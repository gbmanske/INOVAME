//Benchmark atmr_prom1_2672_0.0625

module atmr_prom1(x0, x1, x2, x3, x4, x5, x6, x7, x8, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39;
 wire ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1401_, ori_ori_n1402_, ori_ori_n1403_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, ori_ori_n1407_, ori_ori_n1408_, ori_ori_n1409_, ori_ori_n1410_, ori_ori_n1411_, ori_ori_n1412_, ori_ori_n1413_, ori_ori_n1414_, ori_ori_n1415_, ori_ori_n1416_, ori_ori_n1417_, ori_ori_n1418_, ori_ori_n1419_, ori_ori_n1420_, ori_ori_n1421_, ori_ori_n1422_, ori_ori_n1423_, ori_ori_n1424_, ori_ori_n1425_, ori_ori_n1426_, ori_ori_n1427_, ori_ori_n1428_, ori_ori_n1429_, ori_ori_n1430_, ori_ori_n1431_, ori_ori_n1432_, ori_ori_n1433_, ori_ori_n1434_, ori_ori_n1435_, ori_ori_n1436_, ori_ori_n1437_, ori_ori_n1438_, ori_ori_n1439_, ori_ori_n1440_, ori_ori_n1441_, ori_ori_n1442_, ori_ori_n1443_, ori_ori_n1444_, ori_ori_n1445_, ori_ori_n1446_, ori_ori_n1447_, ori_ori_n1448_, ori_ori_n1449_, ori_ori_n1450_, ori_ori_n1451_, ori_ori_n1452_, ori_ori_n1453_, ori_ori_n1454_, ori_ori_n1455_, ori_ori_n1456_, ori_ori_n1457_, ori_ori_n1458_, ori_ori_n1459_, ori_ori_n1460_, ori_ori_n1461_, ori_ori_n1462_, ori_ori_n1463_, ori_ori_n1464_, ori_ori_n1465_, ori_ori_n1467_, ori_ori_n1468_, ori_ori_n1469_, ori_ori_n1470_, ori_ori_n1471_, ori_ori_n1472_, ori_ori_n1473_, ori_ori_n1474_, ori_ori_n1475_, ori_ori_n1476_, ori_ori_n1477_, ori_ori_n1478_, ori_ori_n1479_, ori_ori_n1480_, ori_ori_n1481_, ori_ori_n1482_, ori_ori_n1483_, ori_ori_n1484_, ori_ori_n1485_, ori_ori_n1486_, ori_ori_n1487_, ori_ori_n1488_, ori_ori_n1489_, ori_ori_n1490_, ori_ori_n1491_, ori_ori_n1492_, ori_ori_n1493_, ori_ori_n1495_, ori_ori_n1496_, ori_ori_n1497_, ori_ori_n1498_, ori_ori_n1499_, ori_ori_n1500_, ori_ori_n1501_, ori_ori_n1502_, ori_ori_n1503_, ori_ori_n1504_, ori_ori_n1505_, ori_ori_n1506_, ori_ori_n1507_, ori_ori_n1508_, ori_ori_n1509_, ori_ori_n1510_, ori_ori_n1511_, ori_ori_n1512_, ori_ori_n1513_, ori_ori_n1514_, ori_ori_n1515_, ori_ori_n1516_, ori_ori_n1517_, ori_ori_n1518_, ori_ori_n1519_, ori_ori_n1520_, ori_ori_n1521_, ori_ori_n1522_, ori_ori_n1523_, ori_ori_n1524_, ori_ori_n1525_, ori_ori_n1526_, ori_ori_n1527_, ori_ori_n1528_, ori_ori_n1529_, ori_ori_n1530_, ori_ori_n1531_, ori_ori_n1532_, ori_ori_n1533_, ori_ori_n1534_, ori_ori_n1535_, ori_ori_n1536_, ori_ori_n1537_, ori_ori_n1538_, ori_ori_n1539_, ori_ori_n1540_, ori_ori_n1541_, ori_ori_n1542_, ori_ori_n1543_, ori_ori_n1544_, ori_ori_n1545_, ori_ori_n1546_, ori_ori_n1547_, ori_ori_n1548_, ori_ori_n1549_, ori_ori_n1550_, ori_ori_n1551_, ori_ori_n1552_, ori_ori_n1553_, ori_ori_n1554_, ori_ori_n1555_, ori_ori_n1556_, ori_ori_n1557_, ori_ori_n1558_, ori_ori_n1559_, ori_ori_n1560_, ori_ori_n1562_, ori_ori_n1563_, ori_ori_n1564_, ori_ori_n1565_, ori_ori_n1566_, ori_ori_n1567_, ori_ori_n1568_, ori_ori_n1569_, ori_ori_n1570_, ori_ori_n1571_, ori_ori_n1572_, ori_ori_n1573_, ori_ori_n1574_, ori_ori_n1575_, ori_ori_n1576_, ori_ori_n1577_, ori_ori_n1578_, ori_ori_n1579_, ori_ori_n1580_, ori_ori_n1581_, ori_ori_n1582_, ori_ori_n1583_, ori_ori_n1584_, ori_ori_n1585_, ori_ori_n1586_, ori_ori_n1587_, ori_ori_n1588_, ori_ori_n1589_, ori_ori_n1590_, ori_ori_n1591_, ori_ori_n1592_, ori_ori_n1593_, ori_ori_n1594_, ori_ori_n1595_, ori_ori_n1596_, ori_ori_n1597_, ori_ori_n1598_, ori_ori_n1599_, ori_ori_n1600_, ori_ori_n1601_, ori_ori_n1602_, ori_ori_n1603_, ori_ori_n1604_, ori_ori_n1605_, ori_ori_n1606_, ori_ori_n1607_, ori_ori_n1608_, ori_ori_n1609_, ori_ori_n1610_, ori_ori_n1611_, ori_ori_n1612_, ori_ori_n1613_, ori_ori_n1614_, ori_ori_n1615_, ori_ori_n1616_, ori_ori_n1617_, ori_ori_n1618_, ori_ori_n1620_, ori_ori_n1621_, ori_ori_n1622_, ori_ori_n1623_, ori_ori_n1624_, ori_ori_n1625_, ori_ori_n1626_, ori_ori_n1627_, ori_ori_n1628_, ori_ori_n1629_, ori_ori_n1630_, ori_ori_n1631_, ori_ori_n1632_, ori_ori_n1633_, ori_ori_n1634_, ori_ori_n1635_, ori_ori_n1636_, ori_ori_n1637_, ori_ori_n1638_, ori_ori_n1639_, ori_ori_n1640_, ori_ori_n1641_, ori_ori_n1642_, ori_ori_n1643_, ori_ori_n1644_, ori_ori_n1645_, ori_ori_n1647_, ori_ori_n1648_, ori_ori_n1649_, ori_ori_n1650_, ori_ori_n1651_, ori_ori_n1652_, ori_ori_n1653_, ori_ori_n1654_, ori_ori_n1655_, ori_ori_n1656_, ori_ori_n1657_, ori_ori_n1658_, ori_ori_n1659_, ori_ori_n1660_, ori_ori_n1661_, ori_ori_n1662_, ori_ori_n1663_, ori_ori_n1664_, ori_ori_n1665_, ori_ori_n1666_, ori_ori_n1667_, ori_ori_n1668_, ori_ori_n1669_, ori_ori_n1670_, ori_ori_n1671_, ori_ori_n1672_, ori_ori_n1673_, ori_ori_n1674_, ori_ori_n1675_, ori_ori_n1676_, ori_ori_n1677_, ori_ori_n1678_, ori_ori_n1679_, ori_ori_n1680_, ori_ori_n1681_, ori_ori_n1682_, ori_ori_n1683_, ori_ori_n1684_, ori_ori_n1685_, ori_ori_n1686_, ori_ori_n1687_, ori_ori_n1688_, ori_ori_n1689_, ori_ori_n1690_, ori_ori_n1691_, ori_ori_n1692_, ori_ori_n1693_, ori_ori_n1694_, ori_ori_n1695_, ori_ori_n1696_, ori_ori_n1697_, ori_ori_n1698_, ori_ori_n1699_, ori_ori_n1700_, ori_ori_n1701_, ori_ori_n1702_, ori_ori_n1703_, ori_ori_n1704_, ori_ori_n1705_, ori_ori_n1706_, ori_ori_n1707_, ori_ori_n1708_, ori_ori_n1709_, ori_ori_n1710_, ori_ori_n1711_, ori_ori_n1712_, ori_ori_n1713_, ori_ori_n1714_, ori_ori_n1715_, ori_ori_n1716_, ori_ori_n1717_, ori_ori_n1718_, ori_ori_n1719_, ori_ori_n1720_, ori_ori_n1721_, ori_ori_n1722_, ori_ori_n1723_, ori_ori_n1724_, ori_ori_n1725_, ori_ori_n1726_, ori_ori_n1727_, ori_ori_n1728_, ori_ori_n1729_, ori_ori_n1730_, ori_ori_n1731_, ori_ori_n1732_, ori_ori_n1734_, ori_ori_n1735_, ori_ori_n1736_, ori_ori_n1737_, ori_ori_n1738_, ori_ori_n1739_, ori_ori_n1740_, ori_ori_n1741_, ori_ori_n1742_, ori_ori_n1743_, ori_ori_n1744_, ori_ori_n1745_, ori_ori_n1746_, ori_ori_n1747_, ori_ori_n1748_, ori_ori_n1749_, ori_ori_n1750_, ori_ori_n1751_, ori_ori_n1752_, ori_ori_n1753_, ori_ori_n1754_, ori_ori_n1755_, ori_ori_n1756_, ori_ori_n1757_, ori_ori_n1758_, ori_ori_n1759_, ori_ori_n1760_, ori_ori_n1761_, ori_ori_n1762_, ori_ori_n1763_, ori_ori_n1764_, ori_ori_n1765_, ori_ori_n1766_, ori_ori_n1767_, ori_ori_n1768_, ori_ori_n1769_, ori_ori_n1770_, ori_ori_n1771_, ori_ori_n1772_, ori_ori_n1773_, ori_ori_n1774_, ori_ori_n1775_, ori_ori_n1776_, ori_ori_n1777_, ori_ori_n1778_, ori_ori_n1779_, ori_ori_n1780_, ori_ori_n1781_, ori_ori_n1782_, ori_ori_n1783_, ori_ori_n1784_, ori_ori_n1785_, ori_ori_n1786_, ori_ori_n1787_, ori_ori_n1788_, ori_ori_n1790_, ori_ori_n1791_, ori_ori_n1792_, ori_ori_n1793_, ori_ori_n1794_, ori_ori_n1795_, ori_ori_n1796_, ori_ori_n1797_, ori_ori_n1798_, ori_ori_n1799_, ori_ori_n1800_, ori_ori_n1801_, ori_ori_n1802_, ori_ori_n1803_, ori_ori_n1804_, ori_ori_n1805_, ori_ori_n1806_, ori_ori_n1808_, ori_ori_n1809_, ori_ori_n1810_, ori_ori_n1811_, ori_ori_n1812_, ori_ori_n1813_, ori_ori_n1814_, ori_ori_n1815_, ori_ori_n1816_, ori_ori_n1817_, ori_ori_n1818_, ori_ori_n1819_, ori_ori_n1820_, ori_ori_n1822_, ori_ori_n1823_, ori_ori_n1824_, ori_ori_n1825_, ori_ori_n1826_, ori_ori_n1827_, ori_ori_n1828_, ori_ori_n1829_, ori_ori_n1830_, ori_ori_n1831_, ori_ori_n1832_, ori_ori_n1833_, ori_ori_n1834_, ori_ori_n1835_, ori_ori_n1836_, ori_ori_n1837_, ori_ori_n1838_, ori_ori_n1840_, ori_ori_n1841_, ori_ori_n1842_, ori_ori_n1843_, ori_ori_n1844_, ori_ori_n1845_, ori_ori_n1846_, ori_ori_n1847_, ori_ori_n1848_, ori_ori_n1849_, ori_ori_n1850_, ori_ori_n1851_, ori_ori_n1852_, ori_ori_n1853_, ori_ori_n1854_, ori_ori_n1855_, ori_ori_n1856_, ori_ori_n1857_, ori_ori_n1858_, ori_ori_n1859_, ori_ori_n1860_, ori_ori_n1861_, ori_ori_n1862_, ori_ori_n1863_, ori_ori_n1864_, ori_ori_n1865_, ori_ori_n1866_, ori_ori_n1867_, ori_ori_n1868_, ori_ori_n1869_, ori_ori_n1870_, ori_ori_n1871_, ori_ori_n1872_, ori_ori_n1873_, ori_ori_n1874_, ori_ori_n1875_, ori_ori_n1876_, ori_ori_n1877_, ori_ori_n1878_, ori_ori_n1879_, ori_ori_n1880_, ori_ori_n1881_, ori_ori_n1882_, ori_ori_n1883_, ori_ori_n1884_, ori_ori_n1885_, ori_ori_n1886_, ori_ori_n1888_, ori_ori_n1889_, ori_ori_n1890_, ori_ori_n1891_, ori_ori_n1892_, ori_ori_n1893_, ori_ori_n1894_, ori_ori_n1895_, ori_ori_n1896_, ori_ori_n1897_, ori_ori_n1898_, ori_ori_n1899_, ori_ori_n1900_, ori_ori_n1901_, ori_ori_n1903_, ori_ori_n1904_, ori_ori_n1905_, ori_ori_n1906_, ori_ori_n1907_, ori_ori_n1908_, ori_ori_n1909_, ori_ori_n1910_, ori_ori_n1911_, ori_ori_n1912_, ori_ori_n1913_, ori_ori_n1914_, ori_ori_n1915_, ori_ori_n1916_, ori_ori_n1917_, ori_ori_n1918_, ori_ori_n1919_, ori_ori_n1920_, ori_ori_n1921_, ori_ori_n1922_, ori_ori_n1923_, ori_ori_n1924_, ori_ori_n1925_, ori_ori_n1926_, ori_ori_n1927_, ori_ori_n1928_, ori_ori_n1929_, ori_ori_n1930_, ori_ori_n1931_, ori_ori_n1932_, ori_ori_n1933_, ori_ori_n1934_, ori_ori_n1935_, ori_ori_n1936_, ori_ori_n1937_, ori_ori_n1938_, ori_ori_n1939_, ori_ori_n1940_, ori_ori_n1941_, ori_ori_n1942_, ori_ori_n1943_, ori_ori_n1944_, ori_ori_n1945_, ori_ori_n1946_, ori_ori_n1947_, ori_ori_n1948_, ori_ori_n1949_, ori_ori_n1950_, ori_ori_n1951_, ori_ori_n1952_, ori_ori_n1953_, ori_ori_n1955_, ori_ori_n1956_, ori_ori_n1957_, ori_ori_n1958_, ori_ori_n1959_, ori_ori_n1960_, ori_ori_n1961_, ori_ori_n1962_, ori_ori_n1963_, ori_ori_n1964_, ori_ori_n1965_, ori_ori_n1966_, ori_ori_n1967_, ori_ori_n1968_, ori_ori_n1969_, ori_ori_n1970_, ori_ori_n1971_, ori_ori_n1972_, ori_ori_n1973_, ori_ori_n1974_, ori_ori_n1975_, ori_ori_n1976_, ori_ori_n1977_, ori_ori_n1978_, ori_ori_n1979_, ori_ori_n1980_, ori_ori_n1981_, ori_ori_n1982_, ori_ori_n1983_, ori_ori_n1984_, ori_ori_n1985_, ori_ori_n1986_, ori_ori_n1987_, ori_ori_n1988_, ori_ori_n1989_, ori_ori_n1990_, ori_ori_n1991_, ori_ori_n1992_, ori_ori_n1993_, ori_ori_n1994_, ori_ori_n1995_, ori_ori_n1996_, ori_ori_n1997_, ori_ori_n1998_, ori_ori_n1999_, ori_ori_n2000_, ori_ori_n2001_, ori_ori_n2002_, ori_ori_n2003_, ori_ori_n2004_, ori_ori_n2005_, ori_ori_n2006_, ori_ori_n2007_, ori_ori_n2008_, ori_ori_n2009_, ori_ori_n2010_, ori_ori_n2011_, ori_ori_n2012_, ori_ori_n2013_, ori_ori_n2014_, ori_ori_n2015_, ori_ori_n2016_, ori_ori_n2017_, ori_ori_n2018_, ori_ori_n2019_, ori_ori_n2020_, ori_ori_n2022_, ori_ori_n2023_, ori_ori_n2024_, ori_ori_n2025_, ori_ori_n2026_, ori_ori_n2027_, ori_ori_n2028_, ori_ori_n2029_, ori_ori_n2030_, ori_ori_n2031_, ori_ori_n2032_, ori_ori_n2033_, ori_ori_n2034_, ori_ori_n2035_, ori_ori_n2036_, ori_ori_n2037_, ori_ori_n2038_, ori_ori_n2039_, ori_ori_n2040_, ori_ori_n2041_, ori_ori_n2042_, ori_ori_n2043_, ori_ori_n2044_, ori_ori_n2045_, ori_ori_n2046_, ori_ori_n2047_, ori_ori_n2048_, ori_ori_n2049_, ori_ori_n2050_, ori_ori_n2051_, ori_ori_n2052_, ori_ori_n2053_, ori_ori_n2054_, ori_ori_n2055_, ori_ori_n2056_, ori_ori_n2057_, ori_ori_n2058_, ori_ori_n2059_, ori_ori_n2060_, ori_ori_n2061_, ori_ori_n2062_, ori_ori_n2063_, ori_ori_n2064_, ori_ori_n2065_, ori_ori_n2066_, ori_ori_n2067_, ori_ori_n2068_, ori_ori_n2069_, ori_ori_n2070_, ori_ori_n2071_, ori_ori_n2072_, ori_ori_n2073_, ori_ori_n2074_, ori_ori_n2075_, ori_ori_n2076_, ori_ori_n2077_, ori_ori_n2078_, ori_ori_n2079_, ori_ori_n2080_, ori_ori_n2081_, ori_ori_n2082_, ori_ori_n2083_, ori_ori_n2084_, ori_ori_n2085_, ori_ori_n2086_, ori_ori_n2087_, ori_ori_n2088_, ori_ori_n2089_, ori_ori_n2090_, ori_ori_n2091_, ori_ori_n2092_, ori_ori_n2093_, ori_ori_n2094_, ori_ori_n2095_, ori_ori_n2096_, ori_ori_n2098_, ori_ori_n2099_, ori_ori_n2100_, ori_ori_n2101_, ori_ori_n2102_, ori_ori_n2103_, ori_ori_n2104_, ori_ori_n2105_, ori_ori_n2106_, ori_ori_n2107_, ori_ori_n2108_, ori_ori_n2109_, ori_ori_n2110_, ori_ori_n2111_, ori_ori_n2112_, ori_ori_n2113_, ori_ori_n2114_, ori_ori_n2115_, ori_ori_n2116_, ori_ori_n2117_, ori_ori_n2118_, ori_ori_n2119_, ori_ori_n2120_, ori_ori_n2121_, ori_ori_n2122_, ori_ori_n2123_, ori_ori_n2124_, ori_ori_n2125_, ori_ori_n2126_, ori_ori_n2127_, ori_ori_n2128_, ori_ori_n2129_, ori_ori_n2130_, ori_ori_n2131_, ori_ori_n2132_, ori_ori_n2133_, ori_ori_n2134_, ori_ori_n2135_, ori_ori_n2136_, ori_ori_n2137_, ori_ori_n2138_, ori_ori_n2139_, ori_ori_n2140_, ori_ori_n2141_, ori_ori_n2142_, ori_ori_n2143_, ori_ori_n2144_, ori_ori_n2145_, ori_ori_n2146_, ori_ori_n2147_, ori_ori_n2148_, ori_ori_n2149_, ori_ori_n2150_, ori_ori_n2151_, ori_ori_n2152_, ori_ori_n2153_, ori_ori_n2154_, ori_ori_n2155_, ori_ori_n2156_, ori_ori_n2157_, ori_ori_n2158_, ori_ori_n2159_, ori_ori_n2160_, ori_ori_n2161_, ori_ori_n2162_, ori_ori_n2163_, ori_ori_n2164_, ori_ori_n2165_, ori_ori_n2166_, ori_ori_n2167_, ori_ori_n2168_, ori_ori_n2169_, ori_ori_n2170_, ori_ori_n2171_, ori_ori_n2172_, ori_ori_n2174_, ori_ori_n2175_, ori_ori_n2176_, ori_ori_n2177_, ori_ori_n2178_, ori_ori_n2179_, ori_ori_n2180_, ori_ori_n2181_, ori_ori_n2182_, ori_ori_n2183_, ori_ori_n2184_, ori_ori_n2185_, ori_ori_n2186_, ori_ori_n2187_, ori_ori_n2188_, ori_ori_n2189_, ori_ori_n2190_, ori_ori_n2191_, ori_ori_n2192_, ori_ori_n2193_, ori_ori_n2194_, ori_ori_n2195_, ori_ori_n2196_, ori_ori_n2197_, ori_ori_n2198_, ori_ori_n2199_, ori_ori_n2200_, ori_ori_n2201_, ori_ori_n2202_, ori_ori_n2203_, ori_ori_n2204_, ori_ori_n2205_, ori_ori_n2206_, ori_ori_n2207_, ori_ori_n2208_, ori_ori_n2209_, ori_ori_n2210_, ori_ori_n2211_, ori_ori_n2212_, ori_ori_n2213_, ori_ori_n2214_, ori_ori_n2215_, ori_ori_n2216_, ori_ori_n2217_, ori_ori_n2218_, ori_ori_n2219_, ori_ori_n2220_, ori_ori_n2221_, ori_ori_n2222_, ori_ori_n2223_, ori_ori_n2224_, ori_ori_n2225_, ori_ori_n2226_, ori_ori_n2227_, ori_ori_n2228_, ori_ori_n2229_, ori_ori_n2230_, ori_ori_n2231_, ori_ori_n2232_, ori_ori_n2233_, ori_ori_n2234_, ori_ori_n2235_, ori_ori_n2236_, ori_ori_n2237_, ori_ori_n2238_, ori_ori_n2239_, ori_ori_n2240_, ori_ori_n2241_, ori_ori_n2242_, ori_ori_n2243_, ori_ori_n2244_, ori_ori_n2245_, ori_ori_n2246_, ori_ori_n2247_, ori_ori_n2248_, ori_ori_n2249_, ori_ori_n2250_, ori_ori_n2251_, ori_ori_n2253_, ori_ori_n2254_, ori_ori_n2255_, ori_ori_n2256_, ori_ori_n2257_, ori_ori_n2258_, ori_ori_n2259_, ori_ori_n2260_, ori_ori_n2261_, ori_ori_n2262_, ori_ori_n2263_, ori_ori_n2264_, ori_ori_n2265_, ori_ori_n2266_, ori_ori_n2267_, ori_ori_n2268_, ori_ori_n2269_, ori_ori_n2270_, ori_ori_n2271_, ori_ori_n2272_, ori_ori_n2273_, ori_ori_n2274_, ori_ori_n2275_, ori_ori_n2276_, ori_ori_n2277_, ori_ori_n2278_, ori_ori_n2279_, ori_ori_n2280_, ori_ori_n2281_, ori_ori_n2282_, ori_ori_n2283_, ori_ori_n2284_, ori_ori_n2285_, ori_ori_n2286_, ori_ori_n2287_, ori_ori_n2288_, ori_ori_n2289_, ori_ori_n2290_, ori_ori_n2291_, ori_ori_n2292_, ori_ori_n2293_, ori_ori_n2294_, ori_ori_n2295_, ori_ori_n2296_, ori_ori_n2297_, ori_ori_n2298_, ori_ori_n2299_, ori_ori_n2300_, ori_ori_n2301_, ori_ori_n2302_, ori_ori_n2303_, ori_ori_n2304_, ori_ori_n2305_, ori_ori_n2306_, ori_ori_n2307_, ori_ori_n2308_, ori_ori_n2309_, ori_ori_n2310_, ori_ori_n2311_, ori_ori_n2312_, ori_ori_n2313_, ori_ori_n2314_, ori_ori_n2315_, ori_ori_n2316_, ori_ori_n2317_, ori_ori_n2318_, ori_ori_n2319_, ori_ori_n2321_, ori_ori_n2322_, ori_ori_n2323_, ori_ori_n2324_, ori_ori_n2325_, ori_ori_n2326_, ori_ori_n2327_, ori_ori_n2328_, ori_ori_n2329_, ori_ori_n2330_, ori_ori_n2331_, ori_ori_n2332_, ori_ori_n2333_, ori_ori_n2334_, ori_ori_n2335_, ori_ori_n2336_, ori_ori_n2337_, ori_ori_n2338_, ori_ori_n2339_, ori_ori_n2340_, ori_ori_n2341_, ori_ori_n2342_, ori_ori_n2343_, ori_ori_n2344_, ori_ori_n2345_, ori_ori_n2346_, ori_ori_n2347_, ori_ori_n2348_, ori_ori_n2349_, ori_ori_n2350_, ori_ori_n2351_, ori_ori_n2352_, ori_ori_n2353_, ori_ori_n2354_, ori_ori_n2355_, ori_ori_n2356_, ori_ori_n2357_, ori_ori_n2358_, ori_ori_n2359_, ori_ori_n2360_, ori_ori_n2361_, ori_ori_n2362_, ori_ori_n2363_, ori_ori_n2364_, ori_ori_n2365_, ori_ori_n2366_, ori_ori_n2367_, ori_ori_n2368_, ori_ori_n2369_, ori_ori_n2370_, ori_ori_n2371_, ori_ori_n2372_, ori_ori_n2373_, ori_ori_n2374_, ori_ori_n2375_, ori_ori_n2376_, ori_ori_n2377_, ori_ori_n2378_, ori_ori_n2379_, ori_ori_n2380_, ori_ori_n2381_, ori_ori_n2383_, ori_ori_n2384_, ori_ori_n2385_, ori_ori_n2386_, ori_ori_n2387_, ori_ori_n2388_, ori_ori_n2389_, ori_ori_n2390_, ori_ori_n2391_, ori_ori_n2392_, ori_ori_n2393_, ori_ori_n2394_, ori_ori_n2395_, ori_ori_n2396_, ori_ori_n2397_, ori_ori_n2398_, ori_ori_n2399_, ori_ori_n2400_, ori_ori_n2401_, ori_ori_n2402_, ori_ori_n2403_, ori_ori_n2404_, ori_ori_n2405_, ori_ori_n2406_, ori_ori_n2407_, ori_ori_n2408_, ori_ori_n2409_, ori_ori_n2410_, ori_ori_n2411_, ori_ori_n2412_, ori_ori_n2413_, ori_ori_n2414_, ori_ori_n2415_, ori_ori_n2416_, ori_ori_n2417_, ori_ori_n2418_, ori_ori_n2419_, ori_ori_n2420_, ori_ori_n2421_, ori_ori_n2422_, ori_ori_n2423_, ori_ori_n2424_, ori_ori_n2425_, ori_ori_n2426_, ori_ori_n2427_, ori_ori_n2428_, ori_ori_n2429_, ori_ori_n2430_, ori_ori_n2431_, ori_ori_n2432_, ori_ori_n2433_, ori_ori_n2434_, ori_ori_n2435_, ori_ori_n2436_, ori_ori_n2437_, ori_ori_n2438_, ori_ori_n2439_, ori_ori_n2440_, ori_ori_n2441_, ori_ori_n2442_, ori_ori_n2443_, ori_ori_n2444_, ori_ori_n2445_, ori_ori_n2446_, ori_ori_n2447_, ori_ori_n2448_, ori_ori_n2449_, ori_ori_n2450_, ori_ori_n2451_, ori_ori_n2452_, ori_ori_n2453_, ori_ori_n2454_, ori_ori_n2455_, ori_ori_n2456_, ori_ori_n2457_, ori_ori_n2458_, ori_ori_n2459_, ori_ori_n2461_, ori_ori_n2462_, ori_ori_n2463_, ori_ori_n2464_, ori_ori_n2465_, ori_ori_n2466_, ori_ori_n2467_, ori_ori_n2468_, ori_ori_n2469_, ori_ori_n2470_, ori_ori_n2471_, ori_ori_n2472_, ori_ori_n2473_, ori_ori_n2474_, ori_ori_n2475_, ori_ori_n2476_, ori_ori_n2477_, ori_ori_n2478_, ori_ori_n2479_, ori_ori_n2480_, ori_ori_n2481_, ori_ori_n2482_, ori_ori_n2483_, ori_ori_n2484_, ori_ori_n2485_, ori_ori_n2486_, ori_ori_n2487_, ori_ori_n2488_, ori_ori_n2489_, ori_ori_n2490_, ori_ori_n2491_, ori_ori_n2492_, ori_ori_n2493_, ori_ori_n2494_, ori_ori_n2495_, ori_ori_n2496_, ori_ori_n2497_, ori_ori_n2498_, ori_ori_n2499_, ori_ori_n2500_, ori_ori_n2501_, ori_ori_n2502_, ori_ori_n2503_, ori_ori_n2504_, ori_ori_n2505_, ori_ori_n2506_, ori_ori_n2507_, ori_ori_n2508_, ori_ori_n2509_, ori_ori_n2510_, ori_ori_n2511_, ori_ori_n2512_, ori_ori_n2513_, ori_ori_n2514_, ori_ori_n2515_, ori_ori_n2516_, ori_ori_n2517_, ori_ori_n2518_, ori_ori_n2519_, ori_ori_n2520_, ori_ori_n2521_, ori_ori_n2522_, ori_ori_n2524_, ori_ori_n2525_, ori_ori_n2526_, ori_ori_n2527_, ori_ori_n2528_, ori_ori_n2529_, ori_ori_n2530_, ori_ori_n2531_, ori_ori_n2532_, ori_ori_n2533_, ori_ori_n2534_, ori_ori_n2535_, ori_ori_n2536_, ori_ori_n2537_, ori_ori_n2538_, ori_ori_n2539_, ori_ori_n2540_, ori_ori_n2541_, ori_ori_n2542_, ori_ori_n2543_, ori_ori_n2544_, ori_ori_n2545_, ori_ori_n2546_, ori_ori_n2547_, ori_ori_n2548_, ori_ori_n2549_, ori_ori_n2550_, ori_ori_n2551_, ori_ori_n2552_, ori_ori_n2553_, ori_ori_n2554_, ori_ori_n2555_, ori_ori_n2556_, ori_ori_n2557_, ori_ori_n2558_, ori_ori_n2559_, ori_ori_n2560_, ori_ori_n2561_, ori_ori_n2562_, ori_ori_n2563_, ori_ori_n2564_, ori_ori_n2565_, ori_ori_n2566_, ori_ori_n2567_, ori_ori_n2568_, ori_ori_n2569_, ori_ori_n2570_, ori_ori_n2571_, ori_ori_n2572_, ori_ori_n2573_, ori_ori_n2574_, ori_ori_n2575_, ori_ori_n2576_, ori_ori_n2577_, ori_ori_n2578_, ori_ori_n2579_, ori_ori_n2580_, ori_ori_n2581_, ori_ori_n2582_, ori_ori_n2583_, ori_ori_n2584_, ori_ori_n2585_, ori_ori_n2586_, ori_ori_n2587_, ori_ori_n2588_, ori_ori_n2589_, ori_ori_n2590_, ori_ori_n2591_, ori_ori_n2592_, ori_ori_n2593_, ori_ori_n2595_, ori_ori_n2596_, ori_ori_n2597_, ori_ori_n2598_, ori_ori_n2599_, ori_ori_n2600_, ori_ori_n2601_, ori_ori_n2602_, ori_ori_n2603_, ori_ori_n2604_, ori_ori_n2605_, ori_ori_n2606_, ori_ori_n2607_, ori_ori_n2608_, ori_ori_n2609_, ori_ori_n2610_, ori_ori_n2611_, ori_ori_n2612_, ori_ori_n2613_, ori_ori_n2614_, ori_ori_n2615_, ori_ori_n2616_, ori_ori_n2617_, ori_ori_n2618_, ori_ori_n2619_, ori_ori_n2620_, ori_ori_n2621_, ori_ori_n2622_, ori_ori_n2623_, ori_ori_n2624_, ori_ori_n2625_, ori_ori_n2626_, ori_ori_n2627_, ori_ori_n2628_, ori_ori_n2629_, ori_ori_n2630_, ori_ori_n2631_, ori_ori_n2632_, ori_ori_n2633_, ori_ori_n2634_, ori_ori_n2635_, ori_ori_n2636_, ori_ori_n2637_, ori_ori_n2638_, ori_ori_n2639_, ori_ori_n2640_, ori_ori_n2641_, ori_ori_n2642_, ori_ori_n2643_, ori_ori_n2644_, ori_ori_n2645_, ori_ori_n2646_, ori_ori_n2647_, ori_ori_n2648_, ori_ori_n2649_, ori_ori_n2650_, ori_ori_n2651_, ori_ori_n2652_, ori_ori_n2653_, ori_ori_n2654_, ori_ori_n2655_, ori_ori_n2656_, ori_ori_n2657_, ori_ori_n2658_, ori_ori_n2659_, ori_ori_n2660_, ori_ori_n2661_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, mai_mai_n1552_, mai_mai_n1553_, mai_mai_n1554_, mai_mai_n1555_, mai_mai_n1556_, mai_mai_n1557_, mai_mai_n1558_, mai_mai_n1559_, mai_mai_n1560_, mai_mai_n1561_, mai_mai_n1562_, mai_mai_n1563_, mai_mai_n1564_, mai_mai_n1565_, mai_mai_n1566_, mai_mai_n1567_, mai_mai_n1568_, mai_mai_n1569_, mai_mai_n1570_, mai_mai_n1571_, mai_mai_n1572_, mai_mai_n1573_, mai_mai_n1575_, mai_mai_n1576_, mai_mai_n1577_, mai_mai_n1578_, mai_mai_n1579_, mai_mai_n1580_, mai_mai_n1581_, mai_mai_n1582_, mai_mai_n1583_, mai_mai_n1584_, mai_mai_n1585_, mai_mai_n1586_, mai_mai_n1587_, mai_mai_n1588_, mai_mai_n1589_, mai_mai_n1590_, mai_mai_n1591_, mai_mai_n1592_, mai_mai_n1593_, mai_mai_n1594_, mai_mai_n1595_, mai_mai_n1596_, mai_mai_n1597_, mai_mai_n1598_, mai_mai_n1599_, mai_mai_n1600_, mai_mai_n1601_, mai_mai_n1602_, mai_mai_n1603_, mai_mai_n1604_, mai_mai_n1605_, mai_mai_n1606_, mai_mai_n1607_, mai_mai_n1608_, mai_mai_n1609_, mai_mai_n1610_, mai_mai_n1611_, mai_mai_n1612_, mai_mai_n1613_, mai_mai_n1614_, mai_mai_n1615_, mai_mai_n1616_, mai_mai_n1617_, mai_mai_n1618_, mai_mai_n1619_, mai_mai_n1620_, mai_mai_n1621_, mai_mai_n1622_, mai_mai_n1623_, mai_mai_n1624_, mai_mai_n1625_, mai_mai_n1626_, mai_mai_n1627_, mai_mai_n1628_, mai_mai_n1629_, mai_mai_n1630_, mai_mai_n1631_, mai_mai_n1633_, mai_mai_n1634_, mai_mai_n1635_, mai_mai_n1636_, mai_mai_n1637_, mai_mai_n1638_, mai_mai_n1639_, mai_mai_n1640_, mai_mai_n1641_, mai_mai_n1642_, mai_mai_n1643_, mai_mai_n1644_, mai_mai_n1645_, mai_mai_n1646_, mai_mai_n1647_, mai_mai_n1648_, mai_mai_n1649_, mai_mai_n1650_, mai_mai_n1651_, mai_mai_n1652_, mai_mai_n1653_, mai_mai_n1654_, mai_mai_n1655_, mai_mai_n1656_, mai_mai_n1657_, mai_mai_n1659_, mai_mai_n1660_, mai_mai_n1661_, mai_mai_n1662_, mai_mai_n1663_, mai_mai_n1664_, mai_mai_n1665_, mai_mai_n1666_, mai_mai_n1667_, mai_mai_n1668_, mai_mai_n1669_, mai_mai_n1670_, mai_mai_n1671_, mai_mai_n1672_, mai_mai_n1673_, mai_mai_n1674_, mai_mai_n1675_, mai_mai_n1676_, mai_mai_n1677_, mai_mai_n1678_, mai_mai_n1679_, mai_mai_n1680_, mai_mai_n1681_, mai_mai_n1682_, mai_mai_n1683_, mai_mai_n1684_, mai_mai_n1685_, mai_mai_n1686_, mai_mai_n1687_, mai_mai_n1688_, mai_mai_n1689_, mai_mai_n1690_, mai_mai_n1691_, mai_mai_n1692_, mai_mai_n1693_, mai_mai_n1694_, mai_mai_n1695_, mai_mai_n1696_, mai_mai_n1697_, mai_mai_n1698_, mai_mai_n1699_, mai_mai_n1700_, mai_mai_n1701_, mai_mai_n1702_, mai_mai_n1703_, mai_mai_n1704_, mai_mai_n1705_, mai_mai_n1706_, mai_mai_n1707_, mai_mai_n1708_, mai_mai_n1709_, mai_mai_n1710_, mai_mai_n1711_, mai_mai_n1712_, mai_mai_n1713_, mai_mai_n1714_, mai_mai_n1715_, mai_mai_n1716_, mai_mai_n1717_, mai_mai_n1718_, mai_mai_n1719_, mai_mai_n1720_, mai_mai_n1721_, mai_mai_n1722_, mai_mai_n1723_, mai_mai_n1724_, mai_mai_n1725_, mai_mai_n1726_, mai_mai_n1727_, mai_mai_n1728_, mai_mai_n1729_, mai_mai_n1730_, mai_mai_n1731_, mai_mai_n1732_, mai_mai_n1733_, mai_mai_n1734_, mai_mai_n1735_, mai_mai_n1736_, mai_mai_n1737_, mai_mai_n1738_, mai_mai_n1739_, mai_mai_n1740_, mai_mai_n1741_, mai_mai_n1742_, mai_mai_n1743_, mai_mai_n1745_, mai_mai_n1746_, mai_mai_n1747_, mai_mai_n1748_, mai_mai_n1749_, mai_mai_n1750_, mai_mai_n1751_, mai_mai_n1752_, mai_mai_n1753_, mai_mai_n1754_, mai_mai_n1755_, mai_mai_n1756_, mai_mai_n1757_, mai_mai_n1758_, mai_mai_n1759_, mai_mai_n1760_, mai_mai_n1761_, mai_mai_n1762_, mai_mai_n1763_, mai_mai_n1764_, mai_mai_n1765_, mai_mai_n1766_, mai_mai_n1767_, mai_mai_n1768_, mai_mai_n1769_, mai_mai_n1770_, mai_mai_n1771_, mai_mai_n1772_, mai_mai_n1773_, mai_mai_n1774_, mai_mai_n1775_, mai_mai_n1776_, mai_mai_n1777_, mai_mai_n1778_, mai_mai_n1779_, mai_mai_n1780_, mai_mai_n1781_, mai_mai_n1782_, mai_mai_n1783_, mai_mai_n1784_, mai_mai_n1785_, mai_mai_n1786_, mai_mai_n1787_, mai_mai_n1788_, mai_mai_n1789_, mai_mai_n1790_, mai_mai_n1791_, mai_mai_n1792_, mai_mai_n1793_, mai_mai_n1794_, mai_mai_n1795_, mai_mai_n1796_, mai_mai_n1797_, mai_mai_n1798_, mai_mai_n1799_, mai_mai_n1800_, mai_mai_n1801_, mai_mai_n1803_, mai_mai_n1804_, mai_mai_n1805_, mai_mai_n1806_, mai_mai_n1807_, mai_mai_n1808_, mai_mai_n1809_, mai_mai_n1810_, mai_mai_n1811_, mai_mai_n1812_, mai_mai_n1813_, mai_mai_n1814_, mai_mai_n1815_, mai_mai_n1816_, mai_mai_n1817_, mai_mai_n1818_, mai_mai_n1819_, mai_mai_n1820_, mai_mai_n1821_, mai_mai_n1823_, mai_mai_n1824_, mai_mai_n1825_, mai_mai_n1826_, mai_mai_n1827_, mai_mai_n1828_, mai_mai_n1829_, mai_mai_n1830_, mai_mai_n1831_, mai_mai_n1832_, mai_mai_n1833_, mai_mai_n1835_, mai_mai_n1836_, mai_mai_n1837_, mai_mai_n1838_, mai_mai_n1839_, mai_mai_n1840_, mai_mai_n1841_, mai_mai_n1842_, mai_mai_n1843_, mai_mai_n1844_, mai_mai_n1845_, mai_mai_n1846_, mai_mai_n1847_, mai_mai_n1848_, mai_mai_n1849_, mai_mai_n1851_, mai_mai_n1852_, mai_mai_n1853_, mai_mai_n1854_, mai_mai_n1855_, mai_mai_n1856_, mai_mai_n1857_, mai_mai_n1858_, mai_mai_n1859_, mai_mai_n1860_, mai_mai_n1861_, mai_mai_n1862_, mai_mai_n1863_, mai_mai_n1864_, mai_mai_n1865_, mai_mai_n1866_, mai_mai_n1867_, mai_mai_n1868_, mai_mai_n1869_, mai_mai_n1870_, mai_mai_n1871_, mai_mai_n1872_, mai_mai_n1873_, mai_mai_n1874_, mai_mai_n1875_, mai_mai_n1876_, mai_mai_n1877_, mai_mai_n1878_, mai_mai_n1879_, mai_mai_n1880_, mai_mai_n1881_, mai_mai_n1882_, mai_mai_n1883_, mai_mai_n1884_, mai_mai_n1885_, mai_mai_n1886_, mai_mai_n1887_, mai_mai_n1888_, mai_mai_n1889_, mai_mai_n1890_, mai_mai_n1891_, mai_mai_n1892_, mai_mai_n1893_, mai_mai_n1894_, mai_mai_n1895_, mai_mai_n1897_, mai_mai_n1898_, mai_mai_n1899_, mai_mai_n1900_, mai_mai_n1901_, mai_mai_n1902_, mai_mai_n1903_, mai_mai_n1904_, mai_mai_n1905_, mai_mai_n1906_, mai_mai_n1907_, mai_mai_n1908_, mai_mai_n1909_, mai_mai_n1910_, mai_mai_n1911_, mai_mai_n1912_, mai_mai_n1914_, mai_mai_n1915_, mai_mai_n1916_, mai_mai_n1917_, mai_mai_n1918_, mai_mai_n1919_, mai_mai_n1920_, mai_mai_n1921_, mai_mai_n1922_, mai_mai_n1923_, mai_mai_n1924_, mai_mai_n1925_, mai_mai_n1926_, mai_mai_n1927_, mai_mai_n1928_, mai_mai_n1929_, mai_mai_n1930_, mai_mai_n1931_, mai_mai_n1932_, mai_mai_n1933_, mai_mai_n1934_, mai_mai_n1935_, mai_mai_n1936_, mai_mai_n1937_, mai_mai_n1938_, mai_mai_n1939_, mai_mai_n1940_, mai_mai_n1941_, mai_mai_n1942_, mai_mai_n1943_, mai_mai_n1944_, mai_mai_n1945_, mai_mai_n1946_, mai_mai_n1947_, mai_mai_n1948_, mai_mai_n1949_, mai_mai_n1950_, mai_mai_n1951_, mai_mai_n1952_, mai_mai_n1953_, mai_mai_n1954_, mai_mai_n1955_, mai_mai_n1956_, mai_mai_n1957_, mai_mai_n1958_, mai_mai_n1959_, mai_mai_n1960_, mai_mai_n1961_, mai_mai_n1962_, mai_mai_n1964_, mai_mai_n1965_, mai_mai_n1966_, mai_mai_n1967_, mai_mai_n1968_, mai_mai_n1969_, mai_mai_n1970_, mai_mai_n1971_, mai_mai_n1972_, mai_mai_n1973_, mai_mai_n1974_, mai_mai_n1975_, mai_mai_n1976_, mai_mai_n1977_, mai_mai_n1978_, mai_mai_n1979_, mai_mai_n1980_, mai_mai_n1981_, mai_mai_n1982_, mai_mai_n1983_, mai_mai_n1984_, mai_mai_n1985_, mai_mai_n1986_, mai_mai_n1987_, mai_mai_n1988_, mai_mai_n1989_, mai_mai_n1990_, mai_mai_n1991_, mai_mai_n1992_, mai_mai_n1993_, mai_mai_n1994_, mai_mai_n1995_, mai_mai_n1996_, mai_mai_n1997_, mai_mai_n1998_, mai_mai_n1999_, mai_mai_n2000_, mai_mai_n2001_, mai_mai_n2002_, mai_mai_n2003_, mai_mai_n2004_, mai_mai_n2005_, mai_mai_n2006_, mai_mai_n2007_, mai_mai_n2008_, mai_mai_n2009_, mai_mai_n2010_, mai_mai_n2011_, mai_mai_n2012_, mai_mai_n2013_, mai_mai_n2014_, mai_mai_n2015_, mai_mai_n2016_, mai_mai_n2017_, mai_mai_n2018_, mai_mai_n2019_, mai_mai_n2020_, mai_mai_n2021_, mai_mai_n2022_, mai_mai_n2023_, mai_mai_n2024_, mai_mai_n2025_, mai_mai_n2026_, mai_mai_n2027_, mai_mai_n2028_, mai_mai_n2029_, mai_mai_n2031_, mai_mai_n2032_, mai_mai_n2033_, mai_mai_n2034_, mai_mai_n2035_, mai_mai_n2036_, mai_mai_n2037_, mai_mai_n2038_, mai_mai_n2039_, mai_mai_n2040_, mai_mai_n2041_, mai_mai_n2042_, mai_mai_n2043_, mai_mai_n2044_, mai_mai_n2045_, mai_mai_n2046_, mai_mai_n2047_, mai_mai_n2048_, mai_mai_n2049_, mai_mai_n2050_, mai_mai_n2051_, mai_mai_n2052_, mai_mai_n2053_, mai_mai_n2054_, mai_mai_n2055_, mai_mai_n2056_, mai_mai_n2057_, mai_mai_n2058_, mai_mai_n2059_, mai_mai_n2060_, mai_mai_n2061_, mai_mai_n2062_, mai_mai_n2063_, mai_mai_n2064_, mai_mai_n2065_, mai_mai_n2066_, mai_mai_n2067_, mai_mai_n2068_, mai_mai_n2069_, mai_mai_n2070_, mai_mai_n2071_, mai_mai_n2072_, mai_mai_n2073_, mai_mai_n2074_, mai_mai_n2075_, mai_mai_n2076_, mai_mai_n2077_, mai_mai_n2078_, mai_mai_n2079_, mai_mai_n2080_, mai_mai_n2081_, mai_mai_n2082_, mai_mai_n2083_, mai_mai_n2084_, mai_mai_n2085_, mai_mai_n2086_, mai_mai_n2087_, mai_mai_n2088_, mai_mai_n2089_, mai_mai_n2090_, mai_mai_n2091_, mai_mai_n2092_, mai_mai_n2093_, mai_mai_n2094_, mai_mai_n2095_, mai_mai_n2096_, mai_mai_n2097_, mai_mai_n2098_, mai_mai_n2099_, mai_mai_n2100_, mai_mai_n2101_, mai_mai_n2102_, mai_mai_n2103_, mai_mai_n2104_, mai_mai_n2105_, mai_mai_n2106_, mai_mai_n2108_, mai_mai_n2109_, mai_mai_n2110_, mai_mai_n2111_, mai_mai_n2112_, mai_mai_n2113_, mai_mai_n2114_, mai_mai_n2115_, mai_mai_n2116_, mai_mai_n2117_, mai_mai_n2118_, mai_mai_n2119_, mai_mai_n2120_, mai_mai_n2121_, mai_mai_n2122_, mai_mai_n2123_, mai_mai_n2124_, mai_mai_n2125_, mai_mai_n2126_, mai_mai_n2127_, mai_mai_n2128_, mai_mai_n2129_, mai_mai_n2130_, mai_mai_n2131_, mai_mai_n2132_, mai_mai_n2133_, mai_mai_n2134_, mai_mai_n2135_, mai_mai_n2136_, mai_mai_n2137_, mai_mai_n2138_, mai_mai_n2139_, mai_mai_n2140_, mai_mai_n2141_, mai_mai_n2142_, mai_mai_n2143_, mai_mai_n2144_, mai_mai_n2145_, mai_mai_n2146_, mai_mai_n2147_, mai_mai_n2148_, mai_mai_n2149_, mai_mai_n2150_, mai_mai_n2151_, mai_mai_n2152_, mai_mai_n2153_, mai_mai_n2154_, mai_mai_n2155_, mai_mai_n2156_, mai_mai_n2157_, mai_mai_n2158_, mai_mai_n2159_, mai_mai_n2160_, mai_mai_n2161_, mai_mai_n2162_, mai_mai_n2163_, mai_mai_n2164_, mai_mai_n2165_, mai_mai_n2166_, mai_mai_n2167_, mai_mai_n2168_, mai_mai_n2169_, mai_mai_n2170_, mai_mai_n2171_, mai_mai_n2172_, mai_mai_n2173_, mai_mai_n2174_, mai_mai_n2175_, mai_mai_n2176_, mai_mai_n2177_, mai_mai_n2178_, mai_mai_n2180_, mai_mai_n2181_, mai_mai_n2182_, mai_mai_n2183_, mai_mai_n2184_, mai_mai_n2185_, mai_mai_n2186_, mai_mai_n2187_, mai_mai_n2188_, mai_mai_n2189_, mai_mai_n2190_, mai_mai_n2191_, mai_mai_n2192_, mai_mai_n2193_, mai_mai_n2194_, mai_mai_n2195_, mai_mai_n2196_, mai_mai_n2197_, mai_mai_n2198_, mai_mai_n2199_, mai_mai_n2200_, mai_mai_n2201_, mai_mai_n2202_, mai_mai_n2203_, mai_mai_n2204_, mai_mai_n2205_, mai_mai_n2206_, mai_mai_n2207_, mai_mai_n2208_, mai_mai_n2209_, mai_mai_n2210_, mai_mai_n2211_, mai_mai_n2212_, mai_mai_n2213_, mai_mai_n2214_, mai_mai_n2215_, mai_mai_n2216_, mai_mai_n2217_, mai_mai_n2218_, mai_mai_n2219_, mai_mai_n2220_, mai_mai_n2221_, mai_mai_n2222_, mai_mai_n2223_, mai_mai_n2224_, mai_mai_n2225_, mai_mai_n2226_, mai_mai_n2227_, mai_mai_n2228_, mai_mai_n2229_, mai_mai_n2230_, mai_mai_n2231_, mai_mai_n2232_, mai_mai_n2233_, mai_mai_n2234_, mai_mai_n2235_, mai_mai_n2236_, mai_mai_n2237_, mai_mai_n2238_, mai_mai_n2239_, mai_mai_n2240_, mai_mai_n2241_, mai_mai_n2242_, mai_mai_n2243_, mai_mai_n2244_, mai_mai_n2245_, mai_mai_n2246_, mai_mai_n2247_, mai_mai_n2248_, mai_mai_n2249_, mai_mai_n2250_, mai_mai_n2251_, mai_mai_n2252_, mai_mai_n2253_, mai_mai_n2254_, mai_mai_n2255_, mai_mai_n2256_, mai_mai_n2258_, mai_mai_n2259_, mai_mai_n2260_, mai_mai_n2261_, mai_mai_n2262_, mai_mai_n2263_, mai_mai_n2264_, mai_mai_n2265_, mai_mai_n2266_, mai_mai_n2267_, mai_mai_n2268_, mai_mai_n2269_, mai_mai_n2270_, mai_mai_n2271_, mai_mai_n2272_, mai_mai_n2273_, mai_mai_n2274_, mai_mai_n2275_, mai_mai_n2276_, mai_mai_n2277_, mai_mai_n2278_, mai_mai_n2279_, mai_mai_n2280_, mai_mai_n2281_, mai_mai_n2282_, mai_mai_n2283_, mai_mai_n2284_, mai_mai_n2285_, mai_mai_n2286_, mai_mai_n2287_, mai_mai_n2288_, mai_mai_n2289_, mai_mai_n2290_, mai_mai_n2291_, mai_mai_n2292_, mai_mai_n2293_, mai_mai_n2294_, mai_mai_n2295_, mai_mai_n2296_, mai_mai_n2297_, mai_mai_n2298_, mai_mai_n2299_, mai_mai_n2300_, mai_mai_n2301_, mai_mai_n2302_, mai_mai_n2303_, mai_mai_n2304_, mai_mai_n2305_, mai_mai_n2306_, mai_mai_n2307_, mai_mai_n2308_, mai_mai_n2309_, mai_mai_n2310_, mai_mai_n2311_, mai_mai_n2312_, mai_mai_n2313_, mai_mai_n2314_, mai_mai_n2315_, mai_mai_n2316_, mai_mai_n2317_, mai_mai_n2318_, mai_mai_n2319_, mai_mai_n2320_, mai_mai_n2321_, mai_mai_n2322_, mai_mai_n2323_, mai_mai_n2324_, mai_mai_n2325_, mai_mai_n2327_, mai_mai_n2328_, mai_mai_n2329_, mai_mai_n2330_, mai_mai_n2331_, mai_mai_n2332_, mai_mai_n2333_, mai_mai_n2334_, mai_mai_n2335_, mai_mai_n2336_, mai_mai_n2337_, mai_mai_n2338_, mai_mai_n2339_, mai_mai_n2340_, mai_mai_n2341_, mai_mai_n2342_, mai_mai_n2343_, mai_mai_n2344_, mai_mai_n2345_, mai_mai_n2346_, mai_mai_n2347_, mai_mai_n2348_, mai_mai_n2349_, mai_mai_n2350_, mai_mai_n2351_, mai_mai_n2352_, mai_mai_n2353_, mai_mai_n2354_, mai_mai_n2355_, mai_mai_n2356_, mai_mai_n2357_, mai_mai_n2358_, mai_mai_n2359_, mai_mai_n2360_, mai_mai_n2361_, mai_mai_n2362_, mai_mai_n2363_, mai_mai_n2364_, mai_mai_n2365_, mai_mai_n2366_, mai_mai_n2367_, mai_mai_n2368_, mai_mai_n2369_, mai_mai_n2370_, mai_mai_n2371_, mai_mai_n2372_, mai_mai_n2373_, mai_mai_n2374_, mai_mai_n2375_, mai_mai_n2376_, mai_mai_n2377_, mai_mai_n2378_, mai_mai_n2379_, mai_mai_n2380_, mai_mai_n2381_, mai_mai_n2382_, mai_mai_n2383_, mai_mai_n2384_, mai_mai_n2385_, mai_mai_n2386_, mai_mai_n2387_, mai_mai_n2388_, mai_mai_n2390_, mai_mai_n2391_, mai_mai_n2392_, mai_mai_n2393_, mai_mai_n2394_, mai_mai_n2395_, mai_mai_n2396_, mai_mai_n2397_, mai_mai_n2398_, mai_mai_n2399_, mai_mai_n2400_, mai_mai_n2401_, mai_mai_n2402_, mai_mai_n2403_, mai_mai_n2404_, mai_mai_n2405_, mai_mai_n2406_, mai_mai_n2407_, mai_mai_n2408_, mai_mai_n2409_, mai_mai_n2410_, mai_mai_n2411_, mai_mai_n2412_, mai_mai_n2413_, mai_mai_n2414_, mai_mai_n2415_, mai_mai_n2416_, mai_mai_n2417_, mai_mai_n2418_, mai_mai_n2419_, mai_mai_n2420_, mai_mai_n2421_, mai_mai_n2422_, mai_mai_n2423_, mai_mai_n2424_, mai_mai_n2425_, mai_mai_n2426_, mai_mai_n2427_, mai_mai_n2428_, mai_mai_n2429_, mai_mai_n2430_, mai_mai_n2431_, mai_mai_n2432_, mai_mai_n2433_, mai_mai_n2434_, mai_mai_n2435_, mai_mai_n2436_, mai_mai_n2437_, mai_mai_n2438_, mai_mai_n2439_, mai_mai_n2440_, mai_mai_n2441_, mai_mai_n2442_, mai_mai_n2443_, mai_mai_n2444_, mai_mai_n2445_, mai_mai_n2446_, mai_mai_n2447_, mai_mai_n2448_, mai_mai_n2449_, mai_mai_n2450_, mai_mai_n2451_, mai_mai_n2452_, mai_mai_n2453_, mai_mai_n2454_, mai_mai_n2455_, mai_mai_n2456_, mai_mai_n2457_, mai_mai_n2458_, mai_mai_n2459_, mai_mai_n2460_, mai_mai_n2461_, mai_mai_n2462_, mai_mai_n2463_, mai_mai_n2464_, mai_mai_n2465_, mai_mai_n2467_, mai_mai_n2468_, mai_mai_n2469_, mai_mai_n2470_, mai_mai_n2471_, mai_mai_n2472_, mai_mai_n2473_, mai_mai_n2474_, mai_mai_n2475_, mai_mai_n2476_, mai_mai_n2477_, mai_mai_n2478_, mai_mai_n2479_, mai_mai_n2480_, mai_mai_n2481_, mai_mai_n2482_, mai_mai_n2483_, mai_mai_n2484_, mai_mai_n2485_, mai_mai_n2486_, mai_mai_n2487_, mai_mai_n2488_, mai_mai_n2489_, mai_mai_n2490_, mai_mai_n2491_, mai_mai_n2492_, mai_mai_n2493_, mai_mai_n2494_, mai_mai_n2495_, mai_mai_n2496_, mai_mai_n2497_, mai_mai_n2498_, mai_mai_n2499_, mai_mai_n2500_, mai_mai_n2501_, mai_mai_n2502_, mai_mai_n2503_, mai_mai_n2504_, mai_mai_n2505_, mai_mai_n2506_, mai_mai_n2507_, mai_mai_n2508_, mai_mai_n2509_, mai_mai_n2510_, mai_mai_n2511_, mai_mai_n2512_, mai_mai_n2513_, mai_mai_n2514_, mai_mai_n2515_, mai_mai_n2516_, mai_mai_n2517_, mai_mai_n2518_, mai_mai_n2519_, mai_mai_n2520_, mai_mai_n2521_, mai_mai_n2522_, mai_mai_n2523_, mai_mai_n2524_, mai_mai_n2525_, mai_mai_n2526_, mai_mai_n2527_, mai_mai_n2529_, mai_mai_n2530_, mai_mai_n2531_, mai_mai_n2532_, mai_mai_n2533_, mai_mai_n2534_, mai_mai_n2535_, mai_mai_n2536_, mai_mai_n2537_, mai_mai_n2538_, mai_mai_n2539_, mai_mai_n2540_, mai_mai_n2541_, mai_mai_n2542_, mai_mai_n2543_, mai_mai_n2544_, mai_mai_n2545_, mai_mai_n2546_, mai_mai_n2547_, mai_mai_n2548_, mai_mai_n2549_, mai_mai_n2550_, mai_mai_n2551_, mai_mai_n2552_, mai_mai_n2553_, mai_mai_n2554_, mai_mai_n2555_, mai_mai_n2556_, mai_mai_n2557_, mai_mai_n2558_, mai_mai_n2559_, mai_mai_n2560_, mai_mai_n2561_, mai_mai_n2562_, mai_mai_n2563_, mai_mai_n2564_, mai_mai_n2565_, mai_mai_n2566_, mai_mai_n2567_, mai_mai_n2568_, mai_mai_n2569_, mai_mai_n2570_, mai_mai_n2571_, mai_mai_n2572_, mai_mai_n2573_, mai_mai_n2574_, mai_mai_n2575_, mai_mai_n2576_, mai_mai_n2577_, mai_mai_n2578_, mai_mai_n2579_, mai_mai_n2580_, mai_mai_n2581_, mai_mai_n2582_, mai_mai_n2583_, mai_mai_n2584_, mai_mai_n2585_, mai_mai_n2586_, mai_mai_n2587_, mai_mai_n2588_, mai_mai_n2589_, mai_mai_n2590_, mai_mai_n2591_, mai_mai_n2592_, mai_mai_n2593_, mai_mai_n2594_, mai_mai_n2595_, mai_mai_n2597_, mai_mai_n2598_, mai_mai_n2599_, mai_mai_n2600_, mai_mai_n2601_, mai_mai_n2602_, mai_mai_n2603_, mai_mai_n2604_, mai_mai_n2605_, mai_mai_n2606_, mai_mai_n2607_, mai_mai_n2608_, mai_mai_n2609_, mai_mai_n2610_, mai_mai_n2611_, mai_mai_n2612_, mai_mai_n2613_, mai_mai_n2614_, mai_mai_n2615_, mai_mai_n2616_, mai_mai_n2617_, mai_mai_n2618_, mai_mai_n2619_, mai_mai_n2620_, mai_mai_n2621_, mai_mai_n2622_, mai_mai_n2623_, mai_mai_n2624_, mai_mai_n2625_, mai_mai_n2626_, mai_mai_n2627_, mai_mai_n2628_, mai_mai_n2629_, mai_mai_n2630_, mai_mai_n2631_, mai_mai_n2632_, mai_mai_n2633_, mai_mai_n2634_, mai_mai_n2635_, mai_mai_n2636_, mai_mai_n2637_, mai_mai_n2638_, mai_mai_n2639_, mai_mai_n2640_, mai_mai_n2641_, mai_mai_n2642_, mai_mai_n2643_, mai_mai_n2644_, mai_mai_n2645_, mai_mai_n2646_, mai_mai_n2647_, mai_mai_n2648_, mai_mai_n2649_, mai_mai_n2650_, mai_mai_n2651_, mai_mai_n2652_, mai_mai_n2653_, mai_mai_n2654_, mai_mai_n2655_, mai_mai_n2656_, mai_mai_n2657_, mai_mai_n2658_, mai_mai_n2659_, mai_mai_n2660_, mai_mai_n2661_, mai_mai_n2662_, mai_mai_n2663_, mai_mai_n2667_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1618_, men_men_n1619_, men_men_n1620_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, men_men_n1632_, men_men_n1633_, men_men_n1635_, men_men_n1636_, men_men_n1637_, men_men_n1638_, men_men_n1639_, men_men_n1640_, men_men_n1641_, men_men_n1642_, men_men_n1643_, men_men_n1644_, men_men_n1645_, men_men_n1646_, men_men_n1647_, men_men_n1648_, men_men_n1649_, men_men_n1650_, men_men_n1651_, men_men_n1652_, men_men_n1653_, men_men_n1654_, men_men_n1655_, men_men_n1656_, men_men_n1657_, men_men_n1658_, men_men_n1660_, men_men_n1661_, men_men_n1662_, men_men_n1663_, men_men_n1664_, men_men_n1665_, men_men_n1666_, men_men_n1667_, men_men_n1668_, men_men_n1669_, men_men_n1670_, men_men_n1671_, men_men_n1672_, men_men_n1673_, men_men_n1674_, men_men_n1675_, men_men_n1676_, men_men_n1677_, men_men_n1678_, men_men_n1679_, men_men_n1680_, men_men_n1681_, men_men_n1682_, men_men_n1683_, men_men_n1684_, men_men_n1685_, men_men_n1686_, men_men_n1687_, men_men_n1688_, men_men_n1689_, men_men_n1690_, men_men_n1691_, men_men_n1692_, men_men_n1693_, men_men_n1694_, men_men_n1695_, men_men_n1696_, men_men_n1697_, men_men_n1698_, men_men_n1699_, men_men_n1700_, men_men_n1701_, men_men_n1702_, men_men_n1703_, men_men_n1704_, men_men_n1705_, men_men_n1706_, men_men_n1707_, men_men_n1708_, men_men_n1709_, men_men_n1710_, men_men_n1711_, men_men_n1712_, men_men_n1713_, men_men_n1714_, men_men_n1715_, men_men_n1716_, men_men_n1717_, men_men_n1718_, men_men_n1719_, men_men_n1720_, men_men_n1721_, men_men_n1722_, men_men_n1723_, men_men_n1724_, men_men_n1725_, men_men_n1726_, men_men_n1727_, men_men_n1728_, men_men_n1729_, men_men_n1730_, men_men_n1731_, men_men_n1732_, men_men_n1733_, men_men_n1734_, men_men_n1735_, men_men_n1736_, men_men_n1737_, men_men_n1738_, men_men_n1739_, men_men_n1740_, men_men_n1741_, men_men_n1742_, men_men_n1743_, men_men_n1744_, men_men_n1745_, men_men_n1747_, men_men_n1748_, men_men_n1749_, men_men_n1750_, men_men_n1751_, men_men_n1752_, men_men_n1753_, men_men_n1754_, men_men_n1755_, men_men_n1756_, men_men_n1757_, men_men_n1758_, men_men_n1759_, men_men_n1760_, men_men_n1761_, men_men_n1762_, men_men_n1763_, men_men_n1764_, men_men_n1765_, men_men_n1766_, men_men_n1767_, men_men_n1768_, men_men_n1769_, men_men_n1770_, men_men_n1771_, men_men_n1772_, men_men_n1773_, men_men_n1774_, men_men_n1775_, men_men_n1776_, men_men_n1777_, men_men_n1778_, men_men_n1779_, men_men_n1780_, men_men_n1781_, men_men_n1782_, men_men_n1783_, men_men_n1784_, men_men_n1785_, men_men_n1786_, men_men_n1787_, men_men_n1788_, men_men_n1789_, men_men_n1790_, men_men_n1791_, men_men_n1792_, men_men_n1793_, men_men_n1794_, men_men_n1795_, men_men_n1796_, men_men_n1797_, men_men_n1798_, men_men_n1799_, men_men_n1800_, men_men_n1801_, men_men_n1802_, men_men_n1804_, men_men_n1805_, men_men_n1806_, men_men_n1807_, men_men_n1808_, men_men_n1809_, men_men_n1810_, men_men_n1811_, men_men_n1812_, men_men_n1813_, men_men_n1814_, men_men_n1815_, men_men_n1816_, men_men_n1817_, men_men_n1818_, men_men_n1819_, men_men_n1820_, men_men_n1821_, men_men_n1822_, men_men_n1824_, men_men_n1825_, men_men_n1826_, men_men_n1827_, men_men_n1828_, men_men_n1829_, men_men_n1830_, men_men_n1831_, men_men_n1832_, men_men_n1833_, men_men_n1834_, men_men_n1835_, men_men_n1836_, men_men_n1838_, men_men_n1839_, men_men_n1840_, men_men_n1841_, men_men_n1842_, men_men_n1843_, men_men_n1844_, men_men_n1845_, men_men_n1846_, men_men_n1847_, men_men_n1848_, men_men_n1849_, men_men_n1850_, men_men_n1851_, men_men_n1852_, men_men_n1853_, men_men_n1854_, men_men_n1856_, men_men_n1857_, men_men_n1858_, men_men_n1859_, men_men_n1860_, men_men_n1861_, men_men_n1862_, men_men_n1863_, men_men_n1864_, men_men_n1865_, men_men_n1866_, men_men_n1867_, men_men_n1868_, men_men_n1869_, men_men_n1870_, men_men_n1871_, men_men_n1872_, men_men_n1873_, men_men_n1874_, men_men_n1875_, men_men_n1876_, men_men_n1877_, men_men_n1878_, men_men_n1879_, men_men_n1880_, men_men_n1881_, men_men_n1882_, men_men_n1883_, men_men_n1884_, men_men_n1885_, men_men_n1886_, men_men_n1887_, men_men_n1888_, men_men_n1889_, men_men_n1890_, men_men_n1891_, men_men_n1892_, men_men_n1893_, men_men_n1894_, men_men_n1895_, men_men_n1896_, men_men_n1897_, men_men_n1898_, men_men_n1899_, men_men_n1900_, men_men_n1901_, men_men_n1902_, men_men_n1904_, men_men_n1905_, men_men_n1906_, men_men_n1907_, men_men_n1908_, men_men_n1909_, men_men_n1910_, men_men_n1911_, men_men_n1912_, men_men_n1913_, men_men_n1914_, men_men_n1915_, men_men_n1916_, men_men_n1917_, men_men_n1918_, men_men_n1919_, men_men_n1921_, men_men_n1922_, men_men_n1923_, men_men_n1924_, men_men_n1925_, men_men_n1926_, men_men_n1927_, men_men_n1928_, men_men_n1929_, men_men_n1930_, men_men_n1931_, men_men_n1932_, men_men_n1933_, men_men_n1934_, men_men_n1935_, men_men_n1936_, men_men_n1937_, men_men_n1938_, men_men_n1939_, men_men_n1940_, men_men_n1941_, men_men_n1942_, men_men_n1943_, men_men_n1944_, men_men_n1945_, men_men_n1946_, men_men_n1947_, men_men_n1948_, men_men_n1949_, men_men_n1950_, men_men_n1951_, men_men_n1952_, men_men_n1953_, men_men_n1954_, men_men_n1955_, men_men_n1956_, men_men_n1957_, men_men_n1958_, men_men_n1959_, men_men_n1960_, men_men_n1961_, men_men_n1962_, men_men_n1963_, men_men_n1964_, men_men_n1965_, men_men_n1966_, men_men_n1967_, men_men_n1968_, men_men_n1969_, men_men_n1970_, men_men_n1971_, men_men_n1973_, men_men_n1974_, men_men_n1975_, men_men_n1976_, men_men_n1977_, men_men_n1978_, men_men_n1979_, men_men_n1980_, men_men_n1981_, men_men_n1982_, men_men_n1983_, men_men_n1984_, men_men_n1985_, men_men_n1986_, men_men_n1987_, men_men_n1988_, men_men_n1989_, men_men_n1990_, men_men_n1991_, men_men_n1992_, men_men_n1993_, men_men_n1994_, men_men_n1995_, men_men_n1996_, men_men_n1997_, men_men_n1998_, men_men_n1999_, men_men_n2000_, men_men_n2001_, men_men_n2002_, men_men_n2003_, men_men_n2004_, men_men_n2005_, men_men_n2006_, men_men_n2007_, men_men_n2008_, men_men_n2009_, men_men_n2010_, men_men_n2011_, men_men_n2012_, men_men_n2013_, men_men_n2014_, men_men_n2015_, men_men_n2016_, men_men_n2017_, men_men_n2018_, men_men_n2019_, men_men_n2020_, men_men_n2021_, men_men_n2022_, men_men_n2023_, men_men_n2024_, men_men_n2025_, men_men_n2026_, men_men_n2027_, men_men_n2028_, men_men_n2029_, men_men_n2030_, men_men_n2031_, men_men_n2032_, men_men_n2033_, men_men_n2034_, men_men_n2035_, men_men_n2036_, men_men_n2037_, men_men_n2038_, men_men_n2040_, men_men_n2041_, men_men_n2042_, men_men_n2043_, men_men_n2044_, men_men_n2045_, men_men_n2046_, men_men_n2047_, men_men_n2048_, men_men_n2049_, men_men_n2050_, men_men_n2051_, men_men_n2052_, men_men_n2053_, men_men_n2054_, men_men_n2055_, men_men_n2056_, men_men_n2057_, men_men_n2058_, men_men_n2059_, men_men_n2060_, men_men_n2061_, men_men_n2062_, men_men_n2063_, men_men_n2064_, men_men_n2065_, men_men_n2066_, men_men_n2067_, men_men_n2068_, men_men_n2069_, men_men_n2070_, men_men_n2071_, men_men_n2072_, men_men_n2073_, men_men_n2074_, men_men_n2075_, men_men_n2076_, men_men_n2077_, men_men_n2078_, men_men_n2079_, men_men_n2080_, men_men_n2081_, men_men_n2082_, men_men_n2083_, men_men_n2084_, men_men_n2085_, men_men_n2086_, men_men_n2087_, men_men_n2088_, men_men_n2089_, men_men_n2090_, men_men_n2091_, men_men_n2092_, men_men_n2093_, men_men_n2094_, men_men_n2095_, men_men_n2096_, men_men_n2097_, men_men_n2098_, men_men_n2099_, men_men_n2100_, men_men_n2101_, men_men_n2102_, men_men_n2103_, men_men_n2104_, men_men_n2105_, men_men_n2106_, men_men_n2107_, men_men_n2108_, men_men_n2109_, men_men_n2110_, men_men_n2111_, men_men_n2112_, men_men_n2113_, men_men_n2114_, men_men_n2116_, men_men_n2117_, men_men_n2118_, men_men_n2119_, men_men_n2120_, men_men_n2121_, men_men_n2122_, men_men_n2123_, men_men_n2124_, men_men_n2125_, men_men_n2126_, men_men_n2127_, men_men_n2128_, men_men_n2129_, men_men_n2130_, men_men_n2131_, men_men_n2132_, men_men_n2133_, men_men_n2134_, men_men_n2135_, men_men_n2136_, men_men_n2137_, men_men_n2138_, men_men_n2139_, men_men_n2140_, men_men_n2141_, men_men_n2142_, men_men_n2143_, men_men_n2144_, men_men_n2145_, men_men_n2146_, men_men_n2147_, men_men_n2148_, men_men_n2149_, men_men_n2150_, men_men_n2151_, men_men_n2152_, men_men_n2153_, men_men_n2154_, men_men_n2155_, men_men_n2156_, men_men_n2157_, men_men_n2158_, men_men_n2159_, men_men_n2160_, men_men_n2161_, men_men_n2162_, men_men_n2163_, men_men_n2164_, men_men_n2165_, men_men_n2166_, men_men_n2167_, men_men_n2168_, men_men_n2169_, men_men_n2170_, men_men_n2171_, men_men_n2172_, men_men_n2173_, men_men_n2174_, men_men_n2175_, men_men_n2176_, men_men_n2177_, men_men_n2178_, men_men_n2179_, men_men_n2180_, men_men_n2181_, men_men_n2182_, men_men_n2183_, men_men_n2184_, men_men_n2185_, men_men_n2186_, men_men_n2187_, men_men_n2188_, men_men_n2189_, men_men_n2190_, men_men_n2192_, men_men_n2193_, men_men_n2194_, men_men_n2195_, men_men_n2196_, men_men_n2197_, men_men_n2198_, men_men_n2199_, men_men_n2200_, men_men_n2201_, men_men_n2202_, men_men_n2203_, men_men_n2204_, men_men_n2205_, men_men_n2206_, men_men_n2207_, men_men_n2208_, men_men_n2209_, men_men_n2210_, men_men_n2211_, men_men_n2212_, men_men_n2213_, men_men_n2214_, men_men_n2215_, men_men_n2216_, men_men_n2217_, men_men_n2218_, men_men_n2219_, men_men_n2220_, men_men_n2221_, men_men_n2222_, men_men_n2223_, men_men_n2224_, men_men_n2225_, men_men_n2226_, men_men_n2227_, men_men_n2228_, men_men_n2229_, men_men_n2230_, men_men_n2231_, men_men_n2232_, men_men_n2233_, men_men_n2234_, men_men_n2235_, men_men_n2236_, men_men_n2237_, men_men_n2238_, men_men_n2239_, men_men_n2240_, men_men_n2241_, men_men_n2242_, men_men_n2243_, men_men_n2244_, men_men_n2245_, men_men_n2246_, men_men_n2247_, men_men_n2248_, men_men_n2249_, men_men_n2250_, men_men_n2251_, men_men_n2252_, men_men_n2253_, men_men_n2254_, men_men_n2255_, men_men_n2256_, men_men_n2257_, men_men_n2258_, men_men_n2259_, men_men_n2260_, men_men_n2261_, men_men_n2262_, men_men_n2263_, men_men_n2264_, men_men_n2265_, men_men_n2266_, men_men_n2267_, men_men_n2268_, men_men_n2269_, men_men_n2271_, men_men_n2272_, men_men_n2273_, men_men_n2274_, men_men_n2275_, men_men_n2276_, men_men_n2277_, men_men_n2278_, men_men_n2279_, men_men_n2280_, men_men_n2281_, men_men_n2282_, men_men_n2283_, men_men_n2284_, men_men_n2285_, men_men_n2286_, men_men_n2287_, men_men_n2288_, men_men_n2289_, men_men_n2290_, men_men_n2291_, men_men_n2292_, men_men_n2293_, men_men_n2294_, men_men_n2295_, men_men_n2296_, men_men_n2297_, men_men_n2298_, men_men_n2299_, men_men_n2300_, men_men_n2301_, men_men_n2302_, men_men_n2303_, men_men_n2304_, men_men_n2305_, men_men_n2306_, men_men_n2307_, men_men_n2308_, men_men_n2309_, men_men_n2310_, men_men_n2311_, men_men_n2312_, men_men_n2313_, men_men_n2314_, men_men_n2315_, men_men_n2316_, men_men_n2317_, men_men_n2318_, men_men_n2319_, men_men_n2320_, men_men_n2321_, men_men_n2322_, men_men_n2323_, men_men_n2324_, men_men_n2325_, men_men_n2326_, men_men_n2327_, men_men_n2328_, men_men_n2329_, men_men_n2330_, men_men_n2331_, men_men_n2332_, men_men_n2333_, men_men_n2334_, men_men_n2335_, men_men_n2336_, men_men_n2338_, men_men_n2339_, men_men_n2340_, men_men_n2341_, men_men_n2342_, men_men_n2343_, men_men_n2344_, men_men_n2345_, men_men_n2346_, men_men_n2347_, men_men_n2348_, men_men_n2349_, men_men_n2350_, men_men_n2351_, men_men_n2352_, men_men_n2353_, men_men_n2354_, men_men_n2355_, men_men_n2356_, men_men_n2357_, men_men_n2358_, men_men_n2359_, men_men_n2360_, men_men_n2361_, men_men_n2362_, men_men_n2363_, men_men_n2364_, men_men_n2365_, men_men_n2366_, men_men_n2367_, men_men_n2368_, men_men_n2369_, men_men_n2370_, men_men_n2371_, men_men_n2372_, men_men_n2373_, men_men_n2374_, men_men_n2375_, men_men_n2376_, men_men_n2377_, men_men_n2378_, men_men_n2379_, men_men_n2380_, men_men_n2381_, men_men_n2382_, men_men_n2383_, men_men_n2384_, men_men_n2385_, men_men_n2386_, men_men_n2387_, men_men_n2388_, men_men_n2389_, men_men_n2390_, men_men_n2391_, men_men_n2392_, men_men_n2393_, men_men_n2394_, men_men_n2395_, men_men_n2396_, men_men_n2397_, men_men_n2399_, men_men_n2400_, men_men_n2401_, men_men_n2402_, men_men_n2403_, men_men_n2404_, men_men_n2405_, men_men_n2406_, men_men_n2407_, men_men_n2408_, men_men_n2409_, men_men_n2410_, men_men_n2411_, men_men_n2412_, men_men_n2413_, men_men_n2414_, men_men_n2415_, men_men_n2416_, men_men_n2417_, men_men_n2418_, men_men_n2419_, men_men_n2420_, men_men_n2421_, men_men_n2422_, men_men_n2423_, men_men_n2424_, men_men_n2425_, men_men_n2426_, men_men_n2427_, men_men_n2428_, men_men_n2429_, men_men_n2430_, men_men_n2431_, men_men_n2432_, men_men_n2433_, men_men_n2434_, men_men_n2435_, men_men_n2436_, men_men_n2437_, men_men_n2438_, men_men_n2439_, men_men_n2440_, men_men_n2441_, men_men_n2442_, men_men_n2443_, men_men_n2444_, men_men_n2445_, men_men_n2446_, men_men_n2447_, men_men_n2448_, men_men_n2449_, men_men_n2450_, men_men_n2451_, men_men_n2452_, men_men_n2453_, men_men_n2454_, men_men_n2455_, men_men_n2456_, men_men_n2457_, men_men_n2458_, men_men_n2459_, men_men_n2460_, men_men_n2461_, men_men_n2462_, men_men_n2463_, men_men_n2464_, men_men_n2465_, men_men_n2466_, men_men_n2467_, men_men_n2468_, men_men_n2469_, men_men_n2470_, men_men_n2471_, men_men_n2472_, men_men_n2473_, men_men_n2474_, men_men_n2475_, men_men_n2477_, men_men_n2478_, men_men_n2479_, men_men_n2480_, men_men_n2481_, men_men_n2482_, men_men_n2483_, men_men_n2484_, men_men_n2485_, men_men_n2486_, men_men_n2487_, men_men_n2488_, men_men_n2489_, men_men_n2490_, men_men_n2491_, men_men_n2492_, men_men_n2493_, men_men_n2494_, men_men_n2495_, men_men_n2496_, men_men_n2497_, men_men_n2498_, men_men_n2499_, men_men_n2500_, men_men_n2501_, men_men_n2502_, men_men_n2503_, men_men_n2504_, men_men_n2505_, men_men_n2506_, men_men_n2507_, men_men_n2508_, men_men_n2509_, men_men_n2510_, men_men_n2511_, men_men_n2512_, men_men_n2513_, men_men_n2514_, men_men_n2515_, men_men_n2516_, men_men_n2517_, men_men_n2518_, men_men_n2519_, men_men_n2520_, men_men_n2521_, men_men_n2522_, men_men_n2523_, men_men_n2524_, men_men_n2525_, men_men_n2526_, men_men_n2527_, men_men_n2528_, men_men_n2529_, men_men_n2530_, men_men_n2531_, men_men_n2532_, men_men_n2533_, men_men_n2534_, men_men_n2535_, men_men_n2536_, men_men_n2537_, men_men_n2538_, men_men_n2539_, men_men_n2541_, men_men_n2542_, men_men_n2543_, men_men_n2544_, men_men_n2545_, men_men_n2546_, men_men_n2547_, men_men_n2548_, men_men_n2549_, men_men_n2550_, men_men_n2551_, men_men_n2552_, men_men_n2553_, men_men_n2554_, men_men_n2555_, men_men_n2556_, men_men_n2557_, men_men_n2558_, men_men_n2559_, men_men_n2560_, men_men_n2561_, men_men_n2562_, men_men_n2563_, men_men_n2564_, men_men_n2565_, men_men_n2566_, men_men_n2567_, men_men_n2568_, men_men_n2569_, men_men_n2570_, men_men_n2571_, men_men_n2572_, men_men_n2573_, men_men_n2574_, men_men_n2575_, men_men_n2576_, men_men_n2577_, men_men_n2578_, men_men_n2579_, men_men_n2580_, men_men_n2581_, men_men_n2582_, men_men_n2583_, men_men_n2584_, men_men_n2585_, men_men_n2586_, men_men_n2587_, men_men_n2588_, men_men_n2589_, men_men_n2590_, men_men_n2591_, men_men_n2592_, men_men_n2593_, men_men_n2594_, men_men_n2595_, men_men_n2596_, men_men_n2597_, men_men_n2598_, men_men_n2599_, men_men_n2600_, men_men_n2601_, men_men_n2602_, men_men_n2603_, men_men_n2604_, men_men_n2605_, men_men_n2607_, men_men_n2608_, men_men_n2609_, men_men_n2610_, men_men_n2611_, men_men_n2612_, men_men_n2613_, men_men_n2614_, men_men_n2615_, men_men_n2616_, men_men_n2617_, men_men_n2618_, men_men_n2619_, men_men_n2620_, men_men_n2621_, men_men_n2622_, men_men_n2623_, men_men_n2624_, men_men_n2625_, men_men_n2626_, men_men_n2627_, men_men_n2628_, men_men_n2629_, men_men_n2630_, men_men_n2631_, men_men_n2632_, men_men_n2633_, men_men_n2634_, men_men_n2635_, men_men_n2636_, men_men_n2637_, men_men_n2638_, men_men_n2639_, men_men_n2640_, men_men_n2641_, men_men_n2642_, men_men_n2643_, men_men_n2644_, men_men_n2645_, men_men_n2646_, men_men_n2647_, men_men_n2648_, men_men_n2649_, men_men_n2650_, men_men_n2651_, men_men_n2652_, men_men_n2653_, men_men_n2654_, men_men_n2655_, men_men_n2656_, men_men_n2657_, men_men_n2658_, men_men_n2659_, men_men_n2660_, men_men_n2661_, men_men_n2662_, men_men_n2663_, men_men_n2664_, men_men_n2665_, men_men_n2666_, men_men_n2667_, men_men_n2668_, men_men_n2669_, men_men_n2670_, men_men_n2671_, men_men_n2672_, men_men_n2676_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13, ori14, mai14, men14, ori15, mai15, men15, ori16, mai16, men16, ori17, mai17, men17, ori18, mai18, men18, ori19, mai19, men19, ori20, mai20, men20, ori21, mai21, men21, ori22, mai22, men22, ori23, mai23, men23, ori24, mai24, men24, ori25, mai25, men25, ori26, mai26, men26, ori27, mai27, men27, ori28, mai28, men28, ori29, mai29, men29, ori30, mai30, men30, ori31, mai31, men31, ori32, mai32, men32, ori33, mai33, men33, ori34, mai34, men34, ori35, mai35, men35, ori36, mai36, men36, ori37, mai37, men37, ori38, mai38, men38, ori39, mai39, men39;
  INV        o0000(.A(x3), .Y(ori_ori_n50_));
  NA2        o0001(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n51_));
  NA2        o0002(.A(x7), .B(x0), .Y(ori_ori_n52_));
  INV        o0003(.A(x1), .Y(ori_ori_n53_));
  NA2        o0004(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o0005(.A(x8), .Y(ori_ori_n55_));
  INV        o0006(.A(x4), .Y(ori_ori_n56_));
  INV        o0007(.A(x7), .Y(ori_ori_n57_));
  NA2        o0008(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0009(.A(x0), .Y(ori_ori_n59_));
  NA2        o0010(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NA4        o0011(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n55_), .D(x6), .Y(ori_ori_n61_));
  NA2        o0012(.A(ori_ori_n56_), .B(ori_ori_n59_), .Y(ori_ori_n62_));
  NO2        o0013(.A(ori_ori_n55_), .B(x6), .Y(ori_ori_n63_));
  NA2        o0014(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n64_));
  NA3        o0015(.A(ori_ori_n64_), .B(ori_ori_n63_), .C(ori_ori_n62_), .Y(ori_ori_n65_));
  AOI210     o0016(.A0(ori_ori_n65_), .A1(ori_ori_n61_), .B0(ori_ori_n54_), .Y(ori_ori_n66_));
  NO2        o0017(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n67_));
  NO2        o0018(.A(x7), .B(ori_ori_n59_), .Y(ori_ori_n68_));
  NO2        o0019(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  NAi21      o0020(.An(x5), .B(x1), .Y(ori_ori_n70_));
  INV        o0021(.A(x6), .Y(ori_ori_n71_));
  NA2        o0022(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NO3        o0023(.A(ori_ori_n72_), .B(ori_ori_n70_), .C(ori_ori_n69_), .Y(ori_ori_n73_));
  OAI210     o0024(.A0(ori_ori_n73_), .A1(ori_ori_n66_), .B0(ori_ori_n52_), .Y(ori_ori_n74_));
  NA2        o0025(.A(x7), .B(x4), .Y(ori_ori_n75_));
  NO2        o0026(.A(ori_ori_n75_), .B(x1), .Y(ori_ori_n76_));
  NO2        o0027(.A(ori_ori_n71_), .B(x5), .Y(ori_ori_n77_));
  NO2        o0028(.A(x8), .B(ori_ori_n59_), .Y(ori_ori_n78_));
  NA3        o0029(.A(ori_ori_n78_), .B(ori_ori_n77_), .C(ori_ori_n76_), .Y(ori_ori_n79_));
  AOI210     o0030(.A0(ori_ori_n79_), .A1(ori_ori_n74_), .B0(ori_ori_n51_), .Y(ori_ori_n80_));
  NA2        o0031(.A(x5), .B(x3), .Y(ori_ori_n81_));
  NO2        o0032(.A(x6), .B(x0), .Y(ori_ori_n82_));
  NO2        o0033(.A(ori_ori_n82_), .B(x4), .Y(ori_ori_n83_));
  NO2        o0034(.A(x4), .B(x2), .Y(ori_ori_n84_));
  NO2        o0035(.A(ori_ori_n71_), .B(ori_ori_n59_), .Y(ori_ori_n85_));
  NO2        o0036(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  NA2        o0037(.A(x8), .B(x1), .Y(ori_ori_n87_));
  NO2        o0038(.A(ori_ori_n87_), .B(x7), .Y(ori_ori_n88_));
  NO3        o0039(.A(x8), .B(ori_ori_n57_), .C(x6), .Y(ori_ori_n89_));
  NO2        o0040(.A(x1), .B(ori_ori_n59_), .Y(ori_ori_n90_));
  NO2        o0041(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n91_));
  XO2        o0042(.A(x7), .B(x1), .Y(ori_ori_n92_));
  INV        o0043(.A(ori_ori_n92_), .Y(ori_ori_n93_));
  NO2        o0044(.A(ori_ori_n93_), .B(x6), .Y(ori_ori_n94_));
  NO2        o0045(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n95_));
  NA2        o0046(.A(ori_ori_n95_), .B(ori_ori_n55_), .Y(ori_ori_n96_));
  NO2        o0047(.A(x6), .B(x5), .Y(ori_ori_n97_));
  NO2        o0048(.A(ori_ori_n57_), .B(x5), .Y(ori_ori_n98_));
  NO2        o0049(.A(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  NA2        o0050(.A(x6), .B(x1), .Y(ori_ori_n100_));
  NA2        o0051(.A(ori_ori_n100_), .B(ori_ori_n84_), .Y(ori_ori_n101_));
  NO4        o0052(.A(ori_ori_n101_), .B(ori_ori_n99_), .C(ori_ori_n96_), .D(ori_ori_n94_), .Y(ori_ori_n102_));
  NA2        o0053(.A(x3), .B(x0), .Y(ori_ori_n103_));
  INV        o0054(.A(x5), .Y(ori_ori_n104_));
  NA2        o0055(.A(ori_ori_n71_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  INV        o0056(.A(x2), .Y(ori_ori_n106_));
  NO2        o0057(.A(ori_ori_n56_), .B(ori_ori_n106_), .Y(ori_ori_n107_));
  NA2        o0058(.A(ori_ori_n57_), .B(ori_ori_n104_), .Y(ori_ori_n108_));
  NA3        o0059(.A(ori_ori_n108_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n109_));
  NO3        o0060(.A(ori_ori_n109_), .B(ori_ori_n103_), .C(ori_ori_n53_), .Y(ori_ori_n110_));
  NO3        o0061(.A(ori_ori_n110_), .B(ori_ori_n102_), .C(ori_ori_n80_), .Y(ori00));
  NO2        o0062(.A(x7), .B(x6), .Y(ori_ori_n112_));
  INV        o0063(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NO2        o0064(.A(ori_ori_n55_), .B(ori_ori_n53_), .Y(ori_ori_n114_));
  NA2        o0065(.A(ori_ori_n114_), .B(ori_ori_n56_), .Y(ori_ori_n115_));
  NO2        o0066(.A(ori_ori_n115_), .B(ori_ori_n113_), .Y(ori_ori_n116_));
  XN2        o0067(.A(x6), .B(x1), .Y(ori_ori_n117_));
  INV        o0068(.A(ori_ori_n117_), .Y(ori_ori_n118_));
  NO2        o0069(.A(x6), .B(x4), .Y(ori_ori_n119_));
  NA2        o0070(.A(x6), .B(x4), .Y(ori_ori_n120_));
  NAi21      o0071(.An(ori_ori_n119_), .B(ori_ori_n120_), .Y(ori_ori_n121_));
  XN2        o0072(.A(x7), .B(x6), .Y(ori_ori_n122_));
  NO4        o0073(.A(ori_ori_n122_), .B(ori_ori_n121_), .C(ori_ori_n118_), .D(x8), .Y(ori_ori_n123_));
  NO2        o0074(.A(x3), .B(ori_ori_n106_), .Y(ori_ori_n124_));
  NA2        o0075(.A(ori_ori_n124_), .B(ori_ori_n104_), .Y(ori_ori_n125_));
  NO2        o0076(.A(ori_ori_n125_), .B(ori_ori_n59_), .Y(ori_ori_n126_));
  OAI210     o0077(.A0(ori_ori_n123_), .A1(ori_ori_n116_), .B0(ori_ori_n126_), .Y(ori_ori_n127_));
  NA2        o0078(.A(x3), .B(ori_ori_n106_), .Y(ori_ori_n128_));
  NO2        o0079(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n129_));
  NA2        o0080(.A(ori_ori_n129_), .B(ori_ori_n56_), .Y(ori_ori_n130_));
  NA2        o0081(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n131_));
  NA2        o0082(.A(ori_ori_n131_), .B(x2), .Y(ori_ori_n132_));
  NA2        o0083(.A(x8), .B(x3), .Y(ori_ori_n133_));
  NA2        o0084(.A(ori_ori_n133_), .B(ori_ori_n75_), .Y(ori_ori_n134_));
  OAI220     o0085(.A0(ori_ori_n134_), .A1(ori_ori_n132_), .B0(ori_ori_n130_), .B1(ori_ori_n128_), .Y(ori_ori_n135_));
  NO2        o0086(.A(x5), .B(x0), .Y(ori_ori_n136_));
  NO2        o0087(.A(x6), .B(x1), .Y(ori_ori_n137_));
  NA3        o0088(.A(ori_ori_n137_), .B(ori_ori_n136_), .C(ori_ori_n135_), .Y(ori_ori_n138_));
  NA2        o0089(.A(x8), .B(ori_ori_n104_), .Y(ori_ori_n139_));
  NA2        o0090(.A(x4), .B(ori_ori_n50_), .Y(ori_ori_n140_));
  NO3        o0091(.A(ori_ori_n140_), .B(ori_ori_n139_), .C(ori_ori_n100_), .Y(ori_ori_n141_));
  NAi21      o0092(.An(x7), .B(x2), .Y(ori_ori_n142_));
  NO2        o0093(.A(ori_ori_n142_), .B(x0), .Y(ori_ori_n143_));
  XO2        o0094(.A(x8), .B(x7), .Y(ori_ori_n144_));
  NA2        o0095(.A(ori_ori_n144_), .B(ori_ori_n106_), .Y(ori_ori_n145_));
  NA2        o0096(.A(x6), .B(x5), .Y(ori_ori_n146_));
  NO2        o0097(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n147_));
  NO2        o0098(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n148_));
  NA2        o0099(.A(ori_ori_n148_), .B(ori_ori_n147_), .Y(ori_ori_n149_));
  NO3        o0100(.A(ori_ori_n149_), .B(ori_ori_n146_), .C(ori_ori_n145_), .Y(ori_ori_n150_));
  AOI210     o0101(.A0(ori_ori_n143_), .A1(ori_ori_n141_), .B0(ori_ori_n150_), .Y(ori_ori_n151_));
  NA3        o0102(.A(ori_ori_n151_), .B(ori_ori_n138_), .C(ori_ori_n127_), .Y(ori01));
  NA2        o0103(.A(ori_ori_n57_), .B(ori_ori_n59_), .Y(ori_ori_n153_));
  NO2        o0104(.A(x2), .B(x1), .Y(ori_ori_n154_));
  NA2        o0105(.A(x2), .B(x1), .Y(ori_ori_n155_));
  NOi21      o0106(.An(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NA2        o0107(.A(ori_ori_n104_), .B(ori_ori_n53_), .Y(ori_ori_n157_));
  NO2        o0108(.A(ori_ori_n157_), .B(x8), .Y(ori_ori_n158_));
  NAi21      o0109(.An(x8), .B(x1), .Y(ori_ori_n159_));
  NO2        o0110(.A(ori_ori_n159_), .B(x3), .Y(ori_ori_n160_));
  OAI210     o0111(.A0(ori_ori_n160_), .A1(ori_ori_n158_), .B0(ori_ori_n156_), .Y(ori_ori_n161_));
  NO2        o0112(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n162_));
  NO2        o0113(.A(ori_ori_n106_), .B(x1), .Y(ori_ori_n163_));
  NA2        o0114(.A(ori_ori_n163_), .B(ori_ori_n162_), .Y(ori_ori_n164_));
  AOI210     o0115(.A0(ori_ori_n164_), .A1(ori_ori_n161_), .B0(ori_ori_n153_), .Y(ori_ori_n165_));
  NAi21      o0116(.An(x7), .B(x0), .Y(ori_ori_n166_));
  NO2        o0117(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n167_));
  NO2        o0118(.A(ori_ori_n81_), .B(x1), .Y(ori_ori_n168_));
  NA2        o0119(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n169_));
  NO2        o0120(.A(ori_ori_n169_), .B(ori_ori_n159_), .Y(ori_ori_n170_));
  NA2        o0121(.A(x8), .B(x5), .Y(ori_ori_n171_));
  NO3        o0122(.A(x3), .B(ori_ori_n106_), .C(ori_ori_n53_), .Y(ori_ori_n172_));
  NO2        o0123(.A(ori_ori_n172_), .B(ori_ori_n170_), .Y(ori_ori_n173_));
  NO2        o0124(.A(ori_ori_n173_), .B(ori_ori_n166_), .Y(ori_ori_n174_));
  NO2        o0125(.A(ori_ori_n57_), .B(x3), .Y(ori_ori_n175_));
  NO2        o0126(.A(ori_ori_n55_), .B(x0), .Y(ori_ori_n176_));
  NA3        o0127(.A(ori_ori_n104_), .B(ori_ori_n106_), .C(x1), .Y(ori_ori_n177_));
  NO2        o0128(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  NO2        o0129(.A(ori_ori_n87_), .B(ori_ori_n50_), .Y(ori_ori_n179_));
  NA2        o0130(.A(ori_ori_n104_), .B(x0), .Y(ori_ori_n180_));
  NA2        o0131(.A(ori_ori_n178_), .B(ori_ori_n175_), .Y(ori_ori_n181_));
  NA2        o0132(.A(x7), .B(ori_ori_n106_), .Y(ori_ori_n182_));
  NA2        o0133(.A(ori_ori_n162_), .B(x8), .Y(ori_ori_n183_));
  NA4        o0134(.A(x5), .B(x3), .C(x1), .D(x0), .Y(ori_ori_n184_));
  AO210      o0135(.A0(ori_ori_n184_), .A1(ori_ori_n183_), .B0(ori_ori_n182_), .Y(ori_ori_n185_));
  NO2        o0136(.A(ori_ori_n155_), .B(ori_ori_n50_), .Y(ori_ori_n186_));
  NAi21      o0137(.An(x1), .B(x2), .Y(ori_ori_n187_));
  NO2        o0138(.A(ori_ori_n169_), .B(ori_ori_n187_), .Y(ori_ori_n188_));
  NA2        o0139(.A(x8), .B(x7), .Y(ori_ori_n189_));
  NO2        o0140(.A(ori_ori_n189_), .B(x0), .Y(ori_ori_n190_));
  OAI210     o0141(.A0(ori_ori_n188_), .A1(ori_ori_n186_), .B0(ori_ori_n190_), .Y(ori_ori_n191_));
  NA3        o0142(.A(ori_ori_n191_), .B(ori_ori_n185_), .C(ori_ori_n181_), .Y(ori_ori_n192_));
  NO3        o0143(.A(ori_ori_n192_), .B(ori_ori_n174_), .C(ori_ori_n165_), .Y(ori_ori_n193_));
  NA2        o0144(.A(x3), .B(x1), .Y(ori_ori_n194_));
  NA2        o0145(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n195_));
  NO2        o0146(.A(ori_ori_n195_), .B(ori_ori_n70_), .Y(ori_ori_n196_));
  OAI210     o0147(.A0(ori_ori_n196_), .A1(ori_ori_n188_), .B0(ori_ori_n67_), .Y(ori_ori_n197_));
  NA2        o0148(.A(ori_ori_n129_), .B(ori_ori_n106_), .Y(ori_ori_n198_));
  OAI210     o0149(.A0(ori_ori_n198_), .A1(ori_ori_n194_), .B0(ori_ori_n197_), .Y(ori_ori_n199_));
  XO2        o0150(.A(x5), .B(x3), .Y(ori_ori_n200_));
  NA2        o0151(.A(ori_ori_n200_), .B(x8), .Y(ori_ori_n201_));
  NA2        o0152(.A(x8), .B(ori_ori_n59_), .Y(ori_ori_n202_));
  NA2        o0153(.A(ori_ori_n202_), .B(ori_ori_n133_), .Y(ori_ori_n203_));
  NA2        o0154(.A(x7), .B(ori_ori_n71_), .Y(ori_ori_n204_));
  NO2        o0155(.A(ori_ori_n187_), .B(ori_ori_n204_), .Y(ori_ori_n205_));
  OA210      o0156(.A0(ori_ori_n203_), .A1(ori_ori_n200_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  AOI220     o0157(.A0(ori_ori_n206_), .A1(ori_ori_n201_), .B0(ori_ori_n199_), .B1(x0), .Y(ori_ori_n207_));
  OAI210     o0158(.A0(ori_ori_n193_), .A1(ori_ori_n71_), .B0(ori_ori_n207_), .Y(ori_ori_n208_));
  NO2        o0159(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n209_));
  NA4        o0160(.A(ori_ori_n55_), .B(x5), .C(x3), .D(x2), .Y(ori_ori_n210_));
  NA2        o0161(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n211_));
  NA2        o0162(.A(ori_ori_n211_), .B(x2), .Y(ori_ori_n212_));
  NA2        o0163(.A(ori_ori_n55_), .B(x3), .Y(ori_ori_n213_));
  NA4        o0164(.A(ori_ori_n213_), .B(ori_ori_n212_), .C(ori_ori_n200_), .D(ori_ori_n82_), .Y(ori_ori_n214_));
  AOI210     o0165(.A0(ori_ori_n214_), .A1(ori_ori_n210_), .B0(ori_ori_n53_), .Y(ori_ori_n215_));
  NO2        o0166(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n216_));
  NA2        o0167(.A(x5), .B(x1), .Y(ori_ori_n217_));
  NO2        o0168(.A(ori_ori_n217_), .B(x6), .Y(ori_ori_n218_));
  NO2        o0169(.A(x3), .B(x1), .Y(ori_ori_n219_));
  AOI210     o0170(.A0(ori_ori_n219_), .A1(ori_ori_n77_), .B0(ori_ori_n218_), .Y(ori_ori_n220_));
  NO2        o0171(.A(ori_ori_n81_), .B(ori_ori_n55_), .Y(ori_ori_n221_));
  NO2        o0172(.A(ori_ori_n100_), .B(ori_ori_n50_), .Y(ori_ori_n222_));
  NO2        o0173(.A(ori_ori_n222_), .B(ori_ori_n221_), .Y(ori_ori_n223_));
  OAI210     o0174(.A0(ori_ori_n220_), .A1(x8), .B0(ori_ori_n223_), .Y(ori_ori_n224_));
  NO2        o0175(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n225_));
  NA2        o0176(.A(ori_ori_n225_), .B(ori_ori_n71_), .Y(ori_ori_n226_));
  NAi21      o0177(.An(x2), .B(x5), .Y(ori_ori_n227_));
  NA2        o0178(.A(x8), .B(x6), .Y(ori_ori_n228_));
  OAI210     o0179(.A0(ori_ori_n228_), .A1(ori_ori_n227_), .B0(ori_ori_n226_), .Y(ori_ori_n229_));
  NA2        o0180(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n230_));
  NO2        o0181(.A(ori_ori_n230_), .B(ori_ori_n59_), .Y(ori_ori_n231_));
  AO220      o0182(.A0(ori_ori_n231_), .A1(ori_ori_n229_), .B0(ori_ori_n224_), .B1(ori_ori_n216_), .Y(ori_ori_n232_));
  OAI210     o0183(.A0(ori_ori_n232_), .A1(ori_ori_n215_), .B0(ori_ori_n209_), .Y(ori_ori_n233_));
  NA2        o0184(.A(ori_ori_n71_), .B(ori_ori_n56_), .Y(ori_ori_n234_));
  NO2        o0185(.A(ori_ori_n234_), .B(x7), .Y(ori_ori_n235_));
  NO2        o0186(.A(ori_ori_n104_), .B(ori_ori_n53_), .Y(ori_ori_n236_));
  NA2        o0187(.A(ori_ori_n236_), .B(ori_ori_n106_), .Y(ori_ori_n237_));
  AOI210     o0188(.A0(ori_ori_n237_), .A1(ori_ori_n164_), .B0(ori_ori_n59_), .Y(ori_ori_n238_));
  NA2        o0189(.A(x3), .B(ori_ori_n59_), .Y(ori_ori_n239_));
  NO2        o0190(.A(ori_ori_n177_), .B(ori_ori_n239_), .Y(ori_ori_n240_));
  OA210      o0191(.A0(ori_ori_n240_), .A1(ori_ori_n238_), .B0(x8), .Y(ori_ori_n241_));
  NO2        o0192(.A(x1), .B(x0), .Y(ori_ori_n242_));
  NA2        o0193(.A(ori_ori_n242_), .B(ori_ori_n106_), .Y(ori_ori_n243_));
  NA2        o0194(.A(ori_ori_n104_), .B(ori_ori_n50_), .Y(ori_ori_n244_));
  XN2        o0195(.A(x3), .B(x2), .Y(ori_ori_n245_));
  NA2        o0196(.A(ori_ori_n245_), .B(ori_ori_n156_), .Y(ori_ori_n246_));
  NO2        o0197(.A(ori_ori_n104_), .B(x0), .Y(ori_ori_n247_));
  NA2        o0198(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n248_));
  NA2        o0199(.A(ori_ori_n248_), .B(ori_ori_n247_), .Y(ori_ori_n249_));
  OAI220     o0200(.A0(ori_ori_n249_), .A1(ori_ori_n246_), .B0(ori_ori_n244_), .B1(ori_ori_n243_), .Y(ori_ori_n250_));
  OAI210     o0201(.A0(ori_ori_n250_), .A1(ori_ori_n241_), .B0(ori_ori_n235_), .Y(ori_ori_n251_));
  NO2        o0202(.A(x7), .B(x1), .Y(ori_ori_n252_));
  NOi21      o0203(.An(x8), .B(x3), .Y(ori_ori_n253_));
  NA2        o0204(.A(ori_ori_n253_), .B(ori_ori_n59_), .Y(ori_ori_n254_));
  NA2        o0205(.A(x5), .B(x0), .Y(ori_ori_n255_));
  NAi21      o0206(.An(ori_ori_n136_), .B(ori_ori_n255_), .Y(ori_ori_n256_));
  NA2        o0207(.A(ori_ori_n71_), .B(ori_ori_n50_), .Y(ori_ori_n257_));
  OAI210     o0208(.A0(ori_ori_n257_), .A1(ori_ori_n256_), .B0(ori_ori_n254_), .Y(ori_ori_n258_));
  NA3        o0209(.A(ori_ori_n258_), .B(ori_ori_n139_), .C(ori_ori_n252_), .Y(ori_ori_n259_));
  NA2        o0210(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n260_));
  NO2        o0211(.A(ori_ori_n260_), .B(x5), .Y(ori_ori_n261_));
  NO2        o0212(.A(ori_ori_n148_), .B(ori_ori_n71_), .Y(ori_ori_n262_));
  NA2        o0213(.A(x1), .B(x0), .Y(ori_ori_n263_));
  NA2        o0214(.A(ori_ori_n50_), .B(ori_ori_n59_), .Y(ori_ori_n264_));
  NA4        o0215(.A(ori_ori_n264_), .B(ori_ori_n263_), .C(ori_ori_n262_), .D(ori_ori_n261_), .Y(ori_ori_n265_));
  NA3        o0216(.A(ori_ori_n265_), .B(ori_ori_n259_), .C(ori_ori_n184_), .Y(ori_ori_n266_));
  NO2        o0217(.A(ori_ori_n104_), .B(x3), .Y(ori_ori_n267_));
  NO2        o0218(.A(ori_ori_n106_), .B(x0), .Y(ori_ori_n268_));
  NA2        o0219(.A(ori_ori_n268_), .B(ori_ori_n267_), .Y(ori_ori_n269_));
  NO2        o0220(.A(ori_ori_n55_), .B(x7), .Y(ori_ori_n270_));
  NA2        o0221(.A(ori_ori_n270_), .B(ori_ori_n137_), .Y(ori_ori_n271_));
  NO3        o0222(.A(x8), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n272_));
  NAi21      o0223(.An(x8), .B(x0), .Y(ori_ori_n273_));
  NAi21      o0224(.An(x1), .B(x3), .Y(ori_ori_n274_));
  NO2        o0225(.A(ori_ori_n274_), .B(ori_ori_n273_), .Y(ori_ori_n275_));
  NO2        o0226(.A(x2), .B(ori_ori_n53_), .Y(ori_ori_n276_));
  AOI210     o0227(.A0(ori_ori_n276_), .A1(ori_ori_n272_), .B0(ori_ori_n275_), .Y(ori_ori_n277_));
  NOi21      o0228(.An(x5), .B(x6), .Y(ori_ori_n278_));
  NO2        o0229(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n279_));
  NA2        o0230(.A(ori_ori_n279_), .B(ori_ori_n278_), .Y(ori_ori_n280_));
  OAI220     o0231(.A0(ori_ori_n280_), .A1(ori_ori_n277_), .B0(ori_ori_n271_), .B1(ori_ori_n269_), .Y(ori_ori_n281_));
  AOI210     o0232(.A0(ori_ori_n266_), .A1(ori_ori_n107_), .B0(ori_ori_n281_), .Y(ori_ori_n282_));
  NA3        o0233(.A(ori_ori_n282_), .B(ori_ori_n251_), .C(ori_ori_n233_), .Y(ori_ori_n283_));
  AOI210     o0234(.A0(ori_ori_n208_), .A1(ori_ori_n56_), .B0(ori_ori_n283_), .Y(ori02));
  NO2        o0235(.A(x8), .B(ori_ori_n104_), .Y(ori_ori_n285_));
  XN2        o0236(.A(x7), .B(x3), .Y(ori_ori_n286_));
  INV        o0237(.A(ori_ori_n286_), .Y(ori_ori_n287_));
  NO2        o0238(.A(x2), .B(x0), .Y(ori_ori_n288_));
  NA2        o0239(.A(ori_ori_n288_), .B(ori_ori_n71_), .Y(ori_ori_n289_));
  NO2        o0240(.A(ori_ori_n57_), .B(x1), .Y(ori_ori_n290_));
  NO3        o0241(.A(ori_ori_n290_), .B(ori_ori_n289_), .C(ori_ori_n287_), .Y(ori_ori_n291_));
  NA2        o0242(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n292_));
  NO2        o0243(.A(ori_ori_n274_), .B(x6), .Y(ori_ori_n293_));
  XO2        o0244(.A(x7), .B(x0), .Y(ori_ori_n294_));
  NO2        o0245(.A(ori_ori_n294_), .B(ori_ori_n288_), .Y(ori_ori_n295_));
  NA2        o0246(.A(ori_ori_n295_), .B(ori_ori_n293_), .Y(ori_ori_n296_));
  AN2        o0247(.A(x7), .B(x2), .Y(ori_ori_n297_));
  NA2        o0248(.A(ori_ori_n297_), .B(ori_ori_n50_), .Y(ori_ori_n298_));
  OAI210     o0249(.A0(ori_ori_n298_), .A1(ori_ori_n292_), .B0(ori_ori_n296_), .Y(ori_ori_n299_));
  OAI210     o0250(.A0(ori_ori_n299_), .A1(ori_ori_n291_), .B0(ori_ori_n285_), .Y(ori_ori_n300_));
  NAi21      o0251(.An(x8), .B(x6), .Y(ori_ori_n301_));
  NO2        o0252(.A(ori_ori_n104_), .B(ori_ori_n59_), .Y(ori_ori_n302_));
  NA2        o0253(.A(x7), .B(x3), .Y(ori_ori_n303_));
  NO2        o0254(.A(ori_ori_n303_), .B(x2), .Y(ori_ori_n304_));
  NA2        o0255(.A(x2), .B(x0), .Y(ori_ori_n305_));
  NA2        o0256(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n306_));
  NA2        o0257(.A(ori_ori_n306_), .B(ori_ori_n305_), .Y(ori_ori_n307_));
  NAi21      o0258(.An(x7), .B(x1), .Y(ori_ori_n308_));
  NO2        o0259(.A(ori_ori_n308_), .B(x3), .Y(ori_ori_n309_));
  AOI220     o0260(.A0(ori_ori_n309_), .A1(ori_ori_n307_), .B0(ori_ori_n304_), .B1(ori_ori_n302_), .Y(ori_ori_n310_));
  NA2        o0261(.A(ori_ori_n276_), .B(ori_ori_n50_), .Y(ori_ori_n311_));
  NA3        o0262(.A(x7), .B(ori_ori_n104_), .C(x0), .Y(ori_ori_n312_));
  NA2        o0263(.A(ori_ori_n162_), .B(ori_ori_n57_), .Y(ori_ori_n313_));
  NO2        o0264(.A(ori_ori_n310_), .B(ori_ori_n301_), .Y(ori_ori_n314_));
  INV        o0265(.A(ori_ori_n294_), .Y(ori_ori_n315_));
  NO2        o0266(.A(x7), .B(ori_ori_n71_), .Y(ori_ori_n316_));
  NA2        o0267(.A(ori_ori_n104_), .B(x3), .Y(ori_ori_n317_));
  NO2        o0268(.A(ori_ori_n317_), .B(ori_ori_n316_), .Y(ori_ori_n318_));
  NA2        o0269(.A(ori_ori_n318_), .B(ori_ori_n315_), .Y(ori_ori_n319_));
  NA2        o0270(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n320_));
  NO2        o0271(.A(ori_ori_n320_), .B(x7), .Y(ori_ori_n321_));
  NA2        o0272(.A(ori_ori_n321_), .B(ori_ori_n278_), .Y(ori_ori_n322_));
  NA2        o0273(.A(ori_ori_n167_), .B(x1), .Y(ori_ori_n323_));
  AOI210     o0274(.A0(ori_ori_n322_), .A1(ori_ori_n319_), .B0(ori_ori_n323_), .Y(ori_ori_n324_));
  NO2        o0275(.A(ori_ori_n57_), .B(ori_ori_n50_), .Y(ori_ori_n325_));
  NO2        o0276(.A(ori_ori_n55_), .B(ori_ori_n106_), .Y(ori_ori_n326_));
  NA3        o0277(.A(ori_ori_n326_), .B(ori_ori_n325_), .C(ori_ori_n59_), .Y(ori_ori_n327_));
  NO2        o0278(.A(ori_ori_n157_), .B(x6), .Y(ori_ori_n328_));
  NO2        o0279(.A(ori_ori_n100_), .B(ori_ori_n104_), .Y(ori_ori_n329_));
  NA2        o0280(.A(ori_ori_n57_), .B(ori_ori_n106_), .Y(ori_ori_n330_));
  NO2        o0281(.A(ori_ori_n330_), .B(ori_ori_n264_), .Y(ori_ori_n331_));
  OAI210     o0282(.A0(ori_ori_n329_), .A1(ori_ori_n328_), .B0(ori_ori_n331_), .Y(ori_ori_n332_));
  OAI210     o0283(.A0(ori_ori_n327_), .A1(ori_ori_n100_), .B0(ori_ori_n332_), .Y(ori_ori_n333_));
  NO3        o0284(.A(ori_ori_n333_), .B(ori_ori_n324_), .C(ori_ori_n314_), .Y(ori_ori_n334_));
  AOI210     o0285(.A0(ori_ori_n334_), .A1(ori_ori_n300_), .B0(x4), .Y(ori_ori_n335_));
  NA2        o0286(.A(x8), .B(ori_ori_n71_), .Y(ori_ori_n336_));
  NO2        o0287(.A(x3), .B(ori_ori_n59_), .Y(ori_ori_n337_));
  NA3        o0288(.A(ori_ori_n337_), .B(ori_ori_n104_), .C(ori_ori_n53_), .Y(ori_ori_n338_));
  NO2        o0289(.A(x3), .B(x0), .Y(ori_ori_n339_));
  NAi21      o0290(.An(ori_ori_n339_), .B(ori_ori_n103_), .Y(ori_ori_n340_));
  NA2        o0291(.A(x5), .B(x2), .Y(ori_ori_n341_));
  NO2        o0292(.A(ori_ori_n341_), .B(ori_ori_n219_), .Y(ori_ori_n342_));
  AOI210     o0293(.A0(ori_ori_n342_), .A1(ori_ori_n340_), .B0(ori_ori_n240_), .Y(ori_ori_n343_));
  AO210      o0294(.A0(ori_ori_n343_), .A1(ori_ori_n338_), .B0(ori_ori_n336_), .Y(ori_ori_n344_));
  NO2        o0295(.A(ori_ori_n106_), .B(ori_ori_n53_), .Y(ori_ori_n345_));
  NA2        o0296(.A(ori_ori_n345_), .B(x3), .Y(ori_ori_n346_));
  NO2        o0297(.A(ori_ori_n55_), .B(x1), .Y(ori_ori_n347_));
  NA2        o0298(.A(ori_ori_n347_), .B(ori_ori_n106_), .Y(ori_ori_n348_));
  OAI210     o0299(.A0(ori_ori_n348_), .A1(ori_ori_n169_), .B0(ori_ori_n346_), .Y(ori_ori_n349_));
  NAi32      o0300(.An(x3), .Bn(x0), .C(x2), .Y(ori_ori_n350_));
  NO2        o0301(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n351_));
  NAi21      o0302(.An(x6), .B(x5), .Y(ori_ori_n352_));
  NO2        o0303(.A(x2), .B(ori_ori_n59_), .Y(ori_ori_n353_));
  NO4        o0304(.A(ori_ori_n353_), .B(ori_ori_n352_), .C(ori_ori_n159_), .D(ori_ori_n351_), .Y(ori_ori_n354_));
  AOI220     o0305(.A0(ori_ori_n354_), .A1(ori_ori_n350_), .B0(ori_ori_n349_), .B1(ori_ori_n85_), .Y(ori_ori_n355_));
  AOI210     o0306(.A0(ori_ori_n355_), .A1(ori_ori_n344_), .B0(ori_ori_n75_), .Y(ori_ori_n356_));
  NA2        o0307(.A(ori_ori_n347_), .B(ori_ori_n56_), .Y(ori_ori_n357_));
  NO2        o0308(.A(ori_ori_n104_), .B(ori_ori_n50_), .Y(ori_ori_n358_));
  NO2        o0309(.A(ori_ori_n288_), .B(ori_ori_n216_), .Y(ori_ori_n359_));
  XO2        o0310(.A(x7), .B(x2), .Y(ori_ori_n360_));
  INV        o0311(.A(ori_ori_n360_), .Y(ori_ori_n361_));
  XO2        o0312(.A(x6), .B(x2), .Y(ori_ori_n362_));
  NAi21      o0313(.An(x0), .B(x6), .Y(ori_ori_n363_));
  AOI210     o0314(.A0(ori_ori_n363_), .A1(ori_ori_n142_), .B0(ori_ori_n268_), .Y(ori_ori_n364_));
  XN2        o0315(.A(x7), .B(x5), .Y(ori_ori_n365_));
  NA2        o0316(.A(ori_ori_n365_), .B(ori_ori_n71_), .Y(ori_ori_n366_));
  NA2        o0317(.A(x7), .B(x5), .Y(ori_ori_n367_));
  AOI210     o0318(.A0(ori_ori_n367_), .A1(x6), .B0(ori_ori_n350_), .Y(ori_ori_n368_));
  AOI220     o0319(.A0(ori_ori_n368_), .A1(ori_ori_n366_), .B0(ori_ori_n364_), .B1(ori_ori_n318_), .Y(ori_ori_n369_));
  NO2        o0320(.A(ori_ori_n369_), .B(ori_ori_n357_), .Y(ori_ori_n370_));
  NO2        o0321(.A(x8), .B(x6), .Y(ori_ori_n371_));
  NAi21      o0322(.An(ori_ori_n371_), .B(ori_ori_n228_), .Y(ori_ori_n372_));
  AOI210     o0323(.A0(ori_ori_n372_), .A1(ori_ori_n90_), .B0(x3), .Y(ori_ori_n373_));
  NA2        o0324(.A(ori_ori_n104_), .B(x2), .Y(ori_ori_n374_));
  NO2        o0325(.A(ori_ori_n374_), .B(ori_ori_n64_), .Y(ori_ori_n375_));
  NA2        o0326(.A(x1), .B(ori_ori_n59_), .Y(ori_ori_n376_));
  NO2        o0327(.A(ori_ori_n376_), .B(ori_ori_n228_), .Y(ori_ori_n377_));
  OAI210     o0328(.A0(ori_ori_n377_), .A1(ori_ori_n50_), .B0(ori_ori_n375_), .Y(ori_ori_n378_));
  NA2        o0329(.A(x4), .B(x2), .Y(ori_ori_n379_));
  NO2        o0330(.A(ori_ori_n379_), .B(ori_ori_n104_), .Y(ori_ori_n380_));
  NAi21      o0331(.An(x1), .B(x6), .Y(ori_ori_n381_));
  NA2        o0332(.A(ori_ori_n339_), .B(ori_ori_n270_), .Y(ori_ori_n382_));
  OAI220     o0333(.A0(ori_ori_n382_), .A1(ori_ori_n381_), .B0(ori_ori_n103_), .B1(ori_ori_n53_), .Y(ori_ori_n383_));
  NA2        o0334(.A(x8), .B(x2), .Y(ori_ori_n384_));
  NO2        o0335(.A(ori_ori_n384_), .B(ori_ori_n50_), .Y(ori_ori_n385_));
  INV        o0336(.A(ori_ori_n218_), .Y(ori_ori_n386_));
  NO2        o0337(.A(ori_ori_n386_), .B(ori_ori_n52_), .Y(ori_ori_n387_));
  AOI220     o0338(.A0(ori_ori_n387_), .A1(ori_ori_n385_), .B0(ori_ori_n383_), .B1(ori_ori_n380_), .Y(ori_ori_n388_));
  OAI210     o0339(.A0(ori_ori_n378_), .A1(ori_ori_n373_), .B0(ori_ori_n388_), .Y(ori_ori_n389_));
  NO4        o0340(.A(ori_ori_n389_), .B(ori_ori_n370_), .C(ori_ori_n356_), .D(ori_ori_n335_), .Y(ori03));
  NAi21      o0341(.An(x2), .B(x0), .Y(ori_ori_n391_));
  NO3        o0342(.A(x8), .B(x6), .C(x4), .Y(ori_ori_n392_));
  INV        o0343(.A(ori_ori_n392_), .Y(ori_ori_n393_));
  NO2        o0344(.A(ori_ori_n393_), .B(ori_ori_n391_), .Y(ori_ori_n394_));
  NA2        o0345(.A(ori_ori_n107_), .B(ori_ori_n59_), .Y(ori_ori_n395_));
  NO2        o0346(.A(ori_ori_n395_), .B(ori_ori_n55_), .Y(ori_ori_n396_));
  OAI210     o0347(.A0(ori_ori_n396_), .A1(ori_ori_n394_), .B0(ori_ori_n162_), .Y(ori_ori_n397_));
  NA2        o0348(.A(x3), .B(x2), .Y(ori_ori_n398_));
  NO2        o0349(.A(ori_ori_n159_), .B(x0), .Y(ori_ori_n399_));
  NA2        o0350(.A(x8), .B(x0), .Y(ori_ori_n400_));
  NO2        o0351(.A(ori_ori_n400_), .B(x6), .Y(ori_ori_n401_));
  AOI210     o0352(.A0(ori_ori_n401_), .A1(x5), .B0(ori_ori_n399_), .Y(ori_ori_n402_));
  NO2        o0353(.A(ori_ori_n402_), .B(ori_ori_n398_), .Y(ori_ori_n403_));
  NO2        o0354(.A(x5), .B(ori_ori_n59_), .Y(ori_ori_n404_));
  NO2        o0355(.A(x3), .B(x2), .Y(ori_ori_n405_));
  NA2        o0356(.A(ori_ori_n405_), .B(ori_ori_n404_), .Y(ori_ori_n406_));
  NO2        o0357(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n407_));
  NA2        o0358(.A(ori_ori_n407_), .B(x5), .Y(ori_ori_n408_));
  AOI210     o0359(.A0(ori_ori_n408_), .A1(ori_ori_n406_), .B0(ori_ori_n301_), .Y(ori_ori_n409_));
  NA2        o0360(.A(ori_ori_n254_), .B(ori_ori_n171_), .Y(ori_ori_n410_));
  NO2        o0361(.A(ori_ori_n50_), .B(ori_ori_n59_), .Y(ori_ori_n411_));
  NO2        o0362(.A(ori_ori_n71_), .B(x0), .Y(ori_ori_n412_));
  NO4        o0363(.A(ori_ori_n412_), .B(ori_ori_n411_), .C(x2), .D(ori_ori_n53_), .Y(ori_ori_n413_));
  AO210      o0364(.A0(ori_ori_n413_), .A1(ori_ori_n410_), .B0(ori_ori_n409_), .Y(ori_ori_n414_));
  OAI210     o0365(.A0(ori_ori_n414_), .A1(ori_ori_n403_), .B0(x4), .Y(ori_ori_n415_));
  NO2        o0366(.A(x4), .B(ori_ori_n53_), .Y(ori_ori_n416_));
  NA2        o0367(.A(ori_ori_n416_), .B(ori_ori_n59_), .Y(ori_ori_n417_));
  NO3        o0368(.A(ori_ori_n417_), .B(ori_ori_n228_), .C(x5), .Y(ori_ori_n418_));
  NA2        o0369(.A(x7), .B(ori_ori_n104_), .Y(ori_ori_n419_));
  NO3        o0370(.A(x5), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n420_));
  INV        o0371(.A(ori_ori_n420_), .Y(ori_ori_n421_));
  NO2        o0372(.A(x6), .B(ori_ori_n56_), .Y(ori_ori_n422_));
  NO2        o0373(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n423_));
  NA2        o0374(.A(ori_ori_n423_), .B(ori_ori_n422_), .Y(ori_ori_n424_));
  OAI210     o0375(.A0(ori_ori_n424_), .A1(ori_ori_n421_), .B0(ori_ori_n419_), .Y(ori_ori_n425_));
  AOI210     o0376(.A0(ori_ori_n418_), .A1(x2), .B0(ori_ori_n425_), .Y(ori_ori_n426_));
  AOI220     o0377(.A0(ori_ori_n426_), .A1(ori_ori_n415_), .B0(ori_ori_n397_), .B1(x7), .Y(ori_ori_n427_));
  NA2        o0378(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n428_));
  NO2        o0379(.A(ori_ori_n253_), .B(ori_ori_n106_), .Y(ori_ori_n429_));
  NO2        o0380(.A(ori_ori_n55_), .B(ori_ori_n59_), .Y(ori_ori_n430_));
  NO3        o0381(.A(ori_ori_n430_), .B(ori_ori_n429_), .C(ori_ori_n146_), .Y(ori_ori_n431_));
  AOI210     o0382(.A0(ori_ori_n203_), .A1(ori_ori_n97_), .B0(ori_ori_n431_), .Y(ori_ori_n432_));
  NO2        o0383(.A(x5), .B(x2), .Y(ori_ori_n433_));
  NO2        o0384(.A(x8), .B(x3), .Y(ori_ori_n434_));
  NA2        o0385(.A(ori_ori_n434_), .B(ori_ori_n433_), .Y(ori_ori_n435_));
  NO2        o0386(.A(ori_ori_n435_), .B(x6), .Y(ori_ori_n436_));
  NA2        o0387(.A(ori_ori_n202_), .B(x2), .Y(ori_ori_n437_));
  NO3        o0388(.A(ori_ori_n434_), .B(ori_ori_n340_), .C(ori_ori_n352_), .Y(ori_ori_n438_));
  NA2        o0389(.A(ori_ori_n438_), .B(ori_ori_n437_), .Y(ori_ori_n439_));
  OAI210     o0390(.A0(ori_ori_n432_), .A1(ori_ori_n288_), .B0(ori_ori_n439_), .Y(ori_ori_n440_));
  NA2        o0391(.A(ori_ori_n440_), .B(x4), .Y(ori_ori_n441_));
  NA2        o0392(.A(ori_ori_n55_), .B(ori_ori_n59_), .Y(ori_ori_n442_));
  NO2        o0393(.A(ori_ori_n442_), .B(x5), .Y(ori_ori_n443_));
  NAi21      o0394(.An(x4), .B(x6), .Y(ori_ori_n444_));
  NO2        o0395(.A(ori_ori_n444_), .B(ori_ori_n51_), .Y(ori_ori_n445_));
  NO2        o0396(.A(ori_ori_n55_), .B(ori_ori_n71_), .Y(ori_ori_n446_));
  NO2        o0397(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n447_));
  NO2        o0398(.A(ori_ori_n228_), .B(x0), .Y(ori_ori_n448_));
  NO2        o0399(.A(ori_ori_n352_), .B(x8), .Y(ori_ori_n449_));
  OAI210     o0400(.A0(ori_ori_n449_), .A1(ori_ori_n448_), .B0(ori_ori_n447_), .Y(ori_ori_n450_));
  OAI210     o0401(.A0(ori_ori_n406_), .A1(ori_ori_n446_), .B0(ori_ori_n450_), .Y(ori_ori_n451_));
  AOI220     o0402(.A0(ori_ori_n451_), .A1(ori_ori_n56_), .B0(ori_ori_n445_), .B1(ori_ori_n443_), .Y(ori_ori_n452_));
  AOI210     o0403(.A0(ori_ori_n452_), .A1(ori_ori_n441_), .B0(ori_ori_n428_), .Y(ori_ori_n453_));
  NA2        o0404(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n454_));
  NO2        o0405(.A(ori_ori_n71_), .B(ori_ori_n56_), .Y(ori_ori_n455_));
  NA2        o0406(.A(ori_ori_n351_), .B(ori_ori_n59_), .Y(ori_ori_n456_));
  OAI220     o0407(.A0(ori_ori_n456_), .A1(ori_ori_n55_), .B0(ori_ori_n195_), .B1(ori_ori_n273_), .Y(ori_ori_n457_));
  NA2        o0408(.A(ori_ori_n457_), .B(ori_ori_n455_), .Y(ori_ori_n458_));
  NO3        o0409(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n459_));
  NA2        o0410(.A(ori_ori_n430_), .B(x5), .Y(ori_ori_n460_));
  NO2        o0411(.A(x8), .B(x5), .Y(ori_ori_n461_));
  NAi21      o0412(.An(ori_ori_n461_), .B(ori_ori_n171_), .Y(ori_ori_n462_));
  OAI210     o0413(.A0(ori_ori_n462_), .A1(ori_ori_n306_), .B0(ori_ori_n460_), .Y(ori_ori_n463_));
  NA2        o0414(.A(ori_ori_n359_), .B(ori_ori_n77_), .Y(ori_ori_n464_));
  NOi21      o0415(.An(x3), .B(x4), .Y(ori_ori_n465_));
  NA2        o0416(.A(ori_ori_n55_), .B(ori_ori_n106_), .Y(ori_ori_n466_));
  NA2        o0417(.A(ori_ori_n466_), .B(ori_ori_n465_), .Y(ori_ori_n467_));
  NO2        o0418(.A(ori_ori_n51_), .B(x6), .Y(ori_ori_n468_));
  NO2        o0419(.A(ori_ori_n146_), .B(ori_ori_n55_), .Y(ori_ori_n469_));
  NO3        o0420(.A(ori_ori_n56_), .B(x2), .C(x0), .Y(ori_ori_n470_));
  AOI220     o0421(.A0(ori_ori_n470_), .A1(ori_ori_n469_), .B0(ori_ori_n468_), .B1(ori_ori_n443_), .Y(ori_ori_n471_));
  OAI210     o0422(.A0(ori_ori_n467_), .A1(ori_ori_n464_), .B0(ori_ori_n471_), .Y(ori_ori_n472_));
  AOI210     o0423(.A0(ori_ori_n463_), .A1(ori_ori_n459_), .B0(ori_ori_n472_), .Y(ori_ori_n473_));
  AOI210     o0424(.A0(ori_ori_n473_), .A1(ori_ori_n458_), .B0(ori_ori_n454_), .Y(ori_ori_n474_));
  NA2        o0425(.A(x7), .B(x1), .Y(ori_ori_n475_));
  NO3        o0426(.A(x5), .B(x4), .C(x2), .Y(ori_ori_n476_));
  AN2        o0427(.A(ori_ori_n476_), .B(ori_ori_n371_), .Y(ori_ori_n477_));
  NO3        o0428(.A(ori_ori_n477_), .B(ori_ori_n469_), .C(ori_ori_n380_), .Y(ori_ori_n478_));
  OAI210     o0429(.A0(ori_ori_n371_), .A1(ori_ori_n84_), .B0(ori_ori_n339_), .Y(ori_ori_n479_));
  NO2        o0430(.A(ori_ori_n479_), .B(ori_ori_n478_), .Y(ori_ori_n480_));
  NO2        o0431(.A(x4), .B(ori_ori_n106_), .Y(ori_ori_n481_));
  NA2        o0432(.A(ori_ori_n481_), .B(x6), .Y(ori_ori_n482_));
  NA3        o0433(.A(ori_ori_n104_), .B(x4), .C(ori_ori_n106_), .Y(ori_ori_n483_));
  AOI210     o0434(.A0(ori_ori_n483_), .A1(ori_ori_n482_), .B0(ori_ori_n96_), .Y(ori_ori_n484_));
  NA2        o0435(.A(ori_ori_n465_), .B(ori_ori_n71_), .Y(ori_ori_n485_));
  NA2        o0436(.A(ori_ori_n167_), .B(ori_ori_n59_), .Y(ori_ori_n486_));
  NO2        o0437(.A(ori_ori_n486_), .B(ori_ori_n485_), .Y(ori_ori_n487_));
  NA2        o0438(.A(ori_ori_n447_), .B(x4), .Y(ori_ori_n488_));
  NO3        o0439(.A(ori_ori_n488_), .B(ori_ori_n371_), .C(ori_ori_n412_), .Y(ori_ori_n489_));
  NO4        o0440(.A(ori_ori_n489_), .B(ori_ori_n487_), .C(ori_ori_n484_), .D(ori_ori_n480_), .Y(ori_ori_n490_));
  NA2        o0441(.A(x5), .B(x4), .Y(ori_ori_n491_));
  NO2        o0442(.A(ori_ori_n71_), .B(ori_ori_n53_), .Y(ori_ori_n492_));
  NO3        o0443(.A(x8), .B(x3), .C(x2), .Y(ori_ori_n493_));
  NA3        o0444(.A(ori_ori_n493_), .B(ori_ori_n492_), .C(ori_ori_n59_), .Y(ori_ori_n494_));
  NO3        o0445(.A(x6), .B(x5), .C(x2), .Y(ori_ori_n495_));
  NA3        o0446(.A(ori_ori_n495_), .B(ori_ori_n290_), .C(ori_ori_n78_), .Y(ori_ori_n496_));
  OAI210     o0447(.A0(ori_ori_n494_), .A1(ori_ori_n491_), .B0(ori_ori_n496_), .Y(ori_ori_n497_));
  NA2        o0448(.A(ori_ori_n71_), .B(x2), .Y(ori_ori_n498_));
  NO3        o0449(.A(x4), .B(x3), .C(ori_ori_n59_), .Y(ori_ori_n499_));
  NA2        o0450(.A(ori_ori_n499_), .B(ori_ori_n225_), .Y(ori_ori_n500_));
  NO3        o0451(.A(ori_ori_n500_), .B(ori_ori_n498_), .C(ori_ori_n92_), .Y(ori_ori_n501_));
  XO2        o0452(.A(x4), .B(x0), .Y(ori_ori_n502_));
  NA2        o0453(.A(ori_ori_n264_), .B(x5), .Y(ori_ori_n503_));
  NO2        o0454(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n504_));
  NO2        o0455(.A(ori_ori_n504_), .B(ori_ori_n63_), .Y(ori_ori_n505_));
  NO4        o0456(.A(ori_ori_n505_), .B(ori_ori_n503_), .C(ori_ori_n502_), .D(ori_ori_n155_), .Y(ori_ori_n506_));
  NO3        o0457(.A(ori_ori_n506_), .B(ori_ori_n501_), .C(ori_ori_n497_), .Y(ori_ori_n507_));
  OAI210     o0458(.A0(ori_ori_n490_), .A1(ori_ori_n475_), .B0(ori_ori_n507_), .Y(ori_ori_n508_));
  NO4        o0459(.A(ori_ori_n508_), .B(ori_ori_n474_), .C(ori_ori_n453_), .D(ori_ori_n427_), .Y(ori04));
  NO2        o0460(.A(x7), .B(x2), .Y(ori_ori_n510_));
  NO2        o0461(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n511_));
  NO2        o0462(.A(ori_ori_n511_), .B(ori_ori_n148_), .Y(ori_ori_n512_));
  XN2        o0463(.A(x8), .B(x1), .Y(ori_ori_n513_));
  NO2        o0464(.A(ori_ori_n513_), .B(ori_ori_n146_), .Y(ori_ori_n514_));
  NA2        o0465(.A(ori_ori_n514_), .B(ori_ori_n512_), .Y(ori_ori_n515_));
  NA2        o0466(.A(x6), .B(x3), .Y(ori_ori_n516_));
  NO2        o0467(.A(ori_ori_n516_), .B(x5), .Y(ori_ori_n517_));
  NA2        o0468(.A(ori_ori_n71_), .B(x1), .Y(ori_ori_n518_));
  NO2        o0469(.A(ori_ori_n461_), .B(ori_ori_n253_), .Y(ori_ori_n519_));
  NO3        o0470(.A(ori_ori_n519_), .B(ori_ori_n434_), .C(ori_ori_n518_), .Y(ori_ori_n520_));
  AOI210     o0471(.A0(ori_ori_n517_), .A1(ori_ori_n347_), .B0(ori_ori_n520_), .Y(ori_ori_n521_));
  AOI210     o0472(.A0(ori_ori_n521_), .A1(ori_ori_n515_), .B0(x0), .Y(ori_ori_n522_));
  NOi21      o0473(.An(ori_ori_n171_), .B(ori_ori_n461_), .Y(ori_ori_n523_));
  NA2        o0474(.A(ori_ori_n105_), .B(x1), .Y(ori_ori_n524_));
  NO3        o0475(.A(ori_ori_n524_), .B(ori_ori_n523_), .C(ori_ori_n320_), .Y(ori_ori_n525_));
  OAI210     o0476(.A0(ori_ori_n525_), .A1(ori_ori_n522_), .B0(ori_ori_n510_), .Y(ori_ori_n526_));
  NA2        o0477(.A(ori_ori_n133_), .B(ori_ori_n239_), .Y(ori_ori_n527_));
  OR4        o0478(.A(ori_ori_n527_), .B(ori_ori_n372_), .C(ori_ori_n82_), .D(ori_ori_n54_), .Y(ori_ori_n528_));
  OR2        o0479(.A(x6), .B(x0), .Y(ori_ori_n529_));
  NO3        o0480(.A(ori_ori_n529_), .B(x3), .C(x1), .Y(ori_ori_n530_));
  AOI220     o0481(.A0(ori_ori_n530_), .A1(ori_ori_n104_), .B0(ori_ori_n278_), .B1(ori_ori_n272_), .Y(ori_ori_n531_));
  AOI210     o0482(.A0(ori_ori_n531_), .A1(ori_ori_n528_), .B0(ori_ori_n182_), .Y(ori_ori_n532_));
  NA2        o0483(.A(x7), .B(x2), .Y(ori_ori_n533_));
  INV        o0484(.A(ori_ori_n133_), .Y(ori_ori_n534_));
  OAI210     o0485(.A0(ori_ori_n170_), .A1(ori_ori_n534_), .B0(ori_ori_n82_), .Y(ori_ori_n535_));
  NO2        o0486(.A(ori_ori_n317_), .B(ori_ori_n55_), .Y(ori_ori_n536_));
  NO3        o0487(.A(x3), .B(x1), .C(x0), .Y(ori_ori_n537_));
  OR2        o0488(.A(x6), .B(x1), .Y(ori_ori_n538_));
  NA2        o0489(.A(ori_ori_n538_), .B(x0), .Y(ori_ori_n539_));
  AOI220     o0490(.A0(ori_ori_n539_), .A1(ori_ori_n536_), .B0(ori_ori_n537_), .B1(ori_ori_n469_), .Y(ori_ori_n540_));
  AOI210     o0491(.A0(ori_ori_n540_), .A1(ori_ori_n535_), .B0(ori_ori_n533_), .Y(ori_ori_n541_));
  NA2        o0492(.A(ori_ori_n71_), .B(x0), .Y(ori_ori_n542_));
  NOi31      o0493(.An(ori_ori_n342_), .B(ori_ori_n542_), .C(ori_ori_n260_), .Y(ori_ori_n543_));
  NO4        o0494(.A(ori_ori_n543_), .B(ori_ori_n541_), .C(ori_ori_n532_), .D(ori_ori_n56_), .Y(ori_ori_n544_));
  NA2        o0495(.A(ori_ori_n544_), .B(ori_ori_n526_), .Y(ori_ori_n545_));
  NA3        o0496(.A(x8), .B(x7), .C(x0), .Y(ori_ori_n546_));
  INV        o0497(.A(ori_ori_n546_), .Y(ori_ori_n547_));
  AOI210     o0498(.A0(ori_ori_n270_), .A1(ori_ori_n95_), .B0(ori_ori_n547_), .Y(ori_ori_n548_));
  NO2        o0499(.A(ori_ori_n548_), .B(ori_ori_n155_), .Y(ori_ori_n549_));
  NA2        o0500(.A(ori_ori_n430_), .B(ori_ori_n57_), .Y(ori_ori_n550_));
  NO2        o0501(.A(x8), .B(x0), .Y(ori_ori_n551_));
  NA2        o0502(.A(ori_ori_n551_), .B(ori_ori_n361_), .Y(ori_ori_n552_));
  AOI210     o0503(.A0(ori_ori_n552_), .A1(ori_ori_n550_), .B0(ori_ori_n274_), .Y(ori_ori_n553_));
  OAI210     o0504(.A0(ori_ori_n553_), .A1(ori_ori_n549_), .B0(ori_ori_n278_), .Y(ori_ori_n554_));
  NO2        o0505(.A(ori_ori_n71_), .B(ori_ori_n106_), .Y(ori_ori_n555_));
  NO2        o0506(.A(ori_ori_n367_), .B(x8), .Y(ori_ori_n556_));
  NO2        o0507(.A(ori_ori_n556_), .B(ori_ori_n261_), .Y(ori_ori_n557_));
  NO3        o0508(.A(ori_ori_n557_), .B(ori_ori_n376_), .C(ori_ori_n267_), .Y(ori_ori_n558_));
  NO2        o0509(.A(ori_ori_n287_), .B(x8), .Y(ori_ori_n559_));
  OAI210     o0510(.A0(ori_ori_n461_), .A1(ori_ori_n325_), .B0(ori_ori_n242_), .Y(ori_ori_n560_));
  NA2        o0511(.A(ori_ori_n347_), .B(ori_ori_n175_), .Y(ori_ori_n561_));
  OAI220     o0512(.A0(ori_ori_n561_), .A1(ori_ori_n59_), .B0(ori_ori_n560_), .B1(ori_ori_n559_), .Y(ori_ori_n562_));
  OAI210     o0513(.A0(ori_ori_n562_), .A1(ori_ori_n558_), .B0(ori_ori_n555_), .Y(ori_ori_n563_));
  NO2        o0514(.A(x8), .B(x2), .Y(ori_ori_n564_));
  NO2        o0515(.A(ori_ori_n219_), .B(ori_ori_n57_), .Y(ori_ori_n565_));
  NA3        o0516(.A(ori_ori_n565_), .B(ori_ori_n564_), .C(ori_ori_n340_), .Y(ori_ori_n566_));
  NO2        o0517(.A(ori_ori_n243_), .B(ori_ori_n133_), .Y(ori_ori_n567_));
  AOI210     o0518(.A0(ori_ori_n321_), .A1(ori_ori_n163_), .B0(ori_ori_n567_), .Y(ori_ori_n568_));
  AOI210     o0519(.A0(ori_ori_n568_), .A1(ori_ori_n566_), .B0(ori_ori_n105_), .Y(ori_ori_n569_));
  NA2        o0520(.A(ori_ori_n337_), .B(x2), .Y(ori_ori_n570_));
  NO2        o0521(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n571_));
  NA2        o0522(.A(ori_ori_n571_), .B(ori_ori_n63_), .Y(ori_ori_n572_));
  AOI210     o0523(.A0(ori_ori_n570_), .A1(ori_ori_n456_), .B0(ori_ori_n572_), .Y(ori_ori_n573_));
  NA2        o0524(.A(ori_ori_n106_), .B(ori_ori_n53_), .Y(ori_ori_n574_));
  NO2        o0525(.A(ori_ori_n574_), .B(x8), .Y(ori_ori_n575_));
  NA2        o0526(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n576_));
  NO2        o0527(.A(ori_ori_n180_), .B(ori_ori_n576_), .Y(ori_ori_n577_));
  AN2        o0528(.A(ori_ori_n577_), .B(ori_ori_n575_), .Y(ori_ori_n578_));
  NA2        o0529(.A(ori_ori_n404_), .B(ori_ori_n148_), .Y(ori_ori_n579_));
  NO2        o0530(.A(ori_ori_n71_), .B(x2), .Y(ori_ori_n580_));
  NA2        o0531(.A(ori_ori_n580_), .B(ori_ori_n270_), .Y(ori_ori_n581_));
  NO4        o0532(.A(x4), .B(ori_ori_n578_), .C(ori_ori_n573_), .D(ori_ori_n569_), .Y(ori_ori_n582_));
  NA3        o0533(.A(ori_ori_n582_), .B(ori_ori_n563_), .C(ori_ori_n554_), .Y(ori_ori_n583_));
  NA2        o0534(.A(ori_ori_n53_), .B(ori_ori_n59_), .Y(ori_ori_n584_));
  NOi21      o0535(.An(x2), .B(x7), .Y(ori_ori_n585_));
  NO2        o0536(.A(x6), .B(x3), .Y(ori_ori_n586_));
  NA2        o0537(.A(ori_ori_n586_), .B(ori_ori_n585_), .Y(ori_ori_n587_));
  NO2        o0538(.A(x6), .B(ori_ori_n59_), .Y(ori_ori_n588_));
  NO3        o0539(.A(ori_ori_n57_), .B(x2), .C(x1), .Y(ori_ori_n589_));
  NO3        o0540(.A(ori_ori_n57_), .B(x2), .C(x0), .Y(ori_ori_n590_));
  AOI220     o0541(.A0(ori_ori_n590_), .A1(ori_ori_n222_), .B0(ori_ori_n589_), .B1(ori_ori_n588_), .Y(ori_ori_n591_));
  OAI210     o0542(.A0(ori_ori_n587_), .A1(ori_ori_n584_), .B0(ori_ori_n591_), .Y(ori_ori_n592_));
  NO2        o0543(.A(ori_ori_n97_), .B(ori_ori_n53_), .Y(ori_ori_n593_));
  NA2        o0544(.A(ori_ori_n217_), .B(ori_ori_n57_), .Y(ori_ori_n594_));
  OAI210     o0545(.A0(ori_ori_n593_), .A1(ori_ori_n449_), .B0(ori_ori_n594_), .Y(ori_ori_n595_));
  NO3        o0546(.A(ori_ori_n595_), .B(ori_ori_n488_), .C(ori_ori_n59_), .Y(ori_ori_n596_));
  AO210      o0547(.A0(ori_ori_n592_), .A1(ori_ori_n461_), .B0(ori_ori_n596_), .Y(ori_ori_n597_));
  AOI210     o0548(.A0(ori_ori_n583_), .A1(ori_ori_n545_), .B0(ori_ori_n597_), .Y(ori05));
  AOI210     o0549(.A0(ori_ori_n162_), .A1(ori_ori_n55_), .B0(ori_ori_n504_), .Y(ori_ori_n599_));
  OR2        o0550(.A(ori_ori_n599_), .B(ori_ori_n57_), .Y(ori_ori_n600_));
  NO2        o0551(.A(x7), .B(ori_ori_n104_), .Y(ori_ori_n601_));
  NO2        o0552(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n602_));
  NA2        o0553(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n603_));
  NO2        o0554(.A(ori_ori_n603_), .B(ori_ori_n576_), .Y(ori_ori_n604_));
  AOI210     o0555(.A0(ori_ori_n602_), .A1(ori_ori_n601_), .B0(ori_ori_n604_), .Y(ori_ori_n605_));
  AOI210     o0556(.A0(ori_ori_n605_), .A1(ori_ori_n600_), .B0(ori_ori_n106_), .Y(ori_ori_n606_));
  NO2        o0557(.A(x7), .B(x4), .Y(ori_ori_n607_));
  NO2        o0558(.A(ori_ori_n64_), .B(ori_ori_n55_), .Y(ori_ori_n608_));
  NO2        o0559(.A(ori_ori_n195_), .B(x5), .Y(ori_ori_n609_));
  NA2        o0560(.A(ori_ori_n104_), .B(ori_ori_n106_), .Y(ori_ori_n610_));
  NO2        o0561(.A(ori_ori_n610_), .B(ori_ori_n213_), .Y(ori_ori_n611_));
  AN2        o0562(.A(ori_ori_n609_), .B(ori_ori_n608_), .Y(ori_ori_n612_));
  OAI210     o0563(.A0(ori_ori_n612_), .A1(ori_ori_n606_), .B0(ori_ori_n492_), .Y(ori_ori_n613_));
  NO2        o0564(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n614_));
  NA2        o0565(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n615_));
  NO2        o0566(.A(ori_ori_n104_), .B(ori_ori_n106_), .Y(ori_ori_n616_));
  NA2        o0567(.A(ori_ori_n616_), .B(x7), .Y(ori_ori_n617_));
  NA2        o0568(.A(ori_ori_n433_), .B(ori_ori_n252_), .Y(ori_ori_n618_));
  AOI210     o0569(.A0(ori_ori_n618_), .A1(ori_ori_n617_), .B0(ori_ori_n615_), .Y(ori_ori_n619_));
  NA2        o0570(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n620_));
  XO2        o0571(.A(x7), .B(x5), .Y(ori_ori_n621_));
  NO2        o0572(.A(ori_ori_n621_), .B(ori_ori_n53_), .Y(ori_ori_n622_));
  NA3        o0573(.A(ori_ori_n622_), .B(ori_ori_n620_), .C(ori_ori_n326_), .Y(ori_ori_n623_));
  NO2        o0574(.A(ori_ori_n104_), .B(x2), .Y(ori_ori_n624_));
  NO2        o0575(.A(ori_ori_n75_), .B(ori_ori_n55_), .Y(ori_ori_n625_));
  NA2        o0576(.A(ori_ori_n625_), .B(ori_ori_n624_), .Y(ori_ori_n626_));
  NA2        o0577(.A(ori_ori_n626_), .B(ori_ori_n623_), .Y(ori_ori_n627_));
  OAI210     o0578(.A0(ori_ori_n627_), .A1(ori_ori_n619_), .B0(ori_ori_n614_), .Y(ori_ori_n628_));
  NO2        o0579(.A(ori_ori_n71_), .B(ori_ori_n50_), .Y(ori_ori_n629_));
  NO2        o0580(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n630_));
  XO2        o0581(.A(x5), .B(x2), .Y(ori_ori_n631_));
  NO3        o0582(.A(x8), .B(x7), .C(ori_ori_n106_), .Y(ori_ori_n632_));
  NA2        o0583(.A(ori_ori_n267_), .B(ori_ori_n585_), .Y(ori_ori_n633_));
  NOi21      o0584(.An(x4), .B(x1), .Y(ori_ori_n634_));
  NA2        o0585(.A(ori_ori_n634_), .B(ori_ori_n63_), .Y(ori_ori_n635_));
  NA2        o0586(.A(x4), .B(x1), .Y(ori_ori_n636_));
  NO2        o0587(.A(ori_ori_n636_), .B(ori_ori_n50_), .Y(ori_ori_n637_));
  AOI210     o0588(.A0(ori_ori_n637_), .A1(ori_ori_n616_), .B0(ori_ori_n59_), .Y(ori_ori_n638_));
  OA210      o0589(.A0(ori_ori_n635_), .A1(ori_ori_n633_), .B0(ori_ori_n638_), .Y(ori_ori_n639_));
  NA3        o0590(.A(ori_ori_n639_), .B(ori_ori_n628_), .C(ori_ori_n613_), .Y(ori_ori_n640_));
  NA2        o0591(.A(ori_ori_n629_), .B(ori_ori_n56_), .Y(ori_ori_n641_));
  NA2        o0592(.A(ori_ori_n564_), .B(ori_ori_n601_), .Y(ori_ori_n642_));
  NO2        o0593(.A(ori_ori_n642_), .B(ori_ori_n641_), .Y(ori_ori_n643_));
  NA2        o0594(.A(ori_ori_n270_), .B(ori_ori_n119_), .Y(ori_ori_n644_));
  OAI210     o0595(.A0(ori_ori_n644_), .A1(ori_ori_n164_), .B0(ori_ori_n59_), .Y(ori_ori_n645_));
  NA2        o0596(.A(ori_ori_n57_), .B(x6), .Y(ori_ori_n646_));
  NA2        o0597(.A(ori_ori_n646_), .B(x3), .Y(ori_ori_n647_));
  NA2        o0598(.A(ori_ori_n630_), .B(ori_ori_n154_), .Y(ori_ori_n648_));
  NO3        o0599(.A(ori_ori_n648_), .B(ori_ori_n647_), .C(ori_ori_n423_), .Y(ori_ori_n649_));
  NA2        o0600(.A(ori_ori_n279_), .B(ori_ori_n71_), .Y(ori_ori_n650_));
  NO2        o0601(.A(ori_ori_n384_), .B(x3), .Y(ori_ori_n651_));
  NA2        o0602(.A(ori_ori_n651_), .B(ori_ori_n236_), .Y(ori_ori_n652_));
  INV        o0603(.A(ori_ori_n423_), .Y(ori_ori_n653_));
  NO2        o0604(.A(ori_ori_n465_), .B(ori_ori_n104_), .Y(ori_ori_n654_));
  NO2        o0605(.A(ori_ori_n574_), .B(x6), .Y(ori_ori_n655_));
  NA2        o0606(.A(ori_ori_n655_), .B(ori_ori_n654_), .Y(ori_ori_n656_));
  OAI220     o0607(.A0(ori_ori_n656_), .A1(ori_ori_n653_), .B0(ori_ori_n652_), .B1(ori_ori_n650_), .Y(ori_ori_n657_));
  NO4        o0608(.A(ori_ori_n657_), .B(ori_ori_n649_), .C(ori_ori_n645_), .D(ori_ori_n643_), .Y(ori_ori_n658_));
  NA2        o0609(.A(ori_ori_n57_), .B(x5), .Y(ori_ori_n659_));
  NO2        o0610(.A(ori_ori_n659_), .B(x1), .Y(ori_ori_n660_));
  NA2        o0611(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n661_));
  NO2        o0612(.A(ori_ori_n661_), .B(ori_ori_n128_), .Y(ori_ori_n662_));
  NA2        o0613(.A(x8), .B(x4), .Y(ori_ori_n663_));
  NO2        o0614(.A(x8), .B(x4), .Y(ori_ori_n664_));
  NAi21      o0615(.An(ori_ori_n664_), .B(ori_ori_n663_), .Y(ori_ori_n665_));
  NAi21      o0616(.An(ori_ori_n564_), .B(ori_ori_n384_), .Y(ori_ori_n666_));
  NO4        o0617(.A(ori_ori_n666_), .B(ori_ori_n665_), .C(ori_ori_n423_), .D(ori_ori_n71_), .Y(ori_ori_n667_));
  OAI210     o0618(.A0(ori_ori_n667_), .A1(ori_ori_n662_), .B0(ori_ori_n660_), .Y(ori_ori_n668_));
  NO3        o0619(.A(x8), .B(ori_ori_n104_), .C(x4), .Y(ori_ori_n669_));
  INV        o0620(.A(ori_ori_n669_), .Y(ori_ori_n670_));
  NO2        o0621(.A(ori_ori_n670_), .B(ori_ori_n106_), .Y(ori_ori_n671_));
  NO2        o0622(.A(x5), .B(x4), .Y(ori_ori_n672_));
  NA3        o0623(.A(ori_ori_n672_), .B(ori_ori_n63_), .C(ori_ori_n106_), .Y(ori_ori_n673_));
  NO2        o0624(.A(x6), .B(ori_ori_n106_), .Y(ori_ori_n674_));
  NA2        o0625(.A(ori_ori_n661_), .B(ori_ori_n674_), .Y(ori_ori_n675_));
  OAI210     o0626(.A0(ori_ori_n675_), .A1(ori_ori_n523_), .B0(ori_ori_n673_), .Y(ori_ori_n676_));
  OAI210     o0627(.A0(ori_ori_n676_), .A1(ori_ori_n671_), .B0(ori_ori_n309_), .Y(ori_ori_n677_));
  NA3        o0628(.A(ori_ori_n677_), .B(ori_ori_n668_), .C(ori_ori_n658_), .Y(ori_ori_n678_));
  OR2        o0629(.A(x4), .B(x1), .Y(ori_ori_n679_));
  NO2        o0630(.A(ori_ori_n679_), .B(x3), .Y(ori_ori_n680_));
  NA2        o0631(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n681_));
  NO3        o0632(.A(ori_ori_n365_), .B(ori_ori_n681_), .C(x6), .Y(ori_ori_n682_));
  AOI220     o0633(.A0(ori_ori_n682_), .A1(ori_ori_n680_), .B0(ori_ori_n678_), .B1(ori_ori_n640_), .Y(ori06));
  NA2        o0634(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n684_));
  NA2        o0635(.A(x6), .B(ori_ori_n106_), .Y(ori_ori_n685_));
  NA2        o0636(.A(ori_ori_n685_), .B(ori_ori_n55_), .Y(ori_ori_n686_));
  NA2        o0637(.A(x5), .B(ori_ori_n59_), .Y(ori_ori_n687_));
  NO2        o0638(.A(ori_ori_n687_), .B(ori_ori_n114_), .Y(ori_ori_n688_));
  NA3        o0639(.A(ori_ori_n688_), .B(ori_ori_n686_), .C(ori_ori_n498_), .Y(ori_ori_n689_));
  NO2        o0640(.A(ori_ori_n384_), .B(x0), .Y(ori_ori_n690_));
  NA2        o0641(.A(ori_ori_n336_), .B(x2), .Y(ori_ori_n691_));
  NOi21      o0642(.An(x6), .B(x8), .Y(ori_ori_n692_));
  NA2        o0643(.A(ori_ori_n690_), .B(ori_ori_n328_), .Y(ori_ori_n693_));
  AOI210     o0644(.A0(ori_ori_n693_), .A1(ori_ori_n689_), .B0(ori_ori_n684_), .Y(ori_ori_n694_));
  NA2        o0645(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n695_));
  NA2        o0646(.A(ori_ori_n363_), .B(ori_ori_n352_), .Y(ori_ori_n696_));
  NO2        o0647(.A(ori_ori_n71_), .B(ori_ori_n104_), .Y(ori_ori_n697_));
  NO2        o0648(.A(ori_ori_n53_), .B(ori_ori_n59_), .Y(ori_ori_n698_));
  NO4        o0649(.A(ori_ori_n698_), .B(ori_ori_n681_), .C(ori_ori_n697_), .D(ori_ori_n492_), .Y(ori_ori_n699_));
  AOI220     o0650(.A0(ori_ori_n699_), .A1(ori_ori_n696_), .B0(ori_ori_n420_), .B1(ori_ori_n63_), .Y(ori_ori_n700_));
  NO2        o0651(.A(ori_ori_n700_), .B(ori_ori_n695_), .Y(ori_ori_n701_));
  NO2        o0652(.A(ori_ori_n54_), .B(x0), .Y(ori_ori_n702_));
  NA2        o0653(.A(x4), .B(x3), .Y(ori_ori_n703_));
  OAI210     o0654(.A0(ori_ori_n703_), .A1(x8), .B0(ori_ori_n516_), .Y(ori_ori_n704_));
  NA2        o0655(.A(ori_ori_n704_), .B(ori_ori_n702_), .Y(ori_ori_n705_));
  NO2        o0656(.A(ori_ori_n100_), .B(ori_ori_n56_), .Y(ori_ori_n706_));
  NA3        o0657(.A(ori_ori_n706_), .B(ori_ori_n253_), .C(ori_ori_n404_), .Y(ori_ori_n707_));
  AOI210     o0658(.A0(ori_ori_n707_), .A1(ori_ori_n705_), .B0(x2), .Y(ori_ori_n708_));
  INV        o0659(.A(ori_ori_n380_), .Y(ori_ori_n709_));
  NO2        o0660(.A(ori_ori_n407_), .B(x8), .Y(ori_ori_n710_));
  NO2        o0661(.A(ori_ori_n254_), .B(ori_ori_n518_), .Y(ori_ori_n711_));
  AOI210     o0662(.A0(ori_ori_n710_), .A1(ori_ori_n262_), .B0(ori_ori_n711_), .Y(ori_ori_n712_));
  NO2        o0663(.A(x5), .B(x3), .Y(ori_ori_n713_));
  NA3        o0664(.A(ori_ori_n551_), .B(ori_ori_n713_), .C(x1), .Y(ori_ori_n714_));
  OR2        o0665(.A(ori_ori_n714_), .B(ori_ori_n498_), .Y(ori_ori_n715_));
  OAI210     o0666(.A0(ori_ori_n712_), .A1(ori_ori_n709_), .B0(ori_ori_n715_), .Y(ori_ori_n716_));
  OR4        o0667(.A(ori_ori_n716_), .B(ori_ori_n708_), .C(ori_ori_n701_), .D(ori_ori_n694_), .Y(ori_ori_n717_));
  NA2        o0668(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n718_));
  NO2        o0669(.A(ori_ori_n616_), .B(ori_ori_n59_), .Y(ori_ori_n719_));
  NO2        o0670(.A(ori_ori_n169_), .B(x6), .Y(ori_ori_n720_));
  AN2        o0671(.A(ori_ori_n470_), .B(ori_ori_n318_), .Y(ori_ori_n721_));
  NA2        o0672(.A(ori_ori_n721_), .B(ori_ori_n347_), .Y(ori_ori_n722_));
  NO2        o0673(.A(ori_ori_n305_), .B(ori_ori_n104_), .Y(ori_ori_n723_));
  NO2        o0674(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n724_));
  NA2        o0675(.A(ori_ori_n724_), .B(ori_ori_n71_), .Y(ori_ori_n725_));
  NO2        o0676(.A(ori_ori_n725_), .B(ori_ori_n248_), .Y(ori_ori_n726_));
  NO2        o0677(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n727_));
  NA3        o0678(.A(ori_ori_n727_), .B(ori_ori_n571_), .C(ori_ori_n56_), .Y(ori_ori_n728_));
  NO2        o0679(.A(ori_ori_n57_), .B(x6), .Y(ori_ori_n729_));
  NA2        o0680(.A(ori_ori_n179_), .B(ori_ori_n729_), .Y(ori_ori_n730_));
  NA3        o0681(.A(ori_ori_n602_), .B(ori_ori_n325_), .C(ori_ori_n71_), .Y(ori_ori_n731_));
  NA3        o0682(.A(ori_ori_n731_), .B(ori_ori_n730_), .C(ori_ori_n728_), .Y(ori_ori_n732_));
  OR3        o0683(.A(ori_ori_n732_), .B(ori_ori_n726_), .C(ori_ori_n637_), .Y(ori_ori_n733_));
  NA2        o0684(.A(ori_ori_n733_), .B(ori_ori_n723_), .Y(ori_ori_n734_));
  NA2        o0685(.A(ori_ori_n702_), .B(ori_ori_n629_), .Y(ori_ori_n735_));
  NA3        o0686(.A(ori_ori_n586_), .B(ori_ori_n217_), .C(ori_ori_n255_), .Y(ori_ori_n736_));
  NA2        o0687(.A(ori_ori_n481_), .B(ori_ori_n67_), .Y(ori_ori_n737_));
  AOI210     o0688(.A0(ori_ori_n736_), .A1(ori_ori_n735_), .B0(ori_ori_n737_), .Y(ori_ori_n738_));
  NA2        o0689(.A(x7), .B(x6), .Y(ori_ori_n739_));
  NA3        o0690(.A(x2), .B(x1), .C(x0), .Y(ori_ori_n740_));
  NO3        o0691(.A(ori_ori_n740_), .B(ori_ori_n739_), .C(ori_ori_n599_), .Y(ori_ori_n741_));
  NA2        o0692(.A(ori_ori_n493_), .B(ori_ori_n147_), .Y(ori_ori_n742_));
  NO2        o0693(.A(x5), .B(x1), .Y(ori_ori_n743_));
  NA2        o0694(.A(ori_ori_n743_), .B(ori_ori_n729_), .Y(ori_ori_n744_));
  NA2        o0695(.A(x4), .B(x0), .Y(ori_ori_n745_));
  NO3        o0696(.A(ori_ori_n57_), .B(x6), .C(x2), .Y(ori_ori_n746_));
  NA2        o0697(.A(ori_ori_n746_), .B(ori_ori_n221_), .Y(ori_ori_n747_));
  NO2        o0698(.A(ori_ori_n747_), .B(ori_ori_n745_), .Y(ori_ori_n748_));
  NO3        o0699(.A(ori_ori_n748_), .B(ori_ori_n741_), .C(ori_ori_n738_), .Y(ori_ori_n749_));
  NA3        o0700(.A(ori_ori_n749_), .B(ori_ori_n734_), .C(ori_ori_n722_), .Y(ori_ori_n750_));
  AOI210     o0701(.A0(ori_ori_n717_), .A1(ori_ori_n57_), .B0(ori_ori_n750_), .Y(ori07));
  NA2        o0702(.A(ori_ori_n104_), .B(ori_ori_n59_), .Y(ori_ori_n752_));
  NOi21      o0703(.An(ori_ori_n739_), .B(ori_ori_n112_), .Y(ori_ori_n753_));
  NO4        o0704(.A(ori_ori_n753_), .B(ori_ori_n629_), .C(ori_ori_n248_), .D(ori_ori_n752_), .Y(ori_ori_n754_));
  NO3        o0705(.A(ori_ori_n57_), .B(x5), .C(x1), .Y(ori_ori_n755_));
  NA2        o0706(.A(ori_ori_n755_), .B(ori_ori_n371_), .Y(ori_ori_n756_));
  NO2        o0707(.A(ori_ori_n57_), .B(ori_ori_n71_), .Y(ori_ori_n757_));
  NO2        o0708(.A(ori_ori_n153_), .B(ori_ori_n105_), .Y(ori_ori_n758_));
  INV        o0709(.A(ori_ori_n758_), .Y(ori_ori_n759_));
  NO2        o0710(.A(ori_ori_n759_), .B(ori_ori_n133_), .Y(ori_ori_n760_));
  OAI210     o0711(.A0(ori_ori_n760_), .A1(ori_ori_n754_), .B0(x2), .Y(ori_ori_n761_));
  NAi21      o0712(.An(ori_ori_n154_), .B(ori_ori_n155_), .Y(ori_ori_n762_));
  NA3        o0713(.A(ori_ori_n762_), .B(ori_ori_n89_), .C(x3), .Y(ori_ori_n763_));
  NO3        o0714(.A(ori_ori_n55_), .B(x3), .C(x1), .Y(ori_ori_n764_));
  NO2        o0715(.A(ori_ori_n511_), .B(x2), .Y(ori_ori_n765_));
  AOI210     o0716(.A0(ori_ori_n765_), .A1(ori_ori_n513_), .B0(ori_ori_n764_), .Y(ori_ori_n766_));
  OAI210     o0717(.A0(ori_ori_n766_), .A1(ori_ori_n646_), .B0(ori_ori_n763_), .Y(ori_ori_n767_));
  NO2        o0718(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n768_));
  NA2        o0719(.A(ori_ori_n768_), .B(ori_ori_n59_), .Y(ori_ori_n769_));
  NA2        o0720(.A(ori_ori_n353_), .B(ori_ori_n347_), .Y(ori_ori_n770_));
  NO2        o0721(.A(x7), .B(x3), .Y(ori_ori_n771_));
  NA2        o0722(.A(ori_ori_n771_), .B(ori_ori_n97_), .Y(ori_ori_n772_));
  NO2        o0723(.A(ori_ori_n769_), .B(ori_ori_n772_), .Y(ori_ori_n773_));
  AOI210     o0724(.A0(ori_ori_n767_), .A1(ori_ori_n247_), .B0(ori_ori_n773_), .Y(ori_ori_n774_));
  AOI210     o0725(.A0(ori_ori_n774_), .A1(ori_ori_n761_), .B0(x4), .Y(ori_ori_n775_));
  NO2        o0726(.A(ori_ori_n595_), .B(ori_ori_n106_), .Y(ori_ori_n776_));
  XO2        o0727(.A(x5), .B(x1), .Y(ori_ori_n777_));
  NO4        o0728(.A(ori_ori_n777_), .B(ori_ori_n163_), .C(ori_ori_n204_), .D(ori_ori_n55_), .Y(ori_ori_n778_));
  OAI210     o0729(.A0(ori_ori_n778_), .A1(ori_ori_n776_), .B0(ori_ori_n411_), .Y(ori_ori_n779_));
  NO3        o0730(.A(ori_ori_n50_), .B(x2), .C(x0), .Y(ori_ori_n780_));
  NO2        o0731(.A(ori_ori_n308_), .B(ori_ori_n104_), .Y(ori_ori_n781_));
  NA2        o0732(.A(x6), .B(x0), .Y(ori_ori_n782_));
  NO2        o0733(.A(ori_ori_n681_), .B(ori_ori_n782_), .Y(ori_ori_n783_));
  INV        o0734(.A(ori_ori_n777_), .Y(ori_ori_n784_));
  NA2        o0735(.A(ori_ori_n63_), .B(ori_ori_n57_), .Y(ori_ori_n785_));
  OAI210     o0736(.A0(ori_ori_n785_), .A1(ori_ori_n784_), .B0(ori_ori_n756_), .Y(ori_ori_n786_));
  AOI220     o0737(.A0(ori_ori_n786_), .A1(ori_ori_n780_), .B0(ori_ori_n783_), .B1(ori_ori_n781_), .Y(ori_ori_n787_));
  AOI210     o0738(.A0(ori_ori_n787_), .A1(ori_ori_n779_), .B0(ori_ori_n56_), .Y(ori_ori_n788_));
  NOi21      o0739(.An(ori_ori_n228_), .B(ori_ori_n371_), .Y(ori_ori_n789_));
  NO3        o0740(.A(ori_ori_n789_), .B(ori_ori_n237_), .C(ori_ori_n67_), .Y(ori_ori_n790_));
  NO2        o0741(.A(ori_ori_n187_), .B(ori_ori_n71_), .Y(ori_ori_n791_));
  NO2        o0742(.A(ori_ori_n308_), .B(x6), .Y(ori_ori_n792_));
  AO220      o0743(.A0(ori_ori_n792_), .A1(ori_ori_n326_), .B0(ori_ori_n791_), .B1(ori_ori_n556_), .Y(ori_ori_n793_));
  OAI210     o0744(.A0(ori_ori_n793_), .A1(ori_ori_n790_), .B0(ori_ori_n59_), .Y(ori_ori_n794_));
  NA2        o0745(.A(ori_ori_n90_), .B(ori_ori_n71_), .Y(ori_ori_n795_));
  NO2        o0746(.A(ori_ori_n795_), .B(ori_ori_n642_), .Y(ori_ori_n796_));
  NAi21      o0747(.An(x8), .B(x7), .Y(ori_ori_n797_));
  NA2        o0748(.A(ori_ori_n789_), .B(ori_ori_n797_), .Y(ori_ori_n798_));
  NA2        o0749(.A(ori_ori_n404_), .B(ori_ori_n106_), .Y(ori_ori_n799_));
  NO2        o0750(.A(ori_ori_n692_), .B(x1), .Y(ori_ori_n800_));
  NO3        o0751(.A(ori_ori_n800_), .B(ori_ori_n799_), .C(ori_ori_n571_), .Y(ori_ori_n801_));
  AOI210     o0752(.A0(ori_ori_n801_), .A1(ori_ori_n798_), .B0(ori_ori_n796_), .Y(ori_ori_n802_));
  AOI210     o0753(.A0(ori_ori_n802_), .A1(ori_ori_n794_), .B0(ori_ori_n140_), .Y(ori_ori_n803_));
  NO2        o0754(.A(x8), .B(x7), .Y(ori_ori_n804_));
  NO2        o0755(.A(ori_ori_n804_), .B(x3), .Y(ori_ori_n805_));
  NA3        o0756(.A(ori_ori_n805_), .B(ori_ori_n361_), .C(x1), .Y(ori_ori_n806_));
  NO2        o0757(.A(x8), .B(ori_ori_n106_), .Y(ori_ori_n807_));
  AOI220     o0758(.A0(ori_ori_n325_), .A1(ori_ori_n347_), .B0(ori_ori_n807_), .B1(ori_ori_n252_), .Y(ori_ori_n808_));
  NO2        o0759(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n809_));
  NA2        o0760(.A(ori_ori_n809_), .B(ori_ori_n302_), .Y(ori_ori_n810_));
  AOI210     o0761(.A0(ori_ori_n808_), .A1(ori_ori_n806_), .B0(ori_ori_n810_), .Y(ori_ori_n811_));
  NO4        o0762(.A(ori_ori_n811_), .B(ori_ori_n803_), .C(ori_ori_n788_), .D(ori_ori_n775_), .Y(ori08));
  NA2        o0763(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n813_));
  XN2        o0764(.A(x5), .B(x4), .Y(ori_ori_n814_));
  INV        o0765(.A(ori_ori_n814_), .Y(ori_ori_n815_));
  AOI220     o0766(.A0(ori_ori_n815_), .A1(ori_ori_n353_), .B0(ori_ori_n136_), .B1(ori_ori_n56_), .Y(ori_ori_n816_));
  NO2        o0767(.A(ori_ori_n239_), .B(ori_ori_n104_), .Y(ori_ori_n817_));
  AOI210     o0768(.A0(ori_ori_n817_), .A1(ori_ori_n276_), .B0(ori_ori_n188_), .Y(ori_ori_n818_));
  OAI220     o0769(.A0(ori_ori_n818_), .A1(x4), .B0(ori_ori_n816_), .B1(ori_ori_n813_), .Y(ori_ori_n819_));
  NA2        o0770(.A(ori_ori_n819_), .B(ori_ori_n270_), .Y(ori_ori_n820_));
  AOI210     o0771(.A0(ori_ori_n269_), .A1(ori_ori_n799_), .B0(ori_ori_n615_), .Y(ori_ori_n821_));
  NA2        o0772(.A(ori_ori_n610_), .B(ori_ori_n169_), .Y(ori_ori_n822_));
  OAI220     o0773(.A0(ori_ori_n822_), .A1(ori_ori_n661_), .B0(ori_ori_n483_), .B1(ori_ori_n50_), .Y(ori_ori_n823_));
  AO210      o0774(.A0(ori_ori_n823_), .A1(ori_ori_n340_), .B0(ori_ori_n821_), .Y(ori_ori_n824_));
  NA2        o0775(.A(ori_ori_n276_), .B(ori_ori_n147_), .Y(ori_ori_n825_));
  NA2        o0776(.A(ori_ori_n140_), .B(x7), .Y(ori_ori_n826_));
  OR3        o0777(.A(ori_ori_n740_), .B(ori_ori_n465_), .C(ori_ori_n713_), .Y(ori_ori_n827_));
  OAI220     o0778(.A0(ori_ori_n827_), .A1(ori_ori_n826_), .B0(ori_ori_n825_), .B1(ori_ori_n201_), .Y(ori_ori_n828_));
  AOI210     o0779(.A0(ori_ori_n824_), .A1(ori_ori_n290_), .B0(ori_ori_n828_), .Y(ori_ori_n829_));
  AOI210     o0780(.A0(ori_ori_n829_), .A1(ori_ori_n820_), .B0(ori_ori_n71_), .Y(ori_ori_n830_));
  NO2        o0781(.A(ori_ori_n804_), .B(ori_ori_n106_), .Y(ori_ori_n831_));
  NA2        o0782(.A(ori_ori_n831_), .B(ori_ori_n189_), .Y(ori_ori_n832_));
  OAI210     o0783(.A0(ori_ori_n407_), .A1(ori_ori_n302_), .B0(ori_ori_n340_), .Y(ori_ori_n833_));
  NA2        o0784(.A(ori_ori_n433_), .B(ori_ori_n230_), .Y(ori_ori_n834_));
  NA2        o0785(.A(ori_ori_n710_), .B(ori_ori_n103_), .Y(ori_ori_n835_));
  OAI220     o0786(.A0(ori_ori_n835_), .A1(ori_ori_n834_), .B0(ori_ori_n833_), .B1(ori_ori_n832_), .Y(ori_ori_n836_));
  NA2        o0787(.A(ori_ori_n836_), .B(ori_ori_n286_), .Y(ori_ori_n837_));
  NA2        o0788(.A(ori_ori_n330_), .B(ori_ori_n53_), .Y(ori_ori_n838_));
  NO3        o0789(.A(ori_ori_n407_), .B(ori_ori_n133_), .C(ori_ori_n68_), .Y(ori_ori_n839_));
  NO2        o0790(.A(ori_ori_n698_), .B(ori_ori_n242_), .Y(ori_ori_n840_));
  NO3        o0791(.A(ori_ori_n565_), .B(ori_ori_n466_), .C(ori_ori_n95_), .Y(ori_ori_n841_));
  AO220      o0792(.A0(ori_ori_n841_), .A1(ori_ori_n840_), .B0(ori_ori_n839_), .B1(ori_ori_n838_), .Y(ori_ori_n842_));
  NA2        o0793(.A(x7), .B(ori_ori_n59_), .Y(ori_ori_n843_));
  NO3        o0794(.A(ori_ori_n311_), .B(ori_ori_n843_), .C(ori_ori_n285_), .Y(ori_ori_n844_));
  AOI210     o0795(.A0(ori_ori_n842_), .A1(x5), .B0(ori_ori_n844_), .Y(ori_ori_n845_));
  AOI210     o0796(.A0(ori_ori_n845_), .A1(ori_ori_n837_), .B0(ori_ori_n72_), .Y(ori_ori_n846_));
  NO2        o0797(.A(ori_ori_n70_), .B(x3), .Y(ori_ori_n847_));
  OAI210     o0798(.A0(ori_ori_n847_), .A1(ori_ori_n261_), .B0(ori_ori_n145_), .Y(ori_ori_n848_));
  MUX2       o0799(.S(x3), .A(ori_ori_n163_), .B(ori_ori_n762_), .Y(ori_ori_n849_));
  NA2        o0800(.A(ori_ori_n849_), .B(ori_ori_n556_), .Y(ori_ori_n850_));
  NO3        o0801(.A(x6), .B(x4), .C(x0), .Y(ori_ori_n851_));
  INV        o0802(.A(ori_ori_n851_), .Y(ori_ori_n852_));
  AOI210     o0803(.A0(ori_ori_n850_), .A1(ori_ori_n848_), .B0(ori_ori_n852_), .Y(ori_ori_n853_));
  NO3        o0804(.A(x5), .B(x3), .C(ori_ori_n106_), .Y(ori_ori_n854_));
  AOI220     o0805(.A0(ori_ori_n815_), .A1(ori_ori_n307_), .B0(ori_ori_n854_), .B1(ori_ori_n59_), .Y(ori_ori_n855_));
  OR2        o0806(.A(x8), .B(x1), .Y(ori_ori_n856_));
  NO3        o0807(.A(ori_ori_n856_), .B(ori_ori_n855_), .C(ori_ori_n724_), .Y(ori_ori_n857_));
  NAi21      o0808(.An(x4), .B(x1), .Y(ori_ori_n858_));
  NO2        o0809(.A(ori_ori_n858_), .B(x0), .Y(ori_ori_n859_));
  NA2        o0810(.A(ori_ori_n609_), .B(ori_ori_n859_), .Y(ori_ori_n860_));
  NA3        o0811(.A(ori_ori_n55_), .B(x1), .C(x0), .Y(ori_ori_n861_));
  OAI210     o0812(.A0(ori_ori_n861_), .A1(ori_ori_n709_), .B0(ori_ori_n860_), .Y(ori_ori_n862_));
  OAI210     o0813(.A0(ori_ori_n862_), .A1(ori_ori_n857_), .B0(ori_ori_n316_), .Y(ori_ori_n863_));
  AO210      o0814(.A0(ori_ori_n288_), .A1(ori_ori_n261_), .B0(ori_ori_n723_), .Y(ori_ori_n864_));
  NA2        o0815(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n865_));
  NO2        o0816(.A(ori_ori_n57_), .B(x2), .Y(ori_ori_n866_));
  NA2        o0817(.A(ori_ori_n864_), .B(ori_ori_n637_), .Y(ori_ori_n867_));
  NA2        o0818(.A(ori_ori_n867_), .B(ori_ori_n863_), .Y(ori_ori_n868_));
  NO4        o0819(.A(ori_ori_n868_), .B(ori_ori_n853_), .C(ori_ori_n846_), .D(ori_ori_n830_), .Y(ori09));
  NO3        o0820(.A(ori_ori_n777_), .B(ori_ori_n117_), .C(ori_ori_n92_), .Y(ori_ori_n870_));
  AOI220     o0821(.A0(ori_ori_n297_), .A1(ori_ori_n70_), .B0(ori_ori_n585_), .B1(ori_ori_n538_), .Y(ori_ori_n871_));
  OAI210     o0822(.A0(ori_ori_n870_), .A1(x2), .B0(ori_ori_n871_), .Y(ori_ori_n872_));
  AOI210     o0823(.A0(ori_ori_n872_), .A1(ori_ori_n744_), .B0(ori_ori_n442_), .Y(ori_ori_n873_));
  NO2        o0824(.A(ori_ori_n584_), .B(ori_ori_n260_), .Y(ori_ori_n874_));
  NO2        o0825(.A(ori_ori_n743_), .B(ori_ori_n336_), .Y(ori_ori_n875_));
  NO3        o0826(.A(ori_ori_n601_), .B(ori_ori_n98_), .C(ori_ori_n106_), .Y(ori_ori_n876_));
  AO220      o0827(.A0(ori_ori_n876_), .A1(ori_ori_n875_), .B0(ori_ori_n874_), .B1(ori_ori_n616_), .Y(ori_ori_n877_));
  OAI210     o0828(.A0(ori_ori_n877_), .A1(ori_ori_n873_), .B0(x4), .Y(ori_ori_n878_));
  OAI220     o0829(.A0(ori_ori_n363_), .A1(ori_ori_n142_), .B0(ori_ori_n391_), .B1(ori_ori_n278_), .Y(ori_ori_n879_));
  NO2        o0830(.A(ori_ori_n187_), .B(ori_ori_n104_), .Y(ori_ori_n880_));
  AOI220     o0831(.A0(ori_ori_n880_), .A1(ori_ori_n122_), .B0(ori_ori_n879_), .B1(ori_ori_n622_), .Y(ori_ori_n881_));
  NO2        o0832(.A(ori_ori_n777_), .B(ori_ori_n92_), .Y(ori_ori_n882_));
  NAi21      o0833(.An(x0), .B(x2), .Y(ori_ori_n883_));
  NO2        o0834(.A(ori_ori_n301_), .B(ori_ori_n883_), .Y(ori_ori_n884_));
  OAI210     o0835(.A0(ori_ori_n475_), .A1(ori_ori_n273_), .B0(ori_ori_n187_), .Y(ori_ori_n885_));
  AOI210     o0836(.A0(ori_ori_n166_), .A1(ori_ori_n797_), .B0(ori_ori_n352_), .Y(ori_ori_n886_));
  AOI220     o0837(.A0(ori_ori_n886_), .A1(ori_ori_n885_), .B0(ori_ori_n884_), .B1(ori_ori_n882_), .Y(ori_ori_n887_));
  OAI210     o0838(.A0(ori_ori_n881_), .A1(ori_ori_n55_), .B0(ori_ori_n887_), .Y(ori_ori_n888_));
  NA2        o0839(.A(ori_ori_n888_), .B(ori_ori_n56_), .Y(ori_ori_n889_));
  NO2        o0840(.A(ori_ori_n56_), .B(ori_ori_n59_), .Y(ori_ori_n890_));
  INV        o0841(.A(ori_ori_n122_), .Y(ori_ori_n891_));
  NA2        o0842(.A(ori_ori_n743_), .B(ori_ori_n55_), .Y(ori_ori_n892_));
  AOI210     o0843(.A0(x6), .A1(x1), .B0(x5), .Y(ori_ori_n893_));
  OAI210     o0844(.A0(ori_ori_n893_), .A1(ori_ori_n329_), .B0(x2), .Y(ori_ori_n894_));
  AOI210     o0845(.A0(ori_ori_n894_), .A1(ori_ori_n892_), .B0(ori_ori_n891_), .Y(ori_ori_n895_));
  NA2        o0846(.A(ori_ori_n555_), .B(ori_ori_n55_), .Y(ori_ori_n896_));
  NO2        o0847(.A(ori_ori_n227_), .B(ori_ori_n381_), .Y(ori_ori_n897_));
  NO2        o0848(.A(ori_ori_n308_), .B(ori_ori_n146_), .Y(ori_ori_n898_));
  NO2        o0849(.A(ori_ori_n898_), .B(ori_ori_n897_), .Y(ori_ori_n899_));
  OAI220     o0850(.A0(ori_ori_n899_), .A1(ori_ori_n55_), .B0(ori_ori_n896_), .B1(ori_ori_n454_), .Y(ori_ori_n900_));
  OAI210     o0851(.A0(ori_ori_n900_), .A1(ori_ori_n895_), .B0(ori_ori_n890_), .Y(ori_ori_n901_));
  NO2        o0852(.A(ori_ori_n400_), .B(ori_ori_n104_), .Y(ori_ori_n902_));
  NO2        o0853(.A(ori_ori_n330_), .B(ori_ori_n492_), .Y(ori_ori_n903_));
  AOI220     o0854(.A0(ori_ori_n903_), .A1(ori_ori_n902_), .B0(ori_ori_n205_), .B1(ori_ori_n225_), .Y(ori_ori_n904_));
  NA4        o0855(.A(ori_ori_n904_), .B(ori_ori_n901_), .C(ori_ori_n889_), .D(ori_ori_n878_), .Y(ori_ori_n905_));
  NA2        o0856(.A(ori_ori_n905_), .B(ori_ori_n50_), .Y(ori_ori_n906_));
  NO2        o0857(.A(ori_ori_n374_), .B(ori_ori_n159_), .Y(ori_ori_n907_));
  NA2        o0858(.A(ori_ori_n236_), .B(ori_ori_n585_), .Y(ori_ori_n908_));
  OAI210     o0859(.A0(ori_ori_n428_), .A1(ori_ori_n807_), .B0(ori_ori_n908_), .Y(ori_ori_n909_));
  OAI210     o0860(.A0(ori_ori_n909_), .A1(ori_ori_n907_), .B0(x0), .Y(ori_ori_n910_));
  NO3        o0861(.A(x8), .B(x7), .C(x2), .Y(ori_ori_n911_));
  NO3        o0862(.A(ori_ori_n57_), .B(x5), .C(x2), .Y(ori_ori_n912_));
  OAI210     o0863(.A0(ori_ori_n912_), .A1(ori_ori_n911_), .B0(ori_ori_n513_), .Y(ori_ori_n913_));
  AOI210     o0864(.A0(ori_ori_n913_), .A1(ori_ori_n910_), .B0(x4), .Y(ori_ori_n914_));
  NO2        o0865(.A(ori_ori_n421_), .B(ori_ori_n145_), .Y(ori_ori_n915_));
  NO2        o0866(.A(ori_ori_n52_), .B(x2), .Y(ori_ori_n916_));
  NO2        o0867(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n917_));
  NA2        o0868(.A(ori_ori_n917_), .B(x8), .Y(ori_ori_n918_));
  NA2        o0869(.A(ori_ori_n918_), .B(ori_ori_n892_), .Y(ori_ori_n919_));
  AO210      o0870(.A0(ori_ori_n919_), .A1(ori_ori_n916_), .B0(ori_ori_n915_), .Y(ori_ori_n920_));
  OAI210     o0871(.A0(ori_ori_n920_), .A1(ori_ori_n914_), .B0(ori_ori_n614_), .Y(ori_ori_n921_));
  NO2        o0872(.A(ori_ori_n256_), .B(ori_ori_n115_), .Y(ori_ori_n922_));
  OAI210     o0873(.A0(x4), .A1(x2), .B0(x0), .Y(ori_ori_n923_));
  NA3        o0874(.A(ori_ori_n603_), .B(ori_ori_n615_), .C(ori_ori_n341_), .Y(ori_ori_n924_));
  OAI210     o0875(.A0(ori_ori_n923_), .A1(ori_ori_n285_), .B0(ori_ori_n53_), .Y(ori_ori_n925_));
  AOI210     o0876(.A0(ori_ori_n924_), .A1(ori_ori_n923_), .B0(ori_ori_n925_), .Y(ori_ori_n926_));
  OAI210     o0877(.A0(ori_ori_n926_), .A1(ori_ori_n922_), .B0(ori_ori_n325_), .Y(ori_ori_n927_));
  AOI220     o0878(.A0(ori_ori_n663_), .A1(ori_ori_n345_), .B0(ori_ori_n347_), .B1(ori_ori_n91_), .Y(ori_ori_n928_));
  NA2        o0879(.A(ori_ori_n91_), .B(x5), .Y(ori_ori_n929_));
  OAI220     o0880(.A0(ori_ori_n929_), .A1(ori_ori_n856_), .B0(ori_ori_n928_), .B1(ori_ori_n317_), .Y(ori_ori_n930_));
  NA2        o0881(.A(ori_ori_n930_), .B(ori_ori_n68_), .Y(ori_ori_n931_));
  NA2        o0882(.A(ori_ori_n404_), .B(ori_ori_n762_), .Y(ori_ori_n932_));
  NA2        o0883(.A(ori_ori_n247_), .B(ori_ori_n163_), .Y(ori_ori_n933_));
  AO210      o0884(.A0(ori_ori_n933_), .A1(ori_ori_n932_), .B0(ori_ori_n130_), .Y(ori_ori_n934_));
  NO2        o0885(.A(ori_ori_n434_), .B(x2), .Y(ori_ori_n935_));
  NO2        o0886(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n936_));
  NA2        o0887(.A(ori_ori_n936_), .B(x5), .Y(ori_ori_n937_));
  NO2        o0888(.A(ori_ori_n937_), .B(ori_ori_n60_), .Y(ori_ori_n938_));
  AOI220     o0889(.A0(ori_ori_n938_), .A1(ori_ori_n935_), .B0(ori_ori_n664_), .B1(ori_ori_n240_), .Y(ori_ori_n939_));
  NA4        o0890(.A(ori_ori_n939_), .B(ori_ori_n934_), .C(ori_ori_n931_), .D(ori_ori_n927_), .Y(ori_ori_n940_));
  NO4        o0891(.A(ori_ori_n924_), .B(ori_ori_n630_), .C(ori_ori_n454_), .D(ori_ori_n50_), .Y(ori_ori_n941_));
  AOI220     o0892(.A0(ori_ori_n602_), .A1(ori_ori_n601_), .B0(ori_ori_n279_), .B1(x5), .Y(ori_ori_n942_));
  NO2        o0893(.A(ori_ori_n672_), .B(ori_ori_n187_), .Y(ori_ori_n943_));
  NA3        o0894(.A(ori_ori_n943_), .B(ori_ori_n665_), .C(x7), .Y(ori_ori_n944_));
  OAI210     o0895(.A0(ori_ori_n942_), .A1(ori_ori_n346_), .B0(ori_ori_n944_), .Y(ori_ori_n945_));
  OAI210     o0896(.A0(ori_ori_n945_), .A1(ori_ori_n941_), .B0(ori_ori_n82_), .Y(ori_ori_n946_));
  NA2        o0897(.A(ori_ori_n768_), .B(x2), .Y(ori_ori_n947_));
  NO2        o0898(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n948_));
  NAi21      o0899(.An(x1), .B(x4), .Y(ori_ori_n949_));
  NA2        o0900(.A(ori_ori_n949_), .B(ori_ori_n858_), .Y(ori_ori_n950_));
  NA3        o0901(.A(ori_ori_n394_), .B(ori_ori_n743_), .C(ori_ori_n57_), .Y(ori_ori_n951_));
  NA2        o0902(.A(ori_ori_n951_), .B(ori_ori_n946_), .Y(ori_ori_n952_));
  AOI210     o0903(.A0(ori_ori_n940_), .A1(x6), .B0(ori_ori_n952_), .Y(ori_ori_n953_));
  NA3        o0904(.A(ori_ori_n953_), .B(ori_ori_n921_), .C(ori_ori_n906_), .Y(ori10));
  NO2        o0905(.A(x4), .B(x1), .Y(ori_ori_n955_));
  NO2        o0906(.A(ori_ori_n955_), .B(ori_ori_n147_), .Y(ori_ori_n956_));
  NA3        o0907(.A(x5), .B(x4), .C(x0), .Y(ori_ori_n957_));
  OAI220     o0908(.A0(ori_ori_n957_), .A1(ori_ori_n274_), .B0(ori_ori_n698_), .B1(ori_ori_n244_), .Y(ori_ori_n958_));
  NA2        o0909(.A(ori_ori_n958_), .B(ori_ori_n956_), .Y(ori_ori_n959_));
  NO3        o0910(.A(ori_ori_n353_), .B(ori_ori_n317_), .C(ori_ori_n90_), .Y(ori_ori_n960_));
  NA3        o0911(.A(ori_ori_n960_), .B(ori_ori_n379_), .C(ori_ori_n62_), .Y(ori_ori_n961_));
  AOI210     o0912(.A0(ori_ori_n961_), .A1(ori_ori_n959_), .B0(ori_ori_n301_), .Y(ori_ori_n962_));
  NOi21      o0913(.An(ori_ori_n255_), .B(ori_ori_n136_), .Y(ori_ori_n963_));
  AOI210     o0914(.A0(ori_ori_n499_), .A1(ori_ori_n616_), .B0(ori_ori_n326_), .Y(ori_ori_n964_));
  NO2        o0915(.A(ori_ori_n890_), .B(ori_ori_n339_), .Y(ori_ori_n965_));
  NOi31      o0916(.An(ori_ori_n965_), .B(ori_ori_n964_), .C(ori_ori_n963_), .Y(ori_ori_n966_));
  NA2        o0917(.A(x4), .B(ori_ori_n106_), .Y(ori_ori_n967_));
  NO2        o0918(.A(ori_ori_n320_), .B(ori_ori_n967_), .Y(ori_ori_n968_));
  NA2        o0919(.A(ori_ori_n95_), .B(x5), .Y(ori_ori_n969_));
  NO3        o0920(.A(ori_ori_n969_), .B(ori_ori_n107_), .C(ori_ori_n55_), .Y(ori_ori_n970_));
  NO3        o0921(.A(ori_ori_n970_), .B(ori_ori_n968_), .C(ori_ori_n966_), .Y(ori_ori_n971_));
  NA2        o0922(.A(ori_ori_n948_), .B(ori_ori_n50_), .Y(ori_ori_n972_));
  NA2        o0923(.A(ori_ori_n602_), .B(ori_ori_n268_), .Y(ori_ori_n973_));
  NO2        o0924(.A(ori_ori_n973_), .B(ori_ori_n972_), .Y(ori_ori_n974_));
  OAI220     o0925(.A0(ori_ori_n918_), .A1(ori_ori_n103_), .B0(ori_ori_n865_), .B1(ori_ori_n442_), .Y(ori_ori_n975_));
  AOI210     o0926(.A0(ori_ori_n975_), .A1(ori_ori_n276_), .B0(ori_ori_n974_), .Y(ori_ori_n976_));
  OAI210     o0927(.A0(ori_ori_n971_), .A1(ori_ori_n381_), .B0(ori_ori_n976_), .Y(ori_ori_n977_));
  OAI210     o0928(.A0(ori_ori_n977_), .A1(ori_ori_n962_), .B0(x7), .Y(ori_ori_n978_));
  NA2        o0929(.A(ori_ori_n55_), .B(ori_ori_n71_), .Y(ori_ori_n979_));
  AOI210     o0930(.A0(ori_ori_n442_), .A1(ori_ori_n352_), .B0(ori_ori_n967_), .Y(ori_ori_n980_));
  NO3        o0931(.A(ori_ori_n444_), .B(ori_ori_n883_), .C(x5), .Y(ori_ori_n981_));
  OAI210     o0932(.A0(ori_ori_n981_), .A1(ori_ori_n980_), .B0(ori_ori_n979_), .Y(ori_ori_n982_));
  NO2        o0933(.A(ori_ori_n353_), .B(ori_ori_n139_), .Y(ori_ori_n983_));
  NA2        o0934(.A(ori_ori_n983_), .B(ori_ori_n422_), .Y(ori_ori_n984_));
  AOI210     o0935(.A0(ori_ori_n984_), .A1(ori_ori_n982_), .B0(x3), .Y(ori_ori_n985_));
  NA2        o0936(.A(ori_ori_n692_), .B(ori_ori_n247_), .Y(ori_ori_n986_));
  NO2        o0937(.A(x5), .B(ori_ori_n106_), .Y(ori_ori_n987_));
  OAI210     o0938(.A0(ori_ori_n987_), .A1(ori_ori_n234_), .B0(ori_ori_n929_), .Y(ori_ori_n988_));
  NA3        o0939(.A(ori_ori_n461_), .B(ori_ori_n128_), .C(ori_ori_n422_), .Y(ori_ori_n989_));
  OAI210     o0940(.A0(ori_ori_n444_), .A1(ori_ori_n210_), .B0(ori_ori_n989_), .Y(ori_ori_n990_));
  AOI210     o0941(.A0(ori_ori_n988_), .A1(ori_ori_n253_), .B0(ori_ori_n990_), .Y(ori_ori_n991_));
  OAI220     o0942(.A0(ori_ori_n991_), .A1(ori_ori_n59_), .B0(ori_ori_n986_), .B1(ori_ori_n703_), .Y(ori_ori_n992_));
  OAI210     o0943(.A0(ori_ori_n992_), .A1(ori_ori_n985_), .B0(ori_ori_n936_), .Y(ori_ori_n993_));
  NO2        o0944(.A(x4), .B(x3), .Y(ori_ori_n994_));
  NO3        o0945(.A(ori_ori_n994_), .B(ori_ori_n340_), .C(ori_ori_n87_), .Y(ori_ori_n995_));
  OAI210     o0946(.A0(ori_ori_n995_), .A1(ori_ori_n275_), .B0(ori_ori_n433_), .Y(ori_ori_n996_));
  AOI210     o0947(.A0(ori_ori_n395_), .A1(ori_ori_n125_), .B0(ori_ori_n248_), .Y(ori_ori_n997_));
  NA2        o0948(.A(ori_ori_n955_), .B(ori_ori_n55_), .Y(ori_ori_n998_));
  NO2        o0949(.A(ori_ori_n998_), .B(ori_ori_n969_), .Y(ori_ori_n999_));
  NO2        o0950(.A(ori_ori_n523_), .B(ori_ori_n358_), .Y(ori_ori_n1000_));
  NO3        o0951(.A(x4), .B(ori_ori_n106_), .C(ori_ori_n59_), .Y(ori_ori_n1001_));
  NO2        o0952(.A(ori_ori_n434_), .B(x1), .Y(ori_ori_n1002_));
  NOi31      o0953(.An(ori_ori_n1001_), .B(ori_ori_n1002_), .C(ori_ori_n1000_), .Y(ori_ori_n1003_));
  NA2        o0954(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n1004_));
  NO4        o0955(.A(ori_ori_n956_), .B(ori_ori_n512_), .C(ori_ori_n1004_), .D(x2), .Y(ori_ori_n1005_));
  NO4        o0956(.A(ori_ori_n1005_), .B(ori_ori_n1003_), .C(ori_ori_n999_), .D(ori_ori_n997_), .Y(ori_ori_n1006_));
  AOI210     o0957(.A0(ori_ori_n1006_), .A1(ori_ori_n996_), .B0(ori_ori_n204_), .Y(ori_ori_n1007_));
  NO2        o0958(.A(ori_ori_n661_), .B(ori_ori_n498_), .Y(ori_ori_n1008_));
  NO2        o0959(.A(x6), .B(x2), .Y(ori_ori_n1009_));
  NO3        o0960(.A(ori_ori_n1009_), .B(ori_ori_n692_), .C(ori_ori_n60_), .Y(ori_ori_n1010_));
  OAI210     o0961(.A0(ori_ori_n1010_), .A1(ori_ori_n1008_), .B0(ori_ori_n267_), .Y(ori_ori_n1011_));
  NO2        o0962(.A(ori_ori_n865_), .B(ori_ori_n442_), .Y(ori_ori_n1012_));
  NA3        o0963(.A(x4), .B(x3), .C(ori_ori_n106_), .Y(ori_ori_n1013_));
  NO3        o0964(.A(ori_ori_n1013_), .B(ori_ori_n696_), .C(ori_ori_n461_), .Y(ori_ori_n1014_));
  AOI210     o0965(.A0(ori_ori_n1012_), .A1(ori_ori_n468_), .B0(ori_ori_n1014_), .Y(ori_ori_n1015_));
  AOI210     o0966(.A0(ori_ori_n1015_), .A1(ori_ori_n1011_), .B0(ori_ori_n454_), .Y(ori_ori_n1016_));
  NO2        o0967(.A(ori_ori_n55_), .B(ori_ori_n56_), .Y(ori_ori_n1017_));
  OAI220     o0968(.A0(ori_ori_n815_), .A1(ori_ori_n456_), .B0(ori_ori_n745_), .B1(ori_ori_n125_), .Y(ori_ori_n1018_));
  NOi21      o0969(.An(ori_ori_n120_), .B(ori_ori_n119_), .Y(ori_ori_n1019_));
  NO3        o0970(.A(ori_ori_n341_), .B(ori_ori_n320_), .C(ori_ori_n1019_), .Y(ori_ori_n1020_));
  AOI220     o0971(.A0(ori_ori_n1020_), .A1(ori_ori_n252_), .B0(ori_ori_n1018_), .B1(ori_ori_n112_), .Y(ori_ori_n1021_));
  NO2        o0972(.A(ori_ori_n1021_), .B(ori_ori_n1017_), .Y(ori_ori_n1022_));
  NA2        o0973(.A(ori_ori_n516_), .B(ori_ori_n257_), .Y(ori_ori_n1023_));
  NO2        o0974(.A(ori_ori_n483_), .B(ori_ori_n584_), .Y(ori_ori_n1024_));
  NO2        o0975(.A(ori_ori_n180_), .B(ori_ori_n106_), .Y(ori_ori_n1025_));
  NO3        o0976(.A(ori_ori_n1022_), .B(ori_ori_n1016_), .C(ori_ori_n1007_), .Y(ori_ori_n1026_));
  NA3        o0977(.A(ori_ori_n1026_), .B(ori_ori_n993_), .C(ori_ori_n978_), .Y(ori11));
  NA2        o0978(.A(ori_ori_n372_), .B(ori_ori_n90_), .Y(ori_ori_n1028_));
  INV        o0979(.A(ori_ori_n884_), .Y(ori_ori_n1029_));
  OAI220     o0980(.A0(ori_ori_n1029_), .A1(ori_ori_n53_), .B0(ori_ori_n1028_), .B1(ori_ori_n362_), .Y(ori_ori_n1030_));
  NO2        o0981(.A(ori_ori_n762_), .B(x5), .Y(ori_ori_n1031_));
  NO2        o0982(.A(ori_ori_n167_), .B(ori_ori_n529_), .Y(ori_ori_n1032_));
  AOI220     o0983(.A0(ori_ori_n1032_), .A1(ori_ori_n1031_), .B0(ori_ori_n1030_), .B1(x5), .Y(ori_ori_n1033_));
  OAI220     o0984(.A0(ori_ori_n963_), .A1(ori_ori_n213_), .B0(ori_ori_n211_), .B1(ori_ori_n180_), .Y(ori_ori_n1034_));
  NO2        o0985(.A(ori_ori_n337_), .B(ori_ori_n423_), .Y(ori_ori_n1035_));
  AOI220     o0986(.A0(ori_ori_n1035_), .A1(ori_ori_n178_), .B0(ori_ori_n1034_), .B1(ori_ori_n163_), .Y(ori_ori_n1036_));
  NO2        o0987(.A(ori_ori_n1036_), .B(ori_ori_n444_), .Y(ori_ori_n1037_));
  NO2        o0988(.A(ori_ori_n248_), .B(x2), .Y(ori_ori_n1038_));
  OAI210     o0989(.A0(ori_ori_n907_), .A1(ori_ori_n1038_), .B0(ori_ori_n412_), .Y(ori_ori_n1039_));
  NO2        o0990(.A(ori_ori_n55_), .B(ori_ori_n104_), .Y(ori_ori_n1040_));
  NA2        o0991(.A(ori_ori_n276_), .B(ori_ori_n1040_), .Y(ori_ori_n1041_));
  NO2        o0992(.A(ori_ori_n71_), .B(x1), .Y(ori_ori_n1042_));
  NA2        o0993(.A(ori_ori_n1042_), .B(ori_ori_n78_), .Y(ori_ori_n1043_));
  OA220      o0994(.A0(ori_ori_n1043_), .A1(ori_ori_n610_), .B0(ori_ori_n1041_), .B1(ori_ori_n529_), .Y(ori_ori_n1044_));
  AOI210     o0995(.A0(ori_ori_n1044_), .A1(ori_ori_n1039_), .B0(ori_ori_n703_), .Y(ori_ori_n1045_));
  NO2        o0996(.A(ori_ori_n302_), .B(ori_ori_n53_), .Y(ori_ori_n1046_));
  NO2        o0997(.A(ori_ori_n433_), .B(x3), .Y(ori_ori_n1047_));
  NA3        o0998(.A(ori_ori_n1047_), .B(ori_ori_n1046_), .C(ori_ori_n883_), .Y(ori_ori_n1048_));
  AOI210     o0999(.A0(ori_ori_n1048_), .A1(ori_ori_n933_), .B0(ori_ori_n393_), .Y(ori_ori_n1049_));
  NA2        o1000(.A(ori_ori_n106_), .B(x1), .Y(ori_ori_n1050_));
  NO2        o1001(.A(ori_ori_n616_), .B(ori_ori_n216_), .Y(ori_ori_n1051_));
  NA4        o1002(.A(ori_ori_n1051_), .B(ori_ori_n875_), .C(ori_ori_n465_), .D(ori_ori_n1050_), .Y(ori_ori_n1052_));
  NA3        o1003(.A(x6), .B(x5), .C(ori_ori_n106_), .Y(ori_ori_n1053_));
  NO2        o1004(.A(ori_ori_n1053_), .B(ori_ori_n274_), .Y(ori_ori_n1054_));
  NO2        o1005(.A(ori_ori_n444_), .B(x0), .Y(ori_ori_n1055_));
  NOi31      o1006(.An(ori_ori_n1055_), .B(ori_ori_n171_), .C(ori_ori_n51_), .Y(ori_ori_n1056_));
  AOI210     o1007(.A0(ori_ori_n1054_), .A1(ori_ori_n176_), .B0(ori_ori_n1056_), .Y(ori_ori_n1057_));
  NA2        o1008(.A(ori_ori_n1057_), .B(ori_ori_n1052_), .Y(ori_ori_n1058_));
  NO4        o1009(.A(ori_ori_n1058_), .B(ori_ori_n1049_), .C(ori_ori_n1045_), .D(ori_ori_n1037_), .Y(ori_ori_n1059_));
  OAI210     o1010(.A0(ori_ori_n1033_), .A1(ori_ori_n140_), .B0(ori_ori_n1059_), .Y(ori_ori_n1060_));
  NA2        o1011(.A(ori_ori_n856_), .B(ori_ori_n87_), .Y(ori_ori_n1061_));
  NO3        o1012(.A(ori_ori_n462_), .B(ori_ori_n768_), .C(ori_ori_n120_), .Y(ori_ori_n1062_));
  AOI210     o1013(.A0(ori_ori_n1061_), .A1(ori_ori_n97_), .B0(ori_ori_n1062_), .Y(ori_ori_n1063_));
  NO2        o1014(.A(x8), .B(x1), .Y(ori_ori_n1064_));
  NO3        o1015(.A(ori_ori_n1064_), .B(ori_ori_n684_), .C(ori_ori_n446_), .Y(ori_ori_n1065_));
  OAI210     o1016(.A0(ori_ori_n77_), .A1(ori_ori_n53_), .B0(ori_ori_n1065_), .Y(ori_ori_n1066_));
  OAI210     o1017(.A0(ori_ori_n1063_), .A1(x3), .B0(ori_ori_n1066_), .Y(ori_ori_n1067_));
  NO2        o1018(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n1068_));
  OAI210     o1019(.A0(ori_ori_n1068_), .A1(x2), .B0(ori_ori_n230_), .Y(ori_ori_n1069_));
  NO2        o1020(.A(ori_ori_n603_), .B(ori_ori_n228_), .Y(ori_ori_n1070_));
  NA2        o1021(.A(ori_ori_n1070_), .B(ori_ori_n1069_), .Y(ori_ori_n1071_));
  NO2        o1022(.A(ori_ori_n516_), .B(x4), .Y(ori_ori_n1072_));
  NO3        o1023(.A(ori_ori_n55_), .B(x6), .C(x1), .Y(ori_ori_n1073_));
  NOi21      o1024(.An(ori_ori_n1073_), .B(ori_ori_n483_), .Y(ori_ori_n1074_));
  AOI210     o1025(.A0(ori_ori_n1072_), .A1(ori_ori_n575_), .B0(ori_ori_n1074_), .Y(ori_ori_n1075_));
  NA2        o1026(.A(ori_ori_n1075_), .B(ori_ori_n1071_), .Y(ori_ori_n1076_));
  AOI210     o1027(.A0(ori_ori_n1067_), .A1(x2), .B0(ori_ori_n1076_), .Y(ori_ori_n1077_));
  NO2        o1028(.A(ori_ori_n228_), .B(x2), .Y(ori_ori_n1078_));
  NA2        o1029(.A(ori_ori_n1078_), .B(ori_ori_n994_), .Y(ori_ori_n1079_));
  NOi21      o1030(.An(ori_ori_n384_), .B(ori_ori_n564_), .Y(ori_ori_n1080_));
  NO3        o1031(.A(ori_ori_n1080_), .B(ori_ori_n602_), .C(ori_ori_n320_), .Y(ori_ori_n1081_));
  NA2        o1032(.A(x8), .B(ori_ori_n106_), .Y(ori_ori_n1082_));
  OAI220     o1033(.A0(ori_ori_n703_), .A1(ori_ori_n1082_), .B0(ori_ori_n320_), .B1(ori_ori_n379_), .Y(ori_ori_n1083_));
  OAI210     o1034(.A0(ori_ori_n1083_), .A1(ori_ori_n1081_), .B0(ori_ori_n71_), .Y(ori_ori_n1084_));
  NO2        o1035(.A(ori_ori_n104_), .B(x1), .Y(ori_ori_n1085_));
  NA2        o1036(.A(ori_ori_n1085_), .B(x7), .Y(ori_ori_n1086_));
  AOI210     o1037(.A0(ori_ori_n1084_), .A1(ori_ori_n1079_), .B0(ori_ori_n1086_), .Y(ori_ori_n1087_));
  NA2        o1038(.A(ori_ori_n84_), .B(ori_ori_n71_), .Y(ori_ori_n1088_));
  INV        o1039(.A(ori_ori_n245_), .Y(ori_ori_n1089_));
  NA2        o1040(.A(ori_ori_n1089_), .B(ori_ori_n147_), .Y(ori_ori_n1090_));
  OAI220     o1041(.A0(ori_ori_n1090_), .A1(ori_ori_n362_), .B0(ori_ori_n1088_), .B1(ori_ori_n320_), .Y(ori_ori_n1091_));
  NO2        o1042(.A(ori_ori_n157_), .B(ori_ori_n55_), .Y(ori_ori_n1092_));
  AOI210     o1043(.A0(ori_ori_n1092_), .A1(ori_ori_n1091_), .B0(ori_ori_n1087_), .Y(ori_ori_n1093_));
  OAI210     o1044(.A0(ori_ori_n1077_), .A1(ori_ori_n843_), .B0(ori_ori_n1093_), .Y(ori_ori_n1094_));
  AO210      o1045(.A0(ori_ori_n1060_), .A1(ori_ori_n57_), .B0(ori_ori_n1094_), .Y(ori12));
  NA2        o1046(.A(ori_ori_n874_), .B(ori_ori_n244_), .Y(ori_ori_n1096_));
  NO2        o1047(.A(ori_ori_n620_), .B(x7), .Y(ori_ori_n1097_));
  NA2        o1048(.A(ori_ori_n1097_), .B(ori_ori_n275_), .Y(ori_ori_n1098_));
  NA2        o1049(.A(ori_ori_n695_), .B(ori_ori_n865_), .Y(ori_ori_n1099_));
  AOI210     o1050(.A0(ori_ori_n1098_), .A1(ori_ori_n1096_), .B0(ori_ori_n1099_), .Y(ori_ori_n1100_));
  NOi21      o1051(.An(ori_ori_n400_), .B(ori_ori_n551_), .Y(ori_ori_n1101_));
  NO2        o1052(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n1102_));
  NO2        o1053(.A(ori_ori_n603_), .B(ori_ori_n1102_), .Y(ori_ori_n1103_));
  NO3        o1054(.A(ori_ori_n858_), .B(ori_ori_n108_), .C(ori_ori_n95_), .Y(ori_ori_n1104_));
  AOI210     o1055(.A0(ori_ori_n1103_), .A1(ori_ori_n1002_), .B0(ori_ori_n1104_), .Y(ori_ori_n1105_));
  NA2        o1056(.A(ori_ori_n1040_), .B(ori_ori_n56_), .Y(ori_ori_n1106_));
  OAI220     o1057(.A0(ori_ori_n1106_), .A1(ori_ori_n576_), .B0(ori_ori_n1105_), .B1(ori_ori_n1101_), .Y(ori_ori_n1107_));
  OAI210     o1058(.A0(ori_ori_n1107_), .A1(ori_ori_n1100_), .B0(ori_ori_n580_), .Y(ori_ori_n1108_));
  NA2        o1059(.A(ori_ori_n87_), .B(x5), .Y(ori_ori_n1109_));
  OAI210     o1060(.A0(ori_ori_n1109_), .A1(ori_ori_n320_), .B0(ori_ori_n714_), .Y(ori_ori_n1110_));
  AOI210     o1061(.A0(ori_ori_n817_), .A1(ori_ori_n114_), .B0(ori_ori_n1110_), .Y(ori_ori_n1111_));
  NA2        o1062(.A(ori_ori_n601_), .B(ori_ori_n53_), .Y(ori_ori_n1112_));
  NA2        o1063(.A(ori_ori_n285_), .B(ori_ori_n50_), .Y(ori_ori_n1113_));
  OAI220     o1064(.A0(ori_ori_n1113_), .A1(ori_ori_n308_), .B0(ori_ori_n1112_), .B1(ori_ori_n133_), .Y(ori_ori_n1114_));
  NO2        o1065(.A(ori_ori_n1061_), .B(ori_ori_n511_), .Y(ori_ori_n1115_));
  NO4        o1066(.A(ori_ori_n236_), .B(ori_ori_n267_), .C(ori_ori_n60_), .D(ori_ori_n57_), .Y(ori_ori_n1116_));
  AOI220     o1067(.A0(ori_ori_n1116_), .A1(ori_ori_n1115_), .B0(ori_ori_n1114_), .B1(ori_ori_n56_), .Y(ori_ori_n1117_));
  OAI210     o1068(.A0(ori_ori_n1111_), .A1(ori_ori_n64_), .B0(ori_ori_n1117_), .Y(ori_ori_n1118_));
  NO2        o1069(.A(ori_ori_n57_), .B(x0), .Y(ori_ori_n1119_));
  NO2        o1070(.A(ori_ori_n661_), .B(ori_ori_n317_), .Y(ori_ori_n1120_));
  NO2        o1071(.A(ori_ori_n745_), .B(x3), .Y(ori_ori_n1121_));
  NO2        o1072(.A(ori_ori_n659_), .B(x8), .Y(ori_ori_n1122_));
  AOI220     o1073(.A0(ori_ori_n1122_), .A1(ori_ori_n1121_), .B0(ori_ori_n1120_), .B1(ori_ori_n1119_), .Y(ori_ori_n1123_));
  AOI210     o1074(.A0(ori_ori_n684_), .A1(ori_ori_n244_), .B0(x7), .Y(ori_ori_n1124_));
  NO3        o1075(.A(ori_ori_n1124_), .B(ori_ori_n604_), .C(x8), .Y(ori_ori_n1125_));
  NA4        o1076(.A(ori_ori_n663_), .B(ori_ori_n655_), .C(ori_ori_n201_), .D(x0), .Y(ori_ori_n1126_));
  OAI220     o1077(.A0(ori_ori_n1126_), .A1(ori_ori_n1125_), .B0(ori_ori_n1123_), .B1(ori_ori_n574_), .Y(ori_ori_n1127_));
  AOI210     o1078(.A0(ori_ori_n1118_), .A1(ori_ori_n1009_), .B0(ori_ori_n1127_), .Y(ori_ori_n1128_));
  NO2        o1079(.A(ori_ori_n244_), .B(ori_ori_n55_), .Y(ori_ori_n1129_));
  NO2        o1080(.A(ori_ori_n252_), .B(x8), .Y(ori_ori_n1130_));
  NOi32      o1081(.An(ori_ori_n1130_), .Bn(ori_ori_n200_), .C(ori_ori_n565_), .Y(ori_ori_n1131_));
  NO2        o1082(.A(ori_ori_n88_), .B(ori_ori_n60_), .Y(ori_ori_n1132_));
  OAI210     o1083(.A0(ori_ori_n1131_), .A1(ori_ori_n1129_), .B0(ori_ori_n1132_), .Y(ori_ori_n1133_));
  NO2        o1084(.A(ori_ori_n936_), .B(ori_ori_n96_), .Y(ori_ori_n1134_));
  NO2        o1085(.A(ori_ori_n166_), .B(ori_ori_n53_), .Y(ori_ori_n1135_));
  AOI210     o1086(.A0(ori_ori_n337_), .A1(x8), .B0(ori_ori_n1135_), .Y(ori_ori_n1136_));
  AOI210     o1087(.A0(ori_ori_n213_), .A1(ori_ori_n92_), .B0(ori_ori_n1136_), .Y(ori_ori_n1137_));
  OAI210     o1088(.A0(ori_ori_n1137_), .A1(ori_ori_n1134_), .B0(ori_ori_n672_), .Y(ori_ori_n1138_));
  NO2        o1089(.A(x7), .B(x0), .Y(ori_ori_n1139_));
  NO3        o1090(.A(ori_ori_n157_), .B(ori_ori_n1139_), .C(ori_ori_n144_), .Y(ori_ori_n1140_));
  XN2        o1091(.A(x8), .B(x7), .Y(ori_ori_n1141_));
  NO3        o1092(.A(ori_ori_n1064_), .B(ori_ori_n255_), .C(ori_ori_n1141_), .Y(ori_ori_n1142_));
  OAI210     o1093(.A0(ori_ori_n1142_), .A1(ori_ori_n1140_), .B0(ori_ori_n724_), .Y(ori_ori_n1143_));
  NO2        o1094(.A(ori_ori_n264_), .B(ori_ori_n260_), .Y(ori_ori_n1144_));
  NO2        o1095(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n1145_));
  OAI210     o1096(.A0(ori_ori_n1144_), .A1(ori_ori_n275_), .B0(ori_ori_n1145_), .Y(ori_ori_n1146_));
  NA4        o1097(.A(ori_ori_n1146_), .B(ori_ori_n1143_), .C(ori_ori_n1138_), .D(ori_ori_n1133_), .Y(ori_ori_n1147_));
  NA2        o1098(.A(ori_ori_n1147_), .B(ori_ori_n555_), .Y(ori_ori_n1148_));
  NO2        o1099(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n1149_));
  NA2        o1100(.A(ori_ori_n1149_), .B(ori_ori_n162_), .Y(ori_ori_n1150_));
  NO2        o1101(.A(ori_ori_n665_), .B(ori_ori_n255_), .Y(ori_ori_n1151_));
  OAI210     o1102(.A0(ori_ori_n1151_), .A1(ori_ori_n1012_), .B0(ori_ori_n50_), .Y(ori_ori_n1152_));
  AOI210     o1103(.A0(ori_ori_n1152_), .A1(ori_ori_n1150_), .B0(ori_ori_n428_), .Y(ori_ori_n1153_));
  OAI220     o1104(.A0(ori_ori_n287_), .A1(ori_ori_n273_), .B0(ori_ori_n260_), .B1(ori_ori_n239_), .Y(ori_ori_n1154_));
  NA3        o1105(.A(ori_ori_n1154_), .B(ori_ori_n672_), .C(x1), .Y(ori_ori_n1155_));
  OAI210     o1106(.A0(x8), .A1(x0), .B0(x4), .Y(ori_ori_n1156_));
  NO2        o1107(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n1157_));
  NO2        o1108(.A(ori_ori_n68_), .B(ori_ori_n1157_), .Y(ori_ori_n1158_));
  NOi21      o1109(.An(ori_ori_n1156_), .B(ori_ori_n1158_), .Y(ori_ori_n1159_));
  NO2        o1110(.A(ori_ori_n663_), .B(ori_ori_n320_), .Y(ori_ori_n1160_));
  NO2        o1111(.A(ori_ori_n771_), .B(ori_ori_n217_), .Y(ori_ori_n1161_));
  OAI210     o1112(.A0(ori_ori_n1160_), .A1(ori_ori_n1159_), .B0(ori_ori_n1161_), .Y(ori_ori_n1162_));
  NO2        o1113(.A(ori_ori_n140_), .B(ori_ori_n139_), .Y(ori_ori_n1163_));
  NO2        o1114(.A(ori_ori_n603_), .B(ori_ori_n442_), .Y(ori_ori_n1164_));
  OAI210     o1115(.A0(ori_ori_n1164_), .A1(ori_ori_n1163_), .B0(ori_ori_n252_), .Y(ori_ori_n1165_));
  NA2        o1116(.A(ori_ori_n325_), .B(ori_ori_n59_), .Y(ori_ori_n1166_));
  NO2        o1117(.A(ori_ori_n1106_), .B(ori_ori_n1166_), .Y(ori_ori_n1167_));
  INV        o1118(.A(ori_ori_n1167_), .Y(ori_ori_n1168_));
  NA4        o1119(.A(ori_ori_n1168_), .B(ori_ori_n1165_), .C(ori_ori_n1162_), .D(ori_ori_n1155_), .Y(ori_ori_n1169_));
  OAI210     o1120(.A0(ori_ori_n1169_), .A1(ori_ori_n1153_), .B0(ori_ori_n674_), .Y(ori_ori_n1170_));
  NA4        o1121(.A(ori_ori_n1170_), .B(ori_ori_n1148_), .C(ori_ori_n1128_), .D(ori_ori_n1108_), .Y(ori13));
  NO2        o1122(.A(ori_ori_n461_), .B(ori_ori_n347_), .Y(ori_ori_n1172_));
  NOi41      o1123(.An(ori_ori_n1172_), .B(ori_ori_n672_), .C(ori_ori_n289_), .D(ori_ori_n236_), .Y(ori_ori_n1173_));
  NO2        o1124(.A(ori_ori_n858_), .B(ori_ori_n180_), .Y(ori_ori_n1174_));
  NO2        o1125(.A(ori_ori_n156_), .B(ori_ori_n71_), .Y(ori_ori_n1175_));
  XN2        o1126(.A(x4), .B(x0), .Y(ori_ori_n1176_));
  NO3        o1127(.A(ori_ori_n1176_), .B(ori_ori_n107_), .C(ori_ori_n419_), .Y(ori_ori_n1177_));
  AO220      o1128(.A0(ori_ori_n1177_), .A1(ori_ori_n1175_), .B0(ori_ori_n1174_), .B1(ori_ori_n326_), .Y(ori_ori_n1178_));
  OAI210     o1129(.A0(ori_ori_n1178_), .A1(ori_ori_n1173_), .B0(x3), .Y(ori_ori_n1179_));
  NO2        o1130(.A(ori_ori_n858_), .B(x6), .Y(ori_ori_n1180_));
  NO2        o1131(.A(ori_ori_n1113_), .B(ori_ori_n391_), .Y(ori_ori_n1181_));
  NO3        o1132(.A(x8), .B(x5), .C(ori_ori_n106_), .Y(ori_ori_n1182_));
  NA2        o1133(.A(ori_ori_n1182_), .B(ori_ori_n637_), .Y(ori_ori_n1183_));
  NO2        o1134(.A(ori_ori_n603_), .B(ori_ori_n195_), .Y(ori_ori_n1184_));
  NA2        o1135(.A(ori_ori_n1184_), .B(ori_ori_n1073_), .Y(ori_ori_n1185_));
  NA2        o1136(.A(ori_ori_n446_), .B(ori_ori_n53_), .Y(ori_ori_n1186_));
  NO2        o1137(.A(ori_ori_n1186_), .B(ori_ori_n929_), .Y(ori_ori_n1187_));
  NA2        o1138(.A(ori_ori_n1106_), .B(ori_ori_n466_), .Y(ori_ori_n1188_));
  NA2        o1139(.A(ori_ori_n56_), .B(ori_ori_n106_), .Y(ori_ori_n1189_));
  NA2        o1140(.A(ori_ori_n1189_), .B(x1), .Y(ori_ori_n1190_));
  NO2        o1141(.A(ori_ori_n1190_), .B(ori_ori_n257_), .Y(ori_ori_n1191_));
  NO2        o1142(.A(ori_ori_n317_), .B(x6), .Y(ori_ori_n1192_));
  OAI210     o1143(.A0(ori_ori_n248_), .A1(ori_ori_n967_), .B0(ori_ori_n947_), .Y(ori_ori_n1193_));
  AOI220     o1144(.A0(ori_ori_n1193_), .A1(ori_ori_n1192_), .B0(ori_ori_n1191_), .B1(ori_ori_n1188_), .Y(ori_ori_n1194_));
  NAi41      o1145(.An(ori_ori_n1187_), .B(ori_ori_n1194_), .C(ori_ori_n1185_), .D(ori_ori_n1183_), .Y(ori_ori_n1195_));
  AOI220     o1146(.A0(ori_ori_n1195_), .A1(ori_ori_n68_), .B0(ori_ori_n1181_), .B1(ori_ori_n1180_), .Y(ori_ori_n1196_));
  NA2        o1147(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n1197_));
  NA2        o1148(.A(ori_ori_n1197_), .B(ori_ori_n892_), .Y(ori_ori_n1198_));
  OAI220     o1149(.A0(ori_ori_n301_), .A1(ori_ori_n813_), .B0(ori_ori_n87_), .B1(ori_ori_n77_), .Y(ori_ori_n1199_));
  AOI210     o1150(.A0(ori_ori_n1109_), .A1(ori_ori_n614_), .B0(ori_ori_n967_), .Y(ori_ori_n1200_));
  OA210      o1151(.A0(ori_ori_n1199_), .A1(ori_ori_n1198_), .B0(ori_ori_n1200_), .Y(ori_ori_n1201_));
  NA2        o1152(.A(ori_ori_n616_), .B(ori_ori_n55_), .Y(ori_ori_n1202_));
  NA2        o1153(.A(ori_ori_n504_), .B(ori_ori_n492_), .Y(ori_ori_n1203_));
  NA2        o1154(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n1204_));
  NA2        o1155(.A(ori_ori_n1204_), .B(ori_ori_n538_), .Y(ori_ori_n1205_));
  NO2        o1156(.A(ori_ori_n159_), .B(ori_ori_n128_), .Y(ori_ori_n1206_));
  AOI210     o1157(.A0(ori_ori_n1205_), .A1(ori_ori_n429_), .B0(ori_ori_n1206_), .Y(ori_ori_n1207_));
  OAI220     o1158(.A0(ori_ori_n1207_), .A1(ori_ori_n865_), .B0(ori_ori_n1203_), .B1(ori_ori_n1202_), .Y(ori_ori_n1208_));
  OAI210     o1159(.A0(ori_ori_n1208_), .A1(ori_ori_n1201_), .B0(ori_ori_n1139_), .Y(ori_ori_n1209_));
  NAi21      o1160(.An(ori_ori_n84_), .B(ori_ori_n379_), .Y(ori_ori_n1210_));
  NO2        o1161(.A(ori_ori_n1210_), .B(ori_ori_n71_), .Y(ori_ori_n1211_));
  AOI210     o1162(.A0(ori_ori_n162_), .A1(x4), .B0(ori_ori_n172_), .Y(ori_ori_n1212_));
  NO2        o1163(.A(ori_ori_n1212_), .B(x0), .Y(ori_ori_n1213_));
  NO2        o1164(.A(ori_ori_n169_), .B(ori_ori_n292_), .Y(ori_ori_n1214_));
  OAI210     o1165(.A0(ori_ori_n1214_), .A1(ori_ori_n1213_), .B0(ori_ori_n1211_), .Y(ori_ori_n1215_));
  NA3        o1166(.A(ori_ori_n1145_), .B(ori_ori_n186_), .C(ori_ori_n71_), .Y(ori_ori_n1216_));
  NO2        o1167(.A(x4), .B(x0), .Y(ori_ori_n1217_));
  NO3        o1168(.A(ori_ori_n987_), .B(ori_ori_n245_), .C(ori_ori_n538_), .Y(ori_ori_n1218_));
  OAI210     o1169(.A0(ori_ori_n1218_), .A1(ori_ori_n196_), .B0(ori_ori_n1217_), .Y(ori_ori_n1219_));
  NA3        o1170(.A(ori_ori_n1219_), .B(ori_ori_n1216_), .C(ori_ori_n1215_), .Y(ori_ori_n1220_));
  NA2        o1171(.A(ori_ori_n247_), .B(ori_ori_n724_), .Y(ori_ori_n1221_));
  NA2        o1172(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n1222_));
  NO3        o1173(.A(ori_ori_n1222_), .B(ori_ori_n492_), .C(ori_ori_n81_), .Y(ori_ori_n1223_));
  NA2        o1174(.A(ori_ori_n1223_), .B(x2), .Y(ori_ori_n1224_));
  NO2        o1175(.A(ori_ori_n320_), .B(ori_ori_n379_), .Y(ori_ori_n1225_));
  NO2        o1176(.A(ori_ori_n684_), .B(x0), .Y(ori_ori_n1226_));
  OAI210     o1177(.A0(ori_ori_n1226_), .A1(ori_ori_n1225_), .B0(ori_ori_n329_), .Y(ori_ori_n1227_));
  NO2        o1178(.A(ori_ori_n782_), .B(x1), .Y(ori_ori_n1228_));
  AOI220     o1179(.A0(ori_ori_n1228_), .A1(ori_ori_n609_), .B0(ori_ori_n476_), .B1(ori_ori_n293_), .Y(ori_ori_n1229_));
  NA2        o1180(.A(ori_ori_n498_), .B(ori_ori_n50_), .Y(ori_ori_n1230_));
  AOI220     o1181(.A0(ori_ori_n1230_), .A1(ori_ori_n1174_), .B0(ori_ori_n968_), .B1(ori_ori_n97_), .Y(ori_ori_n1231_));
  NA4        o1182(.A(ori_ori_n1231_), .B(ori_ori_n1229_), .C(ori_ori_n1227_), .D(ori_ori_n1224_), .Y(ori_ori_n1232_));
  AOI220     o1183(.A0(ori_ori_n1232_), .A1(ori_ori_n129_), .B0(ori_ori_n1220_), .B1(ori_ori_n67_), .Y(ori_ori_n1233_));
  NA4        o1184(.A(ori_ori_n1233_), .B(ori_ori_n1209_), .C(ori_ori_n1196_), .D(ori_ori_n1179_), .Y(ori14));
  NO2        o1185(.A(ori_ori_n367_), .B(ori_ori_n71_), .Y(ori_ori_n1235_));
  NO3        o1186(.A(x7), .B(x6), .C(x0), .Y(ori_ori_n1236_));
  OAI210     o1187(.A0(ori_ori_n1236_), .A1(ori_ori_n1235_), .B0(x8), .Y(ori_ori_n1237_));
  NA2        o1188(.A(ori_ori_n1122_), .B(ori_ori_n85_), .Y(ori_ori_n1238_));
  AOI210     o1189(.A0(ori_ori_n1238_), .A1(ori_ori_n1237_), .B0(ori_ori_n155_), .Y(ori_ori_n1239_));
  AOI220     o1190(.A0(ori_ori_n371_), .A1(ori_ori_n843_), .B0(ori_ori_n446_), .B1(ori_ori_n419_), .Y(ori_ori_n1240_));
  NA2        o1191(.A(ori_ori_n276_), .B(ori_ori_n963_), .Y(ori_ori_n1241_));
  OAI220     o1192(.A0(ori_ori_n1241_), .A1(ori_ori_n1240_), .B0(ori_ori_n464_), .B1(ori_ori_n797_), .Y(ori_ori_n1242_));
  OA210      o1193(.A0(ori_ori_n1242_), .A1(ori_ori_n1239_), .B0(x4), .Y(ori_ori_n1243_));
  NO2        o1194(.A(ori_ori_n139_), .B(ori_ori_n607_), .Y(ori_ori_n1244_));
  NA2        o1195(.A(x6), .B(x2), .Y(ori_ori_n1245_));
  NO2        o1196(.A(ori_ori_n625_), .B(ori_ori_n1245_), .Y(ori_ori_n1246_));
  OA210      o1197(.A0(ori_ori_n1244_), .A1(ori_ori_n209_), .B0(ori_ori_n1246_), .Y(ori_ori_n1247_));
  NO4        o1198(.A(ori_ori_n603_), .B(ori_ori_n372_), .C(ori_ori_n297_), .D(ori_ori_n112_), .Y(ori_ori_n1248_));
  OAI210     o1199(.A0(ori_ori_n1248_), .A1(ori_ori_n1247_), .B0(ori_ori_n59_), .Y(ori_ori_n1249_));
  NA2        o1200(.A(x6), .B(ori_ori_n104_), .Y(ori_ori_n1250_));
  NO2        o1201(.A(ori_ori_n661_), .B(ori_ori_n1250_), .Y(ori_ori_n1251_));
  NA2        o1202(.A(ori_ori_n1251_), .B(ori_ori_n916_), .Y(ori_ori_n1252_));
  AOI210     o1203(.A0(ori_ori_n1122_), .A1(ori_ori_n1001_), .B0(x1), .Y(ori_ori_n1253_));
  NO2        o1204(.A(ori_ori_n533_), .B(x5), .Y(ori_ori_n1254_));
  NA3        o1205(.A(ori_ori_n1254_), .B(ori_ori_n119_), .C(x0), .Y(ori_ori_n1255_));
  NA4        o1206(.A(ori_ori_n691_), .B(ori_ori_n917_), .C(ori_ori_n301_), .D(ori_ori_n68_), .Y(ori_ori_n1256_));
  AN4        o1207(.A(ori_ori_n1256_), .B(ori_ori_n1255_), .C(ori_ori_n1253_), .D(ori_ori_n1252_), .Y(ori_ori_n1257_));
  NO2        o1208(.A(ori_ori_n696_), .B(ori_ori_n1082_), .Y(ori_ori_n1258_));
  NO2        o1209(.A(ori_ori_n77_), .B(ori_ori_n58_), .Y(ori_ori_n1259_));
  OAI210     o1210(.A0(ori_ori_n1258_), .A1(ori_ori_n443_), .B0(ori_ori_n1259_), .Y(ori_ori_n1260_));
  AO210      o1211(.A0(ori_ori_n1235_), .A1(ori_ori_n1001_), .B0(ori_ori_n53_), .Y(ori_ori_n1261_));
  AOI210     o1212(.A0(ori_ori_n758_), .A1(ori_ori_n807_), .B0(ori_ori_n1261_), .Y(ori_ori_n1262_));
  AOI220     o1213(.A0(ori_ori_n1262_), .A1(ori_ori_n1260_), .B0(ori_ori_n1257_), .B1(ori_ori_n1249_), .Y(ori_ori_n1263_));
  NO2        o1214(.A(ori_ori_n1263_), .B(ori_ori_n1243_), .Y(ori_ori_n1264_));
  NO2        o1215(.A(ori_ori_n317_), .B(x2), .Y(ori_ori_n1265_));
  XN2        o1216(.A(x4), .B(x1), .Y(ori_ori_n1266_));
  NO2        o1217(.A(ori_ori_n1266_), .B(ori_ori_n301_), .Y(ori_ori_n1267_));
  NO2        o1218(.A(ori_ori_n336_), .B(ori_ori_n60_), .Y(ori_ori_n1268_));
  NA2        o1219(.A(ori_ori_n1268_), .B(ori_ori_n1265_), .Y(ori_ori_n1269_));
  NA2        o1220(.A(ori_ori_n685_), .B(ori_ori_n56_), .Y(ori_ori_n1270_));
  OAI220     o1221(.A0(ori_ori_n1270_), .A1(ori_ori_n156_), .B0(ori_ori_n187_), .B1(ori_ori_n71_), .Y(ori_ori_n1271_));
  NO2        o1222(.A(ori_ori_n213_), .B(ori_ori_n255_), .Y(ori_ori_n1272_));
  AOI220     o1223(.A0(ori_ori_n136_), .A1(ori_ori_n56_), .B0(ori_ori_n91_), .B1(x5), .Y(ori_ori_n1273_));
  NA2        o1224(.A(ori_ori_n1073_), .B(ori_ori_n306_), .Y(ori_ori_n1274_));
  NA2        o1225(.A(ori_ori_n247_), .B(ori_ori_n351_), .Y(ori_ori_n1275_));
  NA2        o1226(.A(ori_ori_n636_), .B(ori_ori_n1019_), .Y(ori_ori_n1276_));
  OAI220     o1227(.A0(ori_ori_n1276_), .A1(ori_ori_n1275_), .B0(ori_ori_n1274_), .B1(ori_ori_n1273_), .Y(ori_ori_n1277_));
  AOI210     o1228(.A0(ori_ori_n1272_), .A1(ori_ori_n1271_), .B0(ori_ori_n1277_), .Y(ori_ori_n1278_));
  AOI210     o1229(.A0(ori_ori_n1278_), .A1(ori_ori_n1269_), .B0(x7), .Y(ori_ori_n1279_));
  NO2        o1230(.A(ori_ori_n491_), .B(x6), .Y(ori_ori_n1280_));
  AOI210     o1231(.A0(ori_ori_n809_), .A1(ori_ori_n948_), .B0(ori_ori_n1280_), .Y(ori_ori_n1281_));
  OAI220     o1232(.A0(ori_ori_n1281_), .A1(ori_ori_n55_), .B0(ori_ori_n491_), .B1(ori_ori_n100_), .Y(ori_ori_n1282_));
  NA2        o1233(.A(ori_ori_n1282_), .B(ori_ori_n353_), .Y(ori_ori_n1283_));
  NA3        o1234(.A(ori_ori_n610_), .B(ori_ori_n1050_), .C(ori_ori_n70_), .Y(ori_ori_n1284_));
  NO4        o1235(.A(ori_ori_n1284_), .B(ori_ori_n1222_), .C(ori_ori_n117_), .D(ori_ori_n55_), .Y(ori_ori_n1285_));
  NO3        o1236(.A(ori_ori_n1043_), .B(ori_ori_n815_), .C(ori_ori_n481_), .Y(ori_ori_n1286_));
  NO3        o1237(.A(ori_ori_n745_), .B(ori_ori_n498_), .C(ori_ori_n54_), .Y(ori_ori_n1287_));
  NO4        o1238(.A(ori_ori_n1287_), .B(ori_ori_n1286_), .C(ori_ori_n1285_), .D(ori_ori_n1024_), .Y(ori_ori_n1288_));
  AOI210     o1239(.A0(ori_ori_n1288_), .A1(ori_ori_n1283_), .B0(ori_ori_n303_), .Y(ori_ori_n1289_));
  NA2        o1240(.A(ori_ori_n890_), .B(ori_ori_n53_), .Y(ori_ori_n1290_));
  OAI210     o1241(.A0(ori_ori_n242_), .A1(ori_ori_n114_), .B0(x2), .Y(ori_ori_n1291_));
  NA2        o1242(.A(ori_ori_n363_), .B(ori_ori_n56_), .Y(ori_ori_n1292_));
  OA220      o1243(.A0(ori_ori_n1292_), .A1(ori_ori_n1291_), .B0(ori_ori_n1290_), .B1(ori_ori_n371_), .Y(ori_ori_n1293_));
  NA2        o1244(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n1294_));
  NO2        o1245(.A(ori_ori_n1294_), .B(ori_ori_n194_), .Y(ori_ori_n1295_));
  NA4        o1246(.A(ori_ori_n1295_), .B(ori_ori_n363_), .C(ori_ori_n255_), .D(ori_ori_n67_), .Y(ori_ori_n1296_));
  OAI210     o1247(.A0(ori_ori_n1293_), .A1(ori_ori_n313_), .B0(ori_ori_n1296_), .Y(ori_ori_n1297_));
  NO3        o1248(.A(ori_ori_n1297_), .B(ori_ori_n1289_), .C(ori_ori_n1279_), .Y(ori_ori_n1298_));
  OAI210     o1249(.A0(ori_ori_n1264_), .A1(x3), .B0(ori_ori_n1298_), .Y(ori15));
  NA2        o1250(.A(ori_ori_n585_), .B(ori_ori_n59_), .Y(ori_ori_n1300_));
  NAi41      o1251(.An(x2), .B(x7), .C(x6), .D(x0), .Y(ori_ori_n1301_));
  AOI210     o1252(.A0(ori_ori_n1301_), .A1(ori_ori_n1300_), .B0(ori_ori_n53_), .Y(ori_ori_n1302_));
  NA3        o1253(.A(ori_ori_n57_), .B(x6), .C(ori_ori_n106_), .Y(ori_ori_n1303_));
  NO2        o1254(.A(ori_ori_n1303_), .B(ori_ori_n292_), .Y(ori_ori_n1304_));
  OAI210     o1255(.A0(ori_ori_n1304_), .A1(ori_ori_n1302_), .B0(ori_ori_n1145_), .Y(ori_ori_n1305_));
  NA2        o1256(.A(ori_ori_n108_), .B(ori_ori_n106_), .Y(ori_ori_n1306_));
  NA4        o1257(.A(ori_ori_n1306_), .B(ori_ori_n634_), .C(ori_ori_n307_), .D(x6), .Y(ori_ori_n1307_));
  AOI210     o1258(.A0(ori_ori_n723_), .A1(ori_ori_n76_), .B0(x3), .Y(ori_ori_n1308_));
  NA3        o1259(.A(ori_ori_n1308_), .B(ori_ori_n1307_), .C(ori_ori_n1305_), .Y(ori_ori_n1309_));
  AOI210     o1260(.A0(ori_ori_n1055_), .A1(ori_ori_n589_), .B0(ori_ori_n50_), .Y(ori_ori_n1310_));
  NO2        o1261(.A(ori_ori_n292_), .B(ori_ori_n106_), .Y(ori_ori_n1311_));
  NO2        o1262(.A(ori_ori_n234_), .B(x5), .Y(ori_ori_n1312_));
  NA2        o1263(.A(ori_ori_n1312_), .B(ori_ori_n1311_), .Y(ori_ori_n1313_));
  NA3        o1264(.A(ori_ori_n1228_), .B(ori_ori_n624_), .C(ori_ori_n1157_), .Y(ori_ori_n1314_));
  NA4        o1265(.A(ori_ori_n1314_), .B(ori_ori_n1313_), .C(ori_ori_n1310_), .D(ori_ori_n1255_), .Y(ori_ori_n1315_));
  NA2        o1266(.A(ori_ori_n330_), .B(ori_ori_n339_), .Y(ori_ori_n1316_));
  AOI210     o1267(.A0(ori_ori_n1190_), .A1(ori_ori_n58_), .B0(ori_ori_n1316_), .Y(ori_ori_n1317_));
  NA4        o1268(.A(ori_ori_n1190_), .B(ori_ori_n695_), .C(ori_ori_n1119_), .D(ori_ori_n379_), .Y(ori_ori_n1318_));
  NA2        o1269(.A(ori_ori_n589_), .B(ori_ori_n465_), .Y(ori_ori_n1319_));
  NO2        o1270(.A(ori_ori_n745_), .B(ori_ori_n53_), .Y(ori_ori_n1320_));
  NO2        o1271(.A(ori_ori_n771_), .B(ori_ori_n297_), .Y(ori_ori_n1321_));
  NA2        o1272(.A(ori_ori_n1321_), .B(ori_ori_n1320_), .Y(ori_ori_n1322_));
  NA3        o1273(.A(ori_ori_n1322_), .B(ori_ori_n1319_), .C(ori_ori_n1318_), .Y(ori_ori_n1323_));
  OAI210     o1274(.A0(ori_ori_n1323_), .A1(ori_ori_n1317_), .B0(ori_ori_n77_), .Y(ori_ori_n1324_));
  NA2        o1275(.A(ori_ori_n365_), .B(ori_ori_n698_), .Y(ori_ori_n1325_));
  NA2        o1276(.A(ori_ori_n571_), .B(ori_ori_n56_), .Y(ori_ori_n1326_));
  NA3        o1277(.A(ori_ori_n1326_), .B(ori_ori_n339_), .C(ori_ori_n108_), .Y(ori_ori_n1327_));
  AOI210     o1278(.A0(ori_ori_n1327_), .A1(ori_ori_n1325_), .B0(ori_ori_n498_), .Y(ori_ori_n1328_));
  NO3        o1279(.A(ori_ori_n795_), .B(ori_ori_n621_), .C(ori_ori_n195_), .Y(ori_ori_n1329_));
  OAI210     o1280(.A0(ori_ori_n1329_), .A1(ori_ori_n1328_), .B0(ori_ori_n491_), .Y(ori_ori_n1330_));
  NO2        o1281(.A(ori_ori_n865_), .B(ori_ori_n50_), .Y(ori_ori_n1331_));
  NO2        o1282(.A(ori_ori_n244_), .B(ori_ori_n64_), .Y(ori_ori_n1332_));
  OA210      o1283(.A0(ori_ori_n1332_), .A1(ori_ori_n1331_), .B0(ori_ori_n407_), .Y(ori_ori_n1333_));
  NA2        o1284(.A(ori_ori_n57_), .B(x3), .Y(ori_ori_n1334_));
  AOI210     o1285(.A0(ori_ori_n969_), .A1(ori_ori_n1334_), .B0(ori_ori_n679_), .Y(ori_ori_n1335_));
  OAI210     o1286(.A0(ori_ori_n1335_), .A1(ori_ori_n1333_), .B0(ori_ori_n1009_), .Y(ori_ori_n1336_));
  NA2        o1287(.A(ori_ori_n1295_), .B(ori_ori_n68_), .Y(ori_ori_n1337_));
  NO2        o1288(.A(ori_ori_n1245_), .B(x0), .Y(ori_ori_n1338_));
  AOI210     o1289(.A0(ori_ori_n1338_), .A1(ori_ori_n604_), .B0(x8), .Y(ori_ori_n1339_));
  NO2        o1290(.A(ori_ori_n428_), .B(ori_ori_n81_), .Y(ori_ori_n1340_));
  NO2        o1291(.A(ori_ori_n923_), .B(ori_ori_n71_), .Y(ori_ori_n1341_));
  NA2        o1292(.A(ori_ori_n1341_), .B(ori_ori_n1340_), .Y(ori_ori_n1342_));
  NO2        o1293(.A(ori_ori_n967_), .B(x6), .Y(ori_ori_n1343_));
  NA4        o1294(.A(ori_ori_n1343_), .B(ori_ori_n594_), .C(ori_ori_n157_), .D(ori_ori_n411_), .Y(ori_ori_n1344_));
  AN4        o1295(.A(ori_ori_n1344_), .B(ori_ori_n1342_), .C(ori_ori_n1339_), .D(ori_ori_n1337_), .Y(ori_ori_n1345_));
  NA4        o1296(.A(ori_ori_n1345_), .B(ori_ori_n1336_), .C(ori_ori_n1330_), .D(ori_ori_n1324_), .Y(ori_ori_n1346_));
  NA2        o1297(.A(ori_ori_n163_), .B(ori_ori_n729_), .Y(ori_ori_n1347_));
  NO2        o1298(.A(ori_ori_n646_), .B(x2), .Y(ori_ori_n1348_));
  OAI210     o1299(.A0(ori_ori_n1348_), .A1(ori_ori_n85_), .B0(x1), .Y(ori_ori_n1349_));
  AOI210     o1300(.A0(ori_ori_n1349_), .A1(ori_ori_n1347_), .B0(ori_ori_n317_), .Y(ori_ori_n1350_));
  NA3        o1301(.A(ori_ori_n57_), .B(x1), .C(x0), .Y(ori_ori_n1351_));
  NA3        o1302(.A(ori_ori_n71_), .B(x5), .C(x2), .Y(ori_ori_n1352_));
  NA4        o1303(.A(x7), .B(x3), .C(ori_ori_n53_), .D(x0), .Y(ori_ori_n1353_));
  OAI220     o1304(.A0(ori_ori_n1353_), .A1(x6), .B0(ori_ori_n1352_), .B1(ori_ori_n1351_), .Y(ori_ori_n1354_));
  INV        o1305(.A(ori_ori_n1354_), .Y(ori_ori_n1355_));
  NAi21      o1306(.An(ori_ori_n112_), .B(ori_ori_n739_), .Y(ori_ori_n1356_));
  NA4        o1307(.A(ori_ori_n1356_), .B(ori_ori_n315_), .C(ori_ori_n287_), .D(ori_ori_n624_), .Y(ori_ori_n1357_));
  OAI220     o1308(.A0(ori_ori_n320_), .A1(x7), .B0(ori_ori_n128_), .B1(ori_ori_n71_), .Y(ori_ori_n1358_));
  NA3        o1309(.A(ori_ori_n1358_), .B(ori_ori_n782_), .C(ori_ori_n1085_), .Y(ori_ori_n1359_));
  NA2        o1310(.A(ori_ori_n82_), .B(ori_ori_n50_), .Y(ori_ori_n1360_));
  AO210      o1311(.A0(ori_ori_n1360_), .A1(ori_ori_n312_), .B0(ori_ori_n155_), .Y(ori_ori_n1361_));
  NA4        o1312(.A(ori_ori_n1361_), .B(ori_ori_n1359_), .C(ori_ori_n1357_), .D(ori_ori_n1355_), .Y(ori_ori_n1362_));
  OAI210     o1313(.A0(ori_ori_n1362_), .A1(ori_ori_n1350_), .B0(ori_ori_n56_), .Y(ori_ori_n1363_));
  AOI210     o1314(.A0(ori_ori_n687_), .A1(x4), .B0(ori_ori_n948_), .Y(ori_ori_n1364_));
  OAI220     o1315(.A0(ori_ori_n1364_), .A1(ori_ori_n298_), .B0(ori_ori_n1013_), .B1(ori_ori_n937_), .Y(ori_ori_n1365_));
  NA2        o1316(.A(ori_ori_n826_), .B(ori_ori_n404_), .Y(ori_ori_n1366_));
  OAI210     o1317(.A0(ori_ori_n1340_), .A1(ori_ori_n1332_), .B0(ori_ori_n288_), .Y(ori_ori_n1367_));
  OAI210     o1318(.A0(ori_ori_n1366_), .A1(ori_ori_n838_), .B0(ori_ori_n1367_), .Y(ori_ori_n1368_));
  OAI210     o1319(.A0(ori_ori_n1368_), .A1(ori_ori_n1365_), .B0(x6), .Y(ori_ori_n1369_));
  NO2        o1320(.A(ori_ori_n57_), .B(ori_ori_n59_), .Y(ori_ori_n1370_));
  NO2        o1321(.A(x7), .B(x5), .Y(ori_ori_n1371_));
  AOI220     o1322(.A0(ori_ori_n847_), .A1(ori_ori_n1370_), .B0(ori_ori_n537_), .B1(ori_ori_n1371_), .Y(ori_ori_n1372_));
  NA2        o1323(.A(ori_ori_n755_), .B(ori_ori_n288_), .Y(ori_ori_n1373_));
  NA3        o1324(.A(ori_ori_n616_), .B(ori_ori_n290_), .C(ori_ori_n239_), .Y(ori_ori_n1374_));
  NA3        o1325(.A(ori_ori_n1374_), .B(ori_ori_n1373_), .C(ori_ori_n1372_), .Y(ori_ori_n1375_));
  NA2        o1326(.A(ori_ori_n1375_), .B(ori_ori_n422_), .Y(ori_ori_n1376_));
  AOI210     o1327(.A0(ori_ori_n375_), .A1(ori_ori_n337_), .B0(ori_ori_n55_), .Y(ori_ori_n1377_));
  NA4        o1328(.A(ori_ori_n1377_), .B(ori_ori_n1376_), .C(ori_ori_n1369_), .D(ori_ori_n1363_), .Y(ori_ori_n1378_));
  AO220      o1329(.A0(ori_ori_n1378_), .A1(ori_ori_n1346_), .B0(ori_ori_n1315_), .B1(ori_ori_n1309_), .Y(ori16));
  NO2        o1330(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n1380_));
  NA2        o1331(.A(ori_ori_n660_), .B(ori_ori_n534_), .Y(ori_ori_n1381_));
  NA3        o1332(.A(ori_ori_n228_), .B(ori_ori_n429_), .C(ori_ori_n948_), .Y(ori_ori_n1382_));
  NA2        o1333(.A(ori_ori_n131_), .B(ori_ori_n204_), .Y(ori_ori_n1383_));
  AOI210     o1334(.A0(ori_ori_n1382_), .A1(ori_ori_n1381_), .B0(ori_ori_n1383_), .Y(ori_ori_n1384_));
  NO3        o1335(.A(x8), .B(x6), .C(ori_ori_n50_), .Y(ori_ori_n1385_));
  NO2        o1336(.A(ori_ori_n727_), .B(ori_ori_n182_), .Y(ori_ori_n1386_));
  OAI210     o1337(.A0(ori_ori_n1385_), .A1(ori_ori_n236_), .B0(ori_ori_n1386_), .Y(ori_ori_n1387_));
  NO2        o1338(.A(ori_ori_n159_), .B(x5), .Y(ori_ori_n1388_));
  INV        o1339(.A(ori_ori_n1387_), .Y(ori_ori_n1389_));
  OAI210     o1340(.A0(ori_ori_n1389_), .A1(ori_ori_n1384_), .B0(ori_ori_n1380_), .Y(ori_ori_n1390_));
  OAI210     o1341(.A0(ori_ori_n1265_), .A1(ori_ori_n916_), .B0(ori_ori_n419_), .Y(ori_ori_n1391_));
  NO2        o1342(.A(ori_ori_n317_), .B(x7), .Y(ori_ori_n1392_));
  NA2        o1343(.A(ori_ori_n1392_), .B(x0), .Y(ori_ori_n1393_));
  AOI210     o1344(.A0(ori_ori_n1393_), .A1(ori_ori_n1391_), .B0(ori_ori_n635_), .Y(ori_ori_n1394_));
  NA2        o1345(.A(ori_ori_n1064_), .B(ori_ori_n195_), .Y(ori_ori_n1395_));
  NA2        o1346(.A(ori_ori_n55_), .B(ori_ori_n104_), .Y(ori_ori_n1396_));
  NA2        o1347(.A(ori_ori_n1396_), .B(ori_ori_n681_), .Y(ori_ori_n1397_));
  NA2        o1348(.A(ori_ori_n374_), .B(ori_ori_n1068_), .Y(ori_ori_n1398_));
  OA220      o1349(.A0(ori_ori_n1398_), .A1(ori_ori_n1397_), .B0(ori_ori_n1395_), .B1(ori_ori_n631_), .Y(ori_ori_n1399_));
  OAI210     o1350(.A0(ori_ori_n1399_), .A1(ori_ori_n650_), .B0(ori_ori_n496_), .Y(ori_ori_n1400_));
  INV        o1351(.A(ori_ori_n1009_), .Y(ori_ori_n1401_));
  NO2        o1352(.A(ori_ori_n1401_), .B(ori_ori_n62_), .Y(ori_ori_n1402_));
  AOI220     o1353(.A0(ori_ori_n1402_), .A1(ori_ori_n267_), .B0(ori_ori_n1251_), .B1(ori_ori_n124_), .Y(ori_ori_n1403_));
  AOI220     o1354(.A0(ori_ori_n634_), .A1(ori_ori_n360_), .B0(ori_ori_n624_), .B1(ori_ori_n88_), .Y(ori_ori_n1404_));
  NA3        o1355(.A(ori_ori_n462_), .B(ori_ori_n586_), .C(ori_ori_n189_), .Y(ori_ori_n1405_));
  OAI220     o1356(.A0(ori_ori_n1405_), .A1(ori_ori_n1404_), .B0(ori_ori_n1403_), .B1(ori_ori_n308_), .Y(ori_ori_n1406_));
  NO3        o1357(.A(ori_ori_n1406_), .B(ori_ori_n1400_), .C(ori_ori_n1394_), .Y(ori_ori_n1407_));
  NO3        o1358(.A(x6), .B(x4), .C(x3), .Y(ori_ori_n1408_));
  NA2        o1359(.A(ori_ori_n1408_), .B(ori_ori_n533_), .Y(ori_ori_n1409_));
  NA4        o1360(.A(ori_ori_n703_), .B(ori_ori_n182_), .C(ori_ori_n58_), .D(x6), .Y(ori_ori_n1410_));
  AOI210     o1361(.A0(ori_ori_n1410_), .A1(ori_ori_n1409_), .B0(ori_ori_n54_), .Y(ori_ori_n1411_));
  NO2        o1362(.A(ori_ori_n718_), .B(x3), .Y(ori_ori_n1412_));
  AOI210     o1363(.A0(ori_ori_n659_), .A1(ori_ori_n146_), .B0(ori_ori_n1050_), .Y(ori_ori_n1413_));
  OA210      o1364(.A0(ori_ori_n1412_), .A1(ori_ori_n422_), .B0(ori_ori_n1413_), .Y(ori_ori_n1414_));
  NO2        o1365(.A(ori_ori_n755_), .B(ori_ori_n510_), .Y(ori_ori_n1415_));
  NO3        o1366(.A(ori_ori_n1415_), .B(ori_ori_n257_), .C(ori_ori_n154_), .Y(ori_ori_n1416_));
  NO3        o1367(.A(ori_ori_n1416_), .B(ori_ori_n1414_), .C(ori_ori_n1411_), .Y(ori_ori_n1417_));
  NA2        o1368(.A(ori_ori_n405_), .B(ori_ori_n948_), .Y(ori_ori_n1418_));
  NA4        o1369(.A(ori_ori_n481_), .B(ori_ori_n367_), .C(ori_ori_n219_), .D(x6), .Y(ori_ori_n1419_));
  OAI210     o1370(.A0(ori_ori_n718_), .A1(ori_ori_n1418_), .B0(ori_ori_n1419_), .Y(ori_ori_n1420_));
  NA2        o1371(.A(ori_ori_n898_), .B(ori_ori_n1294_), .Y(ori_ori_n1421_));
  NA2        o1372(.A(ori_ori_n724_), .B(x7), .Y(ori_ori_n1422_));
  OAI210     o1373(.A0(ori_ori_n1422_), .A1(ori_ori_n386_), .B0(ori_ori_n1421_), .Y(ori_ori_n1423_));
  NA2        o1374(.A(ori_ori_n274_), .B(x2), .Y(ori_ori_n1424_));
  NO3        o1375(.A(ori_ori_n1424_), .B(ori_ori_n594_), .C(ori_ori_n72_), .Y(ori_ori_n1425_));
  AOI210     o1376(.A0(ori_ori_n580_), .A1(ori_ori_n50_), .B0(ori_ori_n589_), .Y(ori_ori_n1426_));
  OAI210     o1377(.A0(ori_ori_n917_), .A1(ori_ori_n936_), .B0(ori_ori_n381_), .Y(ori_ori_n1427_));
  OAI220     o1378(.A0(ori_ori_n1427_), .A1(ori_ori_n1426_), .B0(ori_ori_n772_), .B1(ori_ori_n187_), .Y(ori_ori_n1428_));
  NO4        o1379(.A(ori_ori_n1428_), .B(ori_ori_n1425_), .C(ori_ori_n1423_), .D(ori_ori_n1420_), .Y(ori_ori_n1429_));
  OA220      o1380(.A0(ori_ori_n1429_), .A1(ori_ori_n442_), .B0(ori_ori_n1417_), .B1(ori_ori_n202_), .Y(ori_ori_n1430_));
  NO2        o1381(.A(ori_ori_n912_), .B(ori_ori_n55_), .Y(ori_ori_n1431_));
  NA2        o1382(.A(ori_ori_n416_), .B(ori_ori_n797_), .Y(ori_ori_n1432_));
  NO2        o1383(.A(ori_ori_n1432_), .B(ori_ori_n1431_), .Y(ori_ori_n1433_));
  NO3        o1384(.A(ori_ori_n949_), .B(ori_ori_n330_), .C(x8), .Y(ori_ori_n1434_));
  OAI210     o1385(.A0(ori_ori_n1434_), .A1(ori_ori_n1433_), .B0(x6), .Y(ori_ori_n1435_));
  NO2        o1386(.A(ori_ori_n1080_), .B(ori_ori_n1042_), .Y(ori_ori_n1436_));
  NA2        o1387(.A(ori_ori_n187_), .B(x7), .Y(ori_ori_n1437_));
  OAI220     o1388(.A0(ori_ori_n1437_), .A1(ori_ori_n1436_), .B0(ori_ori_n757_), .B1(ori_ori_n87_), .Y(ori_ori_n1438_));
  NA2        o1389(.A(ori_ori_n1438_), .B(ori_ori_n917_), .Y(ori_ori_n1439_));
  NA2        o1390(.A(ori_ori_n866_), .B(ori_ori_n71_), .Y(ori_ori_n1440_));
  OAI210     o1391(.A0(ori_ori_n1440_), .A1(ori_ori_n157_), .B0(ori_ori_n998_), .Y(ori_ori_n1441_));
  AOI210     o1392(.A0(ori_ori_n498_), .A1(ori_ori_n57_), .B0(ori_ori_n631_), .Y(ori_ori_n1442_));
  NA3        o1393(.A(ori_ori_n225_), .B(ori_ori_n76_), .C(ori_ori_n71_), .Y(ori_ori_n1443_));
  OAI210     o1394(.A0(ori_ori_n908_), .A1(ori_ori_n228_), .B0(ori_ori_n1443_), .Y(ori_ori_n1444_));
  AOI210     o1395(.A0(ori_ori_n1442_), .A1(ori_ori_n1441_), .B0(ori_ori_n1444_), .Y(ori_ori_n1445_));
  NA3        o1396(.A(ori_ori_n1445_), .B(ori_ori_n1439_), .C(ori_ori_n1435_), .Y(ori_ori_n1446_));
  NO2        o1397(.A(ori_ori_n636_), .B(x6), .Y(ori_ori_n1447_));
  OAI210     o1398(.A0(ori_ori_n381_), .A1(ori_ori_n84_), .B0(ori_ori_n379_), .Y(ori_ori_n1448_));
  OA210      o1399(.A0(ori_ori_n1448_), .A1(ori_ori_n1447_), .B0(ori_ori_n129_), .Y(ori_ori_n1449_));
  NO3        o1400(.A(ori_ori_n444_), .B(ori_ori_n384_), .C(x7), .Y(ori_ori_n1450_));
  NO3        o1401(.A(ori_ori_n159_), .B(ori_ori_n75_), .C(x2), .Y(ori_ori_n1451_));
  NO3        o1402(.A(ori_ori_n1451_), .B(ori_ori_n1450_), .C(ori_ori_n1449_), .Y(ori_ori_n1452_));
  NO2        o1403(.A(ori_ori_n228_), .B(x1), .Y(ori_ori_n1453_));
  OAI210     o1404(.A0(ori_ori_n1453_), .A1(ori_ori_n449_), .B0(ori_ori_n510_), .Y(ori_ori_n1454_));
  NO2        o1405(.A(ori_ori_n57_), .B(ori_ori_n104_), .Y(ori_ori_n1455_));
  NA2        o1406(.A(ori_ori_n1073_), .B(ori_ori_n1455_), .Y(ori_ori_n1456_));
  AOI210     o1407(.A0(ori_ori_n1456_), .A1(ori_ori_n1454_), .B0(ori_ori_n56_), .Y(ori_ori_n1457_));
  AOI220     o1408(.A0(ori_ori_n757_), .A1(ori_ori_n768_), .B0(ori_ori_n513_), .B1(ori_ori_n278_), .Y(ori_ori_n1458_));
  NO2        o1409(.A(ori_ori_n1458_), .B(ori_ori_n1294_), .Y(ori_ori_n1459_));
  NO3        o1410(.A(ori_ori_n533_), .B(ori_ori_n171_), .C(ori_ori_n1042_), .Y(ori_ori_n1460_));
  NA2        o1411(.A(ori_ori_n936_), .B(x4), .Y(ori_ori_n1461_));
  OAI220     o1412(.A0(ori_ori_n1461_), .A1(ori_ori_n686_), .B0(ori_ori_n644_), .B1(ori_ori_n610_), .Y(ori_ori_n1462_));
  NO4        o1413(.A(ori_ori_n1462_), .B(ori_ori_n1460_), .C(ori_ori_n1459_), .D(ori_ori_n1457_), .Y(ori_ori_n1463_));
  OAI210     o1414(.A0(ori_ori_n1452_), .A1(x5), .B0(ori_ori_n1463_), .Y(ori_ori_n1464_));
  AOI220     o1415(.A0(ori_ori_n1464_), .A1(ori_ori_n95_), .B0(ori_ori_n1446_), .B1(ori_ori_n337_), .Y(ori_ori_n1465_));
  NA4        o1416(.A(ori_ori_n1465_), .B(ori_ori_n1430_), .C(ori_ori_n1407_), .D(ori_ori_n1390_), .Y(ori17));
  NO4        o1417(.A(ori_ori_n601_), .B(ori_ori_n697_), .C(ori_ori_n98_), .D(ori_ori_n97_), .Y(ori_ori_n1467_));
  NO2        o1418(.A(ori_ori_n122_), .B(ori_ori_n1157_), .Y(ori_ori_n1468_));
  AOI220     o1419(.A0(ori_ori_n1468_), .A1(ori_ori_n713_), .B0(ori_ori_n1467_), .B1(ori_ori_n504_), .Y(ori_ori_n1469_));
  NA2        o1420(.A(ori_ori_n163_), .B(ori_ori_n78_), .Y(ori_ori_n1470_));
  NOi21      o1421(.An(ori_ori_n379_), .B(ori_ori_n84_), .Y(ori_ori_n1471_));
  OAI210     o1422(.A0(ori_ori_n624_), .A1(ori_ori_n55_), .B0(ori_ori_n1471_), .Y(ori_ori_n1472_));
  NA2        o1423(.A(ori_ori_n1210_), .B(ori_ori_n1004_), .Y(ori_ori_n1473_));
  NA4        o1424(.A(ori_ori_n1473_), .B(ori_ori_n1472_), .C(ori_ori_n727_), .D(ori_ori_n57_), .Y(ori_ori_n1474_));
  OAI210     o1425(.A0(ori_ori_n703_), .A1(x8), .B0(ori_ori_n1294_), .Y(ori_ori_n1475_));
  NA3        o1426(.A(ori_ori_n1475_), .B(ori_ori_n1235_), .C(ori_ori_n398_), .Y(ori_ori_n1476_));
  NA3        o1427(.A(ori_ori_n392_), .B(ori_ori_n267_), .C(ori_ori_n585_), .Y(ori_ori_n1477_));
  BUFFER     o1428(.A(ori_ori_n747_), .Y(ori_ori_n1478_));
  NA4        o1429(.A(ori_ori_n1478_), .B(ori_ori_n1477_), .C(ori_ori_n1476_), .D(ori_ori_n1474_), .Y(ori_ori_n1479_));
  AOI210     o1430(.A0(ori_ori_n1070_), .A1(ori_ori_n304_), .B0(ori_ori_n59_), .Y(ori_ori_n1480_));
  INV        o1431(.A(ori_ori_n1480_), .Y(ori_ori_n1481_));
  AOI210     o1432(.A0(ori_ori_n1479_), .A1(x1), .B0(ori_ori_n1481_), .Y(ori_ori_n1482_));
  NO2        o1433(.A(ori_ori_n972_), .B(ori_ori_n498_), .Y(ori_ori_n1483_));
  OAI210     o1434(.A0(ori_ori_n1483_), .A1(ori_ori_n1054_), .B0(ori_ori_n607_), .Y(ori_ori_n1484_));
  NO3        o1435(.A(ori_ori_n631_), .B(ori_ori_n555_), .C(ori_ori_n524_), .Y(ori_ori_n1485_));
  OAI210     o1436(.A0(ori_ori_n1485_), .A1(ori_ori_n897_), .B0(ori_ori_n1412_), .Y(ori_ori_n1486_));
  AOI210     o1437(.A0(ori_ori_n1486_), .A1(ori_ori_n1484_), .B0(x8), .Y(ori_ori_n1487_));
  NA3        o1438(.A(ori_ori_n631_), .B(ori_ori_n270_), .C(ori_ori_n119_), .Y(ori_ori_n1488_));
  NO2        o1439(.A(ori_ori_n142_), .B(ori_ori_n140_), .Y(ori_ori_n1489_));
  NO3        o1440(.A(ori_ori_n893_), .B(ori_ori_n768_), .C(ori_ori_n697_), .Y(ori_ori_n1490_));
  AOI210     o1441(.A0(ori_ori_n1490_), .A1(ori_ori_n1489_), .B0(x0), .Y(ori_ori_n1491_));
  OAI210     o1442(.A0(ori_ori_n1488_), .A1(ori_ori_n246_), .B0(ori_ori_n1491_), .Y(ori_ori_n1492_));
  NO2        o1443(.A(ori_ori_n1492_), .B(ori_ori_n1487_), .Y(ori_ori_n1493_));
  OAI220     o1444(.A0(ori_ori_n1493_), .A1(ori_ori_n1482_), .B0(ori_ori_n1470_), .B1(ori_ori_n1469_), .Y(ori18));
  AOI210     o1445(.A0(x8), .A1(x0), .B0(x5), .Y(ori_ori_n1495_));
  NOi31      o1446(.An(ori_ori_n304_), .B(ori_ori_n1495_), .C(ori_ori_n1040_), .Y(ori_ori_n1496_));
  NA2        o1447(.A(ori_ori_n601_), .B(ori_ori_n59_), .Y(ori_ori_n1497_));
  AOI210     o1448(.A0(ori_ori_n1395_), .A1(ori_ori_n348_), .B0(ori_ori_n1497_), .Y(ori_ori_n1498_));
  NO2        o1449(.A(ori_ori_n617_), .B(ori_ori_n769_), .Y(ori_ori_n1499_));
  NO4        o1450(.A(ori_ori_n253_), .B(ori_ori_n807_), .C(ori_ori_n153_), .D(ori_ori_n70_), .Y(ori_ori_n1500_));
  NO4        o1451(.A(ori_ori_n1500_), .B(ori_ori_n1499_), .C(ori_ori_n1498_), .D(ori_ori_n1496_), .Y(ori_ori_n1501_));
  NA3        o1452(.A(ori_ori_n519_), .B(ori_ori_n213_), .C(x0), .Y(ori_ori_n1502_));
  NAi21      o1453(.An(ori_ori_n385_), .B(ori_ori_n1502_), .Y(ori_ori_n1503_));
  NO2        o1454(.A(ori_ori_n883_), .B(x5), .Y(ori_ori_n1504_));
  AOI210     o1455(.A0(ori_ori_n1135_), .A1(x5), .B0(ori_ori_n1504_), .Y(ori_ori_n1505_));
  OA220      o1456(.A0(ori_ori_n519_), .A1(ori_ori_n330_), .B0(ori_ori_n398_), .B1(x5), .Y(ori_ori_n1506_));
  OAI220     o1457(.A0(ori_ori_n1506_), .A1(ori_ori_n292_), .B0(ori_ori_n1505_), .B1(ori_ori_n211_), .Y(ori_ori_n1507_));
  AOI210     o1458(.A0(ori_ori_n1503_), .A1(ori_ori_n290_), .B0(ori_ori_n1507_), .Y(ori_ori_n1508_));
  AOI210     o1459(.A0(ori_ori_n1508_), .A1(ori_ori_n1501_), .B0(x6), .Y(ori_ori_n1509_));
  NA3        o1460(.A(ori_ori_n523_), .B(ori_ori_n419_), .C(x2), .Y(ori_ori_n1510_));
  NA3        o1461(.A(ori_ori_n1040_), .B(ori_ori_n51_), .C(ori_ori_n57_), .Y(ori_ori_n1511_));
  AOI210     o1462(.A0(ori_ori_n1511_), .A1(ori_ori_n1510_), .B0(ori_ori_n782_), .Y(ori_ori_n1512_));
  AOI210     o1463(.A0(ori_ori_n423_), .A1(ori_ori_n136_), .B0(ori_ori_n780_), .Y(ori_ori_n1513_));
  NA2        o1464(.A(ori_ori_n267_), .B(x6), .Y(ori_ori_n1514_));
  OAI210     o1465(.A0(ori_ori_n176_), .A1(ori_ori_n106_), .B0(ori_ori_n1141_), .Y(ori_ori_n1515_));
  OAI220     o1466(.A0(ori_ori_n1515_), .A1(ori_ori_n1514_), .B0(ori_ori_n1513_), .B1(ori_ori_n739_), .Y(ori_ori_n1516_));
  OAI210     o1467(.A0(ori_ori_n1516_), .A1(ori_ori_n1512_), .B0(ori_ori_n53_), .Y(ori_ori_n1517_));
  NO2        o1468(.A(ori_ori_n685_), .B(ori_ori_n260_), .Y(ori_ori_n1518_));
  NO2        o1469(.A(ori_ori_n263_), .B(x3), .Y(ori_ori_n1519_));
  NO3        o1470(.A(ori_ori_n433_), .B(ori_ori_n601_), .C(ori_ori_n831_), .Y(ori_ori_n1520_));
  OAI210     o1471(.A0(ori_ori_n1520_), .A1(ori_ori_n1518_), .B0(ori_ori_n1519_), .Y(ori_ori_n1521_));
  AOI210     o1472(.A0(ori_ori_n1144_), .A1(ori_ori_n616_), .B0(x4), .Y(ori_ori_n1522_));
  OAI210     o1473(.A0(ori_ori_n555_), .A1(ori_ori_n601_), .B0(ori_ori_n59_), .Y(ori_ori_n1523_));
  OAI210     o1474(.A0(ori_ori_n624_), .A1(ori_ori_n646_), .B0(ori_ori_n1523_), .Y(ori_ori_n1524_));
  AO220      o1475(.A0(ori_ori_n1254_), .A1(ori_ori_n727_), .B0(ori_ori_n556_), .B1(ori_ori_n353_), .Y(ori_ori_n1525_));
  AOI220     o1476(.A0(ori_ori_n1525_), .A1(x1), .B0(ori_ori_n1524_), .B1(ori_ori_n160_), .Y(ori_ori_n1526_));
  NA4        o1477(.A(ori_ori_n1526_), .B(ori_ori_n1522_), .C(ori_ori_n1521_), .D(ori_ori_n1517_), .Y(ori_ori_n1527_));
  NO3        o1478(.A(ori_ori_n1061_), .B(ori_ori_n129_), .C(ori_ori_n128_), .Y(ori_ori_n1528_));
  OAI210     o1479(.A0(ori_ori_n1528_), .A1(ori_ori_n651_), .B0(ori_ori_n104_), .Y(ori_ori_n1529_));
  AOI210     o1480(.A0(ori_ori_n1529_), .A1(ori_ori_n561_), .B0(ori_ori_n782_), .Y(ori_ori_n1530_));
  NA3        o1481(.A(ori_ori_n1202_), .B(ori_ori_n187_), .C(ori_ori_n139_), .Y(ori_ori_n1531_));
  NA3        o1482(.A(ori_ori_n1064_), .B(ori_ori_n771_), .C(ori_ori_n341_), .Y(ori_ori_n1532_));
  NA2        o1483(.A(ori_ori_n169_), .B(ori_ori_n768_), .Y(ori_ori_n1533_));
  OAI210     o1484(.A0(ori_ori_n1533_), .A1(ori_ori_n1306_), .B0(ori_ori_n1532_), .Y(ori_ori_n1534_));
  AOI210     o1485(.A0(ori_ori_n1531_), .A1(ori_ori_n175_), .B0(ori_ori_n1534_), .Y(ori_ori_n1535_));
  OAI210     o1486(.A0(ori_ori_n1535_), .A1(ori_ori_n542_), .B0(x4), .Y(ori_ori_n1536_));
  OAI220     o1487(.A0(ori_ori_n1536_), .A1(ori_ori_n1530_), .B0(ori_ori_n1527_), .B1(ori_ori_n1509_), .Y(ori_ori_n1537_));
  NO2        o1488(.A(ori_ori_n145_), .B(ori_ori_n120_), .Y(ori_ori_n1538_));
  NO2        o1489(.A(ori_ori_n187_), .B(ori_ori_n797_), .Y(ori_ori_n1539_));
  AOI210     o1490(.A0(ori_ori_n602_), .A1(ori_ori_n510_), .B0(ori_ori_n1539_), .Y(ori_ori_n1540_));
  NO2        o1491(.A(ori_ori_n1540_), .B(x6), .Y(ori_ori_n1541_));
  NO2        o1492(.A(ori_ori_n384_), .B(ori_ori_n252_), .Y(ori_ori_n1542_));
  NO2        o1493(.A(ori_ori_n129_), .B(ori_ori_n729_), .Y(ori_ori_n1543_));
  NO2        o1494(.A(ori_ori_n949_), .B(ori_ori_n585_), .Y(ori_ori_n1544_));
  AO220      o1495(.A0(ori_ori_n1544_), .A1(ori_ori_n1543_), .B0(ori_ori_n1542_), .B1(ori_ori_n122_), .Y(ori_ori_n1545_));
  NO3        o1496(.A(ori_ori_n1545_), .B(ori_ori_n1541_), .C(ori_ori_n1538_), .Y(ori_ori_n1546_));
  NA2        o1497(.A(ori_ori_n1061_), .B(x3), .Y(ori_ori_n1547_));
  NA2        o1498(.A(ori_ori_n1343_), .B(ori_ori_n131_), .Y(ori_ori_n1548_));
  OAI220     o1499(.A0(ori_ori_n1548_), .A1(ori_ori_n1547_), .B0(ori_ori_n1546_), .B1(x3), .Y(ori_ori_n1549_));
  NO3        o1500(.A(ori_ori_n994_), .B(ori_ori_n685_), .C(ori_ori_n325_), .Y(ori_ori_n1550_));
  AO210      o1501(.A0(ori_ori_n1023_), .A1(ori_ori_n297_), .B0(ori_ori_n1550_), .Y(ori_ori_n1551_));
  AOI220     o1502(.A0(ori_ori_n1551_), .A1(x8), .B0(ori_ori_n1343_), .B1(ori_ori_n434_), .Y(ori_ori_n1552_));
  NA2        o1503(.A(ori_ori_n743_), .B(ori_ori_n316_), .Y(ori_ori_n1553_));
  NO4        o1504(.A(ori_ori_n365_), .B(ori_ori_n200_), .C(ori_ori_n336_), .D(x2), .Y(ori_ori_n1554_));
  NA2        o1505(.A(ori_ori_n1396_), .B(ori_ori_n106_), .Y(ori_ori_n1555_));
  NO3        o1506(.A(ori_ori_n1204_), .B(ori_ori_n987_), .C(ori_ori_n1141_), .Y(ori_ori_n1556_));
  AOI210     o1507(.A0(ori_ori_n1556_), .A1(ori_ori_n1555_), .B0(ori_ori_n1554_), .Y(ori_ori_n1557_));
  OA220      o1508(.A0(ori_ori_n1557_), .A1(ori_ori_n949_), .B0(ori_ori_n1553_), .B1(ori_ori_n570_), .Y(ori_ori_n1558_));
  OAI210     o1509(.A0(ori_ori_n1552_), .A1(ori_ori_n408_), .B0(ori_ori_n1558_), .Y(ori_ori_n1559_));
  AOI210     o1510(.A0(ori_ori_n1549_), .A1(ori_ori_n136_), .B0(ori_ori_n1559_), .Y(ori_ori_n1560_));
  NA2        o1511(.A(ori_ori_n1560_), .B(ori_ori_n1537_), .Y(ori19));
  NO2        o1512(.A(ori_ori_n1440_), .B(ori_ori_n256_), .Y(ori_ori_n1562_));
  NA2        o1513(.A(ori_ori_n646_), .B(x3), .Y(ori_ori_n1563_));
  OAI210     o1514(.A0(ori_ori_n153_), .A1(ori_ori_n105_), .B0(ori_ori_n81_), .Y(ori_ori_n1564_));
  NA3        o1515(.A(ori_ori_n1564_), .B(ori_ori_n1563_), .C(ori_ori_n239_), .Y(ori_ori_n1565_));
  NO2        o1516(.A(ori_ori_n1301_), .B(ori_ori_n169_), .Y(ori_ori_n1566_));
  AOI210     o1517(.A0(ori_ori_n1467_), .A1(ori_ori_n351_), .B0(ori_ori_n1566_), .Y(ori_ori_n1567_));
  AOI210     o1518(.A0(ori_ori_n1567_), .A1(ori_ori_n1565_), .B0(ori_ori_n56_), .Y(ori_ori_n1568_));
  NO2        o1519(.A(ori_ori_n856_), .B(ori_ori_n1217_), .Y(ori_ori_n1569_));
  OAI210     o1520(.A0(ori_ori_n1568_), .A1(ori_ori_n1562_), .B0(ori_ori_n1569_), .Y(ori_ori_n1570_));
  NOi21      o1521(.An(ori_ori_n611_), .B(ori_ori_n650_), .Y(ori_ori_n1571_));
  AOI210     o1522(.A0(ori_ori_n351_), .A1(x6), .B0(ori_ori_n119_), .Y(ori_ori_n1572_));
  NO3        o1523(.A(ori_ori_n1572_), .B(ori_ori_n752_), .C(ori_ori_n124_), .Y(ori_ori_n1573_));
  NA2        o1524(.A(ori_ori_n1197_), .B(ori_ori_n120_), .Y(ori_ori_n1574_));
  NO4        o1525(.A(ori_ori_n1574_), .B(ori_ori_n994_), .C(ori_ori_n883_), .D(ori_ori_n77_), .Y(ori_ori_n1575_));
  NO3        o1526(.A(ori_ori_n1575_), .B(ori_ori_n1573_), .C(ori_ori_n1020_), .Y(ori_ori_n1576_));
  NO2        o1527(.A(ori_ori_n542_), .B(ori_ori_n620_), .Y(ori_ori_n1577_));
  NA2        o1528(.A(ori_ori_n1250_), .B(ori_ori_n50_), .Y(ori_ori_n1578_));
  NO3        o1529(.A(ori_ori_n517_), .B(ori_ori_n306_), .C(ori_ori_n64_), .Y(ori_ori_n1579_));
  AOI220     o1530(.A0(ori_ori_n1579_), .A1(ori_ori_n1578_), .B0(ori_ori_n1577_), .B1(ori_ori_n771_), .Y(ori_ori_n1580_));
  OAI210     o1531(.A0(ori_ori_n1576_), .A1(ori_ori_n57_), .B0(ori_ori_n1580_), .Y(ori_ori_n1581_));
  AOI210     o1532(.A0(ori_ori_n1581_), .A1(ori_ori_n768_), .B0(ori_ori_n1571_), .Y(ori_ori_n1582_));
  AOI210     o1533(.A0(ori_ori_n817_), .A1(ori_ori_n729_), .B0(ori_ori_n758_), .Y(ori_ori_n1583_));
  NO2        o1534(.A(ori_ori_n1583_), .B(x4), .Y(ori_ori_n1584_));
  NA3        o1535(.A(ori_ori_n727_), .B(ori_ori_n255_), .C(x7), .Y(ori_ori_n1585_));
  AOI220     o1536(.A0(ori_ori_n1392_), .A1(ori_ori_n782_), .B0(ori_ori_n697_), .B1(ori_ori_n1157_), .Y(ori_ori_n1586_));
  AOI210     o1537(.A0(ori_ori_n1586_), .A1(ori_ori_n1585_), .B0(ori_ori_n502_), .Y(ori_ori_n1587_));
  OAI210     o1538(.A0(ori_ori_n1587_), .A1(ori_ori_n1584_), .B0(ori_ori_n807_), .Y(ori_ori_n1588_));
  NO2        o1539(.A(ori_ori_n739_), .B(ori_ori_n320_), .Y(ori_ori_n1589_));
  NO2        o1540(.A(ori_ori_n153_), .B(ori_ori_n1019_), .Y(ori_ori_n1590_));
  AOI220     o1541(.A0(ori_ori_n1590_), .A1(ori_ori_n1265_), .B0(ori_ori_n1589_), .B1(ori_ori_n476_), .Y(ori_ori_n1591_));
  AO210      o1542(.A0(ori_ori_n1591_), .A1(ori_ori_n1588_), .B0(x1), .Y(ori_ori_n1592_));
  NA3        o1543(.A(ori_ori_n631_), .B(ori_ori_n1042_), .C(ori_ori_n1189_), .Y(ori_ori_n1593_));
  NA2        o1544(.A(ori_ori_n146_), .B(ori_ori_n107_), .Y(ori_ori_n1594_));
  NOi21      o1545(.An(x1), .B(x6), .Y(ori_ori_n1595_));
  NA2        o1546(.A(ori_ori_n1595_), .B(ori_ori_n84_), .Y(ori_ori_n1596_));
  NA3        o1547(.A(ori_ori_n1596_), .B(ori_ori_n1594_), .C(ori_ori_n1593_), .Y(ori_ori_n1597_));
  AOI220     o1548(.A0(ori_ori_n1597_), .A1(x3), .B0(ori_ori_n1205_), .B1(ori_ori_n380_), .Y(ori_ori_n1598_));
  NA3        o1549(.A(ori_ori_n1210_), .B(ori_ori_n792_), .C(ori_ori_n603_), .Y(ori_ori_n1599_));
  AOI220     o1550(.A0(ori_ori_n1254_), .A1(ori_ori_n119_), .B0(ori_ori_n912_), .B1(ori_ori_n809_), .Y(ori_ori_n1600_));
  AOI210     o1551(.A0(ori_ori_n1600_), .A1(ori_ori_n1599_), .B0(ori_ori_n320_), .Y(ori_ori_n1601_));
  NA2        o1552(.A(ori_ori_n936_), .B(ori_ori_n50_), .Y(ori_ori_n1602_));
  NA3        o1553(.A(ori_ori_n1197_), .B(ori_ori_n381_), .C(ori_ori_n106_), .Y(ori_ori_n1603_));
  AOI210     o1554(.A0(ori_ori_n1603_), .A1(ori_ori_n1602_), .B0(ori_ori_n957_), .Y(ori_ori_n1604_));
  NO2        o1555(.A(ori_ori_n1604_), .B(ori_ori_n1601_), .Y(ori_ori_n1605_));
  OAI210     o1556(.A0(ori_ori_n1598_), .A1(ori_ori_n843_), .B0(ori_ori_n1605_), .Y(ori_ori_n1606_));
  NO2        o1557(.A(ori_ori_n555_), .B(ori_ori_n68_), .Y(ori_ori_n1607_));
  OAI220     o1558(.A0(ori_ori_n1607_), .A1(ori_ori_n1563_), .B0(ori_ori_n305_), .B1(ori_ori_n891_), .Y(ori_ori_n1608_));
  AOI220     o1559(.A0(ori_ori_n1608_), .A1(ori_ori_n56_), .B0(ori_ori_n1348_), .B1(ori_ori_n724_), .Y(ori_ori_n1609_));
  NO2        o1560(.A(ori_ori_n54_), .B(ori_ori_n71_), .Y(ori_ori_n1610_));
  AO220      o1561(.A0(ori_ori_n1610_), .A1(ori_ori_n994_), .B0(ori_ori_n809_), .B1(ori_ori_n948_), .Y(ori_ori_n1611_));
  NA2        o1562(.A(ori_ori_n1180_), .B(ori_ori_n358_), .Y(ori_ori_n1612_));
  NO2        o1563(.A(ori_ori_n987_), .B(ori_ori_n1595_), .Y(ori_ori_n1613_));
  NA2        o1564(.A(ori_ori_n498_), .B(ori_ori_n724_), .Y(ori_ori_n1614_));
  OAI210     o1565(.A0(ori_ori_n1614_), .A1(ori_ori_n1613_), .B0(ori_ori_n1612_), .Y(ori_ori_n1615_));
  AOI210     o1566(.A0(ori_ori_n1611_), .A1(x2), .B0(ori_ori_n1615_), .Y(ori_ori_n1616_));
  OAI220     o1567(.A0(ori_ori_n1616_), .A1(ori_ori_n153_), .B0(ori_ori_n1609_), .B1(ori_ori_n54_), .Y(ori_ori_n1617_));
  OAI210     o1568(.A0(ori_ori_n1617_), .A1(ori_ori_n1606_), .B0(x8), .Y(ori_ori_n1618_));
  NA4        o1569(.A(ori_ori_n1618_), .B(ori_ori_n1592_), .C(ori_ori_n1582_), .D(ori_ori_n1570_), .Y(ori20));
  NA4        o1570(.A(ori_ori_n391_), .B(ori_ori_n278_), .C(ori_ori_n379_), .D(ori_ori_n62_), .Y(ori_ori_n1620_));
  NA2        o1571(.A(ori_ori_n476_), .B(ori_ori_n412_), .Y(ori_ori_n1621_));
  AOI210     o1572(.A0(ori_ori_n1621_), .A1(ori_ori_n1620_), .B0(ori_ori_n87_), .Y(ori_ori_n1622_));
  AOI210     o1573(.A0(ori_ori_n1046_), .A1(ori_ori_n62_), .B0(ori_ori_n1577_), .Y(ori_ori_n1623_));
  AOI210     o1574(.A0(ori_ori_n981_), .A1(ori_ori_n347_), .B0(ori_ori_n1187_), .Y(ori_ori_n1624_));
  OAI210     o1575(.A0(ori_ori_n1623_), .A1(ori_ori_n681_), .B0(ori_ori_n1624_), .Y(ori_ori_n1625_));
  OAI210     o1576(.A0(ori_ori_n1625_), .A1(ori_ori_n1622_), .B0(ori_ori_n1102_), .Y(ori_ori_n1626_));
  NAi21      o1577(.An(ori_ori_n551_), .B(ori_ori_n400_), .Y(ori_ori_n1627_));
  NA3        o1578(.A(ori_ori_n1627_), .B(ori_ori_n979_), .C(ori_ori_n948_), .Y(ori_ori_n1628_));
  NA2        o1579(.A(ori_ori_n1101_), .B(ori_ori_n278_), .Y(ori_ori_n1629_));
  AOI210     o1580(.A0(ori_ori_n1629_), .A1(ori_ori_n1628_), .B0(ori_ori_n1294_), .Y(ori_ori_n1630_));
  NO2        o1581(.A(ori_ori_n743_), .B(ori_ori_n967_), .Y(ori_ori_n1631_));
  NOi31      o1582(.An(ori_ori_n1631_), .B(ori_ori_n1172_), .C(ori_ori_n529_), .Y(ori_ori_n1632_));
  OAI210     o1583(.A0(ori_ori_n1632_), .A1(ori_ori_n1630_), .B0(ori_ori_n325_), .Y(ori_ori_n1633_));
  NO4        o1584(.A(ori_ori_n546_), .B(ori_ori_n234_), .C(x5), .D(x2), .Y(ori_ori_n1634_));
  NA2        o1585(.A(ori_ori_n316_), .B(ori_ori_n91_), .Y(ori_ori_n1635_));
  NA2        o1586(.A(ori_ori_n326_), .B(ori_ori_n104_), .Y(ori_ori_n1636_));
  NA2        o1587(.A(ori_ori_n422_), .B(ori_ori_n52_), .Y(ori_ori_n1637_));
  OAI220     o1588(.A0(ori_ori_n1637_), .A1(ori_ori_n1636_), .B0(ori_ori_n1635_), .B1(ori_ori_n273_), .Y(ori_ori_n1638_));
  OAI210     o1589(.A0(ori_ori_n1638_), .A1(ori_ori_n1634_), .B0(ori_ori_n219_), .Y(ori_ori_n1639_));
  NO2        o1590(.A(ori_ori_n665_), .B(ori_ori_n607_), .Y(ori_ori_n1640_));
  NA2        o1591(.A(ori_ori_n949_), .B(ori_ori_n50_), .Y(ori_ori_n1641_));
  NO3        o1592(.A(ori_ori_n1641_), .B(ori_ori_n363_), .C(ori_ori_n227_), .Y(ori_ori_n1642_));
  NA4        o1593(.A(ori_ori_n337_), .B(ori_ori_n236_), .C(ori_ori_n797_), .D(ori_ori_n64_), .Y(ori_ori_n1643_));
  OAI220     o1594(.A0(ori_ori_n1643_), .A1(ori_ori_n675_), .B0(ori_ori_n1461_), .B1(ori_ori_n1029_), .Y(ori_ori_n1644_));
  AOI210     o1595(.A0(ori_ori_n1642_), .A1(ori_ori_n1640_), .B0(ori_ori_n1644_), .Y(ori_ori_n1645_));
  NA4        o1596(.A(ori_ori_n1645_), .B(ori_ori_n1639_), .C(ori_ori_n1633_), .D(ori_ori_n1626_), .Y(ori21));
  OAI210     o1597(.A0(ori_ori_n405_), .A1(ori_ori_n54_), .B0(x7), .Y(ori_ori_n1647_));
  OAI220     o1598(.A0(ori_ori_n1647_), .A1(ori_ori_n1284_), .B0(ori_ori_n1047_), .B1(ori_ori_n92_), .Y(ori_ori_n1648_));
  NA2        o1599(.A(ori_ori_n1648_), .B(ori_ori_n78_), .Y(ori_ori_n1649_));
  NA2        o1600(.A(ori_ori_n290_), .B(ori_ori_n854_), .Y(ori_ori_n1650_));
  AOI220     o1601(.A0(ori_ori_n1650_), .A1(ori_ori_n308_), .B0(ori_ori_n570_), .B1(ori_ori_n460_), .Y(ori_ori_n1651_));
  NA2        o1602(.A(ori_ori_n936_), .B(ori_ori_n272_), .Y(ori_ori_n1652_));
  NA2        o1603(.A(ori_ori_n537_), .B(ori_ori_n461_), .Y(ori_ori_n1653_));
  NA4        o1604(.A(ori_ori_n1653_), .B(ori_ori_n1652_), .C(ori_ori_n1373_), .D(ori_ori_n56_), .Y(ori_ori_n1654_));
  NO2        o1605(.A(ori_ori_n771_), .B(ori_ori_n433_), .Y(ori_ori_n1655_));
  NO3        o1606(.A(ori_ori_n1655_), .B(ori_ori_n719_), .C(ori_ori_n248_), .Y(ori_ori_n1656_));
  NOi31      o1607(.An(ori_ori_n190_), .B(ori_ori_n631_), .C(ori_ori_n1085_), .Y(ori_ori_n1657_));
  NO4        o1608(.A(ori_ori_n1657_), .B(ori_ori_n1656_), .C(ori_ori_n1654_), .D(ori_ori_n1651_), .Y(ori_ori_n1658_));
  NO3        o1609(.A(ori_ori_n433_), .B(ori_ori_n276_), .C(ori_ori_n52_), .Y(ori_ori_n1659_));
  OA210      o1610(.A0(ori_ori_n1659_), .A1(ori_ori_n880_), .B0(x3), .Y(ori_ori_n1660_));
  OAI210     o1611(.A0(ori_ori_n781_), .A1(ori_ori_n589_), .B0(ori_ori_n339_), .Y(ori_ori_n1661_));
  NO2        o1612(.A(ori_ori_n70_), .B(x2), .Y(ori_ori_n1662_));
  OAI210     o1613(.A0(ori_ori_n175_), .A1(x0), .B0(ori_ori_n1662_), .Y(ori_ori_n1663_));
  NA2        o1614(.A(ori_ori_n143_), .B(ori_ori_n104_), .Y(ori_ori_n1664_));
  NA3        o1615(.A(ori_ori_n1664_), .B(ori_ori_n1663_), .C(ori_ori_n1661_), .Y(ori_ori_n1665_));
  OAI210     o1616(.A0(ori_ori_n1665_), .A1(ori_ori_n1660_), .B0(x8), .Y(ori_ori_n1666_));
  NO3        o1617(.A(ori_ori_n769_), .B(ori_ori_n621_), .C(ori_ori_n585_), .Y(ori_ori_n1667_));
  NA2        o1618(.A(ori_ori_n55_), .B(ori_ori_n50_), .Y(ori_ori_n1668_));
  MUX2       o1619(.S(ori_ori_n601_), .A(ori_ori_n1668_), .B(ori_ori_n103_), .Y(ori_ori_n1669_));
  AOI210     o1620(.A0(ori_ori_n1351_), .A1(ori_ori_n237_), .B0(ori_ori_n1669_), .Y(ori_ori_n1670_));
  OAI210     o1621(.A0(ori_ori_n642_), .A1(ori_ori_n584_), .B0(x4), .Y(ori_ori_n1671_));
  NO3        o1622(.A(ori_ori_n1671_), .B(ori_ori_n1670_), .C(ori_ori_n1667_), .Y(ori_ori_n1672_));
  AO220      o1623(.A0(ori_ori_n1672_), .A1(ori_ori_n1666_), .B0(ori_ori_n1658_), .B1(ori_ori_n1649_), .Y(ori_ori_n1673_));
  AO220      o1624(.A0(ori_ori_n632_), .A1(ori_ori_n320_), .B0(ori_ori_n590_), .B1(x8), .Y(ori_ori_n1674_));
  NO2        o1625(.A(ori_ori_n856_), .B(x0), .Y(ori_ori_n1675_));
  NO3        o1626(.A(ori_ori_n1675_), .B(ori_ori_n547_), .C(ori_ori_n88_), .Y(ori_ori_n1676_));
  NO2        o1627(.A(ori_ori_n159_), .B(x2), .Y(ori_ori_n1677_));
  NO3        o1628(.A(ori_ori_n376_), .B(ori_ori_n253_), .C(ori_ori_n182_), .Y(ori_ori_n1678_));
  AOI210     o1629(.A0(ori_ori_n1677_), .A1(ori_ori_n68_), .B0(ori_ori_n1678_), .Y(ori_ori_n1679_));
  OAI210     o1630(.A0(ori_ori_n1676_), .A1(ori_ori_n398_), .B0(ori_ori_n1679_), .Y(ori_ori_n1680_));
  AOI220     o1631(.A0(ori_ori_n1680_), .A1(x5), .B0(ori_ori_n1674_), .B1(ori_ori_n743_), .Y(ori_ori_n1681_));
  AOI210     o1632(.A0(ori_ori_n1681_), .A1(ori_ori_n1673_), .B0(ori_ori_n71_), .Y(ori_ori_n1682_));
  NO2        o1633(.A(ori_ori_n902_), .B(ori_ori_n168_), .Y(ori_ori_n1683_));
  NOi41      o1634(.An(ori_ori_n1424_), .B(ori_ori_n1495_), .C(ori_ori_n1156_), .D(ori_ori_n847_), .Y(ori_ori_n1684_));
  NA2        o1635(.A(ori_ori_n1684_), .B(ori_ori_n1683_), .Y(ori_ori_n1685_));
  NO2        o1636(.A(ori_ori_n78_), .B(x4), .Y(ori_ori_n1686_));
  OAI210     o1637(.A0(ori_ori_n288_), .A1(ori_ori_n157_), .B0(ori_ori_n1686_), .Y(ori_ori_n1687_));
  OAI210     o1638(.A0(ori_ori_n407_), .A1(ori_ori_n423_), .B0(ori_ori_n227_), .Y(ori_ori_n1688_));
  NO2        o1639(.A(ori_ori_n255_), .B(ori_ori_n50_), .Y(ori_ori_n1689_));
  NO2        o1640(.A(ori_ori_n1689_), .B(ori_ori_n57_), .Y(ori_ori_n1690_));
  NA2        o1641(.A(ori_ori_n1690_), .B(ori_ori_n1688_), .Y(ori_ori_n1691_));
  AOI210     o1642(.A0(ori_ori_n1687_), .A1(ori_ori_n1685_), .B0(ori_ori_n1691_), .Y(ori_ori_n1692_));
  NA2        o1643(.A(ori_ori_n755_), .B(ori_ori_n551_), .Y(ori_ori_n1693_));
  AO210      o1644(.A0(ori_ori_n1693_), .A1(ori_ori_n957_), .B0(ori_ori_n50_), .Y(ori_ori_n1694_));
  NA2        o1645(.A(ori_ori_n1320_), .B(ori_ori_n1040_), .Y(ori_ori_n1695_));
  AOI210     o1646(.A0(ori_ori_n1695_), .A1(ori_ori_n1694_), .B0(ori_ori_n106_), .Y(ori_ori_n1696_));
  NA2        o1647(.A(ori_ori_n297_), .B(ori_ori_n104_), .Y(ori_ori_n1697_));
  NA2        o1648(.A(ori_ori_n890_), .B(ori_ori_n55_), .Y(ori_ori_n1698_));
  NO2        o1649(.A(ori_ori_n1698_), .B(ori_ori_n1697_), .Y(ori_ori_n1699_));
  NO2        o1650(.A(ori_ori_n670_), .B(ori_ori_n1050_), .Y(ori_ori_n1700_));
  NO4        o1651(.A(ori_ori_n1700_), .B(ori_ori_n1699_), .C(ori_ori_n1696_), .D(ori_ori_n1692_), .Y(ori_ori_n1701_));
  NO2        o1652(.A(ori_ori_n1701_), .B(x6), .Y(ori_ori_n1702_));
  NO2        o1653(.A(ori_ori_n610_), .B(ori_ori_n1495_), .Y(ori_ori_n1703_));
  OAI210     o1654(.A0(ori_ori_n1703_), .A1(ori_ori_n688_), .B0(ori_ori_n56_), .Y(ori_ori_n1704_));
  NO2        o1655(.A(ori_ori_n745_), .B(ori_ori_n54_), .Y(ori_ori_n1705_));
  NO4        o1656(.A(ori_ori_n955_), .B(ori_ori_n276_), .C(ori_ori_n768_), .D(ori_ori_n752_), .Y(ori_ori_n1706_));
  NO2        o1657(.A(ori_ori_n861_), .B(x5), .Y(ori_ori_n1707_));
  NO4        o1658(.A(ori_ori_n1707_), .B(ori_ori_n1706_), .C(ori_ori_n1705_), .D(ori_ori_n943_), .Y(ori_ori_n1708_));
  AOI210     o1659(.A0(ori_ori_n1708_), .A1(ori_ori_n1704_), .B0(ori_ori_n50_), .Y(ori_ori_n1709_));
  NA2        o1660(.A(ori_ori_n159_), .B(ori_ori_n104_), .Y(ori_ori_n1710_));
  OA220      o1661(.A0(ori_ori_n1710_), .A1(ori_ori_n437_), .B0(ori_ori_n466_), .B1(ori_ori_n743_), .Y(ori_ori_n1711_));
  NA3        o1662(.A(ori_ori_n55_), .B(x2), .C(x0), .Y(ori_ori_n1712_));
  AOI220     o1663(.A0(ori_ori_n1712_), .A1(ori_ori_n169_), .B0(ori_ori_n861_), .B1(ori_ori_n155_), .Y(ori_ori_n1713_));
  NO2        o1664(.A(ori_ori_n681_), .B(ori_ori_n255_), .Y(ori_ori_n1714_));
  NO3        o1665(.A(ori_ori_n243_), .B(ori_ori_n225_), .C(ori_ori_n358_), .Y(ori_ori_n1715_));
  NO3        o1666(.A(ori_ori_n1715_), .B(ori_ori_n1714_), .C(ori_ori_n1713_), .Y(ori_ori_n1716_));
  OAI220     o1667(.A0(ori_ori_n1716_), .A1(ori_ori_n56_), .B0(ori_ori_n1711_), .B1(ori_ori_n695_), .Y(ori_ori_n1717_));
  OAI210     o1668(.A0(ori_ori_n1717_), .A1(ori_ori_n1709_), .B0(ori_ori_n112_), .Y(ori_ori_n1718_));
  NO2        o1669(.A(ori_ori_n615_), .B(ori_ori_n303_), .Y(ori_ori_n1719_));
  AOI210     o1670(.A0(ori_ori_n608_), .A1(x5), .B0(ori_ori_n1719_), .Y(ori_ori_n1720_));
  NO2        o1671(.A(ori_ori_n1720_), .B(ori_ori_n106_), .Y(ori_ori_n1721_));
  NA2        o1672(.A(ori_ori_n703_), .B(ori_ori_n81_), .Y(ori_ori_n1722_));
  NA3        o1673(.A(ori_ori_n1722_), .B(ori_ori_n430_), .C(ori_ori_n57_), .Y(ori_ori_n1723_));
  OAI210     o1674(.A0(ori_ori_n1698_), .A1(ori_ori_n1697_), .B0(ori_ori_n1723_), .Y(ori_ori_n1724_));
  OAI210     o1675(.A0(ori_ori_n1724_), .A1(ori_ori_n1721_), .B0(x1), .Y(ori_ori_n1725_));
  NO4        o1676(.A(ori_ori_n416_), .B(ori_ori_n78_), .C(ori_ori_n147_), .D(x3), .Y(ori_ori_n1726_));
  NO2        o1677(.A(ori_ori_n326_), .B(ori_ori_n108_), .Y(ori_ori_n1727_));
  OAI210     o1678(.A0(ori_ori_n1726_), .A1(ori_ori_n1295_), .B0(ori_ori_n1727_), .Y(ori_ori_n1728_));
  NO2        o1679(.A(ori_ori_n60_), .B(ori_ori_n104_), .Y(ori_ori_n1729_));
  NO4        o1680(.A(ori_ori_n1697_), .B(ori_ori_n955_), .C(ori_ori_n665_), .D(ori_ori_n50_), .Y(ori_ori_n1730_));
  AOI210     o1681(.A0(ori_ori_n1729_), .A1(ori_ori_n1539_), .B0(ori_ori_n1730_), .Y(ori_ori_n1731_));
  NA4        o1682(.A(ori_ori_n1731_), .B(ori_ori_n1728_), .C(ori_ori_n1725_), .D(ori_ori_n1718_), .Y(ori_ori_n1732_));
  NO3        o1683(.A(ori_ori_n1732_), .B(ori_ori_n1702_), .C(ori_ori_n1682_), .Y(ori22));
  AOI210     o1684(.A0(ori_ori_n523_), .A1(ori_ori_n71_), .B0(ori_ori_n469_), .Y(ori_ori_n1734_));
  NO3        o1685(.A(ori_ori_n1192_), .B(ori_ori_n555_), .C(ori_ori_n697_), .Y(ori_ori_n1735_));
  AOI210     o1686(.A0(x5), .A1(x2), .B0(x8), .Y(ori_ori_n1736_));
  NA2        o1687(.A(ori_ori_n1736_), .B(ori_ori_n59_), .Y(ori_ori_n1737_));
  OAI220     o1688(.A0(ori_ori_n1737_), .A1(ori_ori_n1735_), .B0(ori_ori_n1734_), .B1(ori_ori_n398_), .Y(ori_ori_n1738_));
  NA2        o1689(.A(ori_ori_n584_), .B(ori_ori_n87_), .Y(ori_ori_n1739_));
  NA2        o1690(.A(ori_ori_n273_), .B(ori_ori_n77_), .Y(ori_ori_n1740_));
  OA220      o1691(.A0(ori_ori_n1740_), .A1(ori_ori_n1739_), .B0(ori_ori_n840_), .B1(ori_ori_n1004_), .Y(ori_ori_n1741_));
  NO4        o1692(.A(ori_ori_n384_), .B(ori_ori_n217_), .C(ori_ori_n71_), .D(x3), .Y(ori_ori_n1742_));
  NO3        o1693(.A(ori_ori_n1245_), .B(ori_ori_n87_), .C(x0), .Y(ori_ori_n1743_));
  OAI210     o1694(.A0(ori_ori_n398_), .A1(ori_ori_n202_), .B0(x4), .Y(ori_ori_n1744_));
  NO3        o1695(.A(ori_ori_n1744_), .B(ori_ori_n1743_), .C(ori_ori_n1742_), .Y(ori_ori_n1745_));
  OAI210     o1696(.A0(ori_ori_n1741_), .A1(ori_ori_n195_), .B0(ori_ori_n1745_), .Y(ori_ori_n1746_));
  AOI210     o1697(.A0(ori_ori_n1738_), .A1(ori_ori_n53_), .B0(ori_ori_n1746_), .Y(ori_ori_n1747_));
  NA2        o1698(.A(ori_ori_n301_), .B(ori_ori_n306_), .Y(ori_ori_n1748_));
  NA3        o1699(.A(ori_ori_n1748_), .B(ori_ori_n219_), .C(ori_ori_n305_), .Y(ori_ori_n1749_));
  NA2        o1700(.A(ori_ori_n580_), .B(ori_ori_n242_), .Y(ori_ori_n1750_));
  NO3        o1701(.A(ori_ori_n498_), .B(ori_ori_n263_), .C(ori_ori_n211_), .Y(ori_ori_n1751_));
  NAi31      o1702(.An(ori_ori_n1751_), .B(ori_ori_n1750_), .C(ori_ori_n1749_), .Y(ori_ori_n1752_));
  NO2        o1703(.A(ori_ori_n466_), .B(ori_ori_n257_), .Y(ori_ori_n1753_));
  INV        o1704(.A(ori_ori_n1753_), .Y(ori_ori_n1754_));
  OAI210     o1705(.A0(ori_ori_n1080_), .A1(ori_ori_n184_), .B0(ori_ori_n56_), .Y(ori_ori_n1755_));
  NA3        o1706(.A(ori_ori_n55_), .B(ori_ori_n71_), .C(x0), .Y(ori_ori_n1756_));
  OAI220     o1707(.A0(ori_ori_n1756_), .A1(ori_ori_n1050_), .B0(ori_ori_n363_), .B1(ori_ori_n210_), .Y(ori_ori_n1757_));
  NO2        o1708(.A(ori_ori_n1757_), .B(ori_ori_n1755_), .Y(ori_ori_n1758_));
  OAI210     o1709(.A0(ori_ori_n1754_), .A1(ori_ori_n255_), .B0(ori_ori_n1758_), .Y(ori_ori_n1759_));
  AOI210     o1710(.A0(ori_ori_n1752_), .A1(ori_ori_n104_), .B0(ori_ori_n1759_), .Y(ori_ori_n1760_));
  AOI210     o1711(.A0(ori_ori_n947_), .A1(ori_ori_n770_), .B0(ori_ori_n865_), .Y(ori_ori_n1761_));
  OAI210     o1712(.A0(ori_ori_n799_), .A1(ori_ori_n159_), .B0(ori_ori_n933_), .Y(ori_ori_n1762_));
  OAI210     o1713(.A0(ori_ori_n1762_), .A1(ori_ori_n1761_), .B0(ori_ori_n614_), .Y(ori_ori_n1763_));
  OA210      o1714(.A0(ori_ori_n1760_), .A1(ori_ori_n1747_), .B0(ori_ori_n1763_), .Y(ori_ori_n1764_));
  OAI210     o1715(.A0(ori_ori_n1174_), .A1(ori_ori_n702_), .B0(ori_ori_n692_), .Y(ori_ori_n1765_));
  NO2        o1716(.A(ori_ori_n352_), .B(x0), .Y(ori_ori_n1766_));
  NO2        o1717(.A(ori_ori_n1765_), .B(ori_ori_n398_), .Y(ori_ori_n1767_));
  NO3        o1718(.A(ori_ori_n169_), .B(ori_ori_n159_), .C(ori_ori_n62_), .Y(ori_ori_n1768_));
  OAI210     o1719(.A0(ori_ori_n1768_), .A1(ori_ori_n418_), .B0(ori_ori_n106_), .Y(ori_ori_n1769_));
  NA2        o1720(.A(ori_ori_n139_), .B(ori_ori_n782_), .Y(ori_ori_n1770_));
  NA2        o1721(.A(ori_ori_n416_), .B(x3), .Y(ori_ori_n1771_));
  NAi31      o1722(.An(ori_ori_n1771_), .B(ori_ori_n1770_), .C(ori_ori_n1555_), .Y(ori_ori_n1772_));
  NO3        o1723(.A(ori_ori_n856_), .B(ori_ori_n465_), .C(ori_ori_n106_), .Y(ori_ori_n1773_));
  NO2        o1724(.A(ori_ori_n1082_), .B(ori_ori_n140_), .Y(ori_ori_n1774_));
  NO3        o1725(.A(ori_ori_n893_), .B(ori_ori_n412_), .C(ori_ori_n302_), .Y(ori_ori_n1775_));
  AOI220     o1726(.A0(ori_ori_n1775_), .A1(ori_ori_n1774_), .B0(ori_ori_n1773_), .B1(ori_ori_n1766_), .Y(ori_ori_n1776_));
  NA3        o1727(.A(ori_ori_n412_), .B(ori_ori_n91_), .C(ori_ori_n81_), .Y(ori_ori_n1777_));
  AOI210     o1728(.A0(ori_ori_n610_), .A1(ori_ori_n455_), .B0(ori_ori_n495_), .Y(ori_ori_n1778_));
  NA2        o1729(.A(ori_ori_n1176_), .B(x3), .Y(ori_ori_n1779_));
  OAI210     o1730(.A0(ori_ori_n1779_), .A1(ori_ori_n1778_), .B0(ori_ori_n1777_), .Y(ori_ori_n1780_));
  NA3        o1731(.A(ori_ori_n56_), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n1781_));
  NOi21      o1732(.An(ori_ori_n83_), .B(ori_ori_n727_), .Y(ori_ori_n1782_));
  NA3        o1733(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n1783_));
  NA3        o1734(.A(ori_ori_n1783_), .B(ori_ori_n987_), .C(ori_ori_n264_), .Y(ori_ori_n1784_));
  OAI220     o1735(.A0(ori_ori_n1784_), .A1(ori_ori_n1782_), .B0(ori_ori_n1053_), .B1(ori_ori_n1781_), .Y(ori_ori_n1785_));
  AOI220     o1736(.A0(ori_ori_n1785_), .A1(ori_ori_n1064_), .B0(ori_ori_n1780_), .B1(ori_ori_n347_), .Y(ori_ori_n1786_));
  NA4        o1737(.A(ori_ori_n1786_), .B(ori_ori_n1776_), .C(ori_ori_n1772_), .D(ori_ori_n1769_), .Y(ori_ori_n1787_));
  AOI210     o1738(.A0(ori_ori_n1787_), .A1(x7), .B0(ori_ori_n1767_), .Y(ori_ori_n1788_));
  OAI210     o1739(.A0(ori_ori_n1764_), .A1(x7), .B0(ori_ori_n1788_), .Y(ori23));
  OR2        o1740(.A(ori_ori_n517_), .B(ori_ori_n219_), .Y(ori_ori_n1790_));
  AOI220     o1741(.A0(ori_ori_n1790_), .A1(ori_ori_n1631_), .B0(ori_ori_n616_), .B1(ori_ori_n293_), .Y(ori_ori_n1791_));
  NO3        o1742(.A(ori_ori_n840_), .B(ori_ori_n593_), .C(ori_ori_n488_), .Y(ori_ori_n1792_));
  NO3        o1743(.A(ori_ori_n950_), .B(ori_ori_n148_), .C(ori_ori_n113_), .Y(ori_ori_n1793_));
  AOI210     o1744(.A0(ori_ori_n1793_), .A1(ori_ori_n1025_), .B0(ori_ori_n1792_), .Y(ori_ori_n1794_));
  OAI210     o1745(.A0(ori_ori_n1791_), .A1(ori_ori_n153_), .B0(ori_ori_n1794_), .Y(ori_ori_n1795_));
  NA2        o1746(.A(ori_ori_n1795_), .B(ori_ori_n55_), .Y(ori_ori_n1796_));
  NO2        o1747(.A(ori_ori_n955_), .B(ori_ori_n515_), .Y(ori_ori_n1797_));
  AO220      o1748(.A0(ori_ori_n1280_), .A1(ori_ori_n179_), .B0(ori_ori_n994_), .B1(ori_ori_n743_), .Y(ori_ori_n1798_));
  OAI210     o1749(.A0(ori_ori_n1798_), .A1(ori_ori_n1797_), .B0(ori_ori_n590_), .Y(ori_ori_n1799_));
  NA2        o1750(.A(ori_ori_n176_), .B(ori_ori_n168_), .Y(ori_ori_n1800_));
  NA3        o1751(.A(ori_ori_n865_), .B(ori_ori_n423_), .C(ori_ori_n255_), .Y(ori_ori_n1801_));
  AOI210     o1752(.A0(ori_ori_n1801_), .A1(ori_ori_n500_), .B0(ori_ori_n381_), .Y(ori_ori_n1802_));
  NA2        o1753(.A(ori_ori_n1802_), .B(ori_ori_n297_), .Y(ori_ori_n1803_));
  NA3        o1754(.A(ori_ori_n57_), .B(x4), .C(x3), .Y(ori_ori_n1804_));
  NO3        o1755(.A(ori_ori_n1804_), .B(ori_ori_n740_), .C(ori_ori_n139_), .Y(ori_ori_n1805_));
  AOI210     o1756(.A0(ori_ori_n916_), .A1(ori_ori_n141_), .B0(ori_ori_n1805_), .Y(ori_ori_n1806_));
  NA4        o1757(.A(ori_ori_n1806_), .B(ori_ori_n1803_), .C(ori_ori_n1799_), .D(ori_ori_n1796_), .Y(ori24));
  NO2        o1758(.A(ori_ori_n239_), .B(x1), .Y(ori_ori_n1808_));
  NA2        o1759(.A(ori_ori_n337_), .B(ori_ori_n492_), .Y(ori_ori_n1809_));
  NAi21      o1760(.An(ori_ori_n1808_), .B(ori_ori_n1809_), .Y(ori_ori_n1810_));
  NO3        o1761(.A(ori_ori_n542_), .B(ori_ori_n684_), .C(ori_ori_n155_), .Y(ori_ori_n1811_));
  AOI210     o1762(.A0(ori_ori_n1810_), .A1(ori_ori_n91_), .B0(ori_ori_n1811_), .Y(ori_ori_n1812_));
  NA2        o1763(.A(ori_ori_n98_), .B(x8), .Y(ori_ori_n1813_));
  NO3        o1764(.A(ori_ori_n1061_), .B(ori_ori_n1334_), .C(ori_ori_n1042_), .Y(ori_ori_n1814_));
  AOI210     o1765(.A0(ori_ori_n979_), .A1(ori_ori_n56_), .B0(ori_ori_n1447_), .Y(ori_ori_n1815_));
  AO220      o1766(.A0(ori_ori_n1815_), .A1(ori_ori_n1814_), .B0(ori_ori_n1267_), .B1(ori_ori_n325_), .Y(ori_ori_n1816_));
  NA2        o1767(.A(ori_ori_n455_), .B(x8), .Y(ori_ori_n1817_));
  NA2        o1768(.A(ori_ori_n666_), .B(ori_ori_n122_), .Y(ori_ori_n1818_));
  OAI220     o1769(.A0(ori_ori_n1818_), .A1(ori_ori_n1432_), .B0(ori_ori_n1817_), .B1(ori_ori_n838_), .Y(ori_ori_n1819_));
  AOI220     o1770(.A0(ori_ori_n1819_), .A1(ori_ori_n1689_), .B0(ori_ori_n1816_), .B1(ori_ori_n1025_), .Y(ori_ori_n1820_));
  OAI210     o1771(.A0(ori_ori_n1813_), .A1(ori_ori_n1812_), .B0(ori_ori_n1820_), .Y(ori25));
  NA2        o1772(.A(ori_ori_n326_), .B(ori_ori_n59_), .Y(ori_ori_n1822_));
  NO2        o1773(.A(ori_ori_n1822_), .B(ori_ori_n317_), .Y(ori_ori_n1823_));
  OAI210     o1774(.A0(ori_ori_n1823_), .A1(ori_ori_n1181_), .B0(ori_ori_n112_), .Y(ori_ori_n1824_));
  INV        o1775(.A(ori_ori_n1275_), .Y(ori_ori_n1825_));
  NO2        o1776(.A(ori_ori_n739_), .B(ori_ori_n55_), .Y(ori_ori_n1826_));
  AOI220     o1777(.A0(ori_ori_n1826_), .A1(ori_ori_n1825_), .B0(ori_ori_n1589_), .B1(ori_ori_n1182_), .Y(ori_ori_n1827_));
  AOI210     o1778(.A0(ori_ori_n1827_), .A1(ori_ori_n1824_), .B0(ori_ori_n679_), .Y(ori_ori_n1828_));
  NO3        o1779(.A(ori_ori_n1035_), .B(ori_ori_n142_), .C(ori_ori_n78_), .Y(ori_ori_n1829_));
  OAI210     o1780(.A0(ori_ori_n195_), .A1(ori_ori_n273_), .B0(ori_ori_n327_), .Y(ori_ori_n1830_));
  OAI210     o1781(.A0(ori_ori_n1830_), .A1(ori_ori_n1829_), .B0(ori_ori_n1180_), .Y(ori_ori_n1831_));
  NO2        o1782(.A(ori_ori_n1385_), .B(ori_ori_n448_), .Y(ori_ori_n1832_));
  NO3        o1783(.A(ori_ori_n1832_), .B(ori_ori_n533_), .C(ori_ori_n95_), .Y(ori_ori_n1833_));
  NA2        o1784(.A(ori_ori_n510_), .B(ori_ori_n55_), .Y(ori_ori_n1834_));
  OAI220     o1785(.A0(ori_ori_n1834_), .A1(ori_ori_n239_), .B0(ori_ori_n587_), .B1(ori_ori_n273_), .Y(ori_ori_n1835_));
  OAI210     o1786(.A0(ori_ori_n1835_), .A1(ori_ori_n1833_), .B0(ori_ori_n634_), .Y(ori_ori_n1836_));
  AOI220     o1787(.A0(ori_ori_n1753_), .A1(ori_ori_n1135_), .B0(ori_ori_n1489_), .B1(ori_ori_n377_), .Y(ori_ori_n1837_));
  NA3        o1788(.A(ori_ori_n1837_), .B(ori_ori_n1836_), .C(ori_ori_n1831_), .Y(ori_ori_n1838_));
  AO210      o1789(.A0(ori_ori_n1838_), .A1(ori_ori_n104_), .B0(ori_ori_n1828_), .Y(ori26));
  NA2        o1790(.A(ori_ori_n768_), .B(ori_ori_n50_), .Y(ori_ori_n1840_));
  OAI220     o1791(.A0(ori_ori_n303_), .A1(ori_ori_n248_), .B0(ori_ori_n1840_), .B1(x7), .Y(ori_ori_n1841_));
  AOI220     o1792(.A0(ori_ori_n1841_), .A1(ori_ori_n91_), .B0(ori_ori_n1295_), .B1(ori_ori_n1141_), .Y(ori_ori_n1842_));
  NA2        o1793(.A(ori_ori_n625_), .B(ori_ori_n580_), .Y(ori_ori_n1843_));
  OAI210     o1794(.A0(ori_ori_n632_), .A1(ori_ori_n625_), .B0(ori_ori_n743_), .Y(ori_ori_n1844_));
  AOI210     o1795(.A0(ori_ori_n1843_), .A1(ori_ori_n1204_), .B0(ori_ori_n1844_), .Y(ori_ori_n1845_));
  NA2        o1796(.A(ori_ori_n1017_), .B(ori_ori_n585_), .Y(ori_ori_n1846_));
  NO2        o1797(.A(ori_ori_n1846_), .B(ori_ori_n1250_), .Y(ori_ori_n1847_));
  AOI210     o1798(.A0(ori_ori_n1774_), .A1(ori_ori_n1455_), .B0(ori_ori_n1847_), .Y(ori_ori_n1848_));
  NO2        o1799(.A(ori_ori_n1082_), .B(ori_ori_n75_), .Y(ori_ori_n1849_));
  NA2        o1800(.A(ori_ori_n807_), .B(ori_ori_n175_), .Y(ori_ori_n1850_));
  NO2        o1801(.A(ori_ori_n1850_), .B(ori_ori_n538_), .Y(ori_ori_n1851_));
  AOI210     o1802(.A0(ori_ori_n1849_), .A1(ori_ori_n586_), .B0(ori_ori_n1851_), .Y(ori_ori_n1852_));
  OAI220     o1803(.A0(ori_ori_n1852_), .A1(ori_ori_n104_), .B0(ori_ori_n1848_), .B1(ori_ori_n53_), .Y(ori_ori_n1853_));
  NA2        o1804(.A(ori_ori_n602_), .B(ori_ori_n510_), .Y(ori_ori_n1854_));
  NO2        o1805(.A(ori_ori_n132_), .B(ori_ori_n129_), .Y(ori_ori_n1855_));
  NA2        o1806(.A(ori_ori_n1855_), .B(ori_ori_n119_), .Y(ori_ori_n1856_));
  NA2        o1807(.A(ori_ori_n743_), .B(x3), .Y(ori_ori_n1857_));
  AOI210     o1808(.A0(ori_ori_n1856_), .A1(ori_ori_n1854_), .B0(ori_ori_n1857_), .Y(ori_ori_n1858_));
  NO2        o1809(.A(ori_ori_n1004_), .B(x3), .Y(ori_ori_n1859_));
  AOI210     o1810(.A0(ori_ori_n446_), .A1(ori_ori_n104_), .B0(ori_ori_n1859_), .Y(ori_ori_n1860_));
  NA3        o1811(.A(ori_ori_n571_), .B(ori_ori_n51_), .C(ori_ori_n56_), .Y(ori_ori_n1861_));
  AOI210     o1812(.A0(ori_ori_n1640_), .A1(ori_ori_n1054_), .B0(x0), .Y(ori_ori_n1862_));
  OAI210     o1813(.A0(ori_ori_n1861_), .A1(ori_ori_n1860_), .B0(ori_ori_n1862_), .Y(ori_ori_n1863_));
  NO4        o1814(.A(ori_ori_n1863_), .B(ori_ori_n1858_), .C(ori_ori_n1853_), .D(ori_ori_n1845_), .Y(ori_ori_n1864_));
  AOI210     o1815(.A0(x8), .A1(x6), .B0(x5), .Y(ori_ori_n1865_));
  AO220      o1816(.A0(ori_ori_n1865_), .A1(ori_ori_n144_), .B0(ori_ori_n593_), .B1(ori_ori_n139_), .Y(ori_ori_n1866_));
  NA2        o1817(.A(ori_ori_n1866_), .B(ori_ori_n447_), .Y(ori_ori_n1867_));
  NO2        o1818(.A(ori_ori_n753_), .B(ori_ori_n144_), .Y(ori_ori_n1868_));
  NA3        o1819(.A(ori_ori_n1868_), .B(ori_ori_n1662_), .C(ori_ori_n133_), .Y(ori_ori_n1869_));
  NO2        o1820(.A(ori_ori_n398_), .B(ori_ori_n1371_), .Y(ori_ori_n1870_));
  OAI210     o1821(.A0(ori_ori_n1870_), .A1(ori_ori_n1340_), .B0(ori_ori_n446_), .Y(ori_ori_n1871_));
  NA3        o1822(.A(ori_ori_n371_), .B(ori_ori_n854_), .C(ori_ori_n252_), .Y(ori_ori_n1872_));
  NA4        o1823(.A(ori_ori_n1872_), .B(ori_ori_n1871_), .C(ori_ori_n1869_), .D(ori_ori_n1867_), .Y(ori_ori_n1873_));
  AOI210     o1824(.A0(ori_ori_n221_), .A1(x2), .B0(ori_ori_n493_), .Y(ori_ori_n1874_));
  NO2        o1825(.A(ori_ori_n1874_), .B(ori_ori_n113_), .Y(ori_ori_n1875_));
  NA3        o1826(.A(ori_ori_n809_), .B(ori_ori_n1004_), .C(x7), .Y(ori_ori_n1876_));
  AOI210     o1827(.A0(ori_ori_n341_), .A1(ori_ori_n213_), .B0(ori_ori_n1876_), .Y(ori_ori_n1877_));
  OAI220     o1828(.A0(ori_ori_n896_), .A1(ori_ori_n303_), .B0(ori_ori_n642_), .B1(ori_ori_n684_), .Y(ori_ori_n1878_));
  NO3        o1829(.A(ori_ori_n1878_), .B(ori_ori_n1877_), .C(ori_ori_n1875_), .Y(ori_ori_n1879_));
  NA3        o1830(.A(ori_ori_n666_), .B(ori_ori_n189_), .C(ori_ori_n948_), .Y(ori_ori_n1880_));
  NA2        o1831(.A(ori_ori_n1880_), .B(ori_ori_n642_), .Y(ori_ori_n1881_));
  NA2        o1832(.A(ori_ori_n139_), .B(ori_ori_n131_), .Y(ori_ori_n1882_));
  OAI210     o1833(.A0(ori_ori_n1882_), .A1(ori_ori_n1419_), .B0(x0), .Y(ori_ori_n1883_));
  AOI210     o1834(.A0(ori_ori_n1881_), .A1(ori_ori_n1408_), .B0(ori_ori_n1883_), .Y(ori_ori_n1884_));
  OAI210     o1835(.A0(ori_ori_n1879_), .A1(ori_ori_n53_), .B0(ori_ori_n1884_), .Y(ori_ori_n1885_));
  AOI210     o1836(.A0(ori_ori_n1873_), .A1(x4), .B0(ori_ori_n1885_), .Y(ori_ori_n1886_));
  OA220      o1837(.A0(ori_ori_n1886_), .A1(ori_ori_n1864_), .B0(ori_ori_n1842_), .B1(ori_ori_n105_), .Y(ori27));
  NA2        o1838(.A(ori_ori_n1145_), .B(ori_ori_n446_), .Y(ori_ori_n1888_));
  NO2        o1839(.A(ori_ori_n1888_), .B(ori_ori_n298_), .Y(ori_ori_n1889_));
  NA2        o1840(.A(ori_ori_n912_), .B(ori_ori_n809_), .Y(ori_ori_n1890_));
  NA3        o1841(.A(ori_ori_n815_), .B(ori_ori_n361_), .C(ori_ori_n1019_), .Y(ori_ori_n1891_));
  AOI210     o1842(.A0(ori_ori_n1891_), .A1(ori_ori_n1890_), .B0(ori_ori_n213_), .Y(ori_ori_n1892_));
  OAI210     o1843(.A0(ori_ori_n1892_), .A1(ori_ori_n1889_), .B0(ori_ori_n698_), .Y(ori_ori_n1893_));
  XO2        o1844(.A(x8), .B(x4), .Y(ori_ori_n1894_));
  NO3        o1845(.A(ori_ori_n1894_), .B(ori_ori_n446_), .C(ori_ori_n169_), .Y(ori_ori_n1895_));
  OA210      o1846(.A0(ori_ori_n1895_), .A1(ori_ori_n1251_), .B0(ori_ori_n276_), .Y(ori_ori_n1896_));
  NO2        o1847(.A(ori_ori_n393_), .B(ori_ori_n164_), .Y(ori_ori_n1897_));
  OAI210     o1848(.A0(ori_ori_n1897_), .A1(ori_ori_n1896_), .B0(ori_ori_n1119_), .Y(ori_ori_n1898_));
  AOI210     o1849(.A0(ori_ori_n632_), .A1(ori_ori_n56_), .B0(ori_ori_n1849_), .Y(ori_ori_n1899_));
  OAI220     o1850(.A0(ori_ori_n1899_), .A1(ori_ori_n1250_), .B0(ori_ori_n1202_), .B1(ori_ori_n204_), .Y(ori_ori_n1900_));
  NA2        o1851(.A(ori_ori_n1900_), .B(ori_ori_n537_), .Y(ori_ori_n1901_));
  NA3        o1852(.A(ori_ori_n1901_), .B(ori_ori_n1898_), .C(ori_ori_n1893_), .Y(ori28));
  NO3        o1853(.A(ori_ori_n1894_), .B(ori_ori_n1380_), .C(ori_ori_n146_), .Y(ori_ori_n1903_));
  OAI210     o1854(.A0(ori_ori_n1903_), .A1(ori_ori_n1268_), .B0(ori_ori_n585_), .Y(ori_ori_n1904_));
  NA3        o1855(.A(ori_ori_n1182_), .B(ori_ori_n890_), .C(x7), .Y(ori_ori_n1905_));
  NA3        o1856(.A(ori_ori_n495_), .B(ori_ori_n78_), .C(ori_ori_n607_), .Y(ori_ori_n1906_));
  NA3        o1857(.A(ori_ori_n1906_), .B(ori_ori_n1905_), .C(ori_ori_n1904_), .Y(ori_ori_n1907_));
  NA2        o1858(.A(ori_ori_n1245_), .B(ori_ori_n444_), .Y(ori_ori_n1908_));
  NA3        o1859(.A(ori_ori_n1908_), .B(ori_ori_n1397_), .C(ori_ori_n411_), .Y(ori_ori_n1909_));
  NO2        o1860(.A(ori_ori_n306_), .B(x4), .Y(ori_ori_n1910_));
  AOI220     o1861(.A0(ori_ori_n1910_), .A1(ori_ori_n1859_), .B0(ori_ori_n1120_), .B1(ori_ori_n674_), .Y(ori_ori_n1911_));
  NA2        o1862(.A(ori_ori_n1911_), .B(ori_ori_n1909_), .Y(ori_ori_n1912_));
  NO2        o1863(.A(ori_ori_n1245_), .B(ori_ori_n1222_), .Y(ori_ori_n1913_));
  NO4        o1864(.A(x6), .B(ori_ori_n56_), .C(x2), .D(x0), .Y(ori_ori_n1914_));
  OAI210     o1865(.A0(ori_ori_n1914_), .A1(ori_ori_n1913_), .B0(ori_ori_n1040_), .Y(ori_ori_n1915_));
  NA2        o1866(.A(ori_ori_n1176_), .B(ori_ori_n104_), .Y(ori_ori_n1916_));
  NA2        o1867(.A(ori_ori_n1078_), .B(ori_ori_n103_), .Y(ori_ori_n1917_));
  OAI210     o1868(.A0(ori_ori_n1917_), .A1(ori_ori_n1916_), .B0(ori_ori_n1915_), .Y(ori_ori_n1918_));
  OAI210     o1869(.A0(ori_ori_n1918_), .A1(ori_ori_n1912_), .B0(x7), .Y(ori_ori_n1919_));
  NO2        o1870(.A(ori_ori_n384_), .B(x7), .Y(ori_ori_n1920_));
  NO3        o1871(.A(ori_ori_n398_), .B(ori_ori_n270_), .C(ori_ori_n120_), .Y(ori_ori_n1921_));
  OAI210     o1872(.A0(ori_ori_n865_), .A1(ori_ori_n257_), .B0(ori_ori_n81_), .Y(ori_ori_n1922_));
  OAI220     o1873(.A0(ori_ori_n1922_), .A1(ori_ori_n1921_), .B0(ori_ori_n1920_), .B1(ori_ori_n107_), .Y(ori_ori_n1923_));
  NA2        o1874(.A(ori_ori_n1783_), .B(ori_ori_n654_), .Y(ori_ori_n1924_));
  NO2        o1875(.A(ori_ori_n1834_), .B(ori_ori_n77_), .Y(ori_ori_n1925_));
  AOI220     o1876(.A0(ori_ori_n1925_), .A1(ori_ori_n1924_), .B0(ori_ori_n477_), .B1(ori_ori_n50_), .Y(ori_ori_n1926_));
  AOI210     o1877(.A0(ori_ori_n1926_), .A1(ori_ori_n1923_), .B0(ori_ori_n59_), .Y(ori_ori_n1927_));
  AOI220     o1878(.A0(ori_ori_n1385_), .A1(ori_ori_n672_), .B0(ori_ori_n410_), .B1(ori_ori_n455_), .Y(ori_ori_n1928_));
  OAI210     o1879(.A0(ori_ori_n1928_), .A1(ori_ori_n142_), .B0(x1), .Y(ori_ori_n1929_));
  NO2        o1880(.A(ori_ori_n1929_), .B(ori_ori_n1927_), .Y(ori_ori_n1930_));
  AOI210     o1881(.A0(ori_ori_n1574_), .A1(ori_ori_n398_), .B0(ori_ori_n664_), .Y(ori_ori_n1931_));
  NO2        o1882(.A(ori_ori_n398_), .B(x5), .Y(ori_ori_n1932_));
  NO2        o1883(.A(ori_ori_n1932_), .B(ori_ori_n225_), .Y(ori_ori_n1933_));
  NO2        o1884(.A(ori_ori_n1933_), .B(ori_ori_n1931_), .Y(ori_ori_n1934_));
  NOi21      o1885(.An(ori_ori_n703_), .B(ori_ori_n994_), .Y(ori_ori_n1935_));
  NA3        o1886(.A(ori_ori_n1935_), .B(ori_ori_n1078_), .C(ori_ori_n865_), .Y(ori_ori_n1936_));
  OAI210     o1887(.A0(ori_ori_n1352_), .A1(ori_ori_n1668_), .B0(ori_ori_n1936_), .Y(ori_ori_n1937_));
  OAI210     o1888(.A0(ori_ori_n1937_), .A1(ori_ori_n1934_), .B0(ori_ori_n1119_), .Y(ori_ori_n1938_));
  OAI210     o1889(.A0(ori_ori_n444_), .A1(ori_ori_n51_), .B0(ori_ori_n1013_), .Y(ori_ori_n1939_));
  AOI220     o1890(.A0(ori_ori_n1939_), .A1(ori_ori_n461_), .B0(ori_ori_n444_), .B1(ori_ori_n385_), .Y(ori_ori_n1940_));
  NO2        o1891(.A(ori_ori_n1940_), .B(ori_ori_n153_), .Y(ori_ori_n1941_));
  NA2        o1892(.A(ori_ori_n162_), .B(ori_ori_n71_), .Y(ori_ori_n1942_));
  OAI210     o1893(.A0(ori_ori_n1846_), .A1(ori_ori_n1942_), .B0(ori_ori_n53_), .Y(ori_ori_n1943_));
  OAI220     o1894(.A0(ori_ori_n685_), .A1(ori_ori_n260_), .B0(ori_ori_n681_), .B1(x6), .Y(ori_ori_n1944_));
  NO2        o1895(.A(ori_ori_n301_), .B(x4), .Y(ori_ori_n1945_));
  AOI220     o1896(.A0(ori_ori_n1945_), .A1(ori_ori_n361_), .B0(ori_ori_n1944_), .B1(x4), .Y(ori_ori_n1946_));
  NO3        o1897(.A(ori_ori_n1946_), .B(ori_ori_n320_), .C(x5), .Y(ori_ori_n1947_));
  NO2        o1898(.A(ori_ori_n703_), .B(ori_ori_n57_), .Y(ori_ori_n1948_));
  NA2        o1899(.A(ori_ori_n1948_), .B(ori_ori_n446_), .Y(ori_ori_n1949_));
  AOI220     o1900(.A0(ori_ori_n662_), .A1(ori_ori_n729_), .B0(ori_ori_n493_), .B1(ori_ori_n235_), .Y(ori_ori_n1950_));
  AOI210     o1901(.A0(ori_ori_n1950_), .A1(ori_ori_n1949_), .B0(ori_ori_n255_), .Y(ori_ori_n1951_));
  NO4        o1902(.A(ori_ori_n1951_), .B(ori_ori_n1947_), .C(ori_ori_n1943_), .D(ori_ori_n1941_), .Y(ori_ori_n1952_));
  AOI220     o1903(.A0(ori_ori_n1952_), .A1(ori_ori_n1938_), .B0(ori_ori_n1930_), .B1(ori_ori_n1919_), .Y(ori_ori_n1953_));
  AOI210     o1904(.A0(ori_ori_n1907_), .A1(x3), .B0(ori_ori_n1953_), .Y(ori29));
  OAI210     o1905(.A0(ori_ori_n556_), .A1(ori_ori_n261_), .B0(ori_ori_n724_), .Y(ori_ori_n1955_));
  NA2        o1906(.A(ori_ori_n745_), .B(ori_ori_n1040_), .Y(ori_ori_n1956_));
  AO210      o1907(.A0(ori_ori_n1158_), .A1(ori_ori_n1166_), .B0(ori_ori_n1956_), .Y(ori_ori_n1957_));
  AOI210     o1908(.A0(ori_ori_n180_), .A1(ori_ori_n166_), .B0(ori_ori_n703_), .Y(ori_ori_n1958_));
  INV        o1909(.A(ori_ori_n1958_), .Y(ori_ori_n1959_));
  NA3        o1910(.A(ori_ori_n1959_), .B(ori_ori_n1957_), .C(ori_ori_n1955_), .Y(ori_ori_n1960_));
  NO3        o1911(.A(ori_ori_n664_), .B(ori_ori_n1141_), .C(ori_ori_n50_), .Y(ori_ori_n1961_));
  NO3        o1912(.A(ori_ori_n1961_), .B(ori_ori_n1244_), .C(ori_ori_n556_), .Y(ori_ori_n1962_));
  NO2        o1913(.A(ori_ori_n442_), .B(ori_ori_n58_), .Y(ori_ori_n1963_));
  AOI220     o1914(.A0(ori_ori_n1963_), .A1(ori_ori_n1204_), .B0(ori_ori_n669_), .B1(ori_ori_n1370_), .Y(ori_ori_n1964_));
  OAI210     o1915(.A0(ori_ori_n1962_), .A1(ori_ori_n542_), .B0(ori_ori_n1964_), .Y(ori_ori_n1965_));
  AOI210     o1916(.A0(ori_ori_n1960_), .A1(x6), .B0(ori_ori_n1965_), .Y(ori_ori_n1966_));
  OAI210     o1917(.A0(x8), .A1(x4), .B0(x5), .Y(ori_ori_n1967_));
  NA2        o1918(.A(ori_ori_n1967_), .B(ori_ori_n108_), .Y(ori_ori_n1968_));
  NA2        o1919(.A(ori_ori_n301_), .B(ori_ori_n146_), .Y(ori_ori_n1969_));
  NA4        o1920(.A(ori_ori_n1969_), .B(ori_ori_n1968_), .C(ori_ori_n663_), .D(ori_ori_n64_), .Y(ori_ori_n1970_));
  AOI210     o1921(.A0(ori_ori_n1312_), .A1(ori_ori_n270_), .B0(ori_ori_n1719_), .Y(ori_ori_n1971_));
  AOI210     o1922(.A0(ori_ori_n1971_), .A1(ori_ori_n1970_), .B0(ori_ori_n883_), .Y(ori_ori_n1972_));
  NA4        o1923(.A(ori_ori_n664_), .B(ori_ori_n306_), .C(ori_ori_n180_), .D(ori_ori_n166_), .Y(ori_ori_n1973_));
  NA3        o1924(.A(ori_ori_n630_), .B(ori_ori_n294_), .C(ori_ori_n797_), .Y(ori_ori_n1974_));
  AOI210     o1925(.A0(ori_ori_n1974_), .A1(ori_ori_n1973_), .B0(ori_ori_n1204_), .Y(ori_ori_n1975_));
  OAI210     o1926(.A0(ori_ori_n890_), .A1(x8), .B0(x7), .Y(ori_ori_n1976_));
  NO2        o1927(.A(ori_ori_n1976_), .B(ori_ori_n125_), .Y(ori_ori_n1977_));
  OA210      o1928(.A0(ori_ori_n865_), .A1(ori_ori_n273_), .B0(ori_ori_n1967_), .Y(ori_ori_n1978_));
  OAI220     o1929(.A0(ori_ori_n1978_), .A1(ori_ori_n587_), .B0(ori_ori_n1497_), .B1(ori_ori_n393_), .Y(ori_ori_n1979_));
  NO4        o1930(.A(ori_ori_n1979_), .B(ori_ori_n1977_), .C(ori_ori_n1975_), .D(ori_ori_n1972_), .Y(ori_ori_n1980_));
  OAI210     o1931(.A0(ori_ori_n1966_), .A1(x2), .B0(ori_ori_n1980_), .Y(ori_ori_n1981_));
  NA3        o1932(.A(x6), .B(ori_ori_n50_), .C(x2), .Y(ori_ori_n1982_));
  OAI210     o1933(.A0(ori_ori_n1222_), .A1(ori_ori_n351_), .B0(ori_ori_n1982_), .Y(ori_ori_n1983_));
  NO3        o1934(.A(ori_ori_n444_), .B(x3), .C(x0), .Y(ori_ori_n1984_));
  AO220      o1935(.A0(ori_ori_n1984_), .A1(x5), .B0(ori_ori_n1914_), .B1(ori_ori_n81_), .Y(ori_ori_n1985_));
  AOI210     o1936(.A0(ori_ori_n1983_), .A1(ori_ori_n341_), .B0(ori_ori_n1985_), .Y(ori_ori_n1986_));
  NO3        o1937(.A(ori_ori_n696_), .B(ori_ori_n362_), .C(ori_ori_n140_), .Y(ori_ori_n1987_));
  AOI210     o1938(.A0(ori_ori_n723_), .A1(ori_ori_n614_), .B0(ori_ori_n1987_), .Y(ori_ori_n1988_));
  OAI210     o1939(.A0(ori_ori_n1986_), .A1(x7), .B0(ori_ori_n1988_), .Y(ori_ori_n1989_));
  AOI210     o1940(.A0(ori_ori_n1088_), .A1(ori_ori_n398_), .B0(ori_ori_n1396_), .Y(ori_ori_n1990_));
  NO2        o1941(.A(ori_ori_n146_), .B(x2), .Y(ori_ori_n1991_));
  OA210      o1942(.A0(ori_ori_n1991_), .A1(ori_ori_n629_), .B0(ori_ori_n664_), .Y(ori_ori_n1992_));
  OAI210     o1943(.A0(ori_ori_n1992_), .A1(ori_ori_n1990_), .B0(ori_ori_n68_), .Y(ori_ori_n1993_));
  NO2        o1944(.A(ori_ori_n195_), .B(ori_ori_n85_), .Y(ori_ori_n1994_));
  OAI210     o1945(.A0(ori_ori_n1994_), .A1(ori_ori_n783_), .B0(ori_ori_n1097_), .Y(ori_ori_n1995_));
  NA3        o1946(.A(ori_ori_n1932_), .B(ori_ori_n228_), .C(ori_ori_n83_), .Y(ori_ori_n1996_));
  NA3        o1947(.A(ori_ori_n1996_), .B(ori_ori_n1995_), .C(ori_ori_n1993_), .Y(ori_ori_n1997_));
  AOI210     o1948(.A0(ori_ori_n1989_), .A1(x8), .B0(ori_ori_n1997_), .Y(ori_ori_n1998_));
  OAI210     o1949(.A0(ori_ori_n442_), .A1(ori_ori_n244_), .B0(ori_ori_n957_), .Y(ori_ori_n1999_));
  OAI210     o1950(.A0(ori_ori_n1999_), .A1(ori_ori_n1120_), .B0(ori_ori_n674_), .Y(ori_ori_n2000_));
  NO3        o1951(.A(ori_ori_n1017_), .B(ori_ori_n352_), .C(ori_ori_n147_), .Y(ori_ori_n2001_));
  NA3        o1952(.A(ori_ori_n2001_), .B(ori_ori_n1294_), .C(ori_ori_n50_), .Y(ori_ori_n2002_));
  NO2        o1953(.A(ori_ori_n133_), .B(ori_ori_n91_), .Y(ori_ori_n2003_));
  AOI220     o1954(.A0(ori_ori_n2003_), .A1(ori_ori_n588_), .B0(ori_ori_n1913_), .B1(ori_ori_n358_), .Y(ori_ori_n2004_));
  NOi31      o1955(.An(ori_ori_n1121_), .B(ori_ori_n1865_), .C(ori_ori_n624_), .Y(ori_ori_n2005_));
  NA2        o1956(.A(ori_ori_n171_), .B(x4), .Y(ori_ori_n2006_));
  NO3        o1957(.A(ori_ori_n1471_), .B(ori_ori_n239_), .C(ori_ori_n71_), .Y(ori_ori_n2007_));
  AOI210     o1958(.A0(ori_ori_n2007_), .A1(ori_ori_n2006_), .B0(ori_ori_n2005_), .Y(ori_ori_n2008_));
  NA4        o1959(.A(ori_ori_n2008_), .B(ori_ori_n2004_), .C(ori_ori_n2002_), .D(ori_ori_n2000_), .Y(ori_ori_n2009_));
  NO4        o1960(.A(ori_ori_n1222_), .B(ori_ori_n169_), .C(ori_ori_n55_), .D(ori_ori_n71_), .Y(ori_ori_n2010_));
  NO4        o1961(.A(ori_ori_n1197_), .B(ori_ori_n502_), .C(ori_ori_n1370_), .D(ori_ori_n104_), .Y(ori_ori_n2011_));
  OAI210     o1962(.A0(ori_ori_n2011_), .A1(ori_ori_n2010_), .B0(ori_ori_n106_), .Y(ori_ori_n2012_));
  AOI210     o1963(.A0(ori_ori_n305_), .A1(x4), .B0(ori_ori_n189_), .Y(ori_ori_n2013_));
  OAI210     o1964(.A0(ori_ori_n2013_), .A1(ori_ori_n1963_), .B0(ori_ori_n720_), .Y(ori_ori_n2014_));
  OR3        o1965(.A(ori_ori_n1740_), .B(ori_ori_n1422_), .C(ori_ori_n1080_), .Y(ori_ori_n2015_));
  NA2        o1966(.A(ori_ori_n1914_), .B(ori_ori_n804_), .Y(ori_ori_n2016_));
  OR2        o1967(.A(ori_ori_n2016_), .B(ori_ori_n244_), .Y(ori_ori_n2017_));
  NA4        o1968(.A(ori_ori_n2017_), .B(ori_ori_n2015_), .C(ori_ori_n2014_), .D(ori_ori_n2012_), .Y(ori_ori_n2018_));
  AOI210     o1969(.A0(ori_ori_n2009_), .A1(ori_ori_n290_), .B0(ori_ori_n2018_), .Y(ori_ori_n2019_));
  OAI210     o1970(.A0(ori_ori_n1998_), .A1(x1), .B0(ori_ori_n2019_), .Y(ori_ori_n2020_));
  AO210      o1971(.A0(ori_ori_n1981_), .A1(x1), .B0(ori_ori_n2020_), .Y(ori30));
  NO3        o1972(.A(ori_ori_n1766_), .B(ori_ori_n577_), .C(ori_ori_n95_), .Y(ori_ori_n2022_));
  NO3        o1973(.A(ori_ori_n1139_), .B(ori_ori_n136_), .C(ori_ori_n381_), .Y(ori_ori_n2023_));
  AOI210     o1974(.A0(ori_ori_n720_), .A1(ori_ori_n252_), .B0(ori_ori_n2023_), .Y(ori_ori_n2024_));
  AOI210     o1975(.A0(ori_ori_n2024_), .A1(ori_ori_n2022_), .B0(ori_ori_n56_), .Y(ori_ori_n2025_));
  NA2        o1976(.A(ori_ori_n809_), .B(ori_ori_n339_), .Y(ori_ori_n2026_));
  NA2        o1977(.A(ori_ori_n2026_), .B(ori_ori_n1353_), .Y(ori_ori_n2027_));
  OAI210     o1978(.A0(ori_ori_n2027_), .A1(ori_ori_n2025_), .B0(ori_ori_n106_), .Y(ori_ori_n2028_));
  OAI210     o1979(.A0(ori_ori_n994_), .A1(ori_ori_n571_), .B0(ori_ori_n674_), .Y(ori_ori_n2029_));
  AOI220     o1980(.A0(ori_ori_n447_), .A1(ori_ori_n936_), .B0(ori_ori_n325_), .B1(ori_ori_n455_), .Y(ori_ori_n2030_));
  AOI210     o1981(.A0(ori_ori_n2030_), .A1(ori_ori_n2029_), .B0(ori_ori_n255_), .Y(ori_ori_n2031_));
  NO3        o1982(.A(ori_ori_n279_), .B(ori_ori_n121_), .C(x0), .Y(ori_ori_n2032_));
  AOI210     o1983(.A0(ori_ori_n504_), .A1(x6), .B0(ori_ori_n2032_), .Y(ori_ori_n2033_));
  AOI220     o1984(.A0(ori_ori_n1135_), .A1(ori_ori_n422_), .B0(ori_ori_n757_), .B1(ori_ori_n90_), .Y(ori_ori_n2034_));
  OAI220     o1985(.A0(ori_ori_n2034_), .A1(ori_ori_n244_), .B0(ori_ori_n2033_), .B1(ori_ori_n54_), .Y(ori_ori_n2035_));
  NA3        o1986(.A(ori_ori_n321_), .B(ori_ori_n163_), .C(ori_ori_n71_), .Y(ori_ori_n2036_));
  AO210      o1987(.A0(ori_ori_n570_), .A1(ori_ori_n518_), .B0(x5), .Y(ori_ori_n2037_));
  AOI210     o1988(.A0(ori_ori_n2036_), .A1(ori_ori_n718_), .B0(ori_ori_n2037_), .Y(ori_ori_n2038_));
  AOI210     o1989(.A0(ori_ori_n1595_), .A1(ori_ori_n50_), .B0(ori_ori_n455_), .Y(ori_ori_n2039_));
  NA2        o1990(.A(ori_ori_n194_), .B(x2), .Y(ori_ori_n2040_));
  OA220      o1991(.A0(ori_ori_n2040_), .A1(ori_ori_n2039_), .B0(ori_ori_n274_), .B1(x6), .Y(ori_ori_n2041_));
  OAI210     o1992(.A0(x7), .A1(x6), .B0(x1), .Y(ori_ori_n2042_));
  NA3        o1993(.A(ori_ori_n57_), .B(x4), .C(ori_ori_n59_), .Y(ori_ori_n2043_));
  AOI220     o1994(.A0(ori_ori_n2043_), .A1(ori_ori_n1360_), .B0(ori_ori_n2042_), .B1(ori_ori_n1804_), .Y(ori_ori_n2044_));
  NO3        o1995(.A(ori_ori_n1356_), .B(ori_ori_n341_), .C(ori_ori_n1019_), .Y(ori_ori_n2045_));
  NO2        o1996(.A(ori_ori_n516_), .B(ori_ori_n858_), .Y(ori_ori_n2046_));
  NOi21      o1997(.An(ori_ori_n2046_), .B(ori_ori_n843_), .Y(ori_ori_n2047_));
  NO3        o1998(.A(ori_ori_n1294_), .B(ori_ori_n230_), .C(ori_ori_n646_), .Y(ori_ori_n2048_));
  NO4        o1999(.A(ori_ori_n2048_), .B(ori_ori_n2047_), .C(ori_ori_n2045_), .D(ori_ori_n2044_), .Y(ori_ori_n2049_));
  OAI210     o2000(.A0(ori_ori_n2041_), .A1(ori_ori_n752_), .B0(ori_ori_n2049_), .Y(ori_ori_n2050_));
  NO4        o2001(.A(ori_ori_n2050_), .B(ori_ori_n2038_), .C(ori_ori_n2035_), .D(ori_ori_n2031_), .Y(ori_ori_n2051_));
  AOI210     o2002(.A0(ori_ori_n2051_), .A1(ori_ori_n2028_), .B0(x8), .Y(ori_ori_n2052_));
  NO3        o2003(.A(ori_ori_n491_), .B(ori_ori_n780_), .C(ori_ori_n53_), .Y(ori_ori_n2053_));
  OAI220     o2004(.A0(ori_ori_n1781_), .A1(ori_ori_n341_), .B0(ori_ori_n483_), .B1(ori_ori_n584_), .Y(ori_ori_n2054_));
  OAI210     o2005(.A0(ori_ori_n2054_), .A1(ori_ori_n2053_), .B0(x6), .Y(ori_ori_n2055_));
  OAI210     o2006(.A0(ori_ori_n1031_), .A1(ori_ori_n537_), .B0(ori_ori_n809_), .Y(ori_ori_n2056_));
  OAI210     o2007(.A0(ori_ori_n1729_), .A1(ori_ori_n328_), .B0(ori_ori_n124_), .Y(ori_ori_n2057_));
  AOI210     o2008(.A0(ori_ori_n376_), .A1(ori_ori_n227_), .B0(ori_ori_n72_), .Y(ori_ori_n2058_));
  AOI210     o2009(.A0(ori_ori_n994_), .A1(ori_ori_n743_), .B0(ori_ori_n2058_), .Y(ori_ori_n2059_));
  NA4        o2010(.A(ori_ori_n2059_), .B(ori_ori_n2057_), .C(ori_ori_n2056_), .D(ori_ori_n2055_), .Y(ori_ori_n2060_));
  NA2        o2011(.A(ori_ori_n1085_), .B(ori_ori_n59_), .Y(ori_ori_n2061_));
  AOI210     o2012(.A0(ori_ori_n917_), .A1(ori_ori_n492_), .B0(ori_ori_n680_), .Y(ori_ori_n2062_));
  OAI220     o2013(.A0(ori_ori_n2062_), .A1(ori_ori_n305_), .B0(ori_ori_n2061_), .B1(ori_ori_n482_), .Y(ori_ori_n2063_));
  AOI210     o2014(.A0(ori_ori_n2060_), .A1(x8), .B0(ori_ori_n2063_), .Y(ori_ori_n2064_));
  NO2        o2015(.A(ori_ori_n2064_), .B(ori_ori_n57_), .Y(ori_ori_n2065_));
  NO2        o2016(.A(ori_ori_n916_), .B(ori_ori_n660_), .Y(ori_ori_n2066_));
  NO2        o2017(.A(ori_ori_n2066_), .B(ori_ori_n444_), .Y(ori_ori_n2067_));
  NO3        o2018(.A(ori_ori_n634_), .B(ori_ori_n407_), .C(ori_ori_n1139_), .Y(ori_ori_n2068_));
  NO3        o2019(.A(ori_ori_n2068_), .B(ori_ori_n1250_), .C(ori_ori_n1370_), .Y(ori_ori_n2069_));
  AOI210     o2020(.A0(ori_ori_n302_), .A1(x1), .B0(ori_ori_n147_), .Y(ori_ori_n2070_));
  NO2        o2021(.A(ori_ori_n308_), .B(x5), .Y(ori_ori_n2071_));
  NO2        o2022(.A(ori_ori_n2071_), .B(ori_ori_n851_), .Y(ori_ori_n2072_));
  OAI220     o2023(.A0(ori_ori_n2072_), .A1(ori_ori_n1051_), .B0(ori_ori_n2070_), .B1(ori_ori_n204_), .Y(ori_ori_n2073_));
  NO3        o2024(.A(ori_ori_n2073_), .B(ori_ori_n2069_), .C(ori_ori_n2067_), .Y(ori_ori_n2074_));
  NA2        o2025(.A(ori_ori_n955_), .B(ori_ori_n82_), .Y(ori_ori_n2075_));
  AO210      o2026(.A0(ori_ori_n2075_), .A1(ori_ori_n1596_), .B0(x3), .Y(ori_ori_n2076_));
  NO2        o2027(.A(ori_ori_n216_), .B(ori_ori_n56_), .Y(ori_ori_n2077_));
  OAI220     o2028(.A0(ori_ori_n376_), .A1(ori_ori_n1250_), .B0(ori_ori_n352_), .B1(ori_ori_n230_), .Y(ori_ori_n2078_));
  AOI220     o2029(.A0(ori_ori_n2078_), .A1(x2), .B0(ori_ori_n2077_), .B1(ori_ori_n1610_), .Y(ori_ori_n2079_));
  AOI210     o2030(.A0(ori_ori_n2079_), .A1(ori_ori_n2076_), .B0(ori_ori_n260_), .Y(ori_ori_n2080_));
  NO2        o2031(.A(ori_ori_n302_), .B(ori_ori_n120_), .Y(ori_ori_n2081_));
  NO3        o2032(.A(ori_ori_n814_), .B(ori_ori_n697_), .C(ori_ori_n166_), .Y(ori_ori_n2082_));
  OAI210     o2033(.A0(ori_ori_n2082_), .A1(ori_ori_n2081_), .B0(ori_ori_n154_), .Y(ori_ori_n2083_));
  NA3        o2034(.A(x5), .B(x4), .C(ori_ori_n59_), .Y(ori_ori_n2084_));
  AOI210     o2035(.A0(ori_ori_n2084_), .A1(ori_ori_n1300_), .B0(ori_ori_n538_), .Y(ori_ori_n2085_));
  AOI210     o2036(.A0(ori_ori_n1320_), .A1(x2), .B0(ori_ori_n2085_), .Y(ori_ori_n2086_));
  AOI210     o2037(.A0(ori_ori_n2086_), .A1(ori_ori_n2083_), .B0(ori_ori_n50_), .Y(ori_ori_n2087_));
  NA3        o2038(.A(ori_ori_n1468_), .B(ori_ori_n1130_), .C(ori_ori_n475_), .Y(ori_ori_n2088_));
  AOI210     o2039(.A0(ori_ori_n2088_), .A1(ori_ori_n2075_), .B0(ori_ori_n610_), .Y(ori_ori_n2089_));
  AOI210     o2040(.A0(ori_ori_n1019_), .A1(x1), .B0(ori_ori_n1312_), .Y(ori_ori_n2090_));
  OAI220     o2041(.A0(ori_ori_n306_), .A1(x4), .B0(ori_ori_n51_), .B1(x6), .Y(ori_ori_n2091_));
  NO2        o2042(.A(ori_ori_n119_), .B(ori_ori_n108_), .Y(ori_ori_n2092_));
  AOI220     o2043(.A0(ori_ori_n2092_), .A1(ori_ori_n2091_), .B0(ori_ori_n1160_), .B1(ori_ori_n624_), .Y(ori_ori_n2093_));
  OAI210     o2044(.A0(ori_ori_n2090_), .A1(ori_ori_n486_), .B0(ori_ori_n2093_), .Y(ori_ori_n2094_));
  NO4        o2045(.A(ori_ori_n2094_), .B(ori_ori_n2089_), .C(ori_ori_n2087_), .D(ori_ori_n2080_), .Y(ori_ori_n2095_));
  OAI210     o2046(.A0(ori_ori_n2074_), .A1(ori_ori_n133_), .B0(ori_ori_n2095_), .Y(ori_ori_n2096_));
  NO3        o2047(.A(ori_ori_n2096_), .B(ori_ori_n2065_), .C(ori_ori_n2052_), .Y(ori31));
  NA2        o2048(.A(ori_ori_n979_), .B(ori_ori_n353_), .Y(ori_ori_n2098_));
  NO2        o2049(.A(ori_ori_n448_), .B(ori_ori_n674_), .Y(ori_ori_n2099_));
  AOI210     o2050(.A0(ori_ori_n2099_), .A1(ori_ori_n2098_), .B0(ori_ori_n58_), .Y(ori_ori_n2100_));
  NO2        o2051(.A(ori_ori_n782_), .B(ori_ori_n56_), .Y(ori_ori_n2101_));
  AOI220     o2052(.A0(ori_ori_n2101_), .A1(x2), .B0(ori_ori_n89_), .B1(x0), .Y(ori_ori_n2102_));
  NA3        o2053(.A(ori_ori_n2102_), .B(ori_ori_n2016_), .C(ori_ori_n1843_), .Y(ori_ori_n2103_));
  OAI210     o2054(.A0(ori_ori_n2103_), .A1(ori_ori_n2100_), .B0(ori_ori_n53_), .Y(ori_ori_n2104_));
  NO2        o2055(.A(ori_ori_n430_), .B(ori_ori_n674_), .Y(ori_ori_n2105_));
  NO3        o2056(.A(ori_ori_n1945_), .B(ori_ori_n1914_), .C(ori_ori_n884_), .Y(ori_ori_n2106_));
  OA220      o2057(.A0(ori_ori_n2106_), .A1(ori_ori_n475_), .B0(ori_ori_n2105_), .B1(ori_ori_n1461_), .Y(ori_ori_n2107_));
  AOI210     o2058(.A0(ori_ori_n2107_), .A1(ori_ori_n2104_), .B0(ori_ori_n104_), .Y(ori_ori_n2108_));
  NO2        o2059(.A(ori_ori_n498_), .B(ori_ori_n75_), .Y(ori_ori_n2109_));
  NA2        o2060(.A(ori_ori_n444_), .B(ori_ori_n57_), .Y(ori_ori_n2110_));
  AOI210     o2061(.A0(ori_ori_n305_), .A1(ori_ori_n86_), .B0(ori_ori_n2110_), .Y(ori_ori_n2111_));
  OAI210     o2062(.A0(ori_ori_n2111_), .A1(ori_ori_n2109_), .B0(ori_ori_n768_), .Y(ori_ori_n2112_));
  NO4        o2063(.A(ori_ori_n1156_), .B(ori_ori_n362_), .C(ori_ori_n1595_), .D(ori_ori_n67_), .Y(ori_ori_n2113_));
  AOI210     o2064(.A0(ori_ori_n1635_), .A1(ori_ori_n1347_), .B0(ori_ori_n442_), .Y(ori_ori_n2114_));
  NO2        o2065(.A(ori_ori_n1301_), .B(ori_ori_n949_), .Y(ori_ori_n2115_));
  NO3        o2066(.A(ori_ori_n2115_), .B(ori_ori_n2114_), .C(ori_ori_n2113_), .Y(ori_ori_n2116_));
  AOI210     o2067(.A0(ori_ori_n2116_), .A1(ori_ori_n2112_), .B0(x5), .Y(ori_ori_n2117_));
  AOI220     o2068(.A0(ori_ori_n446_), .A1(ori_ori_n624_), .B0(ori_ori_n571_), .B1(ori_ori_n63_), .Y(ori_ori_n2118_));
  AOI210     o2069(.A0(ori_ori_n2118_), .A1(ori_ori_n581_), .B0(ori_ori_n1222_), .Y(ori_ori_n2119_));
  AOI220     o2070(.A0(ori_ori_n956_), .A1(ori_ori_n729_), .B0(ori_ori_n1139_), .B1(ori_ori_n118_), .Y(ori_ori_n2120_));
  OAI220     o2071(.A0(ori_ori_n2120_), .A1(ori_ori_n384_), .B0(ori_ori_n482_), .B1(ori_ori_n769_), .Y(ori_ori_n2121_));
  NO4        o2072(.A(ori_ori_n2121_), .B(ori_ori_n2119_), .C(ori_ori_n2117_), .D(ori_ori_n2108_), .Y(ori_ori_n2122_));
  NA2        o2073(.A(ori_ori_n492_), .B(ori_ori_n59_), .Y(ori_ori_n2123_));
  AOI210     o2074(.A0(ori_ori_n542_), .A1(ori_ori_n2123_), .B0(ori_ori_n139_), .Y(ori_ori_n2124_));
  OAI210     o2075(.A0(ori_ori_n100_), .A1(ori_ori_n273_), .B0(ori_ori_n2061_), .Y(ori_ori_n2125_));
  OAI210     o2076(.A0(ori_ori_n2125_), .A1(ori_ori_n2124_), .B0(x7), .Y(ori_ori_n2126_));
  NO3        o2077(.A(ori_ori_n376_), .B(ori_ori_n55_), .C(x7), .Y(ori_ori_n2127_));
  OA210      o2078(.A0(ori_ori_n2127_), .A1(ori_ori_n1311_), .B0(ori_ori_n97_), .Y(ori_ori_n2128_));
  NA2        o2079(.A(ori_ori_n1082_), .B(ori_ori_n90_), .Y(ori_ori_n2129_));
  AOI210     o2080(.A0(ori_ori_n896_), .A1(ori_ori_n108_), .B0(ori_ori_n2129_), .Y(ori_ori_n2130_));
  NA2        o2081(.A(ori_ori_n1542_), .B(x6), .Y(ori_ori_n2131_));
  AOI210     o2082(.A0(ori_ori_n2131_), .A1(ori_ori_n289_), .B0(ori_ori_n104_), .Y(ori_ori_n2132_));
  NA2        o2083(.A(ori_ori_n1182_), .B(ori_ori_n316_), .Y(ori_ori_n2133_));
  AOI210     o2084(.A0(ori_ori_n2133_), .A1(ori_ori_n642_), .B0(ori_ori_n53_), .Y(ori_ori_n2134_));
  NO4        o2085(.A(ori_ori_n2134_), .B(ori_ori_n2132_), .C(ori_ori_n2130_), .D(ori_ori_n2128_), .Y(ori_ori_n2135_));
  AOI210     o2086(.A0(ori_ori_n2135_), .A1(ori_ori_n2126_), .B0(ori_ori_n684_), .Y(ori_ori_n2136_));
  NOi21      o2087(.An(ori_ori_n1756_), .B(ori_ori_n1055_), .Y(ori_ori_n2137_));
  OAI220     o2088(.A0(ori_ori_n2137_), .A1(ori_ori_n1916_), .B0(ori_ori_n918_), .B1(ori_ori_n2123_), .Y(ori_ori_n2138_));
  NA2        o2089(.A(ori_ori_n2138_), .B(x3), .Y(ori_ori_n2139_));
  AOI220     o2090(.A0(ori_ori_n1380_), .A1(x8), .B0(ori_ori_n60_), .B1(x1), .Y(ori_ori_n2140_));
  NO3        o2091(.A(ori_ori_n2140_), .B(ori_ori_n1109_), .C(x6), .Y(ori_ori_n2141_));
  NA2        o2092(.A(ori_ori_n614_), .B(ori_ori_n407_), .Y(ori_ori_n2142_));
  NA2        o2093(.A(ori_ori_n114_), .B(ori_ori_n529_), .Y(ori_ori_n2143_));
  OAI220     o2094(.A0(ori_ori_n2143_), .A1(ori_ori_n1916_), .B0(ori_ori_n2142_), .B1(x4), .Y(ori_ori_n2144_));
  NO2        o2095(.A(ori_ori_n2144_), .B(ori_ori_n2141_), .Y(ori_ori_n2145_));
  AOI210     o2096(.A0(ori_ori_n2145_), .A1(ori_ori_n2139_), .B0(ori_ori_n182_), .Y(ori_ori_n2146_));
  NO4        o2097(.A(ori_ori_n615_), .B(ori_ori_n588_), .C(ori_ori_n698_), .D(ori_ori_n697_), .Y(ori_ori_n2147_));
  OAI210     o2098(.A0(ori_ori_n2147_), .A1(ori_ori_n1073_), .B0(x3), .Y(ori_ori_n2148_));
  NO4        o2099(.A(ori_ori_n800_), .B(ori_ori_n1222_), .C(ori_ori_n768_), .D(x5), .Y(ori_ori_n2149_));
  NO3        o2100(.A(x6), .B(ori_ori_n56_), .C(x1), .Y(ori_ori_n2150_));
  NA2        o2101(.A(ori_ori_n2150_), .B(ori_ori_n285_), .Y(ori_ori_n2151_));
  OAI210     o2102(.A0(ori_ori_n1888_), .A1(ori_ori_n376_), .B0(ori_ori_n2151_), .Y(ori_ori_n2152_));
  NA4        o2103(.A(ori_ori_n634_), .B(ori_ori_n176_), .C(x6), .D(ori_ori_n104_), .Y(ori_ori_n2153_));
  NO2        o2104(.A(ori_ori_n852_), .B(ori_ori_n248_), .Y(ori_ori_n2154_));
  NOi41      o2105(.An(ori_ori_n2153_), .B(ori_ori_n2154_), .C(ori_ori_n2152_), .D(ori_ori_n2149_), .Y(ori_ori_n2155_));
  AOI210     o2106(.A0(ori_ori_n2155_), .A1(ori_ori_n2148_), .B0(ori_ori_n533_), .Y(ori_ori_n2156_));
  OAI210     o2107(.A0(ori_ori_n614_), .A1(ori_ori_n469_), .B0(ori_ori_n936_), .Y(ori_ori_n2157_));
  NO3        o2108(.A(ori_ori_n371_), .B(ori_ori_n77_), .C(ori_ori_n53_), .Y(ori_ori_n2158_));
  NO3        o2109(.A(ori_ori_n461_), .B(ori_ori_n347_), .C(ori_ori_n50_), .Y(ori_ori_n2159_));
  OAI210     o2110(.A0(ori_ori_n2159_), .A1(ori_ori_n2158_), .B0(ori_ori_n1157_), .Y(ori_ori_n2160_));
  AOI210     o2111(.A0(ori_ori_n2160_), .A1(ori_ori_n2157_), .B0(ori_ori_n391_), .Y(ori_ori_n2161_));
  NO2        o2112(.A(ori_ori_n213_), .B(ori_ori_n538_), .Y(ori_ori_n2162_));
  OAI210     o2113(.A0(ori_ori_n136_), .A1(x2), .B0(ori_ori_n2162_), .Y(ori_ori_n2163_));
  NA3        o2114(.A(ori_ori_n407_), .B(ori_ori_n326_), .C(ori_ori_n77_), .Y(ori_ori_n2164_));
  OA210      o2115(.A0(ori_ori_n243_), .A1(ori_ori_n226_), .B0(ori_ori_n2164_), .Y(ori_ori_n2165_));
  AOI210     o2116(.A0(ori_ori_n2165_), .A1(ori_ori_n2163_), .B0(ori_ori_n64_), .Y(ori_ori_n2166_));
  NA2        o2117(.A(ori_ori_n119_), .B(ori_ori_n57_), .Y(ori_ori_n2167_));
  AOI220     o2118(.A0(ori_ori_n1574_), .A1(ori_ori_n902_), .B0(ori_ori_n272_), .B1(x4), .Y(ori_ori_n2168_));
  AOI220     o2119(.A0(ori_ori_n1627_), .A1(ori_ori_n616_), .B0(ori_ori_n719_), .B1(ori_ori_n768_), .Y(ori_ori_n2169_));
  OAI220     o2120(.A0(ori_ori_n2169_), .A1(ori_ori_n2167_), .B0(ori_ori_n2168_), .B1(ori_ori_n187_), .Y(ori_ori_n2170_));
  OR3        o2121(.A(ori_ori_n2170_), .B(ori_ori_n2166_), .C(ori_ori_n2161_), .Y(ori_ori_n2171_));
  NO4        o2122(.A(ori_ori_n2171_), .B(ori_ori_n2156_), .C(ori_ori_n2146_), .D(ori_ori_n2136_), .Y(ori_ori_n2172_));
  OAI210     o2123(.A0(ori_ori_n2122_), .A1(x3), .B0(ori_ori_n2172_), .Y(ori32));
  OAI210     o2124(.A0(ori_ori_n564_), .A1(ori_ori_n53_), .B0(ori_ori_n412_), .Y(ori_ori_n2174_));
  NA2        o2125(.A(ori_ori_n513_), .B(x2), .Y(ori_ori_n2175_));
  AOI210     o2126(.A0(ori_ori_n2175_), .A1(ori_ori_n2174_), .B0(ori_ori_n57_), .Y(ori_ori_n2176_));
  OAI210     o2127(.A0(ori_ori_n2176_), .A1(ori_ori_n783_), .B0(ori_ori_n56_), .Y(ori_ori_n2177_));
  OAI210     o2128(.A0(ori_ori_n1698_), .A1(ori_ori_n1440_), .B0(ori_ori_n1470_), .Y(ori_ori_n2178_));
  AOI210     o2129(.A0(ori_ori_n2101_), .A1(ori_ori_n276_), .B0(ori_ori_n2178_), .Y(ori_ori_n2179_));
  AOI210     o2130(.A0(ori_ori_n2179_), .A1(ori_ori_n2177_), .B0(ori_ori_n50_), .Y(ori_ori_n2180_));
  NA3        o2131(.A(ori_ori_n1543_), .B(ori_ori_n798_), .C(ori_ori_n288_), .Y(ori_ori_n2181_));
  NA2        o2132(.A(ori_ori_n740_), .B(ori_ori_n546_), .Y(ori_ori_n2182_));
  OAI220     o2133(.A0(ori_ori_n1050_), .A1(ori_ori_n228_), .B0(ori_ori_n681_), .B1(ori_ori_n204_), .Y(ori_ori_n2183_));
  NO3        o2134(.A(ori_ori_n372_), .B(ori_ori_n574_), .C(ori_ori_n804_), .Y(ori_ori_n2184_));
  NO3        o2135(.A(ori_ori_n1356_), .B(ori_ori_n584_), .C(ori_ori_n270_), .Y(ori_ori_n2185_));
  NO4        o2136(.A(ori_ori_n2185_), .B(ori_ori_n2184_), .C(ori_ori_n2183_), .D(ori_ori_n2182_), .Y(ori_ori_n2186_));
  AOI210     o2137(.A0(ori_ori_n2186_), .A1(ori_ori_n2181_), .B0(ori_ori_n140_), .Y(ori_ori_n2187_));
  OAI220     o2138(.A0(ori_ori_n400_), .A1(x7), .B0(ori_ori_n301_), .B1(ori_ori_n294_), .Y(ori_ori_n2188_));
  NA2        o2139(.A(ori_ori_n2188_), .B(ori_ori_n955_), .Y(ori_ori_n2189_));
  NO2        o2140(.A(ori_ori_n551_), .B(ori_ori_n858_), .Y(ori_ori_n2190_));
  AOI220     o2141(.A0(ori_ori_n2190_), .A1(ori_ori_n1868_), .B0(ori_ori_n530_), .B1(ori_ori_n129_), .Y(ori_ori_n2191_));
  AOI210     o2142(.A0(ori_ori_n2191_), .A1(ori_ori_n2189_), .B0(ori_ori_n106_), .Y(ori_ori_n2192_));
  NA3        o2143(.A(ori_ori_n1311_), .B(ori_ori_n1141_), .C(ori_ori_n113_), .Y(ori_ori_n2193_));
  AOI220     o2144(.A0(ori_ori_n1348_), .A1(ori_ori_n698_), .B0(ori_ori_n1236_), .B1(ori_ori_n1038_), .Y(ori_ori_n2194_));
  AOI210     o2145(.A0(ori_ori_n2194_), .A1(ori_ori_n2193_), .B0(ori_ori_n56_), .Y(ori_ori_n2195_));
  NA2        o2146(.A(ori_ori_n955_), .B(ori_ori_n57_), .Y(ori_ori_n2196_));
  NOi21      o2147(.An(ori_ori_n2196_), .B(ori_ori_n129_), .Y(ori_ori_n2197_));
  NA2        o2148(.A(ori_ori_n1009_), .B(ori_ori_n248_), .Y(ori_ori_n2198_));
  NO3        o2149(.A(ori_ori_n2198_), .B(ori_ori_n2197_), .C(ori_ori_n59_), .Y(ori_ori_n2199_));
  OR4        o2150(.A(ori_ori_n2199_), .B(ori_ori_n2195_), .C(ori_ori_n2192_), .D(ori_ori_n2187_), .Y(ori_ori_n2200_));
  OAI210     o2151(.A0(ori_ori_n2200_), .A1(ori_ori_n2180_), .B0(ori_ori_n104_), .Y(ori_ori_n2201_));
  NO3        o2152(.A(ori_ori_n1222_), .B(ori_ori_n144_), .C(ori_ori_n122_), .Y(ori_ori_n2202_));
  NO2        o2153(.A(ori_ori_n379_), .B(ori_ori_n55_), .Y(ori_ori_n2203_));
  NA2        o2154(.A(ori_ori_n2203_), .B(ori_ori_n112_), .Y(ori_ori_n2204_));
  OAI210     o2155(.A0(ori_ori_n632_), .A1(ori_ori_n590_), .B0(ori_ori_n809_), .Y(ori_ori_n2205_));
  NA2        o2156(.A(ori_ori_n2205_), .B(ori_ori_n2204_), .Y(ori_ori_n2206_));
  OAI210     o2157(.A0(ori_ori_n2206_), .A1(ori_ori_n2202_), .B0(x3), .Y(ori_ori_n2207_));
  OAI210     o2158(.A0(ori_ori_n890_), .A1(ori_ori_n270_), .B0(ori_ori_n50_), .Y(ori_ori_n2208_));
  AOI210     o2159(.A0(ori_ori_n62_), .A1(ori_ori_n106_), .B0(ori_ori_n2208_), .Y(ori_ori_n2209_));
  OAI210     o2160(.A0(ori_ori_n2209_), .A1(ori_ori_n1849_), .B0(ori_ori_n697_), .Y(ori_ori_n2210_));
  NO3        o2161(.A(ori_ori_n303_), .B(ori_ori_n171_), .C(ori_ori_n120_), .Y(ori_ori_n2211_));
  NO3        o2162(.A(ori_ori_n798_), .B(ori_ori_n360_), .C(ori_ori_n140_), .Y(ori_ori_n2212_));
  OAI210     o2163(.A0(ori_ori_n2212_), .A1(ori_ori_n2211_), .B0(ori_ori_n59_), .Y(ori_ori_n2213_));
  NA2        o2164(.A(ori_ori_n1145_), .B(ori_ori_n71_), .Y(ori_ori_n2214_));
  NO2        o2165(.A(ori_ori_n1920_), .B(ori_ori_n590_), .Y(ori_ori_n2215_));
  AOI210     o2166(.A0(ori_ori_n2215_), .A1(ori_ori_n1850_), .B0(ori_ori_n2214_), .Y(ori_ori_n2216_));
  NO2        o2167(.A(ori_ori_n273_), .B(ori_ori_n57_), .Y(ori_ori_n2217_));
  NO2        o2168(.A(ori_ori_n2217_), .B(ori_ori_n1001_), .Y(ori_ori_n2218_));
  NOi31      o2169(.An(ori_ori_n720_), .B(ori_ori_n2218_), .C(ori_ori_n279_), .Y(ori_ori_n2219_));
  NO3        o2170(.A(ori_ori_n1303_), .B(ori_ori_n213_), .C(ori_ori_n255_), .Y(ori_ori_n2220_));
  NO4        o2171(.A(ori_ori_n2220_), .B(ori_ori_n2219_), .C(ori_ori_n2216_), .D(x1), .Y(ori_ori_n2221_));
  NA4        o2172(.A(ori_ori_n2221_), .B(ori_ori_n2213_), .C(ori_ori_n2210_), .D(ori_ori_n2207_), .Y(ori_ori_n2222_));
  AO210      o2173(.A0(ori_ori_n1088_), .A1(ori_ori_n395_), .B0(ori_ori_n1004_), .Y(ori_ori_n2223_));
  NA3        o2174(.A(ori_ori_n1894_), .B(ori_ori_n555_), .C(ori_ori_n273_), .Y(ori_ori_n2224_));
  AOI210     o2175(.A0(ori_ori_n2224_), .A1(ori_ori_n2223_), .B0(ori_ori_n303_), .Y(ori_ori_n2225_));
  NA4        o2176(.A(ori_ori_n1259_), .B(ori_ori_n527_), .C(ori_ori_n384_), .D(ori_ori_n228_), .Y(ori_ori_n2226_));
  NO3        o2177(.A(ori_ori_n1422_), .B(ori_ori_n1004_), .C(x2), .Y(ori_ori_n2227_));
  NO2        o2178(.A(ori_ori_n1245_), .B(ori_ori_n382_), .Y(ori_ori_n2228_));
  NO2        o2179(.A(ori_ori_n1822_), .B(ori_ori_n64_), .Y(ori_ori_n2229_));
  NO4        o2180(.A(ori_ori_n2229_), .B(ori_ori_n2228_), .C(ori_ori_n2227_), .D(ori_ori_n53_), .Y(ori_ori_n2230_));
  NO3        o2181(.A(ori_ori_n465_), .B(ori_ori_n1082_), .C(ori_ori_n119_), .Y(ori_ori_n2231_));
  OAI220     o2182(.A0(ori_ori_n684_), .A1(ori_ori_n171_), .B0(ori_ori_n352_), .B1(ori_ori_n140_), .Y(ori_ori_n2232_));
  OAI210     o2183(.A0(ori_ori_n2232_), .A1(ori_ori_n2231_), .B0(ori_ori_n68_), .Y(ori_ori_n2233_));
  NO2        o2184(.A(ori_ori_n1967_), .B(ori_ori_n363_), .Y(ori_ori_n2234_));
  OAI210     o2185(.A0(ori_ori_n1855_), .A1(ori_ori_n608_), .B0(ori_ori_n2234_), .Y(ori_ori_n2235_));
  NA4        o2186(.A(ori_ori_n2235_), .B(ori_ori_n2233_), .C(ori_ori_n2230_), .D(ori_ori_n2226_), .Y(ori_ori_n2236_));
  OAI210     o2187(.A0(ori_ori_n2236_), .A1(ori_ori_n2225_), .B0(ori_ori_n2222_), .Y(ori_ori_n2237_));
  NO3        o2188(.A(ori_ori_n1210_), .B(ori_ori_n103_), .C(ori_ori_n71_), .Y(ori_ori_n2238_));
  NO2        o2189(.A(ori_ori_n564_), .B(ori_ori_n367_), .Y(ori_ori_n2239_));
  OAI210     o2190(.A0(ori_ori_n2238_), .A1(ori_ori_n1402_), .B0(ori_ori_n2239_), .Y(ori_ori_n2240_));
  NO3        o2191(.A(x8), .B(ori_ori_n71_), .C(x2), .Y(ori_ori_n2241_));
  OAI220     o2192(.A0(ori_ori_n2241_), .A1(ori_ori_n624_), .B0(ori_ori_n1412_), .B1(ori_ori_n89_), .Y(ori_ori_n2242_));
  AOI220     o2193(.A0(ori_ori_n556_), .A1(ori_ori_n809_), .B0(ori_ori_n674_), .B1(ori_ori_n253_), .Y(ori_ori_n2243_));
  AOI210     o2194(.A0(ori_ori_n2243_), .A1(ori_ori_n2242_), .B0(ori_ori_n263_), .Y(ori_ori_n2244_));
  NA2        o2195(.A(ori_ori_n1009_), .B(ori_ori_n1139_), .Y(ori_ori_n2245_));
  AOI210     o2196(.A0(ori_ori_n670_), .A1(ori_ori_n684_), .B0(ori_ori_n2245_), .Y(ori_ori_n2246_));
  AOI210     o2197(.A0(ori_ori_n588_), .A1(ori_ori_n624_), .B0(ori_ori_n690_), .Y(ori_ori_n2247_));
  NO2        o2198(.A(ori_ori_n2247_), .B(ori_ori_n1804_), .Y(ori_ori_n2248_));
  NO2        o2199(.A(ori_ori_n449_), .B(ori_ori_n430_), .Y(ori_ori_n2249_));
  NOi31      o2200(.An(ori_ori_n1489_), .B(ori_ori_n2249_), .C(ori_ori_n588_), .Y(ori_ori_n2250_));
  NO4        o2201(.A(ori_ori_n2250_), .B(ori_ori_n2248_), .C(ori_ori_n2246_), .D(ori_ori_n2244_), .Y(ori_ori_n2251_));
  NA4        o2202(.A(ori_ori_n2251_), .B(ori_ori_n2240_), .C(ori_ori_n2237_), .D(ori_ori_n2201_), .Y(ori33));
  OAI210     o2203(.A0(ori_ori_n805_), .A1(x1), .B0(ori_ori_n198_), .Y(ori_ori_n2253_));
  OAI210     o2204(.A0(ori_ori_n2071_), .A1(ori_ori_n175_), .B0(ori_ori_n326_), .Y(ori_ori_n2254_));
  OAI220     o2205(.A0(ori_ori_n1068_), .A1(ori_ori_n804_), .B0(ori_ori_n1662_), .B1(ori_ori_n351_), .Y(ori_ori_n2255_));
  NA3        o2206(.A(ori_ori_n2255_), .B(ori_ori_n2254_), .C(ori_ori_n633_), .Y(ori_ori_n2256_));
  AOI210     o2207(.A0(ori_ori_n2253_), .A1(x5), .B0(ori_ori_n2256_), .Y(ori_ori_n2257_));
  NA2        o2208(.A(ori_ori_n227_), .B(ori_ori_n76_), .Y(ori_ori_n2258_));
  NA4        o2209(.A(ori_ori_n1736_), .B(ori_ori_n565_), .C(ori_ori_n244_), .D(x4), .Y(ori_ori_n2259_));
  AOI210     o2210(.A0(ori_ori_n2259_), .A1(ori_ori_n2258_), .B0(ori_ori_n351_), .Y(ori_ori_n2260_));
  OAI210     o2211(.A0(ori_ori_n433_), .A1(ori_ori_n267_), .B0(ori_ori_n53_), .Y(ori_ori_n2261_));
  AOI210     o2212(.A0(ori_ori_n2261_), .A1(ori_ori_n435_), .B0(ori_ori_n64_), .Y(ori_ori_n2262_));
  NA2        o2213(.A(ori_ori_n1650_), .B(ori_ori_n71_), .Y(ori_ori_n2263_));
  NO3        o2214(.A(ori_ori_n2263_), .B(ori_ori_n2262_), .C(ori_ori_n2260_), .Y(ori_ori_n2264_));
  OAI210     o2215(.A0(ori_ori_n2257_), .A1(x4), .B0(ori_ori_n2264_), .Y(ori_ori_n2265_));
  OAI210     o2216(.A0(ori_ori_n142_), .A1(x5), .B0(ori_ori_n237_), .Y(ori_ori_n2266_));
  NA2        o2217(.A(ori_ori_n182_), .B(x4), .Y(ori_ori_n2267_));
  NA2        o2218(.A(ori_ori_n308_), .B(ori_ori_n285_), .Y(ori_ori_n2268_));
  NO2        o2219(.A(ori_ori_n955_), .B(ori_ori_n225_), .Y(ori_ori_n2269_));
  NA2        o2220(.A(ori_ori_n636_), .B(x7), .Y(ori_ori_n2270_));
  OAI220     o2221(.A0(ori_ori_n2270_), .A1(ori_ori_n2269_), .B0(ori_ori_n2268_), .B1(ori_ori_n2267_), .Y(ori_ori_n2271_));
  AOI210     o2222(.A0(ori_ori_n2266_), .A1(ori_ori_n1017_), .B0(ori_ori_n2271_), .Y(ori_ori_n2272_));
  NA2        o2223(.A(ori_ori_n209_), .B(ori_ori_n948_), .Y(ori_ori_n2273_));
  AOI210     o2224(.A0(ori_ori_n2273_), .A1(ori_ori_n2196_), .B0(ori_ori_n211_), .Y(ori_ori_n2274_));
  NO2        o2225(.A(ori_ori_n1636_), .B(ori_ori_n949_), .Y(ori_ori_n2275_));
  OAI210     o2226(.A0(ori_ori_n858_), .A1(ori_ori_n51_), .B0(x6), .Y(ori_ori_n2276_));
  NA3        o2227(.A(ori_ori_n912_), .B(ori_ori_n724_), .C(ori_ori_n55_), .Y(ori_ori_n2277_));
  OAI210     o2228(.A0(ori_ori_n618_), .A1(ori_ori_n504_), .B0(ori_ori_n2277_), .Y(ori_ori_n2278_));
  NO4        o2229(.A(ori_ori_n2278_), .B(ori_ori_n2276_), .C(ori_ori_n2275_), .D(ori_ori_n2274_), .Y(ori_ori_n2279_));
  OAI210     o2230(.A0(ori_ori_n2272_), .A1(ori_ori_n50_), .B0(ori_ori_n2279_), .Y(ori_ori_n2280_));
  NA3        o2231(.A(ori_ori_n2280_), .B(ori_ori_n2265_), .C(ori_ori_n59_), .Y(ori_ori_n2281_));
  NA2        o2232(.A(ori_ori_n534_), .B(ori_ori_n105_), .Y(ori_ori_n2282_));
  NO3        o2233(.A(ori_ori_n1555_), .B(ori_ori_n371_), .C(x4), .Y(ori_ori_n2283_));
  AOI210     o2234(.A0(ori_ori_n2283_), .A1(ori_ori_n2282_), .B0(ori_ori_n436_), .Y(ori_ori_n2284_));
  NA2        o2235(.A(ori_ori_n807_), .B(ori_ori_n104_), .Y(ori_ori_n2285_));
  NA2        o2236(.A(ori_ori_n500_), .B(ori_ori_n53_), .Y(ori_ori_n2286_));
  INV        o2237(.A(ori_ori_n2286_), .Y(ori_ori_n2287_));
  OAI210     o2238(.A0(ori_ori_n2284_), .A1(ori_ori_n59_), .B0(ori_ori_n2287_), .Y(ori_ori_n2288_));
  AOI220     o2239(.A0(ori_ori_n684_), .A1(ori_ori_n234_), .B0(ori_ori_n384_), .B1(ori_ori_n228_), .Y(ori_ori_n2289_));
  NA2        o2240(.A(ori_ori_n725_), .B(ori_ori_n967_), .Y(ori_ori_n2290_));
  OAI210     o2241(.A0(ori_ori_n2290_), .A1(ori_ori_n2289_), .B0(ori_ori_n302_), .Y(ori_ori_n2291_));
  AOI210     o2242(.A0(ori_ori_n2101_), .A1(ori_ori_n212_), .B0(ori_ori_n53_), .Y(ori_ori_n2292_));
  NO2        o2243(.A(ori_ori_n140_), .B(ori_ori_n336_), .Y(ori_ori_n2293_));
  AOI220     o2244(.A0(ori_ori_n2293_), .A1(ori_ori_n987_), .B0(ori_ori_n669_), .B1(ori_ori_n351_), .Y(ori_ori_n2294_));
  NA2        o2245(.A(ori_ori_n444_), .B(ori_ori_n498_), .Y(ori_ori_n2295_));
  NO3        o2246(.A(ori_ori_n2295_), .B(ori_ori_n1023_), .C(ori_ori_n180_), .Y(ori_ori_n2296_));
  AOI210     o2247(.A0(ori_ori_n1782_), .A1(ori_ori_n1182_), .B0(ori_ori_n2296_), .Y(ori_ori_n2297_));
  NA4        o2248(.A(ori_ori_n2297_), .B(ori_ori_n2294_), .C(ori_ori_n2292_), .D(ori_ori_n2291_), .Y(ori_ori_n2298_));
  NA3        o2249(.A(ori_ori_n2298_), .B(ori_ori_n2288_), .C(ori_ori_n57_), .Y(ori_ori_n2299_));
  NAi21      o2250(.An(ori_ori_n1184_), .B(ori_ori_n488_), .Y(ori_ori_n2300_));
  NA4        o2251(.A(ori_ori_n636_), .B(ori_ori_n1294_), .C(ori_ori_n469_), .D(ori_ori_n50_), .Y(ori_ori_n2301_));
  OAI210     o2252(.A0(ori_ori_n2293_), .A1(ori_ori_n2046_), .B0(x2), .Y(ori_ori_n2302_));
  NA4        o2253(.A(ori_ori_n285_), .B(ori_ori_n155_), .C(ori_ori_n274_), .D(ori_ori_n119_), .Y(ori_ori_n2303_));
  NA3        o2254(.A(ori_ori_n2303_), .B(ori_ori_n2302_), .C(ori_ori_n2301_), .Y(ori_ori_n2304_));
  AO220      o2255(.A0(ori_ori_n2304_), .A1(x0), .B0(ori_ori_n2300_), .B1(ori_ori_n137_), .Y(ori_ori_n2305_));
  NA3        o2256(.A(ori_ori_n768_), .B(ori_ori_n351_), .C(ori_ori_n60_), .Y(ori_ori_n2306_));
  NO2        o2257(.A(ori_ori_n2241_), .B(ori_ori_n411_), .Y(ori_ori_n2307_));
  NA2        o2258(.A(ori_ori_n634_), .B(ori_ori_n516_), .Y(ori_ori_n2308_));
  OAI220     o2259(.A0(ori_ori_n2308_), .A1(ori_ori_n2307_), .B0(ori_ori_n2306_), .B1(ori_ori_n71_), .Y(ori_ori_n2309_));
  OAI210     o2260(.A0(ori_ori_n1519_), .A1(ori_ori_n347_), .B0(ori_ori_n107_), .Y(ori_ori_n2310_));
  AOI210     o2261(.A0(ori_ori_n588_), .A1(ori_ori_n465_), .B0(ori_ori_n137_), .Y(ori_ori_n2311_));
  OAI210     o2262(.A0(ori_ori_n2311_), .A1(ori_ori_n384_), .B0(ori_ori_n2310_), .Y(ori_ori_n2312_));
  OAI210     o2263(.A0(ori_ori_n2312_), .A1(ori_ori_n2309_), .B0(ori_ori_n98_), .Y(ori_ori_n2313_));
  NA3        o2264(.A(ori_ori_n1202_), .B(ori_ori_n130_), .C(ori_ori_n379_), .Y(ori_ori_n2314_));
  NA2        o2265(.A(ori_ori_n2314_), .B(ori_ori_n1808_), .Y(ori_ori_n2315_));
  NA2        o2266(.A(ori_ori_n1181_), .B(ori_ori_n706_), .Y(ori_ori_n2316_));
  AOI220     o2267(.A0(ori_ori_n2203_), .A1(ori_ori_n293_), .B0(ori_ori_n1348_), .B1(ori_ori_n1163_), .Y(ori_ori_n2317_));
  NA4        o2268(.A(ori_ori_n2317_), .B(ori_ori_n2316_), .C(ori_ori_n2315_), .D(ori_ori_n2313_), .Y(ori_ori_n2318_));
  AOI210     o2269(.A0(ori_ori_n2305_), .A1(x7), .B0(ori_ori_n2318_), .Y(ori_ori_n2319_));
  NA3        o2270(.A(ori_ori_n2319_), .B(ori_ori_n2299_), .C(ori_ori_n2281_), .Y(ori34));
  NA2        o2271(.A(ori_ori_n430_), .B(x4), .Y(ori_ori_n2321_));
  NO2        o2272(.A(ori_ori_n1945_), .B(ori_ori_n851_), .Y(ori_ori_n2322_));
  AOI210     o2273(.A0(ori_ori_n2322_), .A1(ori_ori_n2321_), .B0(ori_ori_n317_), .Y(ori_ori_n2323_));
  NA2        o2274(.A(ori_ori_n285_), .B(ori_ori_n120_), .Y(ori_ori_n2324_));
  NO2        o2275(.A(ori_ori_n965_), .B(ori_ori_n2324_), .Y(ori_ori_n2325_));
  AOI210     o2276(.A0(ori_ori_n2026_), .A1(ori_ori_n542_), .B0(ori_ori_n139_), .Y(ori_ori_n2326_));
  NO2        o2277(.A(ori_ori_n1817_), .B(ori_ori_n969_), .Y(ori_ori_n2327_));
  NO4        o2278(.A(ori_ori_n2327_), .B(ori_ori_n2326_), .C(ori_ori_n2325_), .D(ori_ori_n2323_), .Y(ori_ori_n2328_));
  NO2        o2279(.A(ori_ori_n2328_), .B(ori_ori_n475_), .Y(ori_ori_n2329_));
  NA2        o2280(.A(ori_ori_n727_), .B(x8), .Y(ori_ori_n2330_));
  AO210      o2281(.A0(ori_ori_n2330_), .A1(ori_ori_n485_), .B0(ori_ori_n659_), .Y(ori_ori_n2331_));
  NA2        o2282(.A(ori_ori_n669_), .B(ori_ori_n629_), .Y(ori_ori_n2332_));
  AOI210     o2283(.A0(ori_ori_n2332_), .A1(ori_ori_n2331_), .B0(ori_ori_n263_), .Y(ori_ori_n2333_));
  OAI210     o2284(.A0(ori_ori_n119_), .A1(ori_ori_n1042_), .B0(ori_ori_n1455_), .Y(ori_ori_n2334_));
  OAI210     o2285(.A0(ori_ori_n1595_), .A1(ori_ori_n58_), .B0(ori_ori_n2334_), .Y(ori_ori_n2335_));
  NA3        o2286(.A(ori_ori_n2335_), .B(ori_ori_n337_), .C(x8), .Y(ori_ori_n2336_));
  NO3        o2287(.A(ori_ori_n986_), .B(ori_ori_n703_), .C(ori_ori_n454_), .Y(ori_ori_n2337_));
  AOI210     o2288(.A0(ori_ori_n1577_), .A1(ori_ori_n325_), .B0(ori_ori_n2337_), .Y(ori_ori_n2338_));
  NA2        o2289(.A(ori_ori_n663_), .B(ori_ori_n317_), .Y(ori_ori_n2339_));
  NA2        o2290(.A(ori_ori_n133_), .B(x0), .Y(ori_ori_n2340_));
  NAi31      o2291(.An(ori_ori_n2340_), .B(ori_ori_n2339_), .C(ori_ori_n792_), .Y(ori_ori_n2341_));
  NA3        o2292(.A(ori_ori_n1590_), .B(ori_ori_n1388_), .C(ori_ori_n50_), .Y(ori_ori_n2342_));
  NA4        o2293(.A(ori_ori_n2342_), .B(ori_ori_n2341_), .C(ori_ori_n2338_), .D(ori_ori_n2336_), .Y(ori_ori_n2343_));
  NA2        o2294(.A(ori_ori_n1101_), .B(ori_ori_n743_), .Y(ori_ori_n2344_));
  NA3        o2295(.A(ori_ori_n1141_), .B(ori_ori_n166_), .C(ori_ori_n1085_), .Y(ori_ori_n2345_));
  AOI210     o2296(.A0(ori_ori_n2345_), .A1(ori_ori_n2344_), .B0(ori_ori_n753_), .Y(ori_ori_n2346_));
  AOI210     o2297(.A0(ori_ori_n1766_), .A1(ori_ori_n129_), .B0(ori_ori_n2346_), .Y(ori_ori_n2347_));
  AOI210     o2298(.A0(ori_ori_n556_), .A1(ori_ori_n809_), .B0(ori_ori_n252_), .Y(ori_ori_n2348_));
  OAI220     o2299(.A0(ori_ori_n2348_), .A1(ori_ori_n59_), .B0(ori_ori_n1112_), .B1(ori_ori_n55_), .Y(ori_ori_n2349_));
  NA3        o2300(.A(ori_ori_n2349_), .B(ori_ori_n727_), .C(ori_ori_n56_), .Y(ori_ori_n2350_));
  OAI210     o2301(.A0(ori_ori_n2347_), .A1(ori_ori_n140_), .B0(ori_ori_n2350_), .Y(ori_ori_n2351_));
  NO4        o2302(.A(ori_ori_n2351_), .B(ori_ori_n2343_), .C(ori_ori_n2333_), .D(ori_ori_n2329_), .Y(ori_ori_n2352_));
  NO2        o2303(.A(ori_ori_n309_), .B(ori_ori_n948_), .Y(ori_ori_n2353_));
  NO3        o2304(.A(ori_ori_n2353_), .B(ori_ori_n442_), .C(ori_ori_n325_), .Y(ori_ori_n2354_));
  NA2        o2305(.A(ori_ori_n777_), .B(ori_ori_n159_), .Y(ori_ori_n2355_));
  NO3        o2306(.A(ori_ori_n2217_), .B(ori_ori_n302_), .C(ori_ori_n1085_), .Y(ori_ori_n2356_));
  OAI220     o2307(.A0(ori_ori_n2356_), .A1(ori_ori_n1547_), .B0(ori_ori_n2355_), .B1(ori_ori_n1166_), .Y(ori_ori_n2357_));
  OAI210     o2308(.A0(ori_ori_n2357_), .A1(ori_ori_n2354_), .B0(x2), .Y(ori_ori_n2358_));
  OAI210     o2309(.A0(ori_ori_n861_), .A1(ori_ori_n367_), .B0(ori_ori_n2358_), .Y(ori_ori_n2359_));
  NA2        o2310(.A(ori_ori_n312_), .B(x4), .Y(ori_ori_n2360_));
  OAI220     o2311(.A0(ori_ori_n739_), .A1(ori_ori_n55_), .B0(ori_ori_n278_), .B1(ori_ori_n103_), .Y(ori_ori_n2361_));
  NO4        o2312(.A(ori_ori_n446_), .B(ori_ori_n77_), .C(x7), .D(x3), .Y(ori_ori_n2362_));
  NO2        o2313(.A(ori_ori_n1101_), .B(ori_ori_n286_), .Y(ori_ori_n2363_));
  NO4        o2314(.A(ori_ori_n2363_), .B(ori_ori_n2362_), .C(ori_ori_n2361_), .D(ori_ori_n2360_), .Y(ori_ori_n2364_));
  NA2        o2315(.A(ori_ori_n1236_), .B(ori_ori_n1040_), .Y(ori_ori_n2365_));
  NA4        o2316(.A(ori_ori_n727_), .B(ori_ori_n176_), .C(ori_ori_n57_), .D(ori_ori_n104_), .Y(ori_ori_n2366_));
  NA3        o2317(.A(ori_ori_n1385_), .B(ori_ori_n255_), .C(x7), .Y(ori_ori_n2367_));
  NA3        o2318(.A(ori_ori_n2367_), .B(ori_ori_n2366_), .C(ori_ori_n2365_), .Y(ori_ori_n2368_));
  OAI210     o2319(.A0(ori_ori_n2368_), .A1(ori_ori_n2364_), .B0(ori_ori_n163_), .Y(ori_ori_n2369_));
  NA3        o2320(.A(ori_ori_n856_), .B(ori_ori_n87_), .C(x0), .Y(ori_ori_n2370_));
  NA4        o2321(.A(ori_ori_n2370_), .B(ori_ori_n1145_), .C(ori_ori_n295_), .D(ori_ori_n586_), .Y(ori_ori_n2371_));
  NA2        o2322(.A(ori_ori_n1149_), .B(ori_ori_n674_), .Y(ori_ori_n2372_));
  OAI210     o2323(.A0(ori_ori_n2372_), .A1(ori_ori_n264_), .B0(ori_ori_n2153_), .Y(ori_ori_n2373_));
  AOI220     o2324(.A0(ori_ori_n2373_), .A1(x7), .B0(ori_ori_n1008_), .B1(ori_ori_n660_), .Y(ori_ori_n2374_));
  OAI210     o2325(.A0(ori_ori_n2039_), .A1(ori_ori_n260_), .B0(ori_ori_n731_), .Y(ori_ori_n2375_));
  AOI220     o2326(.A0(ori_ori_n407_), .A1(x8), .B0(ori_ori_n90_), .B1(x2), .Y(ori_ori_n2376_));
  AOI210     o2327(.A0(ori_ori_n268_), .A1(ori_ori_n53_), .B0(ori_ori_n651_), .Y(ori_ori_n2377_));
  OAI220     o2328(.A0(ori_ori_n2377_), .A1(ori_ori_n93_), .B0(ori_ori_n2376_), .B1(ori_ori_n1334_), .Y(ori_ori_n2378_));
  AOI220     o2329(.A0(ori_ori_n2378_), .A1(ori_ori_n1312_), .B0(ori_ori_n2375_), .B1(ori_ori_n1504_), .Y(ori_ori_n2379_));
  NA4        o2330(.A(ori_ori_n2379_), .B(ori_ori_n2374_), .C(ori_ori_n2371_), .D(ori_ori_n2369_), .Y(ori_ori_n2380_));
  AOI210     o2331(.A0(ori_ori_n2359_), .A1(ori_ori_n809_), .B0(ori_ori_n2380_), .Y(ori_ori_n2381_));
  OAI210     o2332(.A0(ori_ori_n2352_), .A1(x2), .B0(ori_ori_n2381_), .Y(ori35));
  NA2        o2333(.A(ori_ori_n504_), .B(ori_ori_n176_), .Y(ori_ori_n2383_));
  AOI220     o2334(.A0(ori_ori_n634_), .A1(ori_ori_n55_), .B0(ori_ori_n768_), .B1(ori_ori_n1217_), .Y(ori_ori_n2384_));
  AOI210     o2335(.A0(ori_ori_n2384_), .A1(ori_ori_n2383_), .B0(ori_ori_n71_), .Y(ori_ori_n2385_));
  NO3        o2336(.A(ori_ori_n512_), .B(ori_ori_n465_), .C(ori_ori_n336_), .Y(ori_ori_n2386_));
  OAI210     o2337(.A0(ori_ori_n2386_), .A1(ori_ori_n2385_), .B0(x2), .Y(ori_ori_n2387_));
  AOI210     o2338(.A0(ori_ori_n213_), .A1(x0), .B0(ori_ori_n272_), .Y(ori_ori_n2388_));
  OAI220     o2339(.A0(ori_ori_n2388_), .A1(ori_ori_n665_), .B0(ori_ori_n195_), .B1(x4), .Y(ori_ori_n2389_));
  NA2        o2340(.A(ori_ori_n2389_), .B(ori_ori_n137_), .Y(ori_ori_n2390_));
  NA3        o2341(.A(ori_ori_n407_), .B(x8), .C(ori_ori_n71_), .Y(ori_ori_n2391_));
  AOI210     o2342(.A0(ori_ori_n2391_), .A1(ori_ori_n1712_), .B0(ori_ori_n684_), .Y(ori_ori_n2392_));
  OAI210     o2343(.A0(ori_ori_n2306_), .A1(x6), .B0(ori_ori_n742_), .Y(ori_ori_n2393_));
  NO2        o2344(.A(ori_ori_n2393_), .B(ori_ori_n2392_), .Y(ori_ori_n2394_));
  NA3        o2345(.A(ori_ori_n2394_), .B(ori_ori_n2390_), .C(ori_ori_n2387_), .Y(ori_ori_n2395_));
  NAi21      o2346(.An(ori_ori_n1677_), .B(ori_ori_n1291_), .Y(ori_ori_n2396_));
  NA2        o2347(.A(ori_ori_n211_), .B(ori_ori_n574_), .Y(ori_ori_n2397_));
  NO2        o2348(.A(ori_ori_n430_), .B(ori_ori_n423_), .Y(ori_ori_n2398_));
  AOI220     o2349(.A0(ori_ori_n2398_), .A1(ori_ori_n2397_), .B0(ori_ori_n2396_), .B1(ori_ori_n56_), .Y(ori_ori_n2399_));
  NA2        o2350(.A(ori_ori_n757_), .B(ori_ori_n695_), .Y(ori_ori_n2400_));
  NO3        o2351(.A(ori_ori_n679_), .B(ori_ori_n55_), .C(x6), .Y(ori_ori_n2401_));
  OAI210     o2352(.A0(ori_ori_n2401_), .A1(ori_ori_n706_), .B0(ori_ori_n216_), .Y(ori_ori_n2402_));
  NA2        o2353(.A(ori_ori_n1320_), .B(ori_ori_n63_), .Y(ori_ori_n2403_));
  NA2        o2354(.A(x6), .B(ori_ori_n470_), .Y(ori_ori_n2404_));
  NA3        o2355(.A(ori_ori_n2404_), .B(ori_ori_n2403_), .C(ori_ori_n2402_), .Y(ori_ori_n2405_));
  NA3        o2356(.A(ori_ori_n1266_), .B(ori_ori_n745_), .C(x3), .Y(ori_ori_n2406_));
  NO3        o2357(.A(ori_ori_n2406_), .B(ori_ori_n681_), .C(ori_ori_n204_), .Y(ori_ori_n2407_));
  AOI210     o2358(.A0(ori_ori_n2405_), .A1(ori_ori_n50_), .B0(ori_ori_n2407_), .Y(ori_ori_n2408_));
  OAI210     o2359(.A0(ori_ori_n2400_), .A1(ori_ori_n2399_), .B0(ori_ori_n2408_), .Y(ori_ori_n2409_));
  AOI210     o2360(.A0(ori_ori_n2395_), .A1(ori_ori_n57_), .B0(ori_ori_n2409_), .Y(ori_ori_n2410_));
  NO3        o2361(.A(ori_ori_n1064_), .B(ori_ori_n564_), .C(ori_ori_n120_), .Y(ori_ori_n2411_));
  OAI210     o2362(.A0(ori_ori_n156_), .A1(ori_ori_n67_), .B0(ori_ori_n2411_), .Y(ori_ori_n2412_));
  NO2        o2363(.A(ori_ori_n2412_), .B(ori_ori_n50_), .Y(ori_ori_n2413_));
  NA4        o2364(.A(ori_ori_n465_), .B(ori_ori_n228_), .C(ori_ori_n866_), .D(ori_ori_n100_), .Y(ori_ori_n2414_));
  OAI210     o2365(.A0(ori_ori_n955_), .A1(ori_ori_n253_), .B0(ori_ori_n746_), .Y(ori_ori_n2415_));
  OAI210     o2366(.A0(ori_ori_n253_), .A1(ori_ori_n585_), .B0(ori_ori_n2150_), .Y(ori_ori_n2416_));
  NA3        o2367(.A(ori_ori_n2416_), .B(ori_ori_n2415_), .C(ori_ori_n2414_), .Y(ori_ori_n2417_));
  OAI210     o2368(.A0(ori_ori_n2417_), .A1(ori_ori_n2413_), .B0(ori_ori_n59_), .Y(ori_ori_n2418_));
  AOI210     o2369(.A0(ori_ori_n856_), .A1(ori_ori_n533_), .B0(ori_ori_n1894_), .Y(ori_ori_n2419_));
  AOI210     o2370(.A0(ori_ori_n564_), .A1(ori_ori_n607_), .B0(ori_ori_n2419_), .Y(ori_ori_n2420_));
  NO4        o2371(.A(ori_ori_n949_), .B(ori_ori_n564_), .C(ori_ori_n360_), .D(ori_ori_n405_), .Y(ori_ori_n2421_));
  XN2        o2372(.A(x4), .B(x3), .Y(ori_ori_n2422_));
  NO3        o2373(.A(ori_ori_n2422_), .B(ori_ori_n664_), .C(ori_ori_n308_), .Y(ori_ori_n2423_));
  NO3        o2374(.A(ori_ori_n2423_), .B(ori_ori_n2421_), .C(ori_ori_n1451_), .Y(ori_ori_n2424_));
  OAI210     o2375(.A0(ori_ori_n2420_), .A1(x3), .B0(ori_ori_n2424_), .Y(ori_ori_n2425_));
  NO3        o2376(.A(ori_ori_n739_), .B(ori_ori_n858_), .C(ori_ori_n273_), .Y(ori_ori_n2426_));
  OAI210     o2377(.A0(ori_ori_n2426_), .A1(ori_ori_n1451_), .B0(ori_ori_n50_), .Y(ori_ori_n2427_));
  NA3        o2378(.A(ori_ori_n1072_), .B(ori_ori_n807_), .C(ori_ori_n252_), .Y(ori_ori_n2428_));
  NA2        o2379(.A(ori_ori_n2428_), .B(ori_ori_n2427_), .Y(ori_ori_n2429_));
  AOI210     o2380(.A0(ori_ori_n2425_), .A1(ori_ori_n588_), .B0(ori_ori_n2429_), .Y(ori_ori_n2430_));
  AOI210     o2381(.A0(ori_ori_n1422_), .A1(ori_ori_n641_), .B0(ori_ori_n681_), .Y(ori_ori_n2431_));
  NO2        o2382(.A(ori_ori_n866_), .B(ori_ori_n56_), .Y(ori_ori_n2432_));
  OAI210     o2383(.A0(ori_ori_n1948_), .A1(ori_ori_n607_), .B0(ori_ori_n2241_), .Y(ori_ori_n2433_));
  OAI210     o2384(.A0(ori_ori_n2330_), .A1(ori_ori_n2432_), .B0(ori_ori_n2433_), .Y(ori_ori_n2434_));
  OAI210     o2385(.A0(ori_ori_n2434_), .A1(ori_ori_n2431_), .B0(ori_ori_n90_), .Y(ori_ori_n2435_));
  NO2        o2386(.A(ori_ori_n849_), .B(ori_ori_n661_), .Y(ori_ori_n2436_));
  NO2        o2387(.A(ori_ori_n286_), .B(x6), .Y(ori_ori_n2437_));
  OAI210     o2388(.A0(ori_ori_n2436_), .A1(ori_ori_n1773_), .B0(ori_ori_n2437_), .Y(ori_ori_n2438_));
  NA4        o2389(.A(ori_ori_n2438_), .B(ori_ori_n2435_), .C(ori_ori_n2430_), .D(ori_ori_n2418_), .Y(ori_ori_n2439_));
  NA4        o2390(.A(ori_ori_n615_), .B(ori_ori_n684_), .C(ori_ori_n429_), .D(x6), .Y(ori_ori_n2440_));
  AOI210     o2391(.A0(ori_ori_n2440_), .A1(ori_ori_n424_), .B0(x1), .Y(ori_ori_n2441_));
  NO2        o2392(.A(ori_ori_n725_), .B(ori_ori_n681_), .Y(ori_ori_n2442_));
  OAI210     o2393(.A0(ori_ori_n465_), .A1(ori_ori_n167_), .B0(ori_ori_n789_), .Y(ori_ori_n2443_));
  AOI210     o2394(.A0(ori_ori_n2443_), .A1(ori_ori_n1013_), .B0(ori_ori_n53_), .Y(ori_ori_n2444_));
  NO3        o2395(.A(ori_ori_n2444_), .B(ori_ori_n2442_), .C(ori_ori_n2441_), .Y(ori_ori_n2445_));
  NA3        o2396(.A(ori_ori_n1424_), .B(ori_ori_n1267_), .C(ori_ori_n813_), .Y(ori_ori_n2446_));
  AOI220     o2397(.A0(ori_ori_n1935_), .A1(ori_ori_n137_), .B0(ori_ori_n416_), .B1(ori_ori_n124_), .Y(ori_ori_n2447_));
  AOI210     o2398(.A0(ori_ori_n2447_), .A1(ori_ori_n2446_), .B0(ori_ori_n1497_), .Y(ori_ori_n2448_));
  NO2        o2399(.A(ori_ori_n634_), .B(x3), .Y(ori_ori_n2449_));
  NO3        o2400(.A(ori_ori_n692_), .B(ori_ori_n1595_), .C(x2), .Y(ori_ori_n2450_));
  AOI220     o2401(.A0(ori_ori_n2450_), .A1(ori_ori_n2449_), .B0(ori_ori_n1908_), .B1(ori_ori_n764_), .Y(ori_ori_n2451_));
  NA3        o2402(.A(x6), .B(x4), .C(x0), .Y(ori_ori_n2452_));
  OAI220     o2403(.A0(ori_ori_n2452_), .A1(ori_ori_n194_), .B0(ori_ori_n679_), .B1(ori_ori_n529_), .Y(ori_ori_n2453_));
  OAI220     o2404(.A0(ori_ori_n1301_), .A1(x8), .B0(ori_ori_n371_), .B1(ori_ori_n350_), .Y(ori_ori_n2454_));
  AOI220     o2405(.A0(ori_ori_n2454_), .A1(ori_ori_n416_), .B0(ori_ori_n2453_), .B1(ori_ori_n911_), .Y(ori_ori_n2455_));
  OAI210     o2406(.A0(ori_ori_n2451_), .A1(ori_ori_n1158_), .B0(ori_ori_n2455_), .Y(ori_ori_n2456_));
  NO2        o2407(.A(ori_ori_n2456_), .B(ori_ori_n2448_), .Y(ori_ori_n2457_));
  OAI210     o2408(.A0(ori_ori_n2445_), .A1(ori_ori_n312_), .B0(ori_ori_n2457_), .Y(ori_ori_n2458_));
  AOI210     o2409(.A0(ori_ori_n2439_), .A1(x5), .B0(ori_ori_n2458_), .Y(ori_ori_n2459_));
  OAI210     o2410(.A0(ori_ori_n2410_), .A1(x5), .B0(ori_ori_n2459_), .Y(ori36));
  NO2        o2411(.A(ori_ori_n858_), .B(ori_ori_n301_), .Y(ori_ori_n2461_));
  NO3        o2412(.A(ori_ori_n119_), .B(ori_ori_n1042_), .C(ori_ori_n55_), .Y(ori_ori_n2462_));
  NO3        o2413(.A(ori_ori_n2462_), .B(ori_ori_n1967_), .C(ori_ori_n1064_), .Y(ori_ori_n2463_));
  OAI210     o2414(.A0(ori_ori_n2463_), .A1(ori_ori_n2461_), .B0(ori_ori_n106_), .Y(ori_ori_n2464_));
  OR4        o2415(.A(ori_ori_n950_), .B(ori_ori_n800_), .C(ori_ori_n374_), .D(ori_ori_n492_), .Y(ori_ori_n2465_));
  INV        o2416(.A(ori_ori_n998_), .Y(ori_ori_n2466_));
  OAI210     o2417(.A0(ori_ori_n2203_), .A1(ori_ori_n2466_), .B0(ori_ori_n278_), .Y(ori_ori_n2467_));
  NA3        o2418(.A(ori_ori_n444_), .B(ori_ori_n225_), .C(ori_ori_n118_), .Y(ori_ori_n2468_));
  NA4        o2419(.A(ori_ori_n2468_), .B(ori_ori_n2467_), .C(ori_ori_n2465_), .D(ori_ori_n2464_), .Y(ori_ori_n2469_));
  NO2        o2420(.A(ori_ori_n987_), .B(x8), .Y(ori_ori_n2470_));
  NO3        o2421(.A(ori_ori_n2470_), .B(ori_ori_n983_), .C(ori_ori_n538_), .Y(ori_ori_n2471_));
  AOI220     o2422(.A0(ori_ori_n302_), .A1(x1), .B0(ori_ori_n136_), .B1(x6), .Y(ori_ori_n2472_));
  AOI210     o2423(.A0(ori_ori_n1085_), .A1(x6), .B0(ori_ori_n420_), .Y(ori_ori_n2473_));
  OAI220     o2424(.A0(ori_ori_n2473_), .A1(ori_ori_n359_), .B0(ori_ori_n2472_), .B1(ori_ori_n466_), .Y(ori_ori_n2474_));
  OAI210     o2425(.A0(ori_ori_n2474_), .A1(ori_ori_n2471_), .B0(ori_ori_n465_), .Y(ori_ori_n2475_));
  NA2        o2426(.A(ori_ori_n669_), .B(ori_ori_n492_), .Y(ori_ori_n2476_));
  AOI210     o2427(.A0(ori_ori_n2476_), .A1(ori_ori_n648_), .B0(ori_ori_n264_), .Y(ori_ori_n2477_));
  NO3        o2428(.A(ori_ori_n1865_), .B(ori_ori_n1594_), .C(ori_ori_n274_), .Y(ori_ori_n2478_));
  NO3        o2429(.A(ori_ori_n2478_), .B(ori_ori_n2477_), .C(ori_ori_n418_), .Y(ori_ori_n2479_));
  OAI210     o2430(.A0(ori_ori_n636_), .A1(ori_ori_n799_), .B0(ori_ori_n973_), .Y(ori_ori_n2480_));
  OAI220     o2431(.A0(ori_ori_n1641_), .A1(ori_ori_n1636_), .B0(ori_ori_n973_), .B1(ori_ori_n1085_), .Y(ori_ori_n2481_));
  AOI220     o2432(.A0(ori_ori_n2481_), .A1(ori_ori_n117_), .B0(ori_ori_n2480_), .B1(ori_ori_n629_), .Y(ori_ori_n2482_));
  NA3        o2433(.A(ori_ori_n2482_), .B(ori_ori_n2479_), .C(ori_ori_n2475_), .Y(ori_ori_n2483_));
  AOI210     o2434(.A0(ori_ori_n2469_), .A1(ori_ori_n337_), .B0(ori_ori_n2483_), .Y(ori_ori_n2484_));
  OAI210     o2435(.A0(ori_ori_n593_), .A1(ori_ori_n517_), .B0(ori_ori_n167_), .Y(ori_ori_n2485_));
  OAI210     o2436(.A0(ori_ori_n1982_), .A1(ori_ori_n70_), .B0(ori_ori_n2485_), .Y(ori_ori_n2486_));
  OAI210     o2437(.A0(ori_ori_n495_), .A1(ori_ori_n236_), .B0(ori_ori_n253_), .Y(ori_ori_n2487_));
  NO2        o2438(.A(ori_ori_n1991_), .B(ori_ori_n172_), .Y(ori_ori_n2488_));
  NA2        o2439(.A(ori_ori_n1204_), .B(ori_ori_n55_), .Y(ori_ori_n2489_));
  OAI210     o2440(.A0(ori_ori_n2489_), .A1(ori_ori_n2488_), .B0(ori_ori_n2487_), .Y(ori_ori_n2490_));
  OAI210     o2441(.A0(ori_ori_n2490_), .A1(ori_ori_n2486_), .B0(ori_ori_n890_), .Y(ori_ori_n2491_));
  AOI210     o2442(.A0(ori_ori_n103_), .A1(ori_ori_n106_), .B0(ori_ori_n339_), .Y(ori_ori_n2492_));
  NA2        o2443(.A(ori_ori_n669_), .B(ori_ori_n1595_), .Y(ori_ori_n2493_));
  OAI220     o2444(.A0(ori_ori_n2493_), .A1(ori_ori_n2492_), .B0(ori_ori_n742_), .B1(ori_ori_n1250_), .Y(ori_ori_n2494_));
  NO2        o2445(.A(ori_ori_n1388_), .B(ori_ori_n580_), .Y(ori_ori_n2495_));
  NO3        o2446(.A(ori_ori_n2495_), .B(ori_ori_n1781_), .C(ori_ori_n692_), .Y(ori_ori_n2496_));
  NOi31      o2447(.An(ori_ori_n2003_), .B(ori_ori_n2295_), .C(ori_ori_n752_), .Y(ori_ori_n2497_));
  NO3        o2448(.A(ori_ori_n2497_), .B(ori_ori_n2496_), .C(ori_ori_n2494_), .Y(ori_ori_n2498_));
  AOI210     o2449(.A0(ori_ori_n2498_), .A1(ori_ori_n2491_), .B0(x7), .Y(ori_ori_n2499_));
  NA2        o2450(.A(ori_ori_n136_), .B(ori_ori_n63_), .Y(ori_ori_n2500_));
  AOI210     o2451(.A0(ori_ori_n588_), .A1(ori_ori_n624_), .B0(ori_ori_n1182_), .Y(ori_ori_n2501_));
  NA4        o2452(.A(ori_ori_n2501_), .B(ori_ori_n2500_), .C(ori_ori_n986_), .D(ori_ori_n883_), .Y(ori_ori_n2502_));
  NA2        o2453(.A(ori_ori_n2502_), .B(ori_ori_n504_), .Y(ori_ori_n2503_));
  AOI220     o2454(.A0(ori_ori_n1736_), .A1(ori_ori_n256_), .B0(ori_ori_n1040_), .B1(ori_ori_n124_), .Y(ori_ori_n2504_));
  NO2        o2455(.A(ori_ori_n2504_), .B(ori_ori_n444_), .Y(ori_ori_n2505_));
  NO2        o2456(.A(ori_ori_n405_), .B(ori_ori_n225_), .Y(ori_ori_n2506_));
  NO3        o2457(.A(ori_ori_n2506_), .B(ori_ori_n1270_), .C(ori_ori_n59_), .Y(ori_ori_n2507_));
  AOI210     o2458(.A0(ori_ori_n1221_), .A1(ori_ori_n406_), .B0(x6), .Y(ori_ori_n2508_));
  NA3        o2459(.A(ori_ori_n1668_), .B(ori_ori_n278_), .C(ori_ori_n268_), .Y(ori_ori_n2509_));
  NA2        o2460(.A(ori_ori_n2509_), .B(ori_ori_n1621_), .Y(ori_ori_n2510_));
  NO4        o2461(.A(ori_ori_n2510_), .B(ori_ori_n2508_), .C(ori_ori_n2507_), .D(ori_ori_n2505_), .Y(ori_ori_n2511_));
  AOI210     o2462(.A0(ori_ori_n2511_), .A1(ori_ori_n2503_), .B0(ori_ori_n454_), .Y(ori_ori_n2512_));
  NO3        o2463(.A(ori_ori_n2422_), .B(ori_ori_n896_), .C(ori_ori_n503_), .Y(ori_ori_n2513_));
  AOI210     o2464(.A0(ori_ori_n1268_), .A1(ori_ori_n267_), .B0(ori_ori_n2513_), .Y(ori_ori_n2514_));
  OAI210     o2465(.A0(ori_ori_n865_), .A1(ori_ori_n273_), .B0(ori_ori_n395_), .Y(ori_ori_n2515_));
  NA2        o2466(.A(ori_ori_n1204_), .B(ori_ori_n171_), .Y(ori_ori_n2516_));
  NO2        o2467(.A(ori_ori_n614_), .B(ori_ori_n106_), .Y(ori_ori_n2517_));
  AO210      o2468(.A0(ori_ori_n2517_), .A1(ori_ori_n2516_), .B0(ori_ori_n1753_), .Y(ori_ori_n2518_));
  NO2        o2469(.A(ori_ori_n461_), .B(ori_ori_n417_), .Y(ori_ori_n2519_));
  AOI220     o2470(.A0(ori_ori_n2519_), .A1(ori_ori_n2518_), .B0(ori_ori_n2515_), .B1(ori_ori_n293_), .Y(ori_ori_n2520_));
  OAI210     o2471(.A0(ori_ori_n2514_), .A1(x1), .B0(ori_ori_n2520_), .Y(ori_ori_n2521_));
  NO3        o2472(.A(ori_ori_n2521_), .B(ori_ori_n2512_), .C(ori_ori_n2499_), .Y(ori_ori_n2522_));
  OAI210     o2473(.A0(ori_ori_n2484_), .A1(ori_ori_n57_), .B0(ori_ori_n2522_), .Y(ori37));
  NA2        o2474(.A(ori_ori_n1061_), .B(x3), .Y(ori_ori_n2524_));
  NA3        o2475(.A(ori_ori_n777_), .B(ori_ori_n159_), .C(ori_ori_n50_), .Y(ori_ori_n2525_));
  AOI210     o2476(.A0(ori_ori_n2525_), .A1(ori_ori_n2524_), .B0(ori_ori_n685_), .Y(ori_ori_n2526_));
  NO3        o2477(.A(ori_ori_n1061_), .B(ori_ori_n374_), .C(ori_ori_n511_), .Y(ori_ori_n2527_));
  OAI210     o2478(.A0(ori_ori_n2527_), .A1(ori_ori_n2526_), .B0(ori_ori_n56_), .Y(ori_ori_n2528_));
  NA2        o2479(.A(ori_ori_n602_), .B(ori_ori_n743_), .Y(ori_ori_n2529_));
  AOI210     o2480(.A0(ori_ori_n2529_), .A1(ori_ori_n1041_), .B0(x3), .Y(ori_ori_n2530_));
  AOI220     o2481(.A0(ori_ori_n602_), .A1(ori_ori_n743_), .B0(ori_ori_n465_), .B1(ori_ori_n1040_), .Y(ori_ori_n2531_));
  NO2        o2482(.A(ori_ori_n664_), .B(ori_ori_n179_), .Y(ori_ori_n2532_));
  OAI220     o2483(.A0(ori_ori_n2532_), .A1(ori_ori_n834_), .B0(ori_ori_n2531_), .B1(ori_ori_n106_), .Y(ori_ori_n2533_));
  OAI210     o2484(.A0(ori_ori_n2533_), .A1(ori_ori_n2530_), .B0(ori_ori_n71_), .Y(ori_ori_n2534_));
  NA2        o2485(.A(ori_ori_n1184_), .B(ori_ori_n1064_), .Y(ori_ori_n2535_));
  OAI210     o2486(.A0(ori_ori_n1206_), .A1(ori_ori_n188_), .B0(ori_ori_n455_), .Y(ori_ori_n2536_));
  NA4        o2487(.A(ori_ori_n2536_), .B(ori_ori_n2535_), .C(ori_ori_n2534_), .D(ori_ori_n2528_), .Y(ori_ori_n2537_));
  NA2        o2488(.A(ori_ori_n423_), .B(ori_ori_n136_), .Y(ori_ori_n2538_));
  NO2        o2489(.A(ori_ori_n1698_), .B(ori_ori_n105_), .Y(ori_ori_n2539_));
  AOI210     o2490(.A0(ori_ori_n1969_), .A1(ori_ori_n859_), .B0(ori_ori_n2539_), .Y(ori_ori_n2540_));
  OAI220     o2491(.A0(ori_ori_n2540_), .A1(ori_ori_n51_), .B0(ori_ori_n1596_), .B1(ori_ori_n2538_), .Y(ori_ori_n2541_));
  AOI210     o2492(.A0(ori_ori_n2537_), .A1(ori_ori_n68_), .B0(ori_ori_n2541_), .Y(ori_ori_n2542_));
  OAI210     o2493(.A0(ori_ori_n268_), .A1(ori_ori_n1089_), .B0(ori_ori_n486_), .Y(ori_ori_n2543_));
  NA3        o2494(.A(ori_ori_n2543_), .B(ori_ori_n264_), .C(ori_ori_n1042_), .Y(ori_ori_n2544_));
  OAI210     o2495(.A0(ori_ori_n228_), .A1(ori_ori_n216_), .B0(ori_ori_n1712_), .Y(ori_ori_n2545_));
  NA2        o2496(.A(ori_ori_n345_), .B(ori_ori_n272_), .Y(ori_ori_n2546_));
  NA3        o2497(.A(ori_ori_n401_), .B(ori_ori_n813_), .C(ori_ori_n106_), .Y(ori_ori_n2547_));
  NO2        o2498(.A(ori_ori_n530_), .B(ori_ori_n56_), .Y(ori_ori_n2548_));
  NA3        o2499(.A(ori_ori_n2548_), .B(ori_ori_n2547_), .C(ori_ori_n2546_), .Y(ori_ori_n2549_));
  AOI210     o2500(.A0(ori_ori_n2545_), .A1(ori_ori_n511_), .B0(ori_ori_n2549_), .Y(ori_ori_n2550_));
  NO2        o2501(.A(ori_ori_n1175_), .B(ori_ori_n273_), .Y(ori_ori_n2551_));
  OAI210     o2502(.A0(ori_ori_n293_), .A1(ori_ori_n262_), .B0(ori_ori_n2551_), .Y(ori_ori_n2552_));
  OAI210     o2503(.A0(ori_ori_n666_), .A1(ori_ori_n137_), .B0(x3), .Y(ori_ori_n2553_));
  AOI210     o2504(.A0(ori_ori_n666_), .A1(ori_ori_n363_), .B0(ori_ori_n2553_), .Y(ori_ori_n2554_));
  AOI210     o2505(.A0(ori_ori_n1595_), .A1(ori_ori_n50_), .B0(ori_ori_n345_), .Y(ori_ori_n2555_));
  OAI210     o2506(.A0(ori_ori_n2555_), .A1(ori_ori_n400_), .B0(ori_ori_n56_), .Y(ori_ori_n2556_));
  NO2        o2507(.A(ori_ori_n2556_), .B(ori_ori_n2554_), .Y(ori_ori_n2557_));
  AOI220     o2508(.A0(ori_ori_n2557_), .A1(ori_ori_n2552_), .B0(ori_ori_n2550_), .B1(ori_ori_n2544_), .Y(ori_ori_n2558_));
  OAI210     o2509(.A0(ori_ori_n2558_), .A1(ori_ori_n1751_), .B0(ori_ori_n98_), .Y(ori_ori_n2559_));
  NA2        o2510(.A(ori_ori_n692_), .B(ori_ori_n1189_), .Y(ori_ori_n2560_));
  NOi21      o2511(.An(ori_ori_n1352_), .B(ori_ori_n107_), .Y(ori_ori_n2561_));
  NA2        o2512(.A(ori_ori_n2561_), .B(ori_ori_n2560_), .Y(ori_ori_n2562_));
  NO2        o2513(.A(ori_ori_n2214_), .B(ori_ori_n55_), .Y(ori_ori_n2563_));
  OAI210     o2514(.A0(ori_ori_n2563_), .A1(ori_ori_n2562_), .B0(ori_ori_n1808_), .Y(ori_ori_n2564_));
  NA2        o2515(.A(ori_ori_n176_), .B(ori_ori_n104_), .Y(ori_ori_n2565_));
  NA2        o2516(.A(ori_ori_n684_), .B(x6), .Y(ori_ori_n2566_));
  AOI210     o2517(.A0(ori_ori_n2566_), .A1(ori_ori_n485_), .B0(ori_ori_n2565_), .Y(ori_ori_n2567_));
  AOI210     o2518(.A0(ori_ori_n352_), .A1(ori_ori_n139_), .B0(ori_ori_n140_), .Y(ori_ori_n2568_));
  OAI210     o2519(.A0(ori_ori_n2568_), .A1(ori_ori_n2567_), .B0(ori_ori_n345_), .Y(ori_ori_n2569_));
  AOI210     o2520(.A0(ori_ori_n615_), .A1(ori_ori_n433_), .B0(ori_ori_n1280_), .Y(ori_ori_n2570_));
  NO3        o2521(.A(ori_ori_n2570_), .B(ori_ori_n264_), .C(ori_ori_n63_), .Y(ori_ori_n2571_));
  OAI220     o2522(.A0(ori_ori_n2330_), .A1(ori_ori_n483_), .B0(ori_ori_n2084_), .B1(ori_ori_n384_), .Y(ori_ori_n2572_));
  OAI210     o2523(.A0(ori_ori_n2572_), .A1(ori_ori_n2571_), .B0(ori_ori_n53_), .Y(ori_ori_n2573_));
  NO4        o2524(.A(ori_ori_n2340_), .B(ori_ori_n929_), .C(ori_ori_n434_), .D(ori_ori_n219_), .Y(ori_ori_n2574_));
  NO4        o2525(.A(ori_ori_n727_), .B(ori_ori_n603_), .C(ori_ori_n442_), .D(ori_ori_n1050_), .Y(ori_ori_n2575_));
  NO3        o2526(.A(ori_ori_n2575_), .B(ori_ori_n2574_), .C(ori_ori_n1056_), .Y(ori_ori_n2576_));
  NA4        o2527(.A(ori_ori_n2576_), .B(ori_ori_n2573_), .C(ori_ori_n2569_), .D(ori_ori_n2564_), .Y(ori_ori_n2577_));
  NO3        o2528(.A(ori_ori_n248_), .B(ori_ori_n351_), .C(ori_ori_n84_), .Y(ori_ori_n2578_));
  NO2        o2529(.A(ori_ori_n276_), .B(ori_ori_n768_), .Y(ori_ori_n2579_));
  NO3        o2530(.A(ori_ori_n2579_), .B(ori_ori_n1204_), .C(ori_ori_n1222_), .Y(ori_ori_n2580_));
  OAI220     o2531(.A0(ori_ori_n2580_), .A1(ori_ori_n2578_), .B0(ori_ori_n465_), .B1(ori_ori_n85_), .Y(ori_ori_n2581_));
  OR2        o2532(.A(ori_ori_n935_), .B(ori_ori_n745_), .Y(ori_ori_n2582_));
  NA2        o2533(.A(ori_ori_n1217_), .B(ori_ori_n55_), .Y(ori_ori_n2583_));
  NOi21      o2534(.An(ori_ori_n2583_), .B(ori_ori_n385_), .Y(ori_ori_n2584_));
  AOI210     o2535(.A0(ori_ori_n2584_), .A1(ori_ori_n2582_), .B0(x1), .Y(ori_ori_n2585_));
  NA2        o2536(.A(ori_ori_n263_), .B(ori_ori_n84_), .Y(ori_ori_n2586_));
  AOI210     o2537(.A0(ori_ori_n1547_), .A1(ori_ori_n400_), .B0(ori_ori_n2586_), .Y(ori_ori_n2587_));
  NA2        o2538(.A(ori_ori_n1101_), .B(ori_ori_n62_), .Y(ori_ori_n2588_));
  NA2        o2539(.A(ori_ori_n1149_), .B(ori_ori_n172_), .Y(ori_ori_n2589_));
  OAI210     o2540(.A0(ori_ori_n2588_), .A1(ori_ori_n311_), .B0(ori_ori_n2589_), .Y(ori_ori_n2590_));
  NO3        o2541(.A(ori_ori_n2590_), .B(ori_ori_n2587_), .C(ori_ori_n2585_), .Y(ori_ori_n2591_));
  OAI210     o2542(.A0(ori_ori_n2591_), .A1(x6), .B0(ori_ori_n2581_), .Y(ori_ori_n2592_));
  AOI220     o2543(.A0(ori_ori_n2592_), .A1(ori_ori_n1455_), .B0(ori_ori_n2577_), .B1(ori_ori_n57_), .Y(ori_ori_n2593_));
  NA3        o2544(.A(ori_ori_n2593_), .B(ori_ori_n2559_), .C(ori_ori_n2542_), .Y(ori38));
  NO2        o2545(.A(ori_ori_n184_), .B(ori_ori_n967_), .Y(ori_ori_n2595_));
  AOI210     o2546(.A0(ori_ori_n1221_), .A1(ori_ori_n579_), .B0(ori_ori_n1082_), .Y(ori_ori_n2596_));
  AOI210     o2547(.A0(ori_ori_n2583_), .A1(ori_ori_n1840_), .B0(ori_ori_n227_), .Y(ori_ori_n2597_));
  NO3        o2548(.A(ori_ori_n1290_), .B(ori_ori_n317_), .C(x8), .Y(ori_ori_n2598_));
  NO4        o2549(.A(ori_ori_n2598_), .B(ori_ori_n2597_), .C(ori_ori_n2596_), .D(ori_ori_n2595_), .Y(ori_ori_n2599_));
  NO2        o2550(.A(ori_ori_n2599_), .B(x6), .Y(ori_ori_n2600_));
  NA4        o2551(.A(ori_ori_n376_), .B(ori_ori_n255_), .C(ori_ori_n187_), .D(x8), .Y(ori_ori_n2601_));
  NA2        o2552(.A(ori_ori_n399_), .B(ori_ori_n104_), .Y(ori_ori_n2602_));
  AOI210     o2553(.A0(ori_ori_n2602_), .A1(ori_ori_n2601_), .B0(ori_ori_n140_), .Y(ori_ori_n2603_));
  AOI210     o2554(.A0(ori_ori_n434_), .A1(ori_ori_n404_), .B0(ori_ori_n1722_), .Y(ori_ori_n2604_));
  NO2        o2555(.A(ori_ori_n807_), .B(ori_ori_n90_), .Y(ori_ori_n2605_));
  OAI210     o2556(.A0(ori_ori_n1017_), .A1(ori_ori_n147_), .B0(ori_ori_n358_), .Y(ori_ori_n2606_));
  OAI220     o2557(.A0(ori_ori_n2606_), .A1(ori_ori_n2605_), .B0(ori_ori_n2604_), .B1(ori_ori_n187_), .Y(ori_ori_n2607_));
  OAI210     o2558(.A0(ori_ori_n2607_), .A1(ori_ori_n2603_), .B0(x6), .Y(ori_ori_n2608_));
  NO2        o2559(.A(ori_ori_n245_), .B(ori_ori_n768_), .Y(ori_ori_n2609_));
  NO3        o2560(.A(ori_ori_n2609_), .B(ori_ori_n1677_), .C(ori_ori_n255_), .Y(ori_ori_n2610_));
  NO3        o2561(.A(x3), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n2611_));
  OAI210     o2562(.A0(ori_ori_n523_), .A1(x2), .B0(ori_ori_n2611_), .Y(ori_ori_n2612_));
  NA3        o2563(.A(ori_ori_n433_), .B(ori_ori_n423_), .C(ori_ori_n292_), .Y(ori_ori_n2613_));
  NA3        o2564(.A(ori_ori_n2613_), .B(ori_ori_n2612_), .C(ori_ori_n1800_), .Y(ori_ori_n2614_));
  OAI210     o2565(.A0(ori_ori_n2614_), .A1(ori_ori_n2610_), .B0(ori_ori_n809_), .Y(ori_ori_n2615_));
  AN3        o2566(.A(ori_ori_n814_), .B(ori_ori_n777_), .C(x0), .Y(ori_ori_n2616_));
  NA2        o2567(.A(ori_ori_n2616_), .B(ori_ori_n326_), .Y(ori_ori_n2617_));
  OAI220     o2568(.A0(ori_ori_n603_), .A1(ori_ori_n274_), .B0(ori_ori_n813_), .B1(ori_ori_n91_), .Y(ori_ori_n2618_));
  OAI210     o2569(.A0(ori_ori_n684_), .A1(x0), .B0(ori_ori_n51_), .Y(ori_ori_n2619_));
  AOI210     o2570(.A0(ori_ori_n584_), .A1(x4), .B0(ori_ori_n226_), .Y(ori_ori_n2620_));
  AOI220     o2571(.A0(ori_ori_n2620_), .A1(ori_ori_n2619_), .B0(ori_ori_n2618_), .B1(ori_ori_n401_), .Y(ori_ori_n2621_));
  NA4        o2572(.A(ori_ori_n2621_), .B(ori_ori_n2617_), .C(ori_ori_n2615_), .D(ori_ori_n2608_), .Y(ori_ori_n2622_));
  OAI210     o2573(.A0(ori_ori_n2622_), .A1(ori_ori_n2600_), .B0(x7), .Y(ori_ori_n2623_));
  AOI210     o2574(.A0(ori_ori_n372_), .A1(x1), .B0(ori_ori_n1228_), .Y(ori_ori_n2624_));
  NO2        o2575(.A(ori_ori_n2624_), .B(ori_ori_n51_), .Y(ori_ori_n2625_));
  AOI210     o2576(.A0(ori_ori_n90_), .A1(ori_ori_n71_), .B0(ori_ori_n2241_), .Y(ori_ori_n2626_));
  NA2        o2577(.A(ori_ori_n384_), .B(x3), .Y(ori_ori_n2627_));
  NO2        o2578(.A(ori_ori_n1743_), .B(ori_ori_n530_), .Y(ori_ori_n2628_));
  OAI210     o2579(.A0(ori_ori_n2627_), .A1(ori_ori_n2626_), .B0(ori_ori_n2628_), .Y(ori_ori_n2629_));
  OAI210     o2580(.A0(ori_ori_n2629_), .A1(ori_ori_n2625_), .B0(x4), .Y(ori_ori_n2630_));
  INV        o2581(.A(ori_ori_n459_), .Y(ori_ori_n2631_));
  NO3        o2582(.A(ori_ori_n2631_), .B(ori_ori_n400_), .C(ori_ori_n117_), .Y(ori_ori_n2632_));
  AOI210     o2583(.A0(ori_ori_n1050_), .A1(ori_ori_n239_), .B0(ori_ori_n393_), .Y(ori_ori_n2633_));
  AO210      o2584(.A0(ori_ori_n1295_), .A1(x6), .B0(ori_ori_n2633_), .Y(ori_ori_n2634_));
  NO2        o2585(.A(ori_ori_n1408_), .B(ori_ori_n137_), .Y(ori_ori_n2635_));
  NA2        o2586(.A(ori_ori_n1945_), .B(ori_ori_n320_), .Y(ori_ori_n2636_));
  OAI220     o2587(.A0(ori_ori_n2636_), .A1(ori_ori_n1069_), .B0(ori_ori_n2635_), .B1(ori_ori_n1822_), .Y(ori_ori_n2637_));
  NO3        o2588(.A(ori_ori_n2637_), .B(ori_ori_n2634_), .C(ori_ori_n2632_), .Y(ori_ori_n2638_));
  AOI210     o2589(.A0(ori_ori_n2638_), .A1(ori_ori_n2630_), .B0(ori_ori_n104_), .Y(ori_ori_n2639_));
  NA3        o2590(.A(ori_ori_n1935_), .B(ori_ori_n603_), .C(ori_ori_n163_), .Y(ori_ori_n2640_));
  AOI210     o2591(.A0(ori_ori_n2640_), .A1(ori_ori_n1418_), .B0(ori_ori_n228_), .Y(ori_ori_n2641_));
  AOI210     o2592(.A0(ori_ori_n504_), .A1(ori_ori_n492_), .B0(ori_ori_n680_), .Y(ori_ori_n2642_));
  OAI220     o2593(.A0(ori_ori_n2642_), .A1(ori_ori_n466_), .B0(ori_ori_n195_), .B1(ori_ori_n115_), .Y(ori_ori_n2643_));
  OAI210     o2594(.A0(ori_ori_n2643_), .A1(ori_ori_n2641_), .B0(x0), .Y(ori_ori_n2644_));
  NA3        o2595(.A(ori_ori_n404_), .B(ori_ori_n813_), .C(ori_ori_n274_), .Y(ori_ori_n2645_));
  AOI210     o2596(.A0(ori_ori_n2645_), .A1(ori_ori_n714_), .B0(ori_ori_n2198_), .Y(ori_ori_n2646_));
  NA2        o2597(.A(ori_ori_n1121_), .B(ori_ori_n948_), .Y(ori_ori_n2647_));
  NA4        o2598(.A(ori_ori_n679_), .B(ori_ori_n603_), .C(ori_ori_n176_), .D(x3), .Y(ori_ori_n2648_));
  AOI210     o2599(.A0(ori_ori_n2648_), .A1(ori_ori_n2647_), .B0(ori_ori_n498_), .Y(ori_ori_n2649_));
  NO4        o2600(.A(ori_ori_n1401_), .B(ori_ori_n519_), .C(ori_ori_n1222_), .D(ori_ori_n768_), .Y(ori_ori_n2650_));
  OAI220     o2601(.A0(ori_ori_n1771_), .A1(ori_ori_n2285_), .B0(ori_ori_n226_), .B1(ori_ori_n149_), .Y(ori_ori_n2651_));
  NO4        o2602(.A(ori_ori_n2651_), .B(ori_ori_n2650_), .C(ori_ori_n2649_), .D(ori_ori_n2646_), .Y(ori_ori_n2652_));
  NA2        o2603(.A(ori_ori_n2652_), .B(ori_ori_n2644_), .Y(ori_ori_n2653_));
  OAI210     o2604(.A0(ori_ori_n2653_), .A1(ori_ori_n2639_), .B0(ori_ori_n57_), .Y(ori_ori_n2654_));
  NO2        o2605(.A(ori_ori_n1809_), .B(ori_ori_n681_), .Y(ori_ori_n2655_));
  OAI210     o2606(.A0(ori_ori_n1750_), .A1(ori_ori_n211_), .B0(ori_ori_n494_), .Y(ori_ori_n2656_));
  OAI210     o2607(.A0(ori_ori_n2656_), .A1(ori_ori_n2655_), .B0(ori_ori_n630_), .Y(ori_ori_n2657_));
  OAI220     o2608(.A0(ori_ori_n1756_), .A1(ori_ori_n274_), .B0(ori_ori_n254_), .B1(ori_ori_n100_), .Y(ori_ori_n2658_));
  NA2        o2609(.A(ori_ori_n1859_), .B(ori_ori_n353_), .Y(ori_ori_n2659_));
  OAI220     o2610(.A0(ori_ori_n2659_), .A1(ori_ori_n636_), .B0(ori_ori_n691_), .B1(ori_ori_n149_), .Y(ori_ori_n2660_));
  AOI210     o2611(.A0(ori_ori_n2658_), .A1(ori_ori_n987_), .B0(ori_ori_n2660_), .Y(ori_ori_n2661_));
  NA4        o2612(.A(ori_ori_n2661_), .B(ori_ori_n2657_), .C(ori_ori_n2654_), .D(ori_ori_n2623_), .Y(ori39));
  INV        m0000(.A(x3), .Y(mai_mai_n50_));
  NA2        m0001(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n51_));
  NA2        m0002(.A(x7), .B(x0), .Y(mai_mai_n52_));
  INV        m0003(.A(x1), .Y(mai_mai_n53_));
  NA2        m0004(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  INV        m0005(.A(x8), .Y(mai_mai_n55_));
  INV        m0006(.A(x4), .Y(mai_mai_n56_));
  INV        m0007(.A(x7), .Y(mai_mai_n57_));
  NA2        m0008(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0009(.A(x0), .Y(mai_mai_n59_));
  NA2        m0010(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n60_));
  NA4        m0011(.A(mai_mai_n60_), .B(mai_mai_n58_), .C(mai_mai_n55_), .D(x6), .Y(mai_mai_n61_));
  NA2        m0012(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n62_));
  NO2        m0013(.A(mai_mai_n55_), .B(x6), .Y(mai_mai_n63_));
  NA2        m0014(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n64_));
  NA3        m0015(.A(mai_mai_n64_), .B(mai_mai_n63_), .C(mai_mai_n62_), .Y(mai_mai_n65_));
  AOI210     m0016(.A0(mai_mai_n65_), .A1(mai_mai_n61_), .B0(mai_mai_n54_), .Y(mai_mai_n66_));
  NO2        m0017(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n67_));
  NO2        m0018(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n68_));
  NO2        m0019(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NAi21      m0020(.An(x5), .B(x1), .Y(mai_mai_n70_));
  INV        m0021(.A(x6), .Y(mai_mai_n71_));
  NA2        m0022(.A(mai_mai_n71_), .B(x4), .Y(mai_mai_n72_));
  NO3        m0023(.A(mai_mai_n72_), .B(mai_mai_n70_), .C(mai_mai_n69_), .Y(mai_mai_n73_));
  OAI210     m0024(.A0(mai_mai_n73_), .A1(mai_mai_n66_), .B0(mai_mai_n52_), .Y(mai_mai_n74_));
  NA2        m0025(.A(x7), .B(x4), .Y(mai_mai_n75_));
  NO2        m0026(.A(mai_mai_n75_), .B(x1), .Y(mai_mai_n76_));
  NO2        m0027(.A(mai_mai_n71_), .B(x5), .Y(mai_mai_n77_));
  NO2        m0028(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n78_));
  NA3        m0029(.A(mai_mai_n78_), .B(mai_mai_n77_), .C(mai_mai_n76_), .Y(mai_mai_n79_));
  AOI210     m0030(.A0(mai_mai_n79_), .A1(mai_mai_n74_), .B0(mai_mai_n51_), .Y(mai_mai_n80_));
  NA2        m0031(.A(x5), .B(x3), .Y(mai_mai_n81_));
  NO2        m0032(.A(x6), .B(x0), .Y(mai_mai_n82_));
  NO2        m0033(.A(mai_mai_n82_), .B(x4), .Y(mai_mai_n83_));
  NO2        m0034(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m0035(.A(mai_mai_n71_), .B(mai_mai_n59_), .Y(mai_mai_n85_));
  NO2        m0036(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n86_));
  NA2        m0037(.A(x8), .B(x1), .Y(mai_mai_n87_));
  NO2        m0038(.A(mai_mai_n87_), .B(x7), .Y(mai_mai_n88_));
  INV        m0039(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OR3        m0040(.A(mai_mai_n89_), .B(mai_mai_n86_), .C(mai_mai_n83_), .Y(mai_mai_n90_));
  NO3        m0041(.A(x8), .B(mai_mai_n57_), .C(x6), .Y(mai_mai_n91_));
  NO2        m0042(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n92_));
  NO2        m0043(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n93_));
  NA3        m0044(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n94_));
  AOI210     m0045(.A0(mai_mai_n94_), .A1(mai_mai_n90_), .B0(mai_mai_n81_), .Y(mai_mai_n95_));
  XO2        m0046(.A(x7), .B(x1), .Y(mai_mai_n96_));
  INV        m0047(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NO2        m0048(.A(mai_mai_n97_), .B(x6), .Y(mai_mai_n98_));
  NO2        m0049(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n99_));
  NA2        m0050(.A(mai_mai_n99_), .B(mai_mai_n55_), .Y(mai_mai_n100_));
  NO2        m0051(.A(x6), .B(x5), .Y(mai_mai_n101_));
  NO2        m0052(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n102_));
  NO2        m0053(.A(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  NA2        m0054(.A(x6), .B(x1), .Y(mai_mai_n104_));
  NA2        m0055(.A(mai_mai_n104_), .B(mai_mai_n84_), .Y(mai_mai_n105_));
  NO4        m0056(.A(mai_mai_n105_), .B(mai_mai_n103_), .C(mai_mai_n100_), .D(mai_mai_n98_), .Y(mai_mai_n106_));
  NA2        m0057(.A(x3), .B(x0), .Y(mai_mai_n107_));
  INV        m0058(.A(x5), .Y(mai_mai_n108_));
  NA2        m0059(.A(mai_mai_n71_), .B(mai_mai_n108_), .Y(mai_mai_n109_));
  INV        m0060(.A(x2), .Y(mai_mai_n110_));
  NO2        m0061(.A(mai_mai_n56_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  NA2        m0062(.A(mai_mai_n57_), .B(mai_mai_n108_), .Y(mai_mai_n112_));
  NA3        m0063(.A(mai_mai_n112_), .B(mai_mai_n111_), .C(mai_mai_n109_), .Y(mai_mai_n113_));
  NO3        m0064(.A(mai_mai_n113_), .B(mai_mai_n107_), .C(mai_mai_n53_), .Y(mai_mai_n114_));
  NO4        m0065(.A(mai_mai_n114_), .B(mai_mai_n106_), .C(mai_mai_n95_), .D(mai_mai_n80_), .Y(mai00));
  NO2        m0066(.A(x7), .B(x6), .Y(mai_mai_n116_));
  INV        m0067(.A(mai_mai_n116_), .Y(mai_mai_n117_));
  NO2        m0068(.A(mai_mai_n55_), .B(mai_mai_n53_), .Y(mai_mai_n118_));
  NA2        m0069(.A(mai_mai_n118_), .B(mai_mai_n56_), .Y(mai_mai_n119_));
  NO2        m0070(.A(mai_mai_n119_), .B(mai_mai_n117_), .Y(mai_mai_n120_));
  XN2        m0071(.A(x6), .B(x1), .Y(mai_mai_n121_));
  INV        m0072(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  NO2        m0073(.A(x6), .B(x4), .Y(mai_mai_n123_));
  NA2        m0074(.A(x6), .B(x4), .Y(mai_mai_n124_));
  NAi21      m0075(.An(mai_mai_n123_), .B(mai_mai_n124_), .Y(mai_mai_n125_));
  XN2        m0076(.A(x7), .B(x6), .Y(mai_mai_n126_));
  NO4        m0077(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n122_), .D(x8), .Y(mai_mai_n127_));
  NO2        m0078(.A(x3), .B(mai_mai_n110_), .Y(mai_mai_n128_));
  NA2        m0079(.A(mai_mai_n128_), .B(mai_mai_n108_), .Y(mai_mai_n129_));
  NO2        m0080(.A(mai_mai_n129_), .B(mai_mai_n59_), .Y(mai_mai_n130_));
  OAI210     m0081(.A0(mai_mai_n127_), .A1(mai_mai_n120_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NA2        m0082(.A(x3), .B(mai_mai_n110_), .Y(mai_mai_n132_));
  NO2        m0083(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n133_));
  NA2        m0084(.A(mai_mai_n133_), .B(mai_mai_n56_), .Y(mai_mai_n134_));
  NA2        m0085(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n135_));
  NA2        m0086(.A(mai_mai_n135_), .B(x2), .Y(mai_mai_n136_));
  NA2        m0087(.A(x8), .B(x3), .Y(mai_mai_n137_));
  NA2        m0088(.A(mai_mai_n137_), .B(mai_mai_n75_), .Y(mai_mai_n138_));
  OAI220     m0089(.A0(mai_mai_n138_), .A1(mai_mai_n136_), .B0(mai_mai_n134_), .B1(mai_mai_n132_), .Y(mai_mai_n139_));
  NO2        m0090(.A(x5), .B(x0), .Y(mai_mai_n140_));
  NO2        m0091(.A(x6), .B(x1), .Y(mai_mai_n141_));
  NA3        m0092(.A(mai_mai_n141_), .B(mai_mai_n140_), .C(mai_mai_n139_), .Y(mai_mai_n142_));
  NA2        m0093(.A(x8), .B(mai_mai_n108_), .Y(mai_mai_n143_));
  NA2        m0094(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n144_));
  NAi21      m0095(.An(x7), .B(x2), .Y(mai_mai_n145_));
  XO2        m0096(.A(x8), .B(x7), .Y(mai_mai_n146_));
  NA2        m0097(.A(mai_mai_n146_), .B(mai_mai_n110_), .Y(mai_mai_n147_));
  NA2        m0098(.A(x6), .B(x5), .Y(mai_mai_n148_));
  NO2        m0099(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n149_));
  NO2        m0100(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n150_));
  NA2        m0101(.A(mai_mai_n150_), .B(mai_mai_n149_), .Y(mai_mai_n151_));
  NO3        m0102(.A(mai_mai_n151_), .B(mai_mai_n148_), .C(mai_mai_n147_), .Y(mai_mai_n152_));
  INV        m0103(.A(mai_mai_n152_), .Y(mai_mai_n153_));
  NA3        m0104(.A(mai_mai_n153_), .B(mai_mai_n142_), .C(mai_mai_n131_), .Y(mai01));
  NA2        m0105(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n155_));
  NO2        m0106(.A(x2), .B(x1), .Y(mai_mai_n156_));
  NA2        m0107(.A(x2), .B(x1), .Y(mai_mai_n157_));
  NOi21      m0108(.An(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  NA2        m0109(.A(mai_mai_n108_), .B(mai_mai_n53_), .Y(mai_mai_n159_));
  NO2        m0110(.A(mai_mai_n159_), .B(x8), .Y(mai_mai_n160_));
  NAi21      m0111(.An(x8), .B(x1), .Y(mai_mai_n161_));
  NO2        m0112(.A(mai_mai_n161_), .B(x3), .Y(mai_mai_n162_));
  OAI210     m0113(.A0(mai_mai_n162_), .A1(mai_mai_n160_), .B0(mai_mai_n158_), .Y(mai_mai_n163_));
  NO2        m0114(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n164_));
  NO2        m0115(.A(mai_mai_n110_), .B(x1), .Y(mai_mai_n165_));
  NA2        m0116(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  AOI210     m0117(.A0(mai_mai_n166_), .A1(mai_mai_n163_), .B0(mai_mai_n155_), .Y(mai_mai_n167_));
  NAi21      m0118(.An(x7), .B(x0), .Y(mai_mai_n168_));
  NO2        m0119(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n169_));
  NO2        m0120(.A(mai_mai_n81_), .B(x1), .Y(mai_mai_n170_));
  NA2        m0121(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  NA2        m0122(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n172_));
  NO2        m0123(.A(mai_mai_n172_), .B(mai_mai_n161_), .Y(mai_mai_n173_));
  NA2        m0124(.A(x8), .B(x5), .Y(mai_mai_n174_));
  NO2        m0125(.A(mai_mai_n174_), .B(mai_mai_n51_), .Y(mai_mai_n175_));
  NO3        m0126(.A(x3), .B(mai_mai_n110_), .C(mai_mai_n53_), .Y(mai_mai_n176_));
  NO3        m0127(.A(mai_mai_n176_), .B(mai_mai_n175_), .C(mai_mai_n173_), .Y(mai_mai_n177_));
  AOI210     m0128(.A0(mai_mai_n177_), .A1(mai_mai_n171_), .B0(mai_mai_n168_), .Y(mai_mai_n178_));
  NO2        m0129(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n179_));
  NO2        m0130(.A(mai_mai_n55_), .B(x0), .Y(mai_mai_n180_));
  NA3        m0131(.A(mai_mai_n108_), .B(mai_mai_n110_), .C(x1), .Y(mai_mai_n181_));
  NO2        m0132(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NO2        m0133(.A(mai_mai_n87_), .B(mai_mai_n50_), .Y(mai_mai_n183_));
  NA2        m0134(.A(mai_mai_n108_), .B(x0), .Y(mai_mai_n184_));
  NO2        m0135(.A(mai_mai_n184_), .B(x2), .Y(mai_mai_n185_));
  AOI220     m0136(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(mai_mai_n182_), .B1(mai_mai_n179_), .Y(mai_mai_n186_));
  NA2        m0137(.A(x7), .B(mai_mai_n110_), .Y(mai_mai_n187_));
  NA2        m0138(.A(mai_mai_n164_), .B(x8), .Y(mai_mai_n188_));
  NA4        m0139(.A(x5), .B(x3), .C(x1), .D(x0), .Y(mai_mai_n189_));
  AO210      m0140(.A0(mai_mai_n189_), .A1(mai_mai_n188_), .B0(mai_mai_n187_), .Y(mai_mai_n190_));
  NO2        m0141(.A(mai_mai_n157_), .B(mai_mai_n50_), .Y(mai_mai_n191_));
  NAi21      m0142(.An(x1), .B(x2), .Y(mai_mai_n192_));
  NO2        m0143(.A(mai_mai_n172_), .B(mai_mai_n192_), .Y(mai_mai_n193_));
  NA2        m0144(.A(x8), .B(x7), .Y(mai_mai_n194_));
  NO2        m0145(.A(mai_mai_n194_), .B(x0), .Y(mai_mai_n195_));
  OAI210     m0146(.A0(mai_mai_n193_), .A1(mai_mai_n191_), .B0(mai_mai_n195_), .Y(mai_mai_n196_));
  NA3        m0147(.A(mai_mai_n196_), .B(mai_mai_n190_), .C(mai_mai_n186_), .Y(mai_mai_n197_));
  NO3        m0148(.A(mai_mai_n197_), .B(mai_mai_n178_), .C(mai_mai_n167_), .Y(mai_mai_n198_));
  NA2        m0149(.A(x3), .B(x1), .Y(mai_mai_n199_));
  NA2        m0150(.A(mai_mai_n50_), .B(mai_mai_n110_), .Y(mai_mai_n200_));
  NO2        m0151(.A(mai_mai_n200_), .B(mai_mai_n70_), .Y(mai_mai_n201_));
  OAI210     m0152(.A0(mai_mai_n201_), .A1(mai_mai_n193_), .B0(mai_mai_n67_), .Y(mai_mai_n202_));
  NA2        m0153(.A(mai_mai_n133_), .B(mai_mai_n110_), .Y(mai_mai_n203_));
  OAI210     m0154(.A0(mai_mai_n203_), .A1(mai_mai_n199_), .B0(mai_mai_n202_), .Y(mai_mai_n204_));
  XO2        m0155(.A(x5), .B(x3), .Y(mai_mai_n205_));
  NA2        m0156(.A(mai_mai_n205_), .B(x8), .Y(mai_mai_n206_));
  NA2        m0157(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n207_));
  NA2        m0158(.A(mai_mai_n207_), .B(mai_mai_n137_), .Y(mai_mai_n208_));
  NA2        m0159(.A(x7), .B(mai_mai_n71_), .Y(mai_mai_n209_));
  NO2        m0160(.A(mai_mai_n192_), .B(mai_mai_n209_), .Y(mai_mai_n210_));
  OA210      m0161(.A0(mai_mai_n208_), .A1(mai_mai_n205_), .B0(mai_mai_n210_), .Y(mai_mai_n211_));
  AOI220     m0162(.A0(mai_mai_n211_), .A1(mai_mai_n206_), .B0(mai_mai_n204_), .B1(x0), .Y(mai_mai_n212_));
  OAI210     m0163(.A0(mai_mai_n198_), .A1(mai_mai_n71_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  NO2        m0164(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n214_));
  NA4        m0165(.A(mai_mai_n55_), .B(x5), .C(x3), .D(x2), .Y(mai_mai_n215_));
  NA2        m0166(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n216_));
  NA2        m0167(.A(mai_mai_n216_), .B(x2), .Y(mai_mai_n217_));
  NA2        m0168(.A(mai_mai_n55_), .B(x3), .Y(mai_mai_n218_));
  NA4        m0169(.A(mai_mai_n218_), .B(mai_mai_n217_), .C(mai_mai_n205_), .D(mai_mai_n82_), .Y(mai_mai_n219_));
  AOI210     m0170(.A0(mai_mai_n219_), .A1(mai_mai_n215_), .B0(mai_mai_n53_), .Y(mai_mai_n220_));
  NO2        m0171(.A(mai_mai_n110_), .B(mai_mai_n59_), .Y(mai_mai_n221_));
  NA2        m0172(.A(x5), .B(x1), .Y(mai_mai_n222_));
  NO2        m0173(.A(mai_mai_n222_), .B(x6), .Y(mai_mai_n223_));
  NO2        m0174(.A(x3), .B(x1), .Y(mai_mai_n224_));
  AOI210     m0175(.A0(mai_mai_n224_), .A1(mai_mai_n77_), .B0(mai_mai_n223_), .Y(mai_mai_n225_));
  NO2        m0176(.A(mai_mai_n81_), .B(mai_mai_n55_), .Y(mai_mai_n226_));
  NO2        m0177(.A(mai_mai_n104_), .B(mai_mai_n50_), .Y(mai_mai_n227_));
  NO2        m0178(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  OAI210     m0179(.A0(mai_mai_n225_), .A1(x8), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  NO2        m0180(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n230_));
  NA2        m0181(.A(mai_mai_n230_), .B(mai_mai_n71_), .Y(mai_mai_n231_));
  NAi21      m0182(.An(x2), .B(x5), .Y(mai_mai_n232_));
  NA2        m0183(.A(x8), .B(x6), .Y(mai_mai_n233_));
  OAI210     m0184(.A0(mai_mai_n233_), .A1(mai_mai_n232_), .B0(mai_mai_n231_), .Y(mai_mai_n234_));
  NA2        m0185(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n235_));
  NO2        m0186(.A(mai_mai_n235_), .B(mai_mai_n59_), .Y(mai_mai_n236_));
  AO220      m0187(.A0(mai_mai_n236_), .A1(mai_mai_n234_), .B0(mai_mai_n229_), .B1(mai_mai_n221_), .Y(mai_mai_n237_));
  OAI210     m0188(.A0(mai_mai_n237_), .A1(mai_mai_n220_), .B0(mai_mai_n214_), .Y(mai_mai_n238_));
  NA2        m0189(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n239_));
  NO2        m0190(.A(mai_mai_n239_), .B(x7), .Y(mai_mai_n240_));
  NO2        m0191(.A(mai_mai_n108_), .B(mai_mai_n53_), .Y(mai_mai_n241_));
  NA2        m0192(.A(mai_mai_n241_), .B(mai_mai_n110_), .Y(mai_mai_n242_));
  AOI210     m0193(.A0(mai_mai_n242_), .A1(mai_mai_n166_), .B0(mai_mai_n59_), .Y(mai_mai_n243_));
  NA2        m0194(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n244_));
  NO2        m0195(.A(mai_mai_n181_), .B(mai_mai_n244_), .Y(mai_mai_n245_));
  AN2        m0196(.A(mai_mai_n243_), .B(x8), .Y(mai_mai_n246_));
  NO2        m0197(.A(x1), .B(x0), .Y(mai_mai_n247_));
  NA2        m0198(.A(mai_mai_n247_), .B(mai_mai_n110_), .Y(mai_mai_n248_));
  NA2        m0199(.A(mai_mai_n108_), .B(mai_mai_n50_), .Y(mai_mai_n249_));
  XN2        m0200(.A(x3), .B(x2), .Y(mai_mai_n250_));
  NA2        m0201(.A(mai_mai_n250_), .B(mai_mai_n158_), .Y(mai_mai_n251_));
  NO2        m0202(.A(mai_mai_n108_), .B(x0), .Y(mai_mai_n252_));
  NA2        m0203(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n253_));
  NA2        m0204(.A(mai_mai_n253_), .B(mai_mai_n252_), .Y(mai_mai_n254_));
  OAI220     m0205(.A0(mai_mai_n254_), .A1(mai_mai_n251_), .B0(mai_mai_n249_), .B1(mai_mai_n248_), .Y(mai_mai_n255_));
  OAI210     m0206(.A0(mai_mai_n255_), .A1(mai_mai_n246_), .B0(mai_mai_n240_), .Y(mai_mai_n256_));
  NO2        m0207(.A(x7), .B(x1), .Y(mai_mai_n257_));
  NOi21      m0208(.An(x8), .B(x3), .Y(mai_mai_n258_));
  NA2        m0209(.A(mai_mai_n258_), .B(mai_mai_n59_), .Y(mai_mai_n259_));
  NA2        m0210(.A(x5), .B(x0), .Y(mai_mai_n260_));
  NAi21      m0211(.An(mai_mai_n140_), .B(mai_mai_n260_), .Y(mai_mai_n261_));
  NA2        m0212(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n262_));
  OAI210     m0213(.A0(mai_mai_n262_), .A1(mai_mai_n261_), .B0(mai_mai_n259_), .Y(mai_mai_n263_));
  NA3        m0214(.A(mai_mai_n263_), .B(mai_mai_n143_), .C(mai_mai_n257_), .Y(mai_mai_n264_));
  NA2        m0215(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n265_));
  NO2        m0216(.A(mai_mai_n265_), .B(x5), .Y(mai_mai_n266_));
  NO2        m0217(.A(mai_mai_n150_), .B(mai_mai_n71_), .Y(mai_mai_n267_));
  NA2        m0218(.A(x1), .B(x0), .Y(mai_mai_n268_));
  NA2        m0219(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n269_));
  NA3        m0220(.A(mai_mai_n268_), .B(mai_mai_n267_), .C(mai_mai_n266_), .Y(mai_mai_n270_));
  NA3        m0221(.A(mai_mai_n270_), .B(mai_mai_n264_), .C(mai_mai_n189_), .Y(mai_mai_n271_));
  NO2        m0222(.A(mai_mai_n108_), .B(x3), .Y(mai_mai_n272_));
  NO2        m0223(.A(mai_mai_n110_), .B(x0), .Y(mai_mai_n273_));
  NO2        m0224(.A(mai_mai_n55_), .B(x7), .Y(mai_mai_n274_));
  NO3        m0225(.A(x8), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n275_));
  NAi21      m0226(.An(x8), .B(x0), .Y(mai_mai_n276_));
  NAi21      m0227(.An(x1), .B(x3), .Y(mai_mai_n277_));
  NO2        m0228(.A(mai_mai_n277_), .B(mai_mai_n276_), .Y(mai_mai_n278_));
  NO2        m0229(.A(x2), .B(mai_mai_n53_), .Y(mai_mai_n279_));
  AOI210     m0230(.A0(mai_mai_n279_), .A1(mai_mai_n275_), .B0(mai_mai_n278_), .Y(mai_mai_n280_));
  NOi21      m0231(.An(x5), .B(x6), .Y(mai_mai_n281_));
  NO2        m0232(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n282_));
  NA2        m0233(.A(mai_mai_n282_), .B(mai_mai_n281_), .Y(mai_mai_n283_));
  NO2        m0234(.A(mai_mai_n283_), .B(mai_mai_n280_), .Y(mai_mai_n284_));
  AOI210     m0235(.A0(mai_mai_n271_), .A1(mai_mai_n111_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  NA3        m0236(.A(mai_mai_n285_), .B(mai_mai_n256_), .C(mai_mai_n238_), .Y(mai_mai_n286_));
  AOI210     m0237(.A0(mai_mai_n213_), .A1(mai_mai_n56_), .B0(mai_mai_n286_), .Y(mai02));
  NO2        m0238(.A(x8), .B(mai_mai_n108_), .Y(mai_mai_n288_));
  XN2        m0239(.A(x7), .B(x3), .Y(mai_mai_n289_));
  INV        m0240(.A(mai_mai_n289_), .Y(mai_mai_n290_));
  NO2        m0241(.A(x2), .B(x0), .Y(mai_mai_n291_));
  NA2        m0242(.A(mai_mai_n291_), .B(mai_mai_n71_), .Y(mai_mai_n292_));
  NO2        m0243(.A(mai_mai_n57_), .B(x1), .Y(mai_mai_n293_));
  NO3        m0244(.A(mai_mai_n293_), .B(mai_mai_n292_), .C(mai_mai_n290_), .Y(mai_mai_n294_));
  NA2        m0245(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n295_));
  NO2        m0246(.A(mai_mai_n277_), .B(x6), .Y(mai_mai_n296_));
  XO2        m0247(.A(x7), .B(x0), .Y(mai_mai_n297_));
  NO2        m0248(.A(mai_mai_n297_), .B(mai_mai_n291_), .Y(mai_mai_n298_));
  NA2        m0249(.A(mai_mai_n298_), .B(mai_mai_n296_), .Y(mai_mai_n299_));
  AN2        m0250(.A(x7), .B(x2), .Y(mai_mai_n300_));
  NA2        m0251(.A(mai_mai_n300_), .B(mai_mai_n50_), .Y(mai_mai_n301_));
  OAI210     m0252(.A0(mai_mai_n301_), .A1(mai_mai_n295_), .B0(mai_mai_n299_), .Y(mai_mai_n302_));
  OAI210     m0253(.A0(mai_mai_n302_), .A1(mai_mai_n294_), .B0(mai_mai_n288_), .Y(mai_mai_n303_));
  NAi21      m0254(.An(x8), .B(x6), .Y(mai_mai_n304_));
  NO2        m0255(.A(mai_mai_n108_), .B(mai_mai_n59_), .Y(mai_mai_n305_));
  NA2        m0256(.A(x7), .B(x3), .Y(mai_mai_n306_));
  NO2        m0257(.A(mai_mai_n306_), .B(x2), .Y(mai_mai_n307_));
  NA2        m0258(.A(x2), .B(x0), .Y(mai_mai_n308_));
  NA2        m0259(.A(mai_mai_n110_), .B(mai_mai_n59_), .Y(mai_mai_n309_));
  NA2        m0260(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  NAi21      m0261(.An(x7), .B(x1), .Y(mai_mai_n311_));
  NO2        m0262(.A(mai_mai_n311_), .B(x3), .Y(mai_mai_n312_));
  AOI220     m0263(.A0(mai_mai_n312_), .A1(mai_mai_n310_), .B0(mai_mai_n307_), .B1(mai_mai_n305_), .Y(mai_mai_n313_));
  NA2        m0264(.A(mai_mai_n279_), .B(mai_mai_n50_), .Y(mai_mai_n314_));
  NA3        m0265(.A(x7), .B(mai_mai_n108_), .C(x0), .Y(mai_mai_n315_));
  NA2        m0266(.A(mai_mai_n273_), .B(mai_mai_n53_), .Y(mai_mai_n316_));
  NA2        m0267(.A(mai_mai_n164_), .B(mai_mai_n57_), .Y(mai_mai_n317_));
  OA220      m0268(.A0(mai_mai_n317_), .A1(mai_mai_n316_), .B0(mai_mai_n315_), .B1(mai_mai_n314_), .Y(mai_mai_n318_));
  AOI210     m0269(.A0(mai_mai_n318_), .A1(mai_mai_n313_), .B0(mai_mai_n304_), .Y(mai_mai_n319_));
  INV        m0270(.A(mai_mai_n297_), .Y(mai_mai_n320_));
  NO2        m0271(.A(x7), .B(mai_mai_n71_), .Y(mai_mai_n321_));
  NA2        m0272(.A(mai_mai_n108_), .B(x3), .Y(mai_mai_n322_));
  NO2        m0273(.A(mai_mai_n322_), .B(mai_mai_n321_), .Y(mai_mai_n323_));
  NA2        m0274(.A(mai_mai_n323_), .B(mai_mai_n320_), .Y(mai_mai_n324_));
  NA2        m0275(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n325_));
  NO2        m0276(.A(mai_mai_n325_), .B(x7), .Y(mai_mai_n326_));
  NA2        m0277(.A(mai_mai_n326_), .B(mai_mai_n281_), .Y(mai_mai_n327_));
  NA2        m0278(.A(mai_mai_n169_), .B(x1), .Y(mai_mai_n328_));
  AOI210     m0279(.A0(mai_mai_n327_), .A1(mai_mai_n324_), .B0(mai_mai_n328_), .Y(mai_mai_n329_));
  NO2        m0280(.A(mai_mai_n57_), .B(mai_mai_n50_), .Y(mai_mai_n330_));
  NO2        m0281(.A(mai_mai_n55_), .B(mai_mai_n110_), .Y(mai_mai_n331_));
  NA3        m0282(.A(mai_mai_n331_), .B(mai_mai_n330_), .C(mai_mai_n59_), .Y(mai_mai_n332_));
  NO2        m0283(.A(mai_mai_n159_), .B(x6), .Y(mai_mai_n333_));
  NO2        m0284(.A(mai_mai_n104_), .B(mai_mai_n108_), .Y(mai_mai_n334_));
  NA2        m0285(.A(mai_mai_n57_), .B(mai_mai_n110_), .Y(mai_mai_n335_));
  NO2        m0286(.A(mai_mai_n335_), .B(mai_mai_n269_), .Y(mai_mai_n336_));
  OAI210     m0287(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  OAI210     m0288(.A0(mai_mai_n332_), .A1(mai_mai_n104_), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  NO3        m0289(.A(mai_mai_n338_), .B(mai_mai_n329_), .C(mai_mai_n319_), .Y(mai_mai_n339_));
  AOI210     m0290(.A0(mai_mai_n339_), .A1(mai_mai_n303_), .B0(x4), .Y(mai_mai_n340_));
  NA2        m0291(.A(x8), .B(mai_mai_n71_), .Y(mai_mai_n341_));
  NO2        m0292(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n342_));
  NA3        m0293(.A(mai_mai_n342_), .B(mai_mai_n108_), .C(mai_mai_n53_), .Y(mai_mai_n343_));
  NO2        m0294(.A(x3), .B(x0), .Y(mai_mai_n344_));
  NAi21      m0295(.An(mai_mai_n344_), .B(mai_mai_n107_), .Y(mai_mai_n345_));
  NA2        m0296(.A(x5), .B(x2), .Y(mai_mai_n346_));
  NO2        m0297(.A(mai_mai_n346_), .B(mai_mai_n224_), .Y(mai_mai_n347_));
  AOI210     m0298(.A0(mai_mai_n347_), .A1(mai_mai_n345_), .B0(mai_mai_n245_), .Y(mai_mai_n348_));
  AO210      m0299(.A0(mai_mai_n348_), .A1(mai_mai_n343_), .B0(mai_mai_n341_), .Y(mai_mai_n349_));
  NO2        m0300(.A(mai_mai_n110_), .B(mai_mai_n53_), .Y(mai_mai_n350_));
  NA2        m0301(.A(mai_mai_n350_), .B(x3), .Y(mai_mai_n351_));
  NO2        m0302(.A(mai_mai_n55_), .B(x1), .Y(mai_mai_n352_));
  NA2        m0303(.A(mai_mai_n352_), .B(mai_mai_n110_), .Y(mai_mai_n353_));
  OAI210     m0304(.A0(mai_mai_n353_), .A1(mai_mai_n172_), .B0(mai_mai_n351_), .Y(mai_mai_n354_));
  NAi32      m0305(.An(x3), .Bn(x0), .C(x2), .Y(mai_mai_n355_));
  NO2        m0306(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n356_));
  NAi21      m0307(.An(x6), .B(x5), .Y(mai_mai_n357_));
  NO2        m0308(.A(x2), .B(mai_mai_n59_), .Y(mai_mai_n358_));
  NO4        m0309(.A(mai_mai_n358_), .B(mai_mai_n357_), .C(mai_mai_n161_), .D(mai_mai_n356_), .Y(mai_mai_n359_));
  AOI220     m0310(.A0(mai_mai_n359_), .A1(mai_mai_n355_), .B0(mai_mai_n354_), .B1(mai_mai_n85_), .Y(mai_mai_n360_));
  AOI210     m0311(.A0(mai_mai_n360_), .A1(mai_mai_n349_), .B0(mai_mai_n75_), .Y(mai_mai_n361_));
  NA2        m0312(.A(mai_mai_n352_), .B(mai_mai_n56_), .Y(mai_mai_n362_));
  NO2        m0313(.A(mai_mai_n108_), .B(mai_mai_n50_), .Y(mai_mai_n363_));
  NO2        m0314(.A(mai_mai_n291_), .B(mai_mai_n221_), .Y(mai_mai_n364_));
  XO2        m0315(.A(x7), .B(x2), .Y(mai_mai_n365_));
  INV        m0316(.A(mai_mai_n365_), .Y(mai_mai_n366_));
  XO2        m0317(.A(x6), .B(x2), .Y(mai_mai_n367_));
  NA4        m0318(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(mai_mai_n364_), .D(mai_mai_n363_), .Y(mai_mai_n368_));
  NAi21      m0319(.An(x0), .B(x6), .Y(mai_mai_n369_));
  AOI210     m0320(.A0(mai_mai_n369_), .A1(mai_mai_n145_), .B0(mai_mai_n273_), .Y(mai_mai_n370_));
  XN2        m0321(.A(x7), .B(x5), .Y(mai_mai_n371_));
  NA2        m0322(.A(mai_mai_n371_), .B(mai_mai_n71_), .Y(mai_mai_n372_));
  NA2        m0323(.A(x7), .B(x5), .Y(mai_mai_n373_));
  AOI210     m0324(.A0(mai_mai_n373_), .A1(x6), .B0(mai_mai_n355_), .Y(mai_mai_n374_));
  AOI220     m0325(.A0(mai_mai_n374_), .A1(mai_mai_n372_), .B0(mai_mai_n370_), .B1(mai_mai_n323_), .Y(mai_mai_n375_));
  AOI210     m0326(.A0(mai_mai_n375_), .A1(mai_mai_n368_), .B0(mai_mai_n362_), .Y(mai_mai_n376_));
  NO2        m0327(.A(x8), .B(x6), .Y(mai_mai_n377_));
  NAi21      m0328(.An(mai_mai_n377_), .B(mai_mai_n233_), .Y(mai_mai_n378_));
  AOI210     m0329(.A0(mai_mai_n378_), .A1(mai_mai_n92_), .B0(x3), .Y(mai_mai_n379_));
  NA2        m0330(.A(mai_mai_n108_), .B(x2), .Y(mai_mai_n380_));
  NO2        m0331(.A(mai_mai_n380_), .B(mai_mai_n64_), .Y(mai_mai_n381_));
  NA2        m0332(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n382_));
  NA2        m0333(.A(mai_mai_n50_), .B(mai_mai_n381_), .Y(mai_mai_n383_));
  NA2        m0334(.A(x4), .B(x2), .Y(mai_mai_n384_));
  NO2        m0335(.A(mai_mai_n384_), .B(mai_mai_n108_), .Y(mai_mai_n385_));
  NAi21      m0336(.An(x1), .B(x6), .Y(mai_mai_n386_));
  NA2        m0337(.A(mai_mai_n344_), .B(mai_mai_n274_), .Y(mai_mai_n387_));
  OAI220     m0338(.A0(mai_mai_n387_), .A1(mai_mai_n386_), .B0(mai_mai_n107_), .B1(mai_mai_n53_), .Y(mai_mai_n388_));
  NA2        m0339(.A(x8), .B(x2), .Y(mai_mai_n389_));
  NO2        m0340(.A(mai_mai_n389_), .B(mai_mai_n50_), .Y(mai_mai_n390_));
  INV        m0341(.A(mai_mai_n223_), .Y(mai_mai_n391_));
  NO2        m0342(.A(mai_mai_n391_), .B(mai_mai_n52_), .Y(mai_mai_n392_));
  AOI220     m0343(.A0(mai_mai_n392_), .A1(mai_mai_n390_), .B0(mai_mai_n388_), .B1(mai_mai_n385_), .Y(mai_mai_n393_));
  OAI210     m0344(.A0(mai_mai_n383_), .A1(mai_mai_n379_), .B0(mai_mai_n393_), .Y(mai_mai_n394_));
  NO4        m0345(.A(mai_mai_n394_), .B(mai_mai_n376_), .C(mai_mai_n361_), .D(mai_mai_n340_), .Y(mai03));
  NAi21      m0346(.An(x2), .B(x0), .Y(mai_mai_n396_));
  NO3        m0347(.A(x8), .B(x6), .C(x4), .Y(mai_mai_n397_));
  INV        m0348(.A(mai_mai_n397_), .Y(mai_mai_n398_));
  NO2        m0349(.A(mai_mai_n398_), .B(mai_mai_n396_), .Y(mai_mai_n399_));
  NA2        m0350(.A(mai_mai_n111_), .B(mai_mai_n59_), .Y(mai_mai_n400_));
  NO2        m0351(.A(mai_mai_n400_), .B(mai_mai_n55_), .Y(mai_mai_n401_));
  OAI210     m0352(.A0(mai_mai_n401_), .A1(mai_mai_n399_), .B0(mai_mai_n164_), .Y(mai_mai_n402_));
  NA2        m0353(.A(x3), .B(x2), .Y(mai_mai_n403_));
  NO2        m0354(.A(mai_mai_n161_), .B(x0), .Y(mai_mai_n404_));
  NA2        m0355(.A(x8), .B(x0), .Y(mai_mai_n405_));
  NO2        m0356(.A(mai_mai_n405_), .B(x6), .Y(mai_mai_n406_));
  AOI210     m0357(.A0(mai_mai_n406_), .A1(x5), .B0(mai_mai_n404_), .Y(mai_mai_n407_));
  NO2        m0358(.A(mai_mai_n407_), .B(mai_mai_n403_), .Y(mai_mai_n408_));
  NO2        m0359(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n409_));
  NO2        m0360(.A(x3), .B(x2), .Y(mai_mai_n410_));
  NA2        m0361(.A(mai_mai_n410_), .B(mai_mai_n409_), .Y(mai_mai_n411_));
  NO2        m0362(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n412_));
  NA2        m0363(.A(mai_mai_n412_), .B(x5), .Y(mai_mai_n413_));
  AOI210     m0364(.A0(mai_mai_n413_), .A1(mai_mai_n411_), .B0(mai_mai_n304_), .Y(mai_mai_n414_));
  NA2        m0365(.A(mai_mai_n259_), .B(mai_mai_n174_), .Y(mai_mai_n415_));
  NO2        m0366(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n416_));
  NO2        m0367(.A(mai_mai_n71_), .B(x0), .Y(mai_mai_n417_));
  NO4        m0368(.A(mai_mai_n417_), .B(mai_mai_n416_), .C(x2), .D(mai_mai_n53_), .Y(mai_mai_n418_));
  AO210      m0369(.A0(mai_mai_n418_), .A1(mai_mai_n415_), .B0(mai_mai_n414_), .Y(mai_mai_n419_));
  OAI210     m0370(.A0(mai_mai_n419_), .A1(mai_mai_n408_), .B0(x4), .Y(mai_mai_n420_));
  NO2        m0371(.A(x4), .B(mai_mai_n53_), .Y(mai_mai_n421_));
  NA2        m0372(.A(mai_mai_n421_), .B(mai_mai_n59_), .Y(mai_mai_n422_));
  NO3        m0373(.A(mai_mai_n422_), .B(mai_mai_n233_), .C(x5), .Y(mai_mai_n423_));
  NA2        m0374(.A(x7), .B(mai_mai_n108_), .Y(mai_mai_n424_));
  NO3        m0375(.A(x5), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n425_));
  INV        m0376(.A(mai_mai_n425_), .Y(mai_mai_n426_));
  NO2        m0377(.A(x6), .B(mai_mai_n56_), .Y(mai_mai_n427_));
  NO2        m0378(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n428_));
  NA2        m0379(.A(mai_mai_n428_), .B(mai_mai_n427_), .Y(mai_mai_n429_));
  OAI210     m0380(.A0(mai_mai_n429_), .A1(mai_mai_n426_), .B0(mai_mai_n424_), .Y(mai_mai_n430_));
  AOI210     m0381(.A0(mai_mai_n423_), .A1(x2), .B0(mai_mai_n430_), .Y(mai_mai_n431_));
  AOI220     m0382(.A0(mai_mai_n431_), .A1(mai_mai_n420_), .B0(mai_mai_n402_), .B1(x7), .Y(mai_mai_n432_));
  NA2        m0383(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n433_));
  NO2        m0384(.A(mai_mai_n258_), .B(mai_mai_n110_), .Y(mai_mai_n434_));
  NO2        m0385(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n435_));
  NO3        m0386(.A(mai_mai_n435_), .B(mai_mai_n434_), .C(mai_mai_n148_), .Y(mai_mai_n436_));
  AOI210     m0387(.A0(mai_mai_n208_), .A1(mai_mai_n101_), .B0(mai_mai_n436_), .Y(mai_mai_n437_));
  NO2        m0388(.A(x5), .B(x2), .Y(mai_mai_n438_));
  NO2        m0389(.A(x8), .B(x3), .Y(mai_mai_n439_));
  NA2        m0390(.A(mai_mai_n439_), .B(mai_mai_n438_), .Y(mai_mai_n440_));
  NO2        m0391(.A(mai_mai_n440_), .B(x6), .Y(mai_mai_n441_));
  NA2        m0392(.A(mai_mai_n207_), .B(x2), .Y(mai_mai_n442_));
  NO3        m0393(.A(mai_mai_n439_), .B(mai_mai_n345_), .C(mai_mai_n357_), .Y(mai_mai_n443_));
  AOI210     m0394(.A0(mai_mai_n443_), .A1(mai_mai_n442_), .B0(mai_mai_n441_), .Y(mai_mai_n444_));
  OAI210     m0395(.A0(mai_mai_n437_), .A1(mai_mai_n291_), .B0(mai_mai_n444_), .Y(mai_mai_n445_));
  NA2        m0396(.A(mai_mai_n445_), .B(x4), .Y(mai_mai_n446_));
  NA2        m0397(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n447_));
  NO2        m0398(.A(mai_mai_n447_), .B(x5), .Y(mai_mai_n448_));
  NAi21      m0399(.An(x4), .B(x6), .Y(mai_mai_n449_));
  NO2        m0400(.A(mai_mai_n449_), .B(mai_mai_n51_), .Y(mai_mai_n450_));
  NO2        m0401(.A(mai_mai_n55_), .B(mai_mai_n71_), .Y(mai_mai_n451_));
  NO2        m0402(.A(mai_mai_n50_), .B(mai_mai_n110_), .Y(mai_mai_n452_));
  NO2        m0403(.A(mai_mai_n233_), .B(x0), .Y(mai_mai_n453_));
  NO2        m0404(.A(mai_mai_n357_), .B(x8), .Y(mai_mai_n454_));
  OAI210     m0405(.A0(mai_mai_n454_), .A1(mai_mai_n453_), .B0(mai_mai_n452_), .Y(mai_mai_n455_));
  OAI210     m0406(.A0(mai_mai_n411_), .A1(mai_mai_n451_), .B0(mai_mai_n455_), .Y(mai_mai_n456_));
  AOI220     m0407(.A0(mai_mai_n456_), .A1(mai_mai_n56_), .B0(mai_mai_n450_), .B1(mai_mai_n448_), .Y(mai_mai_n457_));
  AOI210     m0408(.A0(mai_mai_n457_), .A1(mai_mai_n446_), .B0(mai_mai_n433_), .Y(mai_mai_n458_));
  NA2        m0409(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n459_));
  NO2        m0410(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n460_));
  NA2        m0411(.A(mai_mai_n356_), .B(mai_mai_n59_), .Y(mai_mai_n461_));
  NO3        m0412(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n462_));
  NA2        m0413(.A(mai_mai_n435_), .B(x5), .Y(mai_mai_n463_));
  NO2        m0414(.A(x8), .B(x5), .Y(mai_mai_n464_));
  NAi21      m0415(.An(mai_mai_n464_), .B(mai_mai_n174_), .Y(mai_mai_n465_));
  OAI210     m0416(.A0(mai_mai_n465_), .A1(mai_mai_n309_), .B0(mai_mai_n463_), .Y(mai_mai_n466_));
  NA2        m0417(.A(mai_mai_n364_), .B(mai_mai_n77_), .Y(mai_mai_n467_));
  NOi21      m0418(.An(x3), .B(x4), .Y(mai_mai_n468_));
  NA2        m0419(.A(mai_mai_n55_), .B(mai_mai_n110_), .Y(mai_mai_n469_));
  NA2        m0420(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  NO2        m0421(.A(mai_mai_n51_), .B(x6), .Y(mai_mai_n471_));
  NO2        m0422(.A(mai_mai_n148_), .B(mai_mai_n55_), .Y(mai_mai_n472_));
  NO3        m0423(.A(mai_mai_n56_), .B(x2), .C(x0), .Y(mai_mai_n473_));
  AOI220     m0424(.A0(mai_mai_n473_), .A1(mai_mai_n472_), .B0(mai_mai_n471_), .B1(mai_mai_n448_), .Y(mai_mai_n474_));
  OAI210     m0425(.A0(mai_mai_n470_), .A1(mai_mai_n467_), .B0(mai_mai_n474_), .Y(mai_mai_n475_));
  AOI210     m0426(.A0(mai_mai_n466_), .A1(mai_mai_n462_), .B0(mai_mai_n475_), .Y(mai_mai_n476_));
  NO2        m0427(.A(mai_mai_n476_), .B(mai_mai_n459_), .Y(mai_mai_n477_));
  NA2        m0428(.A(x7), .B(x1), .Y(mai_mai_n478_));
  NO3        m0429(.A(x5), .B(x4), .C(x2), .Y(mai_mai_n479_));
  AN2        m0430(.A(mai_mai_n479_), .B(mai_mai_n377_), .Y(mai_mai_n480_));
  NO3        m0431(.A(mai_mai_n480_), .B(mai_mai_n472_), .C(mai_mai_n385_), .Y(mai_mai_n481_));
  OAI210     m0432(.A0(mai_mai_n377_), .A1(mai_mai_n84_), .B0(mai_mai_n344_), .Y(mai_mai_n482_));
  NO2        m0433(.A(mai_mai_n482_), .B(mai_mai_n481_), .Y(mai_mai_n483_));
  NO2        m0434(.A(x4), .B(mai_mai_n110_), .Y(mai_mai_n484_));
  NA2        m0435(.A(mai_mai_n484_), .B(x6), .Y(mai_mai_n485_));
  NA3        m0436(.A(mai_mai_n108_), .B(x4), .C(mai_mai_n110_), .Y(mai_mai_n486_));
  AOI210     m0437(.A0(mai_mai_n486_), .A1(mai_mai_n485_), .B0(mai_mai_n100_), .Y(mai_mai_n487_));
  NA2        m0438(.A(mai_mai_n468_), .B(mai_mai_n71_), .Y(mai_mai_n488_));
  NA2        m0439(.A(mai_mai_n169_), .B(mai_mai_n59_), .Y(mai_mai_n489_));
  NO2        m0440(.A(mai_mai_n489_), .B(mai_mai_n488_), .Y(mai_mai_n490_));
  NA2        m0441(.A(mai_mai_n452_), .B(x4), .Y(mai_mai_n491_));
  NO3        m0442(.A(mai_mai_n491_), .B(mai_mai_n377_), .C(mai_mai_n417_), .Y(mai_mai_n492_));
  NO4        m0443(.A(mai_mai_n492_), .B(mai_mai_n490_), .C(mai_mai_n487_), .D(mai_mai_n483_), .Y(mai_mai_n493_));
  NA2        m0444(.A(x5), .B(x4), .Y(mai_mai_n494_));
  NO2        m0445(.A(mai_mai_n71_), .B(mai_mai_n53_), .Y(mai_mai_n495_));
  NO3        m0446(.A(x8), .B(x3), .C(x2), .Y(mai_mai_n496_));
  NA3        m0447(.A(mai_mai_n496_), .B(mai_mai_n495_), .C(mai_mai_n59_), .Y(mai_mai_n497_));
  NO3        m0448(.A(x6), .B(x5), .C(x2), .Y(mai_mai_n498_));
  NO2        m0449(.A(mai_mai_n497_), .B(mai_mai_n494_), .Y(mai_mai_n499_));
  NA2        m0450(.A(mai_mai_n71_), .B(x2), .Y(mai_mai_n500_));
  NO3        m0451(.A(x4), .B(x3), .C(mai_mai_n59_), .Y(mai_mai_n501_));
  NA2        m0452(.A(mai_mai_n501_), .B(mai_mai_n230_), .Y(mai_mai_n502_));
  NO3        m0453(.A(mai_mai_n502_), .B(mai_mai_n500_), .C(mai_mai_n96_), .Y(mai_mai_n503_));
  XO2        m0454(.A(x4), .B(x0), .Y(mai_mai_n504_));
  NA2        m0455(.A(mai_mai_n269_), .B(x5), .Y(mai_mai_n505_));
  NO2        m0456(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n506_));
  NO2        m0457(.A(mai_mai_n506_), .B(mai_mai_n63_), .Y(mai_mai_n507_));
  NO4        m0458(.A(mai_mai_n507_), .B(mai_mai_n505_), .C(mai_mai_n504_), .D(mai_mai_n157_), .Y(mai_mai_n508_));
  NO3        m0459(.A(mai_mai_n508_), .B(mai_mai_n503_), .C(mai_mai_n499_), .Y(mai_mai_n509_));
  OAI210     m0460(.A0(mai_mai_n493_), .A1(mai_mai_n478_), .B0(mai_mai_n509_), .Y(mai_mai_n510_));
  NO4        m0461(.A(mai_mai_n510_), .B(mai_mai_n477_), .C(mai_mai_n458_), .D(mai_mai_n432_), .Y(mai04));
  NO2        m0462(.A(x7), .B(x2), .Y(mai_mai_n512_));
  NO2        m0463(.A(x3), .B(mai_mai_n53_), .Y(mai_mai_n513_));
  NO2        m0464(.A(mai_mai_n513_), .B(mai_mai_n150_), .Y(mai_mai_n514_));
  XN2        m0465(.A(x8), .B(x1), .Y(mai_mai_n515_));
  NO2        m0466(.A(mai_mai_n515_), .B(mai_mai_n148_), .Y(mai_mai_n516_));
  NA2        m0467(.A(mai_mai_n516_), .B(mai_mai_n514_), .Y(mai_mai_n517_));
  NA2        m0468(.A(x6), .B(x3), .Y(mai_mai_n518_));
  NO2        m0469(.A(mai_mai_n518_), .B(x5), .Y(mai_mai_n519_));
  NA2        m0470(.A(mai_mai_n71_), .B(x1), .Y(mai_mai_n520_));
  NO2        m0471(.A(mai_mai_n464_), .B(mai_mai_n258_), .Y(mai_mai_n521_));
  NO3        m0472(.A(mai_mai_n521_), .B(mai_mai_n439_), .C(mai_mai_n520_), .Y(mai_mai_n522_));
  INV        m0473(.A(mai_mai_n522_), .Y(mai_mai_n523_));
  AOI210     m0474(.A0(mai_mai_n523_), .A1(mai_mai_n517_), .B0(x0), .Y(mai_mai_n524_));
  NOi21      m0475(.An(mai_mai_n174_), .B(mai_mai_n464_), .Y(mai_mai_n525_));
  NA2        m0476(.A(mai_mai_n109_), .B(x1), .Y(mai_mai_n526_));
  NO3        m0477(.A(mai_mai_n526_), .B(mai_mai_n525_), .C(mai_mai_n325_), .Y(mai_mai_n527_));
  OAI210     m0478(.A0(mai_mai_n527_), .A1(mai_mai_n524_), .B0(mai_mai_n512_), .Y(mai_mai_n528_));
  NA2        m0479(.A(mai_mai_n137_), .B(mai_mai_n244_), .Y(mai_mai_n529_));
  OR4        m0480(.A(mai_mai_n529_), .B(mai_mai_n378_), .C(mai_mai_n82_), .D(mai_mai_n54_), .Y(mai_mai_n530_));
  OR2        m0481(.A(x6), .B(x0), .Y(mai_mai_n531_));
  NO3        m0482(.A(mai_mai_n531_), .B(x3), .C(x1), .Y(mai_mai_n532_));
  AOI220     m0483(.A0(mai_mai_n532_), .A1(mai_mai_n108_), .B0(mai_mai_n281_), .B1(mai_mai_n275_), .Y(mai_mai_n533_));
  AOI210     m0484(.A0(mai_mai_n533_), .A1(mai_mai_n530_), .B0(mai_mai_n187_), .Y(mai_mai_n534_));
  NA2        m0485(.A(x7), .B(x2), .Y(mai_mai_n535_));
  INV        m0486(.A(mai_mai_n137_), .Y(mai_mai_n536_));
  OAI210     m0487(.A0(mai_mai_n173_), .A1(mai_mai_n536_), .B0(mai_mai_n82_), .Y(mai_mai_n537_));
  NO2        m0488(.A(mai_mai_n322_), .B(mai_mai_n55_), .Y(mai_mai_n538_));
  NO3        m0489(.A(x3), .B(x1), .C(x0), .Y(mai_mai_n539_));
  OR2        m0490(.A(x6), .B(x1), .Y(mai_mai_n540_));
  NA2        m0491(.A(mai_mai_n540_), .B(x0), .Y(mai_mai_n541_));
  AOI220     m0492(.A0(mai_mai_n541_), .A1(mai_mai_n538_), .B0(mai_mai_n539_), .B1(mai_mai_n472_), .Y(mai_mai_n542_));
  AOI210     m0493(.A0(mai_mai_n542_), .A1(mai_mai_n537_), .B0(mai_mai_n535_), .Y(mai_mai_n543_));
  NA2        m0494(.A(mai_mai_n71_), .B(x0), .Y(mai_mai_n544_));
  NOi31      m0495(.An(mai_mai_n347_), .B(mai_mai_n544_), .C(mai_mai_n265_), .Y(mai_mai_n545_));
  NO4        m0496(.A(mai_mai_n545_), .B(mai_mai_n543_), .C(mai_mai_n534_), .D(mai_mai_n56_), .Y(mai_mai_n546_));
  NA2        m0497(.A(mai_mai_n546_), .B(mai_mai_n528_), .Y(mai_mai_n547_));
  NA3        m0498(.A(x8), .B(x7), .C(x0), .Y(mai_mai_n548_));
  INV        m0499(.A(mai_mai_n548_), .Y(mai_mai_n549_));
  AOI210     m0500(.A0(mai_mai_n274_), .A1(mai_mai_n99_), .B0(mai_mai_n549_), .Y(mai_mai_n550_));
  NO2        m0501(.A(mai_mai_n550_), .B(mai_mai_n157_), .Y(mai_mai_n551_));
  NA2        m0502(.A(mai_mai_n435_), .B(mai_mai_n57_), .Y(mai_mai_n552_));
  NO2        m0503(.A(x8), .B(x0), .Y(mai_mai_n553_));
  NA2        m0504(.A(mai_mai_n553_), .B(mai_mai_n366_), .Y(mai_mai_n554_));
  AOI210     m0505(.A0(mai_mai_n554_), .A1(mai_mai_n552_), .B0(mai_mai_n277_), .Y(mai_mai_n555_));
  OAI210     m0506(.A0(mai_mai_n555_), .A1(mai_mai_n551_), .B0(mai_mai_n281_), .Y(mai_mai_n556_));
  NO2        m0507(.A(mai_mai_n71_), .B(mai_mai_n110_), .Y(mai_mai_n557_));
  NO2        m0508(.A(mai_mai_n373_), .B(x8), .Y(mai_mai_n558_));
  NO2        m0509(.A(mai_mai_n558_), .B(mai_mai_n266_), .Y(mai_mai_n559_));
  NO3        m0510(.A(mai_mai_n559_), .B(mai_mai_n382_), .C(mai_mai_n272_), .Y(mai_mai_n560_));
  NO2        m0511(.A(mai_mai_n290_), .B(x8), .Y(mai_mai_n561_));
  OAI210     m0512(.A0(mai_mai_n464_), .A1(mai_mai_n330_), .B0(mai_mai_n247_), .Y(mai_mai_n562_));
  NA2        m0513(.A(mai_mai_n352_), .B(mai_mai_n179_), .Y(mai_mai_n563_));
  OAI220     m0514(.A0(mai_mai_n563_), .A1(mai_mai_n59_), .B0(mai_mai_n562_), .B1(mai_mai_n561_), .Y(mai_mai_n564_));
  OAI210     m0515(.A0(mai_mai_n564_), .A1(mai_mai_n560_), .B0(mai_mai_n557_), .Y(mai_mai_n565_));
  NO2        m0516(.A(x8), .B(x2), .Y(mai_mai_n566_));
  NO2        m0517(.A(mai_mai_n224_), .B(mai_mai_n57_), .Y(mai_mai_n567_));
  NA3        m0518(.A(mai_mai_n567_), .B(mai_mai_n566_), .C(mai_mai_n345_), .Y(mai_mai_n568_));
  NO2        m0519(.A(mai_mai_n248_), .B(mai_mai_n137_), .Y(mai_mai_n569_));
  AOI210     m0520(.A0(mai_mai_n326_), .A1(mai_mai_n165_), .B0(mai_mai_n569_), .Y(mai_mai_n570_));
  AOI210     m0521(.A0(mai_mai_n570_), .A1(mai_mai_n568_), .B0(mai_mai_n109_), .Y(mai_mai_n571_));
  NA2        m0522(.A(mai_mai_n342_), .B(x2), .Y(mai_mai_n572_));
  NO2        m0523(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n573_));
  NA2        m0524(.A(mai_mai_n573_), .B(mai_mai_n63_), .Y(mai_mai_n574_));
  AOI210     m0525(.A0(mai_mai_n572_), .A1(mai_mai_n461_), .B0(mai_mai_n574_), .Y(mai_mai_n575_));
  NA2        m0526(.A(mai_mai_n110_), .B(mai_mai_n53_), .Y(mai_mai_n576_));
  NO2        m0527(.A(mai_mai_n576_), .B(x8), .Y(mai_mai_n577_));
  NA2        m0528(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n578_));
  NO2        m0529(.A(mai_mai_n184_), .B(mai_mai_n578_), .Y(mai_mai_n579_));
  AN2        m0530(.A(mai_mai_n579_), .B(mai_mai_n577_), .Y(mai_mai_n580_));
  NA2        m0531(.A(mai_mai_n409_), .B(mai_mai_n150_), .Y(mai_mai_n581_));
  NO2        m0532(.A(mai_mai_n71_), .B(x2), .Y(mai_mai_n582_));
  NA2        m0533(.A(mai_mai_n582_), .B(mai_mai_n274_), .Y(mai_mai_n583_));
  OAI210     m0534(.A0(mai_mai_n583_), .A1(mai_mai_n581_), .B0(mai_mai_n56_), .Y(mai_mai_n584_));
  NO4        m0535(.A(mai_mai_n584_), .B(mai_mai_n580_), .C(mai_mai_n575_), .D(mai_mai_n571_), .Y(mai_mai_n585_));
  NA3        m0536(.A(mai_mai_n585_), .B(mai_mai_n565_), .C(mai_mai_n556_), .Y(mai_mai_n586_));
  NA2        m0537(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n587_));
  NOi21      m0538(.An(x2), .B(x7), .Y(mai_mai_n588_));
  NO2        m0539(.A(x6), .B(x3), .Y(mai_mai_n589_));
  NA2        m0540(.A(mai_mai_n589_), .B(mai_mai_n588_), .Y(mai_mai_n590_));
  NO2        m0541(.A(x6), .B(mai_mai_n59_), .Y(mai_mai_n591_));
  NO3        m0542(.A(mai_mai_n57_), .B(x2), .C(x1), .Y(mai_mai_n592_));
  NO3        m0543(.A(mai_mai_n57_), .B(x2), .C(x0), .Y(mai_mai_n593_));
  AOI220     m0544(.A0(mai_mai_n593_), .A1(mai_mai_n227_), .B0(mai_mai_n592_), .B1(mai_mai_n591_), .Y(mai_mai_n594_));
  OAI210     m0545(.A0(mai_mai_n590_), .A1(mai_mai_n587_), .B0(mai_mai_n594_), .Y(mai_mai_n595_));
  NO2        m0546(.A(mai_mai_n101_), .B(mai_mai_n53_), .Y(mai_mai_n596_));
  NA2        m0547(.A(mai_mai_n222_), .B(mai_mai_n57_), .Y(mai_mai_n597_));
  OAI210     m0548(.A0(mai_mai_n596_), .A1(mai_mai_n454_), .B0(mai_mai_n597_), .Y(mai_mai_n598_));
  NO3        m0549(.A(mai_mai_n598_), .B(mai_mai_n491_), .C(mai_mai_n59_), .Y(mai_mai_n599_));
  AO210      m0550(.A0(mai_mai_n595_), .A1(mai_mai_n464_), .B0(mai_mai_n599_), .Y(mai_mai_n600_));
  AOI210     m0551(.A0(mai_mai_n586_), .A1(mai_mai_n547_), .B0(mai_mai_n600_), .Y(mai05));
  AOI210     m0552(.A0(mai_mai_n164_), .A1(mai_mai_n55_), .B0(mai_mai_n506_), .Y(mai_mai_n602_));
  OR2        m0553(.A(mai_mai_n602_), .B(mai_mai_n57_), .Y(mai_mai_n603_));
  NO2        m0554(.A(x7), .B(mai_mai_n108_), .Y(mai_mai_n604_));
  NO2        m0555(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n605_));
  NA2        m0556(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n606_));
  NO2        m0557(.A(mai_mai_n606_), .B(mai_mai_n578_), .Y(mai_mai_n607_));
  AOI210     m0558(.A0(mai_mai_n605_), .A1(mai_mai_n604_), .B0(mai_mai_n607_), .Y(mai_mai_n608_));
  AOI210     m0559(.A0(mai_mai_n608_), .A1(mai_mai_n603_), .B0(mai_mai_n110_), .Y(mai_mai_n609_));
  NO2        m0560(.A(x7), .B(x4), .Y(mai_mai_n610_));
  NO2        m0561(.A(mai_mai_n64_), .B(mai_mai_n55_), .Y(mai_mai_n611_));
  NO2        m0562(.A(mai_mai_n200_), .B(x5), .Y(mai_mai_n612_));
  NA2        m0563(.A(mai_mai_n108_), .B(mai_mai_n110_), .Y(mai_mai_n613_));
  NO2        m0564(.A(mai_mai_n613_), .B(mai_mai_n218_), .Y(mai_mai_n614_));
  AO220      m0565(.A0(mai_mai_n614_), .A1(mai_mai_n610_), .B0(mai_mai_n612_), .B1(mai_mai_n611_), .Y(mai_mai_n615_));
  OAI210     m0566(.A0(mai_mai_n615_), .A1(mai_mai_n609_), .B0(mai_mai_n495_), .Y(mai_mai_n616_));
  NO2        m0567(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n617_));
  NA2        m0568(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n618_));
  NO2        m0569(.A(mai_mai_n108_), .B(mai_mai_n110_), .Y(mai_mai_n619_));
  NA2        m0570(.A(mai_mai_n619_), .B(x7), .Y(mai_mai_n620_));
  NA2        m0571(.A(mai_mai_n438_), .B(mai_mai_n257_), .Y(mai_mai_n621_));
  AOI210     m0572(.A0(mai_mai_n621_), .A1(mai_mai_n620_), .B0(mai_mai_n618_), .Y(mai_mai_n622_));
  NA2        m0573(.A(mai_mai_n108_), .B(x4), .Y(mai_mai_n623_));
  XO2        m0574(.A(x7), .B(x5), .Y(mai_mai_n624_));
  NO2        m0575(.A(mai_mai_n624_), .B(mai_mai_n53_), .Y(mai_mai_n625_));
  NA3        m0576(.A(mai_mai_n625_), .B(mai_mai_n623_), .C(mai_mai_n331_), .Y(mai_mai_n626_));
  NO2        m0577(.A(mai_mai_n108_), .B(x2), .Y(mai_mai_n627_));
  NO2        m0578(.A(mai_mai_n75_), .B(mai_mai_n55_), .Y(mai_mai_n628_));
  NA2        m0579(.A(mai_mai_n628_), .B(mai_mai_n627_), .Y(mai_mai_n629_));
  NA2        m0580(.A(mai_mai_n629_), .B(mai_mai_n626_), .Y(mai_mai_n630_));
  OAI210     m0581(.A0(mai_mai_n630_), .A1(mai_mai_n622_), .B0(mai_mai_n617_), .Y(mai_mai_n631_));
  NO2        m0582(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n632_));
  NO2        m0583(.A(mai_mai_n194_), .B(x4), .Y(mai_mai_n633_));
  NO2        m0584(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n634_));
  XO2        m0585(.A(x5), .B(x2), .Y(mai_mai_n635_));
  NO3        m0586(.A(x8), .B(x7), .C(mai_mai_n110_), .Y(mai_mai_n636_));
  AO220      m0587(.A0(mai_mai_n636_), .A1(mai_mai_n634_), .B0(mai_mai_n635_), .B1(mai_mai_n633_), .Y(mai_mai_n637_));
  NA3        m0588(.A(mai_mai_n637_), .B(mai_mai_n632_), .C(mai_mai_n53_), .Y(mai_mai_n638_));
  NA2        m0589(.A(mai_mai_n272_), .B(mai_mai_n588_), .Y(mai_mai_n639_));
  NOi21      m0590(.An(x4), .B(x1), .Y(mai_mai_n640_));
  NA2        m0591(.A(x4), .B(x1), .Y(mai_mai_n641_));
  NO2        m0592(.A(mai_mai_n641_), .B(mai_mai_n50_), .Y(mai_mai_n642_));
  AOI210     m0593(.A0(mai_mai_n642_), .A1(mai_mai_n619_), .B0(mai_mai_n59_), .Y(mai_mai_n643_));
  NA4        m0594(.A(mai_mai_n643_), .B(mai_mai_n638_), .C(mai_mai_n631_), .D(mai_mai_n616_), .Y(mai_mai_n644_));
  NA2        m0595(.A(mai_mai_n632_), .B(mai_mai_n56_), .Y(mai_mai_n645_));
  NA2        m0596(.A(mai_mai_n566_), .B(mai_mai_n604_), .Y(mai_mai_n646_));
  NO2        m0597(.A(mai_mai_n646_), .B(mai_mai_n645_), .Y(mai_mai_n647_));
  NA2        m0598(.A(mai_mai_n274_), .B(mai_mai_n123_), .Y(mai_mai_n648_));
  OAI210     m0599(.A0(mai_mai_n648_), .A1(mai_mai_n166_), .B0(mai_mai_n59_), .Y(mai_mai_n649_));
  NA2        m0600(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n650_));
  NO2        m0601(.A(x3), .B(mai_mai_n91_), .Y(mai_mai_n651_));
  NA2        m0602(.A(mai_mai_n634_), .B(mai_mai_n156_), .Y(mai_mai_n652_));
  NO3        m0603(.A(mai_mai_n652_), .B(mai_mai_n651_), .C(mai_mai_n428_), .Y(mai_mai_n653_));
  NA2        m0604(.A(mai_mai_n282_), .B(mai_mai_n71_), .Y(mai_mai_n654_));
  NO2        m0605(.A(mai_mai_n389_), .B(x3), .Y(mai_mai_n655_));
  NA2        m0606(.A(mai_mai_n655_), .B(mai_mai_n241_), .Y(mai_mai_n656_));
  NO2        m0607(.A(mai_mai_n428_), .B(mai_mai_n633_), .Y(mai_mai_n657_));
  NO2        m0608(.A(mai_mai_n468_), .B(mai_mai_n108_), .Y(mai_mai_n658_));
  NO2        m0609(.A(mai_mai_n576_), .B(x6), .Y(mai_mai_n659_));
  NA2        m0610(.A(mai_mai_n659_), .B(mai_mai_n658_), .Y(mai_mai_n660_));
  OAI220     m0611(.A0(mai_mai_n660_), .A1(mai_mai_n657_), .B0(mai_mai_n656_), .B1(mai_mai_n654_), .Y(mai_mai_n661_));
  NO4        m0612(.A(mai_mai_n661_), .B(mai_mai_n653_), .C(mai_mai_n649_), .D(mai_mai_n647_), .Y(mai_mai_n662_));
  NA2        m0613(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n663_));
  NO2        m0614(.A(mai_mai_n663_), .B(x1), .Y(mai_mai_n664_));
  NA2        m0615(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n665_));
  NO2        m0616(.A(mai_mai_n665_), .B(mai_mai_n132_), .Y(mai_mai_n666_));
  NA2        m0617(.A(x8), .B(x4), .Y(mai_mai_n667_));
  NO2        m0618(.A(x8), .B(x4), .Y(mai_mai_n668_));
  NAi21      m0619(.An(mai_mai_n668_), .B(mai_mai_n667_), .Y(mai_mai_n669_));
  NAi21      m0620(.An(mai_mai_n566_), .B(mai_mai_n389_), .Y(mai_mai_n670_));
  NO4        m0621(.A(mai_mai_n670_), .B(mai_mai_n669_), .C(mai_mai_n428_), .D(mai_mai_n71_), .Y(mai_mai_n671_));
  OAI210     m0622(.A0(mai_mai_n671_), .A1(mai_mai_n666_), .B0(mai_mai_n664_), .Y(mai_mai_n672_));
  NO3        m0623(.A(x8), .B(mai_mai_n108_), .C(x4), .Y(mai_mai_n673_));
  INV        m0624(.A(mai_mai_n673_), .Y(mai_mai_n674_));
  NO2        m0625(.A(mai_mai_n674_), .B(mai_mai_n110_), .Y(mai_mai_n675_));
  NO2        m0626(.A(x5), .B(x4), .Y(mai_mai_n676_));
  NA3        m0627(.A(mai_mai_n676_), .B(mai_mai_n63_), .C(mai_mai_n110_), .Y(mai_mai_n677_));
  NO2        m0628(.A(x6), .B(mai_mai_n110_), .Y(mai_mai_n678_));
  NA2        m0629(.A(mai_mai_n665_), .B(mai_mai_n678_), .Y(mai_mai_n679_));
  OAI210     m0630(.A0(mai_mai_n679_), .A1(mai_mai_n525_), .B0(mai_mai_n677_), .Y(mai_mai_n680_));
  OAI210     m0631(.A0(mai_mai_n680_), .A1(mai_mai_n675_), .B0(mai_mai_n312_), .Y(mai_mai_n681_));
  NA3        m0632(.A(mai_mai_n681_), .B(mai_mai_n672_), .C(mai_mai_n662_), .Y(mai_mai_n682_));
  OR2        m0633(.A(x4), .B(x1), .Y(mai_mai_n683_));
  NO2        m0634(.A(mai_mai_n683_), .B(x3), .Y(mai_mai_n684_));
  NA2        m0635(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n685_));
  NO3        m0636(.A(mai_mai_n371_), .B(mai_mai_n685_), .C(x6), .Y(mai_mai_n686_));
  AOI220     m0637(.A0(mai_mai_n686_), .A1(mai_mai_n684_), .B0(mai_mai_n682_), .B1(mai_mai_n644_), .Y(mai06));
  NA2        m0638(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n688_));
  NA2        m0639(.A(x6), .B(mai_mai_n110_), .Y(mai_mai_n689_));
  NA2        m0640(.A(mai_mai_n689_), .B(mai_mai_n55_), .Y(mai_mai_n690_));
  NA2        m0641(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n691_));
  NO2        m0642(.A(mai_mai_n691_), .B(mai_mai_n118_), .Y(mai_mai_n692_));
  NA3        m0643(.A(mai_mai_n692_), .B(mai_mai_n690_), .C(mai_mai_n500_), .Y(mai_mai_n693_));
  NO2        m0644(.A(mai_mai_n389_), .B(x0), .Y(mai_mai_n694_));
  NA2        m0645(.A(mai_mai_n341_), .B(x2), .Y(mai_mai_n695_));
  NOi21      m0646(.An(x6), .B(x8), .Y(mai_mai_n696_));
  NO2        m0647(.A(mai_mai_n696_), .B(x2), .Y(mai_mai_n697_));
  NO3        m0648(.A(mai_mai_n697_), .B(mai_mai_n70_), .C(mai_mai_n59_), .Y(mai_mai_n698_));
  AOI220     m0649(.A0(mai_mai_n698_), .A1(mai_mai_n695_), .B0(mai_mai_n694_), .B1(mai_mai_n333_), .Y(mai_mai_n699_));
  AOI210     m0650(.A0(mai_mai_n699_), .A1(mai_mai_n693_), .B0(mai_mai_n688_), .Y(mai_mai_n700_));
  NA2        m0651(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n701_));
  NA2        m0652(.A(mai_mai_n369_), .B(mai_mai_n357_), .Y(mai_mai_n702_));
  NO2        m0653(.A(mai_mai_n71_), .B(mai_mai_n108_), .Y(mai_mai_n703_));
  NO2        m0654(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n704_));
  NO4        m0655(.A(mai_mai_n704_), .B(mai_mai_n685_), .C(mai_mai_n703_), .D(mai_mai_n495_), .Y(mai_mai_n705_));
  AOI220     m0656(.A0(mai_mai_n705_), .A1(mai_mai_n702_), .B0(mai_mai_n425_), .B1(mai_mai_n63_), .Y(mai_mai_n706_));
  NO2        m0657(.A(mai_mai_n706_), .B(mai_mai_n701_), .Y(mai_mai_n707_));
  NO2        m0658(.A(mai_mai_n54_), .B(x0), .Y(mai_mai_n708_));
  NA2        m0659(.A(x4), .B(x3), .Y(mai_mai_n709_));
  OAI210     m0660(.A0(mai_mai_n709_), .A1(x8), .B0(mai_mai_n518_), .Y(mai_mai_n710_));
  NA2        m0661(.A(mai_mai_n710_), .B(mai_mai_n708_), .Y(mai_mai_n711_));
  NO2        m0662(.A(mai_mai_n104_), .B(mai_mai_n56_), .Y(mai_mai_n712_));
  NA3        m0663(.A(mai_mai_n712_), .B(mai_mai_n258_), .C(mai_mai_n409_), .Y(mai_mai_n713_));
  AOI210     m0664(.A0(mai_mai_n713_), .A1(mai_mai_n711_), .B0(x2), .Y(mai_mai_n714_));
  INV        m0665(.A(mai_mai_n385_), .Y(mai_mai_n715_));
  NO2        m0666(.A(mai_mai_n412_), .B(x8), .Y(mai_mai_n716_));
  NO2        m0667(.A(mai_mai_n259_), .B(mai_mai_n520_), .Y(mai_mai_n717_));
  AOI210     m0668(.A0(mai_mai_n716_), .A1(mai_mai_n267_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  NO2        m0669(.A(x5), .B(x3), .Y(mai_mai_n719_));
  NA3        m0670(.A(mai_mai_n553_), .B(mai_mai_n719_), .C(x1), .Y(mai_mai_n720_));
  NA2        m0671(.A(mai_mai_n605_), .B(mai_mai_n557_), .Y(mai_mai_n721_));
  OA220      m0672(.A0(mai_mai_n721_), .A1(mai_mai_n581_), .B0(mai_mai_n720_), .B1(mai_mai_n500_), .Y(mai_mai_n722_));
  OAI210     m0673(.A0(mai_mai_n718_), .A1(mai_mai_n715_), .B0(mai_mai_n722_), .Y(mai_mai_n723_));
  OR4        m0674(.A(mai_mai_n723_), .B(mai_mai_n714_), .C(mai_mai_n707_), .D(mai_mai_n700_), .Y(mai_mai_n724_));
  NA2        m0675(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n725_));
  NO2        m0676(.A(mai_mai_n619_), .B(mai_mai_n59_), .Y(mai_mai_n726_));
  NA2        m0677(.A(mai_mai_n726_), .B(mai_mai_n632_), .Y(mai_mai_n727_));
  NO2        m0678(.A(mai_mai_n172_), .B(x6), .Y(mai_mai_n728_));
  NA2        m0679(.A(mai_mai_n728_), .B(mai_mai_n291_), .Y(mai_mai_n729_));
  AOI210     m0680(.A0(mai_mai_n729_), .A1(mai_mai_n727_), .B0(mai_mai_n725_), .Y(mai_mai_n730_));
  AN2        m0681(.A(mai_mai_n473_), .B(mai_mai_n323_), .Y(mai_mai_n731_));
  OAI210     m0682(.A0(mai_mai_n731_), .A1(mai_mai_n730_), .B0(mai_mai_n352_), .Y(mai_mai_n732_));
  NO2        m0683(.A(mai_mai_n308_), .B(mai_mai_n108_), .Y(mai_mai_n733_));
  NO2        m0684(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n734_));
  NA2        m0685(.A(mai_mai_n734_), .B(mai_mai_n71_), .Y(mai_mai_n735_));
  NO2        m0686(.A(mai_mai_n735_), .B(mai_mai_n253_), .Y(mai_mai_n736_));
  NO2        m0687(.A(mai_mai_n71_), .B(x3), .Y(mai_mai_n737_));
  NA3        m0688(.A(mai_mai_n737_), .B(mai_mai_n573_), .C(mai_mai_n56_), .Y(mai_mai_n738_));
  NO2        m0689(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n739_));
  NA2        m0690(.A(mai_mai_n183_), .B(mai_mai_n739_), .Y(mai_mai_n740_));
  NA3        m0691(.A(mai_mai_n605_), .B(mai_mai_n330_), .C(mai_mai_n71_), .Y(mai_mai_n741_));
  NA3        m0692(.A(mai_mai_n741_), .B(mai_mai_n740_), .C(mai_mai_n738_), .Y(mai_mai_n742_));
  OR3        m0693(.A(mai_mai_n742_), .B(mai_mai_n736_), .C(mai_mai_n642_), .Y(mai_mai_n743_));
  NA2        m0694(.A(mai_mai_n743_), .B(mai_mai_n733_), .Y(mai_mai_n744_));
  NA2        m0695(.A(mai_mai_n708_), .B(mai_mai_n632_), .Y(mai_mai_n745_));
  NA4        m0696(.A(mai_mai_n268_), .B(mai_mai_n589_), .C(mai_mai_n222_), .D(mai_mai_n260_), .Y(mai_mai_n746_));
  NA2        m0697(.A(mai_mai_n484_), .B(mai_mai_n67_), .Y(mai_mai_n747_));
  AOI210     m0698(.A0(mai_mai_n746_), .A1(mai_mai_n745_), .B0(mai_mai_n747_), .Y(mai_mai_n748_));
  NA2        m0699(.A(x7), .B(x6), .Y(mai_mai_n749_));
  NA3        m0700(.A(x2), .B(x1), .C(x0), .Y(mai_mai_n750_));
  NO3        m0701(.A(mai_mai_n750_), .B(mai_mai_n749_), .C(mai_mai_n602_), .Y(mai_mai_n751_));
  NA2        m0702(.A(mai_mai_n496_), .B(mai_mai_n149_), .Y(mai_mai_n752_));
  NO2        m0703(.A(x5), .B(x1), .Y(mai_mai_n753_));
  NA2        m0704(.A(mai_mai_n753_), .B(mai_mai_n739_), .Y(mai_mai_n754_));
  NA2        m0705(.A(x4), .B(x0), .Y(mai_mai_n755_));
  NO3        m0706(.A(mai_mai_n57_), .B(x6), .C(x2), .Y(mai_mai_n756_));
  NA2        m0707(.A(mai_mai_n756_), .B(mai_mai_n226_), .Y(mai_mai_n757_));
  OAI220     m0708(.A0(mai_mai_n757_), .A1(mai_mai_n755_), .B0(mai_mai_n754_), .B1(mai_mai_n752_), .Y(mai_mai_n758_));
  NO3        m0709(.A(mai_mai_n758_), .B(mai_mai_n751_), .C(mai_mai_n748_), .Y(mai_mai_n759_));
  NA3        m0710(.A(mai_mai_n759_), .B(mai_mai_n744_), .C(mai_mai_n732_), .Y(mai_mai_n760_));
  AOI210     m0711(.A0(mai_mai_n724_), .A1(mai_mai_n57_), .B0(mai_mai_n760_), .Y(mai07));
  NA2        m0712(.A(mai_mai_n108_), .B(mai_mai_n59_), .Y(mai_mai_n762_));
  NOi21      m0713(.An(mai_mai_n749_), .B(mai_mai_n116_), .Y(mai_mai_n763_));
  NO3        m0714(.A(mai_mai_n57_), .B(x5), .C(x1), .Y(mai_mai_n764_));
  NA2        m0715(.A(mai_mai_n764_), .B(mai_mai_n377_), .Y(mai_mai_n765_));
  NO2        m0716(.A(mai_mai_n57_), .B(mai_mai_n71_), .Y(mai_mai_n766_));
  NO2        m0717(.A(mai_mai_n155_), .B(mai_mai_n109_), .Y(mai_mai_n767_));
  AOI210     m0718(.A0(mai_mai_n766_), .A1(mai_mai_n92_), .B0(mai_mai_n767_), .Y(mai_mai_n768_));
  OAI220     m0719(.A0(mai_mai_n768_), .A1(mai_mai_n137_), .B0(mai_mai_n765_), .B1(mai_mai_n325_), .Y(mai_mai_n769_));
  NA2        m0720(.A(mai_mai_n769_), .B(x2), .Y(mai_mai_n770_));
  NAi21      m0721(.An(mai_mai_n156_), .B(mai_mai_n157_), .Y(mai_mai_n771_));
  NA3        m0722(.A(mai_mai_n771_), .B(mai_mai_n91_), .C(x3), .Y(mai_mai_n772_));
  NO3        m0723(.A(mai_mai_n55_), .B(x3), .C(x1), .Y(mai_mai_n773_));
  NO2        m0724(.A(mai_mai_n513_), .B(x2), .Y(mai_mai_n774_));
  AOI210     m0725(.A0(mai_mai_n774_), .A1(mai_mai_n515_), .B0(mai_mai_n773_), .Y(mai_mai_n775_));
  OAI210     m0726(.A0(mai_mai_n775_), .A1(mai_mai_n650_), .B0(mai_mai_n772_), .Y(mai_mai_n776_));
  NO2        m0727(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n777_));
  NA2        m0728(.A(mai_mai_n777_), .B(mai_mai_n59_), .Y(mai_mai_n778_));
  NA2        m0729(.A(mai_mai_n358_), .B(mai_mai_n352_), .Y(mai_mai_n779_));
  NO2        m0730(.A(x7), .B(x3), .Y(mai_mai_n780_));
  NA2        m0731(.A(mai_mai_n780_), .B(mai_mai_n101_), .Y(mai_mai_n781_));
  AOI210     m0732(.A0(mai_mai_n779_), .A1(mai_mai_n778_), .B0(mai_mai_n781_), .Y(mai_mai_n782_));
  AOI210     m0733(.A0(mai_mai_n776_), .A1(mai_mai_n252_), .B0(mai_mai_n782_), .Y(mai_mai_n783_));
  AOI210     m0734(.A0(mai_mai_n783_), .A1(mai_mai_n770_), .B0(x4), .Y(mai_mai_n784_));
  NA3        m0735(.A(mai_mai_n753_), .B(mai_mai_n321_), .C(mai_mai_n55_), .Y(mai_mai_n785_));
  AOI210     m0736(.A0(mai_mai_n785_), .A1(mai_mai_n598_), .B0(mai_mai_n110_), .Y(mai_mai_n786_));
  XO2        m0737(.A(x5), .B(x1), .Y(mai_mai_n787_));
  NO4        m0738(.A(mai_mai_n787_), .B(mai_mai_n165_), .C(mai_mai_n209_), .D(mai_mai_n55_), .Y(mai_mai_n788_));
  OAI210     m0739(.A0(mai_mai_n788_), .A1(mai_mai_n786_), .B0(mai_mai_n416_), .Y(mai_mai_n789_));
  NO3        m0740(.A(mai_mai_n50_), .B(x2), .C(x0), .Y(mai_mai_n790_));
  NO2        m0741(.A(mai_mai_n311_), .B(mai_mai_n108_), .Y(mai_mai_n791_));
  NA2        m0742(.A(x6), .B(x0), .Y(mai_mai_n792_));
  NO2        m0743(.A(mai_mai_n685_), .B(mai_mai_n792_), .Y(mai_mai_n793_));
  NO2        m0744(.A(mai_mai_n787_), .B(mai_mai_n696_), .Y(mai_mai_n794_));
  OAI210     m0745(.A0(mai_mai_n753_), .A1(mai_mai_n63_), .B0(mai_mai_n57_), .Y(mai_mai_n795_));
  OAI210     m0746(.A0(mai_mai_n795_), .A1(mai_mai_n794_), .B0(mai_mai_n765_), .Y(mai_mai_n796_));
  AOI220     m0747(.A0(mai_mai_n796_), .A1(mai_mai_n790_), .B0(mai_mai_n793_), .B1(mai_mai_n791_), .Y(mai_mai_n797_));
  AOI210     m0748(.A0(mai_mai_n797_), .A1(mai_mai_n789_), .B0(mai_mai_n56_), .Y(mai_mai_n798_));
  NOi21      m0749(.An(mai_mai_n233_), .B(mai_mai_n377_), .Y(mai_mai_n799_));
  NO3        m0750(.A(mai_mai_n799_), .B(mai_mai_n242_), .C(mai_mai_n67_), .Y(mai_mai_n800_));
  NO2        m0751(.A(mai_mai_n311_), .B(x6), .Y(mai_mai_n801_));
  AN2        m0752(.A(mai_mai_n801_), .B(mai_mai_n331_), .Y(mai_mai_n802_));
  OAI210     m0753(.A0(mai_mai_n802_), .A1(mai_mai_n800_), .B0(mai_mai_n59_), .Y(mai_mai_n803_));
  NA2        m0754(.A(mai_mai_n92_), .B(mai_mai_n71_), .Y(mai_mai_n804_));
  NO2        m0755(.A(mai_mai_n804_), .B(mai_mai_n646_), .Y(mai_mai_n805_));
  NAi21      m0756(.An(x8), .B(x7), .Y(mai_mai_n806_));
  NA2        m0757(.A(mai_mai_n799_), .B(mai_mai_n806_), .Y(mai_mai_n807_));
  NA2        m0758(.A(mai_mai_n409_), .B(mai_mai_n110_), .Y(mai_mai_n808_));
  NO2        m0759(.A(mai_mai_n696_), .B(x1), .Y(mai_mai_n809_));
  NO3        m0760(.A(mai_mai_n809_), .B(mai_mai_n808_), .C(mai_mai_n573_), .Y(mai_mai_n810_));
  AOI210     m0761(.A0(mai_mai_n810_), .A1(mai_mai_n807_), .B0(mai_mai_n805_), .Y(mai_mai_n811_));
  AOI210     m0762(.A0(mai_mai_n811_), .A1(mai_mai_n803_), .B0(mai_mai_n144_), .Y(mai_mai_n812_));
  NO2        m0763(.A(x8), .B(x7), .Y(mai_mai_n813_));
  NO2        m0764(.A(mai_mai_n813_), .B(x3), .Y(mai_mai_n814_));
  NA3        m0765(.A(mai_mai_n814_), .B(mai_mai_n366_), .C(x1), .Y(mai_mai_n815_));
  NO2        m0766(.A(x8), .B(mai_mai_n110_), .Y(mai_mai_n816_));
  AOI220     m0767(.A0(mai_mai_n330_), .A1(mai_mai_n352_), .B0(mai_mai_n816_), .B1(mai_mai_n257_), .Y(mai_mai_n817_));
  NO2        m0768(.A(mai_mai_n71_), .B(x4), .Y(mai_mai_n818_));
  NA2        m0769(.A(mai_mai_n818_), .B(mai_mai_n305_), .Y(mai_mai_n819_));
  AOI210     m0770(.A0(mai_mai_n817_), .A1(mai_mai_n815_), .B0(mai_mai_n819_), .Y(mai_mai_n820_));
  NO4        m0771(.A(mai_mai_n820_), .B(mai_mai_n812_), .C(mai_mai_n798_), .D(mai_mai_n784_), .Y(mai08));
  NA2        m0772(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n822_));
  XN2        m0773(.A(x5), .B(x4), .Y(mai_mai_n823_));
  INV        m0774(.A(mai_mai_n823_), .Y(mai_mai_n824_));
  AOI220     m0775(.A0(mai_mai_n824_), .A1(mai_mai_n358_), .B0(mai_mai_n140_), .B1(mai_mai_n56_), .Y(mai_mai_n825_));
  NO2        m0776(.A(mai_mai_n244_), .B(mai_mai_n108_), .Y(mai_mai_n826_));
  AOI210     m0777(.A0(mai_mai_n826_), .A1(mai_mai_n279_), .B0(mai_mai_n193_), .Y(mai_mai_n827_));
  OAI220     m0778(.A0(mai_mai_n827_), .A1(x4), .B0(mai_mai_n825_), .B1(mai_mai_n822_), .Y(mai_mai_n828_));
  NA2        m0779(.A(mai_mai_n828_), .B(mai_mai_n274_), .Y(mai_mai_n829_));
  NO2        m0780(.A(mai_mai_n808_), .B(mai_mai_n618_), .Y(mai_mai_n830_));
  NA2        m0781(.A(mai_mai_n613_), .B(mai_mai_n172_), .Y(mai_mai_n831_));
  OAI220     m0782(.A0(mai_mai_n831_), .A1(mai_mai_n665_), .B0(mai_mai_n486_), .B1(mai_mai_n50_), .Y(mai_mai_n832_));
  AO210      m0783(.A0(mai_mai_n832_), .A1(mai_mai_n345_), .B0(mai_mai_n830_), .Y(mai_mai_n833_));
  NA2        m0784(.A(mai_mai_n279_), .B(mai_mai_n149_), .Y(mai_mai_n834_));
  NA2        m0785(.A(mai_mai_n144_), .B(x7), .Y(mai_mai_n835_));
  OR3        m0786(.A(mai_mai_n750_), .B(mai_mai_n468_), .C(mai_mai_n719_), .Y(mai_mai_n836_));
  OAI220     m0787(.A0(mai_mai_n836_), .A1(mai_mai_n835_), .B0(mai_mai_n834_), .B1(mai_mai_n206_), .Y(mai_mai_n837_));
  AOI210     m0788(.A0(mai_mai_n833_), .A1(mai_mai_n293_), .B0(mai_mai_n837_), .Y(mai_mai_n838_));
  AOI210     m0789(.A0(mai_mai_n838_), .A1(mai_mai_n829_), .B0(mai_mai_n71_), .Y(mai_mai_n839_));
  NO2        m0790(.A(mai_mai_n813_), .B(mai_mai_n110_), .Y(mai_mai_n840_));
  NA2        m0791(.A(mai_mai_n840_), .B(mai_mai_n194_), .Y(mai_mai_n841_));
  OAI210     m0792(.A0(mai_mai_n412_), .A1(mai_mai_n305_), .B0(mai_mai_n345_), .Y(mai_mai_n842_));
  NA2        m0793(.A(mai_mai_n438_), .B(mai_mai_n235_), .Y(mai_mai_n843_));
  NA2        m0794(.A(mai_mai_n716_), .B(mai_mai_n107_), .Y(mai_mai_n844_));
  OAI220     m0795(.A0(mai_mai_n844_), .A1(mai_mai_n843_), .B0(mai_mai_n842_), .B1(mai_mai_n841_), .Y(mai_mai_n845_));
  NA2        m0796(.A(mai_mai_n845_), .B(mai_mai_n289_), .Y(mai_mai_n846_));
  NA2        m0797(.A(mai_mai_n335_), .B(mai_mai_n53_), .Y(mai_mai_n847_));
  NO3        m0798(.A(mai_mai_n412_), .B(mai_mai_n137_), .C(mai_mai_n68_), .Y(mai_mai_n848_));
  NO2        m0799(.A(mai_mai_n704_), .B(mai_mai_n247_), .Y(mai_mai_n849_));
  NO3        m0800(.A(mai_mai_n567_), .B(mai_mai_n469_), .C(mai_mai_n99_), .Y(mai_mai_n850_));
  AO220      m0801(.A0(mai_mai_n850_), .A1(mai_mai_n849_), .B0(mai_mai_n848_), .B1(mai_mai_n847_), .Y(mai_mai_n851_));
  NA2        m0802(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n852_));
  NO3        m0803(.A(mai_mai_n314_), .B(mai_mai_n852_), .C(mai_mai_n288_), .Y(mai_mai_n853_));
  AOI210     m0804(.A0(mai_mai_n851_), .A1(x5), .B0(mai_mai_n853_), .Y(mai_mai_n854_));
  AOI210     m0805(.A0(mai_mai_n854_), .A1(mai_mai_n846_), .B0(mai_mai_n72_), .Y(mai_mai_n855_));
  NO2        m0806(.A(mai_mai_n70_), .B(x3), .Y(mai_mai_n856_));
  OAI210     m0807(.A0(mai_mai_n856_), .A1(mai_mai_n266_), .B0(mai_mai_n147_), .Y(mai_mai_n857_));
  MUX2       m0808(.S(x3), .A(mai_mai_n165_), .B(mai_mai_n771_), .Y(mai_mai_n858_));
  NA2        m0809(.A(mai_mai_n858_), .B(mai_mai_n558_), .Y(mai_mai_n859_));
  NO3        m0810(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n860_));
  INV        m0811(.A(mai_mai_n860_), .Y(mai_mai_n861_));
  AOI210     m0812(.A0(mai_mai_n859_), .A1(mai_mai_n857_), .B0(mai_mai_n861_), .Y(mai_mai_n862_));
  NO3        m0813(.A(x5), .B(x3), .C(mai_mai_n110_), .Y(mai_mai_n863_));
  AOI220     m0814(.A0(mai_mai_n824_), .A1(mai_mai_n310_), .B0(mai_mai_n863_), .B1(mai_mai_n59_), .Y(mai_mai_n864_));
  OR2        m0815(.A(x8), .B(x1), .Y(mai_mai_n865_));
  NO3        m0816(.A(mai_mai_n865_), .B(mai_mai_n864_), .C(mai_mai_n734_), .Y(mai_mai_n866_));
  NAi21      m0817(.An(x4), .B(x1), .Y(mai_mai_n867_));
  NO2        m0818(.A(mai_mai_n867_), .B(x0), .Y(mai_mai_n868_));
  NA2        m0819(.A(mai_mai_n612_), .B(mai_mai_n868_), .Y(mai_mai_n869_));
  NA3        m0820(.A(mai_mai_n55_), .B(x1), .C(x0), .Y(mai_mai_n870_));
  OAI210     m0821(.A0(mai_mai_n870_), .A1(mai_mai_n715_), .B0(mai_mai_n869_), .Y(mai_mai_n871_));
  OAI210     m0822(.A0(mai_mai_n871_), .A1(mai_mai_n866_), .B0(mai_mai_n321_), .Y(mai_mai_n872_));
  AO210      m0823(.A0(mai_mai_n291_), .A1(mai_mai_n266_), .B0(mai_mai_n733_), .Y(mai_mai_n873_));
  NA2        m0824(.A(mai_mai_n108_), .B(mai_mai_n56_), .Y(mai_mai_n874_));
  NO2        m0825(.A(mai_mai_n874_), .B(mai_mai_n262_), .Y(mai_mai_n875_));
  NO2        m0826(.A(mai_mai_n57_), .B(x2), .Y(mai_mai_n876_));
  NO4        m0827(.A(mai_mai_n331_), .B(mai_mai_n876_), .C(mai_mai_n813_), .D(mai_mai_n295_), .Y(mai_mai_n877_));
  AOI220     m0828(.A0(mai_mai_n877_), .A1(mai_mai_n875_), .B0(mai_mai_n873_), .B1(mai_mai_n642_), .Y(mai_mai_n878_));
  NA2        m0829(.A(mai_mai_n878_), .B(mai_mai_n872_), .Y(mai_mai_n879_));
  NO4        m0830(.A(mai_mai_n879_), .B(mai_mai_n862_), .C(mai_mai_n855_), .D(mai_mai_n839_), .Y(mai09));
  NO3        m0831(.A(mai_mai_n787_), .B(mai_mai_n121_), .C(mai_mai_n96_), .Y(mai_mai_n881_));
  AOI220     m0832(.A0(mai_mai_n300_), .A1(mai_mai_n70_), .B0(mai_mai_n588_), .B1(mai_mai_n540_), .Y(mai_mai_n882_));
  OAI210     m0833(.A0(mai_mai_n881_), .A1(x2), .B0(mai_mai_n882_), .Y(mai_mai_n883_));
  AOI210     m0834(.A0(mai_mai_n883_), .A1(mai_mai_n754_), .B0(mai_mai_n447_), .Y(mai_mai_n884_));
  NO2        m0835(.A(mai_mai_n587_), .B(mai_mai_n265_), .Y(mai_mai_n885_));
  NO2        m0836(.A(mai_mai_n753_), .B(mai_mai_n341_), .Y(mai_mai_n886_));
  NO3        m0837(.A(mai_mai_n604_), .B(mai_mai_n102_), .C(mai_mai_n110_), .Y(mai_mai_n887_));
  AO220      m0838(.A0(mai_mai_n887_), .A1(mai_mai_n886_), .B0(mai_mai_n885_), .B1(mai_mai_n619_), .Y(mai_mai_n888_));
  OAI210     m0839(.A0(mai_mai_n888_), .A1(mai_mai_n884_), .B0(x4), .Y(mai_mai_n889_));
  NO2        m0840(.A(mai_mai_n396_), .B(mai_mai_n281_), .Y(mai_mai_n890_));
  NO2        m0841(.A(mai_mai_n192_), .B(mai_mai_n108_), .Y(mai_mai_n891_));
  AOI220     m0842(.A0(mai_mai_n891_), .A1(mai_mai_n126_), .B0(mai_mai_n890_), .B1(mai_mai_n625_), .Y(mai_mai_n892_));
  NO2        m0843(.A(mai_mai_n787_), .B(mai_mai_n96_), .Y(mai_mai_n893_));
  NAi21      m0844(.An(x0), .B(x2), .Y(mai_mai_n894_));
  NO2        m0845(.A(mai_mai_n304_), .B(mai_mai_n894_), .Y(mai_mai_n895_));
  OAI210     m0846(.A0(mai_mai_n478_), .A1(mai_mai_n276_), .B0(mai_mai_n192_), .Y(mai_mai_n896_));
  AOI210     m0847(.A0(mai_mai_n168_), .A1(mai_mai_n806_), .B0(mai_mai_n357_), .Y(mai_mai_n897_));
  AOI220     m0848(.A0(mai_mai_n897_), .A1(mai_mai_n896_), .B0(mai_mai_n895_), .B1(mai_mai_n893_), .Y(mai_mai_n898_));
  OAI210     m0849(.A0(mai_mai_n892_), .A1(mai_mai_n55_), .B0(mai_mai_n898_), .Y(mai_mai_n899_));
  NA2        m0850(.A(mai_mai_n899_), .B(mai_mai_n56_), .Y(mai_mai_n900_));
  NO2        m0851(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n901_));
  INV        m0852(.A(mai_mai_n126_), .Y(mai_mai_n902_));
  NA2        m0853(.A(mai_mai_n753_), .B(mai_mai_n55_), .Y(mai_mai_n903_));
  AOI210     m0854(.A0(x6), .A1(x1), .B0(x5), .Y(mai_mai_n904_));
  OAI210     m0855(.A0(mai_mai_n904_), .A1(mai_mai_n334_), .B0(x2), .Y(mai_mai_n905_));
  AOI210     m0856(.A0(mai_mai_n905_), .A1(mai_mai_n903_), .B0(mai_mai_n902_), .Y(mai_mai_n906_));
  NA2        m0857(.A(mai_mai_n557_), .B(mai_mai_n55_), .Y(mai_mai_n907_));
  NO4        m0858(.A(mai_mai_n57_), .B(x6), .C(x5), .D(x1), .Y(mai_mai_n908_));
  NO2        m0859(.A(mai_mai_n232_), .B(mai_mai_n386_), .Y(mai_mai_n909_));
  NO2        m0860(.A(mai_mai_n311_), .B(mai_mai_n148_), .Y(mai_mai_n910_));
  NO3        m0861(.A(mai_mai_n910_), .B(mai_mai_n909_), .C(mai_mai_n908_), .Y(mai_mai_n911_));
  OAI220     m0862(.A0(mai_mai_n911_), .A1(mai_mai_n55_), .B0(mai_mai_n907_), .B1(mai_mai_n459_), .Y(mai_mai_n912_));
  OAI210     m0863(.A0(mai_mai_n912_), .A1(mai_mai_n906_), .B0(mai_mai_n901_), .Y(mai_mai_n913_));
  NO2        m0864(.A(mai_mai_n405_), .B(mai_mai_n108_), .Y(mai_mai_n914_));
  NO2        m0865(.A(mai_mai_n335_), .B(mai_mai_n495_), .Y(mai_mai_n915_));
  AOI220     m0866(.A0(mai_mai_n915_), .A1(mai_mai_n914_), .B0(mai_mai_n210_), .B1(mai_mai_n230_), .Y(mai_mai_n916_));
  NA4        m0867(.A(mai_mai_n916_), .B(mai_mai_n913_), .C(mai_mai_n900_), .D(mai_mai_n889_), .Y(mai_mai_n917_));
  NA2        m0868(.A(mai_mai_n917_), .B(mai_mai_n50_), .Y(mai_mai_n918_));
  NO2        m0869(.A(mai_mai_n380_), .B(mai_mai_n161_), .Y(mai_mai_n919_));
  NA2        m0870(.A(mai_mai_n241_), .B(mai_mai_n588_), .Y(mai_mai_n920_));
  OAI210     m0871(.A0(mai_mai_n433_), .A1(mai_mai_n816_), .B0(mai_mai_n920_), .Y(mai_mai_n921_));
  OAI210     m0872(.A0(mai_mai_n921_), .A1(mai_mai_n919_), .B0(x0), .Y(mai_mai_n922_));
  NO3        m0873(.A(x8), .B(x7), .C(x2), .Y(mai_mai_n923_));
  NO3        m0874(.A(mai_mai_n57_), .B(x5), .C(x2), .Y(mai_mai_n924_));
  OAI210     m0875(.A0(mai_mai_n924_), .A1(mai_mai_n923_), .B0(mai_mai_n515_), .Y(mai_mai_n925_));
  AOI210     m0876(.A0(mai_mai_n925_), .A1(mai_mai_n922_), .B0(x4), .Y(mai_mai_n926_));
  NO2        m0877(.A(mai_mai_n426_), .B(mai_mai_n147_), .Y(mai_mai_n927_));
  NO2        m0878(.A(mai_mai_n52_), .B(x2), .Y(mai_mai_n928_));
  NO2        m0879(.A(mai_mai_n108_), .B(mai_mai_n56_), .Y(mai_mai_n929_));
  NA2        m0880(.A(mai_mai_n929_), .B(x8), .Y(mai_mai_n930_));
  OAI210     m0881(.A0(mai_mai_n927_), .A1(mai_mai_n926_), .B0(mai_mai_n617_), .Y(mai_mai_n931_));
  NO2        m0882(.A(mai_mai_n261_), .B(mai_mai_n119_), .Y(mai_mai_n932_));
  OAI210     m0883(.A0(x4), .A1(x2), .B0(x0), .Y(mai_mai_n933_));
  NA3        m0884(.A(mai_mai_n606_), .B(mai_mai_n618_), .C(mai_mai_n346_), .Y(mai_mai_n934_));
  OAI210     m0885(.A0(mai_mai_n933_), .A1(mai_mai_n288_), .B0(mai_mai_n53_), .Y(mai_mai_n935_));
  AOI210     m0886(.A0(mai_mai_n934_), .A1(mai_mai_n933_), .B0(mai_mai_n935_), .Y(mai_mai_n936_));
  OAI210     m0887(.A0(mai_mai_n936_), .A1(mai_mai_n932_), .B0(mai_mai_n330_), .Y(mai_mai_n937_));
  AOI220     m0888(.A0(mai_mai_n667_), .A1(mai_mai_n350_), .B0(mai_mai_n352_), .B1(mai_mai_n93_), .Y(mai_mai_n938_));
  NA2        m0889(.A(mai_mai_n93_), .B(x5), .Y(mai_mai_n939_));
  OAI220     m0890(.A0(mai_mai_n939_), .A1(mai_mai_n865_), .B0(mai_mai_n938_), .B1(mai_mai_n322_), .Y(mai_mai_n940_));
  NA2        m0891(.A(mai_mai_n940_), .B(mai_mai_n68_), .Y(mai_mai_n941_));
  NA2        m0892(.A(mai_mai_n409_), .B(mai_mai_n771_), .Y(mai_mai_n942_));
  NA2        m0893(.A(mai_mai_n252_), .B(mai_mai_n165_), .Y(mai_mai_n943_));
  AO210      m0894(.A0(mai_mai_n943_), .A1(mai_mai_n942_), .B0(mai_mai_n134_), .Y(mai_mai_n944_));
  NO2        m0895(.A(mai_mai_n439_), .B(x2), .Y(mai_mai_n945_));
  NO2        m0896(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n946_));
  NA2        m0897(.A(mai_mai_n946_), .B(x5), .Y(mai_mai_n947_));
  NO2        m0898(.A(mai_mai_n947_), .B(mai_mai_n60_), .Y(mai_mai_n948_));
  AOI220     m0899(.A0(mai_mai_n948_), .A1(mai_mai_n945_), .B0(mai_mai_n668_), .B1(mai_mai_n245_), .Y(mai_mai_n949_));
  NA4        m0900(.A(mai_mai_n949_), .B(mai_mai_n944_), .C(mai_mai_n941_), .D(mai_mai_n937_), .Y(mai_mai_n950_));
  NO4        m0901(.A(mai_mai_n934_), .B(mai_mai_n634_), .C(mai_mai_n459_), .D(mai_mai_n50_), .Y(mai_mai_n951_));
  AOI220     m0902(.A0(mai_mai_n605_), .A1(mai_mai_n604_), .B0(mai_mai_n282_), .B1(x5), .Y(mai_mai_n952_));
  NO2        m0903(.A(mai_mai_n676_), .B(mai_mai_n192_), .Y(mai_mai_n953_));
  NA3        m0904(.A(mai_mai_n953_), .B(mai_mai_n669_), .C(x7), .Y(mai_mai_n954_));
  OAI210     m0905(.A0(mai_mai_n952_), .A1(mai_mai_n351_), .B0(mai_mai_n954_), .Y(mai_mai_n955_));
  OAI210     m0906(.A0(mai_mai_n955_), .A1(mai_mai_n951_), .B0(mai_mai_n82_), .Y(mai_mai_n956_));
  NA2        m0907(.A(mai_mai_n777_), .B(x2), .Y(mai_mai_n957_));
  NO2        m0908(.A(mai_mai_n957_), .B(mai_mai_n58_), .Y(mai_mai_n958_));
  NO2        m0909(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n959_));
  NAi21      m0910(.An(x1), .B(x4), .Y(mai_mai_n960_));
  NA2        m0911(.A(mai_mai_n960_), .B(mai_mai_n867_), .Y(mai_mai_n961_));
  NO3        m0912(.A(mai_mai_n961_), .B(mai_mai_n203_), .C(mai_mai_n959_), .Y(mai_mai_n962_));
  OAI210     m0913(.A0(mai_mai_n962_), .A1(mai_mai_n958_), .B0(mai_mai_n416_), .Y(mai_mai_n963_));
  NA3        m0914(.A(mai_mai_n399_), .B(mai_mai_n753_), .C(mai_mai_n57_), .Y(mai_mai_n964_));
  NA3        m0915(.A(mai_mai_n964_), .B(mai_mai_n963_), .C(mai_mai_n956_), .Y(mai_mai_n965_));
  AOI210     m0916(.A0(mai_mai_n950_), .A1(x6), .B0(mai_mai_n965_), .Y(mai_mai_n966_));
  NA3        m0917(.A(mai_mai_n966_), .B(mai_mai_n931_), .C(mai_mai_n918_), .Y(mai10));
  NO2        m0918(.A(x4), .B(x1), .Y(mai_mai_n968_));
  NO2        m0919(.A(mai_mai_n968_), .B(mai_mai_n149_), .Y(mai_mai_n969_));
  NA3        m0920(.A(x5), .B(x4), .C(x0), .Y(mai_mai_n970_));
  OAI220     m0921(.A0(mai_mai_n970_), .A1(mai_mai_n277_), .B0(mai_mai_n704_), .B1(mai_mai_n249_), .Y(mai_mai_n971_));
  NA2        m0922(.A(mai_mai_n971_), .B(mai_mai_n969_), .Y(mai_mai_n972_));
  NO3        m0923(.A(mai_mai_n358_), .B(mai_mai_n322_), .C(mai_mai_n92_), .Y(mai_mai_n973_));
  NA3        m0924(.A(mai_mai_n973_), .B(mai_mai_n384_), .C(mai_mai_n62_), .Y(mai_mai_n974_));
  AOI210     m0925(.A0(mai_mai_n974_), .A1(mai_mai_n972_), .B0(mai_mai_n304_), .Y(mai_mai_n975_));
  NOi21      m0926(.An(mai_mai_n260_), .B(mai_mai_n140_), .Y(mai_mai_n976_));
  AOI210     m0927(.A0(mai_mai_n501_), .A1(mai_mai_n619_), .B0(mai_mai_n331_), .Y(mai_mai_n977_));
  NO2        m0928(.A(mai_mai_n901_), .B(mai_mai_n344_), .Y(mai_mai_n978_));
  NOi31      m0929(.An(mai_mai_n978_), .B(mai_mai_n977_), .C(mai_mai_n976_), .Y(mai_mai_n979_));
  NA2        m0930(.A(x4), .B(mai_mai_n110_), .Y(mai_mai_n980_));
  NO2        m0931(.A(mai_mai_n325_), .B(mai_mai_n980_), .Y(mai_mai_n981_));
  NA2        m0932(.A(mai_mai_n99_), .B(x5), .Y(mai_mai_n982_));
  NO3        m0933(.A(mai_mai_n982_), .B(mai_mai_n111_), .C(mai_mai_n55_), .Y(mai_mai_n983_));
  NO3        m0934(.A(mai_mai_n983_), .B(mai_mai_n981_), .C(mai_mai_n979_), .Y(mai_mai_n984_));
  NA2        m0935(.A(mai_mai_n959_), .B(mai_mai_n50_), .Y(mai_mai_n985_));
  NA2        m0936(.A(mai_mai_n605_), .B(mai_mai_n273_), .Y(mai_mai_n986_));
  NO2        m0937(.A(mai_mai_n986_), .B(mai_mai_n985_), .Y(mai_mai_n987_));
  OAI220     m0938(.A0(mai_mai_n930_), .A1(mai_mai_n107_), .B0(mai_mai_n874_), .B1(mai_mai_n447_), .Y(mai_mai_n988_));
  AOI210     m0939(.A0(mai_mai_n988_), .A1(mai_mai_n279_), .B0(mai_mai_n987_), .Y(mai_mai_n989_));
  OAI210     m0940(.A0(mai_mai_n984_), .A1(mai_mai_n386_), .B0(mai_mai_n989_), .Y(mai_mai_n990_));
  OAI210     m0941(.A0(mai_mai_n990_), .A1(mai_mai_n975_), .B0(x7), .Y(mai_mai_n991_));
  NA2        m0942(.A(mai_mai_n55_), .B(mai_mai_n71_), .Y(mai_mai_n992_));
  AOI210     m0943(.A0(mai_mai_n447_), .A1(mai_mai_n357_), .B0(mai_mai_n980_), .Y(mai_mai_n993_));
  NO3        m0944(.A(mai_mai_n449_), .B(mai_mai_n894_), .C(x5), .Y(mai_mai_n994_));
  OAI210     m0945(.A0(mai_mai_n994_), .A1(mai_mai_n993_), .B0(mai_mai_n992_), .Y(mai_mai_n995_));
  NO2        m0946(.A(mai_mai_n358_), .B(mai_mai_n143_), .Y(mai_mai_n996_));
  NA2        m0947(.A(mai_mai_n996_), .B(mai_mai_n427_), .Y(mai_mai_n997_));
  AOI210     m0948(.A0(mai_mai_n997_), .A1(mai_mai_n995_), .B0(x3), .Y(mai_mai_n998_));
  NA2        m0949(.A(mai_mai_n696_), .B(mai_mai_n252_), .Y(mai_mai_n999_));
  NO2        m0950(.A(x5), .B(mai_mai_n110_), .Y(mai_mai_n1000_));
  OAI210     m0951(.A0(mai_mai_n1000_), .A1(mai_mai_n239_), .B0(mai_mai_n939_), .Y(mai_mai_n1001_));
  NA3        m0952(.A(mai_mai_n464_), .B(mai_mai_n132_), .C(mai_mai_n427_), .Y(mai_mai_n1002_));
  OAI210     m0953(.A0(mai_mai_n449_), .A1(mai_mai_n215_), .B0(mai_mai_n1002_), .Y(mai_mai_n1003_));
  AOI210     m0954(.A0(mai_mai_n1001_), .A1(mai_mai_n258_), .B0(mai_mai_n1003_), .Y(mai_mai_n1004_));
  OAI220     m0955(.A0(mai_mai_n1004_), .A1(mai_mai_n59_), .B0(mai_mai_n999_), .B1(mai_mai_n709_), .Y(mai_mai_n1005_));
  OAI210     m0956(.A0(mai_mai_n1005_), .A1(mai_mai_n998_), .B0(mai_mai_n946_), .Y(mai_mai_n1006_));
  NO2        m0957(.A(x4), .B(x3), .Y(mai_mai_n1007_));
  NO3        m0958(.A(mai_mai_n1007_), .B(mai_mai_n345_), .C(mai_mai_n87_), .Y(mai_mai_n1008_));
  OAI210     m0959(.A0(mai_mai_n1008_), .A1(mai_mai_n278_), .B0(mai_mai_n438_), .Y(mai_mai_n1009_));
  AOI210     m0960(.A0(mai_mai_n400_), .A1(mai_mai_n129_), .B0(mai_mai_n253_), .Y(mai_mai_n1010_));
  NA2        m0961(.A(mai_mai_n968_), .B(mai_mai_n55_), .Y(mai_mai_n1011_));
  NO2        m0962(.A(mai_mai_n1011_), .B(mai_mai_n982_), .Y(mai_mai_n1012_));
  NO2        m0963(.A(mai_mai_n525_), .B(mai_mai_n363_), .Y(mai_mai_n1013_));
  NO3        m0964(.A(x4), .B(mai_mai_n110_), .C(mai_mai_n59_), .Y(mai_mai_n1014_));
  NO2        m0965(.A(mai_mai_n439_), .B(x1), .Y(mai_mai_n1015_));
  NOi31      m0966(.An(mai_mai_n1014_), .B(mai_mai_n1015_), .C(mai_mai_n1013_), .Y(mai_mai_n1016_));
  NA2        m0967(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n1017_));
  NO4        m0968(.A(mai_mai_n969_), .B(mai_mai_n514_), .C(mai_mai_n1017_), .D(x2), .Y(mai_mai_n1018_));
  NO4        m0969(.A(mai_mai_n1018_), .B(mai_mai_n1016_), .C(mai_mai_n1012_), .D(mai_mai_n1010_), .Y(mai_mai_n1019_));
  AOI210     m0970(.A0(mai_mai_n1019_), .A1(mai_mai_n1009_), .B0(mai_mai_n209_), .Y(mai_mai_n1020_));
  NO2        m0971(.A(mai_mai_n665_), .B(mai_mai_n500_), .Y(mai_mai_n1021_));
  NO2        m0972(.A(x6), .B(x2), .Y(mai_mai_n1022_));
  NO3        m0973(.A(mai_mai_n1022_), .B(mai_mai_n696_), .C(mai_mai_n60_), .Y(mai_mai_n1023_));
  NA2        m0974(.A(mai_mai_n1023_), .B(mai_mai_n272_), .Y(mai_mai_n1024_));
  NO2        m0975(.A(mai_mai_n874_), .B(mai_mai_n447_), .Y(mai_mai_n1025_));
  NA3        m0976(.A(x4), .B(x3), .C(mai_mai_n110_), .Y(mai_mai_n1026_));
  NO3        m0977(.A(mai_mai_n1026_), .B(mai_mai_n702_), .C(mai_mai_n464_), .Y(mai_mai_n1027_));
  AOI210     m0978(.A0(mai_mai_n1025_), .A1(mai_mai_n471_), .B0(mai_mai_n1027_), .Y(mai_mai_n1028_));
  AOI210     m0979(.A0(mai_mai_n1028_), .A1(mai_mai_n1024_), .B0(mai_mai_n459_), .Y(mai_mai_n1029_));
  NO2        m0980(.A(mai_mai_n55_), .B(mai_mai_n56_), .Y(mai_mai_n1030_));
  OAI220     m0981(.A0(mai_mai_n824_), .A1(mai_mai_n461_), .B0(mai_mai_n755_), .B1(mai_mai_n129_), .Y(mai_mai_n1031_));
  NOi21      m0982(.An(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n1032_));
  NO3        m0983(.A(mai_mai_n346_), .B(mai_mai_n325_), .C(mai_mai_n1032_), .Y(mai_mai_n1033_));
  AOI220     m0984(.A0(mai_mai_n1033_), .A1(mai_mai_n257_), .B0(mai_mai_n1031_), .B1(mai_mai_n116_), .Y(mai_mai_n1034_));
  NO2        m0985(.A(mai_mai_n1034_), .B(mai_mai_n1030_), .Y(mai_mai_n1035_));
  NA2        m0986(.A(mai_mai_n518_), .B(mai_mai_n262_), .Y(mai_mai_n1036_));
  NO2        m0987(.A(mai_mai_n486_), .B(mai_mai_n587_), .Y(mai_mai_n1037_));
  NA3        m0988(.A(mai_mai_n1037_), .B(mai_mai_n1036_), .C(mai_mai_n55_), .Y(mai_mai_n1038_));
  NO2        m0989(.A(mai_mai_n184_), .B(mai_mai_n110_), .Y(mai_mai_n1039_));
  NA3        m0990(.A(mai_mai_n1039_), .B(mai_mai_n183_), .C(mai_mai_n123_), .Y(mai_mai_n1040_));
  NA2        m0991(.A(mai_mai_n1040_), .B(mai_mai_n1038_), .Y(mai_mai_n1041_));
  NO4        m0992(.A(mai_mai_n1041_), .B(mai_mai_n1035_), .C(mai_mai_n1029_), .D(mai_mai_n1020_), .Y(mai_mai_n1042_));
  NA3        m0993(.A(mai_mai_n1042_), .B(mai_mai_n1006_), .C(mai_mai_n991_), .Y(mai11));
  NA2        m0994(.A(mai_mai_n378_), .B(mai_mai_n92_), .Y(mai_mai_n1044_));
  INV        m0995(.A(mai_mai_n895_), .Y(mai_mai_n1045_));
  NO2        m0996(.A(mai_mai_n1044_), .B(mai_mai_n367_), .Y(mai_mai_n1046_));
  NO2        m0997(.A(mai_mai_n771_), .B(x5), .Y(mai_mai_n1047_));
  NO2        m0998(.A(mai_mai_n169_), .B(mai_mai_n531_), .Y(mai_mai_n1048_));
  AOI220     m0999(.A0(mai_mai_n1048_), .A1(mai_mai_n1047_), .B0(mai_mai_n1046_), .B1(x5), .Y(mai_mai_n1049_));
  OAI220     m1000(.A0(mai_mai_n976_), .A1(mai_mai_n218_), .B0(mai_mai_n216_), .B1(mai_mai_n184_), .Y(mai_mai_n1050_));
  NO2        m1001(.A(mai_mai_n342_), .B(mai_mai_n428_), .Y(mai_mai_n1051_));
  AOI220     m1002(.A0(mai_mai_n1051_), .A1(mai_mai_n182_), .B0(mai_mai_n1050_), .B1(mai_mai_n165_), .Y(mai_mai_n1052_));
  NO2        m1003(.A(mai_mai_n1052_), .B(mai_mai_n449_), .Y(mai_mai_n1053_));
  NO2        m1004(.A(mai_mai_n55_), .B(mai_mai_n108_), .Y(mai_mai_n1054_));
  NA2        m1005(.A(mai_mai_n279_), .B(mai_mai_n1054_), .Y(mai_mai_n1055_));
  NO2        m1006(.A(mai_mai_n71_), .B(x1), .Y(mai_mai_n1056_));
  NA2        m1007(.A(mai_mai_n1056_), .B(mai_mai_n78_), .Y(mai_mai_n1057_));
  OA220      m1008(.A0(mai_mai_n1057_), .A1(mai_mai_n613_), .B0(mai_mai_n1055_), .B1(mai_mai_n531_), .Y(mai_mai_n1058_));
  NO2        m1009(.A(mai_mai_n1058_), .B(mai_mai_n709_), .Y(mai_mai_n1059_));
  NO2        m1010(.A(mai_mai_n305_), .B(mai_mai_n53_), .Y(mai_mai_n1060_));
  NO2        m1011(.A(mai_mai_n438_), .B(x3), .Y(mai_mai_n1061_));
  NA3        m1012(.A(mai_mai_n1061_), .B(mai_mai_n1060_), .C(mai_mai_n894_), .Y(mai_mai_n1062_));
  AOI210     m1013(.A0(mai_mai_n1062_), .A1(mai_mai_n943_), .B0(mai_mai_n398_), .Y(mai_mai_n1063_));
  NA2        m1014(.A(mai_mai_n110_), .B(x1), .Y(mai_mai_n1064_));
  NO2        m1015(.A(mai_mai_n619_), .B(mai_mai_n221_), .Y(mai_mai_n1065_));
  NA4        m1016(.A(mai_mai_n1065_), .B(mai_mai_n886_), .C(mai_mai_n468_), .D(mai_mai_n1064_), .Y(mai_mai_n1066_));
  NA3        m1017(.A(x6), .B(x5), .C(mai_mai_n110_), .Y(mai_mai_n1067_));
  NO2        m1018(.A(mai_mai_n1067_), .B(mai_mai_n277_), .Y(mai_mai_n1068_));
  NO2        m1019(.A(mai_mai_n449_), .B(x0), .Y(mai_mai_n1069_));
  NOi31      m1020(.An(mai_mai_n1069_), .B(mai_mai_n174_), .C(mai_mai_n51_), .Y(mai_mai_n1070_));
  AOI210     m1021(.A0(mai_mai_n1068_), .A1(mai_mai_n180_), .B0(mai_mai_n1070_), .Y(mai_mai_n1071_));
  NA2        m1022(.A(mai_mai_n1071_), .B(mai_mai_n1066_), .Y(mai_mai_n1072_));
  NO4        m1023(.A(mai_mai_n1072_), .B(mai_mai_n1063_), .C(mai_mai_n1059_), .D(mai_mai_n1053_), .Y(mai_mai_n1073_));
  OAI210     m1024(.A0(mai_mai_n1049_), .A1(mai_mai_n144_), .B0(mai_mai_n1073_), .Y(mai_mai_n1074_));
  NA2        m1025(.A(mai_mai_n865_), .B(mai_mai_n87_), .Y(mai_mai_n1075_));
  NO3        m1026(.A(mai_mai_n465_), .B(mai_mai_n777_), .C(mai_mai_n124_), .Y(mai_mai_n1076_));
  AOI210     m1027(.A0(mai_mai_n1075_), .A1(mai_mai_n101_), .B0(mai_mai_n1076_), .Y(mai_mai_n1077_));
  NO2        m1028(.A(x8), .B(x1), .Y(mai_mai_n1078_));
  NO3        m1029(.A(mai_mai_n1078_), .B(mai_mai_n688_), .C(mai_mai_n451_), .Y(mai_mai_n1079_));
  OAI210     m1030(.A0(mai_mai_n77_), .A1(mai_mai_n53_), .B0(mai_mai_n1079_), .Y(mai_mai_n1080_));
  OAI210     m1031(.A0(mai_mai_n1077_), .A1(x3), .B0(mai_mai_n1080_), .Y(mai_mai_n1081_));
  NO2        m1032(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n1082_));
  OAI210     m1033(.A0(mai_mai_n1082_), .A1(x2), .B0(mai_mai_n235_), .Y(mai_mai_n1083_));
  NO2        m1034(.A(mai_mai_n606_), .B(mai_mai_n233_), .Y(mai_mai_n1084_));
  NA2        m1035(.A(mai_mai_n1084_), .B(mai_mai_n1083_), .Y(mai_mai_n1085_));
  NO2        m1036(.A(mai_mai_n518_), .B(x4), .Y(mai_mai_n1086_));
  NO3        m1037(.A(mai_mai_n55_), .B(x6), .C(x1), .Y(mai_mai_n1087_));
  NOi21      m1038(.An(mai_mai_n1087_), .B(mai_mai_n486_), .Y(mai_mai_n1088_));
  AOI210     m1039(.A0(mai_mai_n1086_), .A1(mai_mai_n577_), .B0(mai_mai_n1088_), .Y(mai_mai_n1089_));
  NA2        m1040(.A(mai_mai_n1089_), .B(mai_mai_n1085_), .Y(mai_mai_n1090_));
  AOI210     m1041(.A0(mai_mai_n1081_), .A1(x2), .B0(mai_mai_n1090_), .Y(mai_mai_n1091_));
  NO2        m1042(.A(mai_mai_n233_), .B(x2), .Y(mai_mai_n1092_));
  NA2        m1043(.A(mai_mai_n1092_), .B(mai_mai_n1007_), .Y(mai_mai_n1093_));
  NOi21      m1044(.An(mai_mai_n389_), .B(mai_mai_n566_), .Y(mai_mai_n1094_));
  NO3        m1045(.A(mai_mai_n1094_), .B(mai_mai_n605_), .C(mai_mai_n325_), .Y(mai_mai_n1095_));
  NA2        m1046(.A(x8), .B(mai_mai_n110_), .Y(mai_mai_n1096_));
  OAI220     m1047(.A0(mai_mai_n709_), .A1(mai_mai_n1096_), .B0(mai_mai_n325_), .B1(mai_mai_n384_), .Y(mai_mai_n1097_));
  OAI210     m1048(.A0(mai_mai_n1097_), .A1(mai_mai_n1095_), .B0(mai_mai_n71_), .Y(mai_mai_n1098_));
  NO2        m1049(.A(mai_mai_n108_), .B(x1), .Y(mai_mai_n1099_));
  NA2        m1050(.A(mai_mai_n1099_), .B(x7), .Y(mai_mai_n1100_));
  AOI210     m1051(.A0(mai_mai_n1098_), .A1(mai_mai_n1093_), .B0(mai_mai_n1100_), .Y(mai_mai_n1101_));
  NA2        m1052(.A(mai_mai_n84_), .B(mai_mai_n71_), .Y(mai_mai_n1102_));
  INV        m1053(.A(mai_mai_n250_), .Y(mai_mai_n1103_));
  INV        m1054(.A(mai_mai_n1101_), .Y(mai_mai_n1104_));
  OAI210     m1055(.A0(mai_mai_n1091_), .A1(mai_mai_n852_), .B0(mai_mai_n1104_), .Y(mai_mai_n1105_));
  AO210      m1056(.A0(mai_mai_n1074_), .A1(mai_mai_n57_), .B0(mai_mai_n1105_), .Y(mai12));
  NA2        m1057(.A(mai_mai_n885_), .B(mai_mai_n249_), .Y(mai_mai_n1107_));
  NO2        m1058(.A(mai_mai_n623_), .B(x7), .Y(mai_mai_n1108_));
  NA2        m1059(.A(mai_mai_n1108_), .B(mai_mai_n278_), .Y(mai_mai_n1109_));
  NA2        m1060(.A(mai_mai_n701_), .B(mai_mai_n874_), .Y(mai_mai_n1110_));
  AOI210     m1061(.A0(mai_mai_n1109_), .A1(mai_mai_n1107_), .B0(mai_mai_n1110_), .Y(mai_mai_n1111_));
  NOi21      m1062(.An(mai_mai_n405_), .B(mai_mai_n553_), .Y(mai_mai_n1112_));
  NO2        m1063(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n1113_));
  NO2        m1064(.A(mai_mai_n606_), .B(mai_mai_n1113_), .Y(mai_mai_n1114_));
  NO3        m1065(.A(mai_mai_n867_), .B(mai_mai_n112_), .C(mai_mai_n99_), .Y(mai_mai_n1115_));
  AOI210     m1066(.A0(mai_mai_n1114_), .A1(mai_mai_n1015_), .B0(mai_mai_n1115_), .Y(mai_mai_n1116_));
  NA2        m1067(.A(mai_mai_n1054_), .B(mai_mai_n56_), .Y(mai_mai_n1117_));
  OAI220     m1068(.A0(mai_mai_n1117_), .A1(mai_mai_n578_), .B0(mai_mai_n1116_), .B1(mai_mai_n1112_), .Y(mai_mai_n1118_));
  OAI210     m1069(.A0(mai_mai_n1118_), .A1(mai_mai_n1111_), .B0(mai_mai_n582_), .Y(mai_mai_n1119_));
  NA2        m1070(.A(mai_mai_n87_), .B(x5), .Y(mai_mai_n1120_));
  OAI210     m1071(.A0(mai_mai_n1120_), .A1(mai_mai_n325_), .B0(mai_mai_n720_), .Y(mai_mai_n1121_));
  AOI210     m1072(.A0(mai_mai_n826_), .A1(mai_mai_n118_), .B0(mai_mai_n1121_), .Y(mai_mai_n1122_));
  NA2        m1073(.A(mai_mai_n604_), .B(mai_mai_n53_), .Y(mai_mai_n1123_));
  NA2        m1074(.A(mai_mai_n288_), .B(mai_mai_n50_), .Y(mai_mai_n1124_));
  OAI220     m1075(.A0(mai_mai_n1124_), .A1(mai_mai_n311_), .B0(mai_mai_n1123_), .B1(mai_mai_n137_), .Y(mai_mai_n1125_));
  NO2        m1076(.A(mai_mai_n1075_), .B(mai_mai_n513_), .Y(mai_mai_n1126_));
  NO4        m1077(.A(mai_mai_n241_), .B(mai_mai_n272_), .C(mai_mai_n60_), .D(mai_mai_n57_), .Y(mai_mai_n1127_));
  AOI220     m1078(.A0(mai_mai_n1127_), .A1(mai_mai_n1126_), .B0(mai_mai_n1125_), .B1(mai_mai_n56_), .Y(mai_mai_n1128_));
  OAI210     m1079(.A0(mai_mai_n1122_), .A1(mai_mai_n64_), .B0(mai_mai_n1128_), .Y(mai_mai_n1129_));
  NO2        m1080(.A(mai_mai_n57_), .B(x0), .Y(mai_mai_n1130_));
  NO2        m1081(.A(mai_mai_n665_), .B(mai_mai_n322_), .Y(mai_mai_n1131_));
  NO2        m1082(.A(mai_mai_n755_), .B(x3), .Y(mai_mai_n1132_));
  NO2        m1083(.A(mai_mai_n663_), .B(x8), .Y(mai_mai_n1133_));
  NA2        m1084(.A(mai_mai_n1131_), .B(mai_mai_n1130_), .Y(mai_mai_n1134_));
  AOI210     m1085(.A0(mai_mai_n688_), .A1(mai_mai_n249_), .B0(x7), .Y(mai_mai_n1135_));
  NO3        m1086(.A(mai_mai_n1135_), .B(mai_mai_n607_), .C(x8), .Y(mai_mai_n1136_));
  NA4        m1087(.A(mai_mai_n667_), .B(mai_mai_n659_), .C(mai_mai_n206_), .D(x0), .Y(mai_mai_n1137_));
  OAI220     m1088(.A0(mai_mai_n1137_), .A1(mai_mai_n1136_), .B0(mai_mai_n1134_), .B1(mai_mai_n576_), .Y(mai_mai_n1138_));
  AOI210     m1089(.A0(mai_mai_n1129_), .A1(mai_mai_n1022_), .B0(mai_mai_n1138_), .Y(mai_mai_n1139_));
  NO2        m1090(.A(mai_mai_n257_), .B(x8), .Y(mai_mai_n1140_));
  NO2        m1091(.A(mai_mai_n946_), .B(mai_mai_n100_), .Y(mai_mai_n1141_));
  NO2        m1092(.A(mai_mai_n168_), .B(mai_mai_n53_), .Y(mai_mai_n1142_));
  AOI210     m1093(.A0(mai_mai_n342_), .A1(x8), .B0(mai_mai_n1142_), .Y(mai_mai_n1143_));
  AOI210     m1094(.A0(mai_mai_n218_), .A1(mai_mai_n96_), .B0(mai_mai_n1143_), .Y(mai_mai_n1144_));
  OAI210     m1095(.A0(mai_mai_n1144_), .A1(mai_mai_n1141_), .B0(mai_mai_n676_), .Y(mai_mai_n1145_));
  NO2        m1096(.A(x7), .B(x0), .Y(mai_mai_n1146_));
  NO3        m1097(.A(mai_mai_n159_), .B(mai_mai_n1146_), .C(mai_mai_n146_), .Y(mai_mai_n1147_));
  XN2        m1098(.A(x8), .B(x7), .Y(mai_mai_n1148_));
  NO3        m1099(.A(mai_mai_n1078_), .B(mai_mai_n260_), .C(mai_mai_n1148_), .Y(mai_mai_n1149_));
  OAI210     m1100(.A0(mai_mai_n1149_), .A1(mai_mai_n1147_), .B0(mai_mai_n734_), .Y(mai_mai_n1150_));
  NO2        m1101(.A(mai_mai_n269_), .B(mai_mai_n265_), .Y(mai_mai_n1151_));
  NO2        m1102(.A(mai_mai_n108_), .B(x4), .Y(mai_mai_n1152_));
  OAI210     m1103(.A0(mai_mai_n1151_), .A1(mai_mai_n278_), .B0(mai_mai_n1152_), .Y(mai_mai_n1153_));
  NA3        m1104(.A(mai_mai_n1153_), .B(mai_mai_n1150_), .C(mai_mai_n1145_), .Y(mai_mai_n1154_));
  NA2        m1105(.A(mai_mai_n1154_), .B(mai_mai_n557_), .Y(mai_mai_n1155_));
  NO2        m1106(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n1156_));
  NA2        m1107(.A(mai_mai_n1156_), .B(mai_mai_n164_), .Y(mai_mai_n1157_));
  NO2        m1108(.A(mai_mai_n669_), .B(mai_mai_n260_), .Y(mai_mai_n1158_));
  OAI210     m1109(.A0(mai_mai_n1158_), .A1(mai_mai_n1025_), .B0(mai_mai_n50_), .Y(mai_mai_n1159_));
  AOI210     m1110(.A0(mai_mai_n1159_), .A1(mai_mai_n1157_), .B0(mai_mai_n433_), .Y(mai_mai_n1160_));
  NO2        m1111(.A(mai_mai_n290_), .B(mai_mai_n276_), .Y(mai_mai_n1161_));
  NA3        m1112(.A(mai_mai_n1161_), .B(mai_mai_n676_), .C(x1), .Y(mai_mai_n1162_));
  OAI210     m1113(.A0(x8), .A1(x0), .B0(x4), .Y(mai_mai_n1163_));
  NO2        m1114(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n1164_));
  NO2        m1115(.A(mai_mai_n68_), .B(mai_mai_n1164_), .Y(mai_mai_n1165_));
  NOi21      m1116(.An(mai_mai_n1163_), .B(mai_mai_n1165_), .Y(mai_mai_n1166_));
  NO2        m1117(.A(mai_mai_n667_), .B(mai_mai_n325_), .Y(mai_mai_n1167_));
  NO2        m1118(.A(mai_mai_n780_), .B(mai_mai_n222_), .Y(mai_mai_n1168_));
  OAI210     m1119(.A0(mai_mai_n1167_), .A1(mai_mai_n1166_), .B0(mai_mai_n1168_), .Y(mai_mai_n1169_));
  NO2        m1120(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n1170_));
  NO2        m1121(.A(mai_mai_n606_), .B(mai_mai_n447_), .Y(mai_mai_n1171_));
  OAI210     m1122(.A0(mai_mai_n1171_), .A1(mai_mai_n1170_), .B0(mai_mai_n257_), .Y(mai_mai_n1172_));
  NO2        m1123(.A(mai_mai_n822_), .B(mai_mai_n424_), .Y(mai_mai_n1173_));
  NA2        m1124(.A(mai_mai_n330_), .B(mai_mai_n59_), .Y(mai_mai_n1174_));
  NO2        m1125(.A(mai_mai_n1117_), .B(mai_mai_n1174_), .Y(mai_mai_n1175_));
  AOI210     m1126(.A0(mai_mai_n1173_), .A1(mai_mai_n180_), .B0(mai_mai_n1175_), .Y(mai_mai_n1176_));
  NA4        m1127(.A(mai_mai_n1176_), .B(mai_mai_n1172_), .C(mai_mai_n1169_), .D(mai_mai_n1162_), .Y(mai_mai_n1177_));
  OAI210     m1128(.A0(mai_mai_n1177_), .A1(mai_mai_n1160_), .B0(mai_mai_n678_), .Y(mai_mai_n1178_));
  NA4        m1129(.A(mai_mai_n1178_), .B(mai_mai_n1155_), .C(mai_mai_n1139_), .D(mai_mai_n1119_), .Y(mai13));
  NO2        m1130(.A(mai_mai_n464_), .B(mai_mai_n352_), .Y(mai_mai_n1180_));
  NOi41      m1131(.An(mai_mai_n1180_), .B(mai_mai_n676_), .C(mai_mai_n292_), .D(mai_mai_n241_), .Y(mai_mai_n1181_));
  NO2        m1132(.A(mai_mai_n867_), .B(mai_mai_n184_), .Y(mai_mai_n1182_));
  NO2        m1133(.A(mai_mai_n158_), .B(mai_mai_n71_), .Y(mai_mai_n1183_));
  XN2        m1134(.A(x4), .B(x0), .Y(mai_mai_n1184_));
  NO3        m1135(.A(mai_mai_n1184_), .B(mai_mai_n111_), .C(mai_mai_n424_), .Y(mai_mai_n1185_));
  AO220      m1136(.A0(mai_mai_n1185_), .A1(mai_mai_n1183_), .B0(mai_mai_n1182_), .B1(mai_mai_n331_), .Y(mai_mai_n1186_));
  OAI210     m1137(.A0(mai_mai_n1186_), .A1(mai_mai_n1181_), .B0(x3), .Y(mai_mai_n1187_));
  NO2        m1138(.A(mai_mai_n867_), .B(x6), .Y(mai_mai_n1188_));
  NO2        m1139(.A(mai_mai_n1124_), .B(mai_mai_n396_), .Y(mai_mai_n1189_));
  NO3        m1140(.A(x8), .B(x5), .C(mai_mai_n110_), .Y(mai_mai_n1190_));
  NA2        m1141(.A(mai_mai_n1190_), .B(mai_mai_n642_), .Y(mai_mai_n1191_));
  NO2        m1142(.A(mai_mai_n606_), .B(mai_mai_n200_), .Y(mai_mai_n1192_));
  NA2        m1143(.A(mai_mai_n1192_), .B(mai_mai_n1087_), .Y(mai_mai_n1193_));
  NA2        m1144(.A(mai_mai_n451_), .B(mai_mai_n53_), .Y(mai_mai_n1194_));
  NO2        m1145(.A(mai_mai_n1194_), .B(mai_mai_n939_), .Y(mai_mai_n1195_));
  NA2        m1146(.A(mai_mai_n1117_), .B(mai_mai_n469_), .Y(mai_mai_n1196_));
  NA2        m1147(.A(mai_mai_n56_), .B(mai_mai_n110_), .Y(mai_mai_n1197_));
  NA2        m1148(.A(mai_mai_n1197_), .B(x1), .Y(mai_mai_n1198_));
  NO2        m1149(.A(mai_mai_n1198_), .B(mai_mai_n262_), .Y(mai_mai_n1199_));
  NO2        m1150(.A(mai_mai_n322_), .B(x6), .Y(mai_mai_n1200_));
  NA2        m1151(.A(mai_mai_n1199_), .B(mai_mai_n1196_), .Y(mai_mai_n1201_));
  NAi41      m1152(.An(mai_mai_n1195_), .B(mai_mai_n1201_), .C(mai_mai_n1193_), .D(mai_mai_n1191_), .Y(mai_mai_n1202_));
  AOI220     m1153(.A0(mai_mai_n1202_), .A1(mai_mai_n68_), .B0(mai_mai_n1189_), .B1(mai_mai_n1188_), .Y(mai_mai_n1203_));
  NA2        m1154(.A(mai_mai_n71_), .B(x3), .Y(mai_mai_n1204_));
  NA2        m1155(.A(mai_mai_n1204_), .B(mai_mai_n903_), .Y(mai_mai_n1205_));
  OAI220     m1156(.A0(mai_mai_n304_), .A1(mai_mai_n822_), .B0(mai_mai_n87_), .B1(mai_mai_n77_), .Y(mai_mai_n1206_));
  AOI210     m1157(.A0(mai_mai_n1120_), .A1(mai_mai_n617_), .B0(mai_mai_n980_), .Y(mai_mai_n1207_));
  OA210      m1158(.A0(mai_mai_n1206_), .A1(mai_mai_n1205_), .B0(mai_mai_n1207_), .Y(mai_mai_n1208_));
  NA2        m1159(.A(mai_mai_n619_), .B(mai_mai_n55_), .Y(mai_mai_n1209_));
  NA2        m1160(.A(mai_mai_n506_), .B(mai_mai_n495_), .Y(mai_mai_n1210_));
  NA2        m1161(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n1211_));
  NA2        m1162(.A(mai_mai_n1211_), .B(mai_mai_n540_), .Y(mai_mai_n1212_));
  NO2        m1163(.A(mai_mai_n161_), .B(mai_mai_n132_), .Y(mai_mai_n1213_));
  AOI210     m1164(.A0(mai_mai_n1212_), .A1(mai_mai_n434_), .B0(mai_mai_n1213_), .Y(mai_mai_n1214_));
  OAI220     m1165(.A0(mai_mai_n1214_), .A1(mai_mai_n874_), .B0(mai_mai_n1210_), .B1(mai_mai_n1209_), .Y(mai_mai_n1215_));
  OAI210     m1166(.A0(mai_mai_n1215_), .A1(mai_mai_n1208_), .B0(mai_mai_n1146_), .Y(mai_mai_n1216_));
  NAi21      m1167(.An(mai_mai_n84_), .B(mai_mai_n384_), .Y(mai_mai_n1217_));
  NO2        m1168(.A(mai_mai_n1217_), .B(mai_mai_n71_), .Y(mai_mai_n1218_));
  AOI210     m1169(.A0(mai_mai_n164_), .A1(x4), .B0(mai_mai_n176_), .Y(mai_mai_n1219_));
  NO2        m1170(.A(mai_mai_n1219_), .B(x0), .Y(mai_mai_n1220_));
  NO2        m1171(.A(mai_mai_n172_), .B(mai_mai_n295_), .Y(mai_mai_n1221_));
  OAI210     m1172(.A0(mai_mai_n1221_), .A1(mai_mai_n1220_), .B0(mai_mai_n1218_), .Y(mai_mai_n1222_));
  NA3        m1173(.A(mai_mai_n1152_), .B(mai_mai_n191_), .C(mai_mai_n71_), .Y(mai_mai_n1223_));
  NO2        m1174(.A(x4), .B(x0), .Y(mai_mai_n1224_));
  NO3        m1175(.A(mai_mai_n1000_), .B(mai_mai_n250_), .C(mai_mai_n540_), .Y(mai_mai_n1225_));
  OAI210     m1176(.A0(mai_mai_n1225_), .A1(mai_mai_n201_), .B0(mai_mai_n1224_), .Y(mai_mai_n1226_));
  NA3        m1177(.A(mai_mai_n1226_), .B(mai_mai_n1223_), .C(mai_mai_n1222_), .Y(mai_mai_n1227_));
  NA2        m1178(.A(mai_mai_n252_), .B(mai_mai_n734_), .Y(mai_mai_n1228_));
  NO2        m1179(.A(mai_mai_n1228_), .B(mai_mai_n520_), .Y(mai_mai_n1229_));
  NA2        m1180(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n1230_));
  NO3        m1181(.A(mai_mai_n1230_), .B(mai_mai_n495_), .C(mai_mai_n81_), .Y(mai_mai_n1231_));
  OAI210     m1182(.A0(mai_mai_n1231_), .A1(mai_mai_n1229_), .B0(x2), .Y(mai_mai_n1232_));
  NO2        m1183(.A(mai_mai_n325_), .B(mai_mai_n384_), .Y(mai_mai_n1233_));
  NO2        m1184(.A(mai_mai_n688_), .B(x0), .Y(mai_mai_n1234_));
  OAI210     m1185(.A0(mai_mai_n1234_), .A1(mai_mai_n1233_), .B0(mai_mai_n334_), .Y(mai_mai_n1235_));
  NO2        m1186(.A(mai_mai_n792_), .B(x1), .Y(mai_mai_n1236_));
  AOI220     m1187(.A0(mai_mai_n1236_), .A1(mai_mai_n612_), .B0(mai_mai_n479_), .B1(mai_mai_n296_), .Y(mai_mai_n1237_));
  NA2        m1188(.A(mai_mai_n500_), .B(mai_mai_n50_), .Y(mai_mai_n1238_));
  AOI220     m1189(.A0(mai_mai_n1238_), .A1(mai_mai_n1182_), .B0(mai_mai_n981_), .B1(mai_mai_n101_), .Y(mai_mai_n1239_));
  NA4        m1190(.A(mai_mai_n1239_), .B(mai_mai_n1237_), .C(mai_mai_n1235_), .D(mai_mai_n1232_), .Y(mai_mai_n1240_));
  AOI220     m1191(.A0(mai_mai_n1240_), .A1(mai_mai_n133_), .B0(mai_mai_n1227_), .B1(mai_mai_n67_), .Y(mai_mai_n1241_));
  NA4        m1192(.A(mai_mai_n1241_), .B(mai_mai_n1216_), .C(mai_mai_n1203_), .D(mai_mai_n1187_), .Y(mai14));
  NO2        m1193(.A(mai_mai_n373_), .B(mai_mai_n71_), .Y(mai_mai_n1243_));
  NO3        m1194(.A(x7), .B(x6), .C(x0), .Y(mai_mai_n1244_));
  OAI210     m1195(.A0(mai_mai_n1244_), .A1(mai_mai_n1243_), .B0(x8), .Y(mai_mai_n1245_));
  NA2        m1196(.A(mai_mai_n1133_), .B(mai_mai_n85_), .Y(mai_mai_n1246_));
  AOI210     m1197(.A0(mai_mai_n1246_), .A1(mai_mai_n1245_), .B0(mai_mai_n157_), .Y(mai_mai_n1247_));
  AOI220     m1198(.A0(mai_mai_n377_), .A1(mai_mai_n852_), .B0(mai_mai_n451_), .B1(mai_mai_n424_), .Y(mai_mai_n1248_));
  NA2        m1199(.A(mai_mai_n279_), .B(mai_mai_n976_), .Y(mai_mai_n1249_));
  OAI220     m1200(.A0(mai_mai_n1249_), .A1(mai_mai_n1248_), .B0(mai_mai_n467_), .B1(mai_mai_n806_), .Y(mai_mai_n1250_));
  OA210      m1201(.A0(mai_mai_n1250_), .A1(mai_mai_n1247_), .B0(x4), .Y(mai_mai_n1251_));
  NO2        m1202(.A(mai_mai_n143_), .B(mai_mai_n610_), .Y(mai_mai_n1252_));
  NA2        m1203(.A(x6), .B(x2), .Y(mai_mai_n1253_));
  NO4        m1204(.A(mai_mai_n606_), .B(mai_mai_n378_), .C(mai_mai_n300_), .D(mai_mai_n116_), .Y(mai_mai_n1254_));
  NA2        m1205(.A(mai_mai_n1254_), .B(mai_mai_n59_), .Y(mai_mai_n1255_));
  NA2        m1206(.A(x6), .B(mai_mai_n108_), .Y(mai_mai_n1256_));
  NO2        m1207(.A(mai_mai_n665_), .B(mai_mai_n1256_), .Y(mai_mai_n1257_));
  NA2        m1208(.A(mai_mai_n1257_), .B(mai_mai_n928_), .Y(mai_mai_n1258_));
  AOI210     m1209(.A0(mai_mai_n1133_), .A1(mai_mai_n1014_), .B0(x1), .Y(mai_mai_n1259_));
  NO2        m1210(.A(mai_mai_n535_), .B(x5), .Y(mai_mai_n1260_));
  NA3        m1211(.A(mai_mai_n1260_), .B(mai_mai_n123_), .C(x0), .Y(mai_mai_n1261_));
  NA4        m1212(.A(mai_mai_n695_), .B(mai_mai_n929_), .C(mai_mai_n304_), .D(mai_mai_n68_), .Y(mai_mai_n1262_));
  AN4        m1213(.A(mai_mai_n1262_), .B(mai_mai_n1261_), .C(mai_mai_n1259_), .D(mai_mai_n1258_), .Y(mai_mai_n1263_));
  NO2        m1214(.A(mai_mai_n702_), .B(mai_mai_n1096_), .Y(mai_mai_n1264_));
  NO2        m1215(.A(mai_mai_n77_), .B(mai_mai_n58_), .Y(mai_mai_n1265_));
  OAI210     m1216(.A0(mai_mai_n1264_), .A1(mai_mai_n448_), .B0(mai_mai_n1265_), .Y(mai_mai_n1266_));
  AO210      m1217(.A0(mai_mai_n1243_), .A1(mai_mai_n1014_), .B0(mai_mai_n53_), .Y(mai_mai_n1267_));
  AOI210     m1218(.A0(mai_mai_n767_), .A1(mai_mai_n816_), .B0(mai_mai_n1267_), .Y(mai_mai_n1268_));
  AOI220     m1219(.A0(mai_mai_n1268_), .A1(mai_mai_n1266_), .B0(mai_mai_n1263_), .B1(mai_mai_n1255_), .Y(mai_mai_n1269_));
  NO2        m1220(.A(mai_mai_n677_), .B(mai_mai_n168_), .Y(mai_mai_n1270_));
  NO3        m1221(.A(mai_mai_n1270_), .B(mai_mai_n1269_), .C(mai_mai_n1251_), .Y(mai_mai_n1271_));
  NO2        m1222(.A(mai_mai_n322_), .B(x2), .Y(mai_mai_n1272_));
  XN2        m1223(.A(x4), .B(x1), .Y(mai_mai_n1273_));
  NO2        m1224(.A(mai_mai_n1273_), .B(mai_mai_n304_), .Y(mai_mai_n1274_));
  NOi21      m1225(.An(mai_mai_n1274_), .B(mai_mai_n412_), .Y(mai_mai_n1275_));
  NO2        m1226(.A(mai_mai_n341_), .B(mai_mai_n60_), .Y(mai_mai_n1276_));
  OAI210     m1227(.A0(mai_mai_n1276_), .A1(mai_mai_n1275_), .B0(mai_mai_n1272_), .Y(mai_mai_n1277_));
  NA2        m1228(.A(mai_mai_n689_), .B(mai_mai_n56_), .Y(mai_mai_n1278_));
  OAI220     m1229(.A0(mai_mai_n1278_), .A1(mai_mai_n158_), .B0(mai_mai_n192_), .B1(mai_mai_n71_), .Y(mai_mai_n1279_));
  NO2        m1230(.A(mai_mai_n218_), .B(mai_mai_n260_), .Y(mai_mai_n1280_));
  NA2        m1231(.A(mai_mai_n252_), .B(mai_mai_n356_), .Y(mai_mai_n1281_));
  NA2        m1232(.A(mai_mai_n641_), .B(mai_mai_n1032_), .Y(mai_mai_n1282_));
  NO2        m1233(.A(mai_mai_n1282_), .B(mai_mai_n1281_), .Y(mai_mai_n1283_));
  AOI210     m1234(.A0(mai_mai_n1280_), .A1(mai_mai_n1279_), .B0(mai_mai_n1283_), .Y(mai_mai_n1284_));
  AOI210     m1235(.A0(mai_mai_n1284_), .A1(mai_mai_n1277_), .B0(x7), .Y(mai_mai_n1285_));
  NO2        m1236(.A(mai_mai_n494_), .B(x6), .Y(mai_mai_n1286_));
  AOI210     m1237(.A0(mai_mai_n818_), .A1(mai_mai_n959_), .B0(mai_mai_n1286_), .Y(mai_mai_n1287_));
  OAI220     m1238(.A0(mai_mai_n1287_), .A1(mai_mai_n55_), .B0(mai_mai_n494_), .B1(mai_mai_n104_), .Y(mai_mai_n1288_));
  NA2        m1239(.A(mai_mai_n1288_), .B(mai_mai_n358_), .Y(mai_mai_n1289_));
  NA3        m1240(.A(mai_mai_n613_), .B(mai_mai_n1064_), .C(mai_mai_n70_), .Y(mai_mai_n1290_));
  NO4        m1241(.A(mai_mai_n1290_), .B(mai_mai_n1230_), .C(mai_mai_n121_), .D(mai_mai_n55_), .Y(mai_mai_n1291_));
  NO3        m1242(.A(mai_mai_n1057_), .B(mai_mai_n824_), .C(mai_mai_n484_), .Y(mai_mai_n1292_));
  NO3        m1243(.A(mai_mai_n755_), .B(mai_mai_n500_), .C(mai_mai_n54_), .Y(mai_mai_n1293_));
  NO4        m1244(.A(mai_mai_n1293_), .B(mai_mai_n1292_), .C(mai_mai_n1291_), .D(mai_mai_n1037_), .Y(mai_mai_n1294_));
  AOI210     m1245(.A0(mai_mai_n1294_), .A1(mai_mai_n1289_), .B0(mai_mai_n306_), .Y(mai_mai_n1295_));
  NA2        m1246(.A(mai_mai_n901_), .B(mai_mai_n53_), .Y(mai_mai_n1296_));
  OAI210     m1247(.A0(mai_mai_n247_), .A1(mai_mai_n118_), .B0(x2), .Y(mai_mai_n1297_));
  NA2        m1248(.A(mai_mai_n369_), .B(mai_mai_n56_), .Y(mai_mai_n1298_));
  OA220      m1249(.A0(mai_mai_n1298_), .A1(mai_mai_n1297_), .B0(mai_mai_n1296_), .B1(mai_mai_n377_), .Y(mai_mai_n1299_));
  NA3        m1250(.A(mai_mai_n1037_), .B(mai_mai_n739_), .C(mai_mai_n55_), .Y(mai_mai_n1300_));
  NA2        m1251(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n1301_));
  NO2        m1252(.A(mai_mai_n1301_), .B(mai_mai_n199_), .Y(mai_mai_n1302_));
  NA4        m1253(.A(mai_mai_n1302_), .B(mai_mai_n369_), .C(mai_mai_n260_), .D(mai_mai_n67_), .Y(mai_mai_n1303_));
  NA3        m1254(.A(mai_mai_n1236_), .B(mai_mai_n619_), .C(mai_mai_n633_), .Y(mai_mai_n1304_));
  AN3        m1255(.A(mai_mai_n1304_), .B(mai_mai_n1303_), .C(mai_mai_n1300_), .Y(mai_mai_n1305_));
  OAI210     m1256(.A0(mai_mai_n1299_), .A1(mai_mai_n317_), .B0(mai_mai_n1305_), .Y(mai_mai_n1306_));
  NO3        m1257(.A(mai_mai_n1306_), .B(mai_mai_n1295_), .C(mai_mai_n1285_), .Y(mai_mai_n1307_));
  OAI210     m1258(.A0(mai_mai_n1271_), .A1(x3), .B0(mai_mai_n1307_), .Y(mai15));
  NA2        m1259(.A(mai_mai_n588_), .B(mai_mai_n59_), .Y(mai_mai_n1309_));
  NAi41      m1260(.An(x2), .B(x7), .C(x6), .D(x0), .Y(mai_mai_n1310_));
  AOI210     m1261(.A0(mai_mai_n1310_), .A1(mai_mai_n1309_), .B0(mai_mai_n53_), .Y(mai_mai_n1311_));
  NA3        m1262(.A(mai_mai_n57_), .B(x6), .C(mai_mai_n110_), .Y(mai_mai_n1312_));
  NO2        m1263(.A(mai_mai_n1312_), .B(mai_mai_n295_), .Y(mai_mai_n1313_));
  OAI210     m1264(.A0(mai_mai_n1313_), .A1(mai_mai_n1311_), .B0(mai_mai_n1152_), .Y(mai_mai_n1314_));
  NA2        m1265(.A(mai_mai_n112_), .B(mai_mai_n110_), .Y(mai_mai_n1315_));
  NA4        m1266(.A(mai_mai_n1315_), .B(mai_mai_n640_), .C(mai_mai_n310_), .D(x6), .Y(mai_mai_n1316_));
  AOI210     m1267(.A0(mai_mai_n733_), .A1(mai_mai_n76_), .B0(x3), .Y(mai_mai_n1317_));
  NA3        m1268(.A(mai_mai_n1317_), .B(mai_mai_n1316_), .C(mai_mai_n1314_), .Y(mai_mai_n1318_));
  AOI210     m1269(.A0(mai_mai_n1069_), .A1(mai_mai_n592_), .B0(mai_mai_n50_), .Y(mai_mai_n1319_));
  NO2        m1270(.A(mai_mai_n295_), .B(mai_mai_n110_), .Y(mai_mai_n1320_));
  NO2        m1271(.A(mai_mai_n239_), .B(x5), .Y(mai_mai_n1321_));
  NA2        m1272(.A(mai_mai_n1321_), .B(mai_mai_n1320_), .Y(mai_mai_n1322_));
  NA3        m1273(.A(mai_mai_n1236_), .B(mai_mai_n627_), .C(mai_mai_n1164_), .Y(mai_mai_n1323_));
  NA4        m1274(.A(mai_mai_n1323_), .B(mai_mai_n1322_), .C(mai_mai_n1319_), .D(mai_mai_n1261_), .Y(mai_mai_n1324_));
  NA2        m1275(.A(mai_mai_n335_), .B(mai_mai_n344_), .Y(mai_mai_n1325_));
  AOI210     m1276(.A0(mai_mai_n1198_), .A1(mai_mai_n58_), .B0(mai_mai_n1325_), .Y(mai_mai_n1326_));
  NA4        m1277(.A(mai_mai_n1198_), .B(mai_mai_n701_), .C(mai_mai_n1130_), .D(mai_mai_n384_), .Y(mai_mai_n1327_));
  NA2        m1278(.A(mai_mai_n592_), .B(mai_mai_n468_), .Y(mai_mai_n1328_));
  NO2        m1279(.A(mai_mai_n755_), .B(mai_mai_n53_), .Y(mai_mai_n1329_));
  NO2        m1280(.A(mai_mai_n780_), .B(mai_mai_n300_), .Y(mai_mai_n1330_));
  NA2        m1281(.A(mai_mai_n1330_), .B(mai_mai_n1329_), .Y(mai_mai_n1331_));
  NA3        m1282(.A(mai_mai_n1331_), .B(mai_mai_n1328_), .C(mai_mai_n1327_), .Y(mai_mai_n1332_));
  OAI210     m1283(.A0(mai_mai_n1332_), .A1(mai_mai_n1326_), .B0(mai_mai_n77_), .Y(mai_mai_n1333_));
  NA2        m1284(.A(mai_mai_n371_), .B(mai_mai_n704_), .Y(mai_mai_n1334_));
  NA2        m1285(.A(mai_mai_n573_), .B(mai_mai_n56_), .Y(mai_mai_n1335_));
  NA3        m1286(.A(mai_mai_n1335_), .B(mai_mai_n344_), .C(mai_mai_n112_), .Y(mai_mai_n1336_));
  AOI210     m1287(.A0(mai_mai_n1336_), .A1(mai_mai_n1334_), .B0(mai_mai_n500_), .Y(mai_mai_n1337_));
  NO3        m1288(.A(mai_mai_n804_), .B(mai_mai_n624_), .C(mai_mai_n200_), .Y(mai_mai_n1338_));
  OAI210     m1289(.A0(mai_mai_n1338_), .A1(mai_mai_n1337_), .B0(mai_mai_n494_), .Y(mai_mai_n1339_));
  NO2        m1290(.A(mai_mai_n874_), .B(mai_mai_n50_), .Y(mai_mai_n1340_));
  NO2        m1291(.A(mai_mai_n249_), .B(mai_mai_n64_), .Y(mai_mai_n1341_));
  OA210      m1292(.A0(mai_mai_n1341_), .A1(mai_mai_n1340_), .B0(mai_mai_n412_), .Y(mai_mai_n1342_));
  NA2        m1293(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n1343_));
  AOI210     m1294(.A0(mai_mai_n982_), .A1(mai_mai_n1343_), .B0(mai_mai_n683_), .Y(mai_mai_n1344_));
  OAI210     m1295(.A0(mai_mai_n1344_), .A1(mai_mai_n1342_), .B0(mai_mai_n1022_), .Y(mai_mai_n1345_));
  NA2        m1296(.A(mai_mai_n1302_), .B(mai_mai_n68_), .Y(mai_mai_n1346_));
  NO2        m1297(.A(mai_mai_n1253_), .B(x0), .Y(mai_mai_n1347_));
  AOI210     m1298(.A0(mai_mai_n1347_), .A1(mai_mai_n607_), .B0(x8), .Y(mai_mai_n1348_));
  NO2        m1299(.A(mai_mai_n433_), .B(mai_mai_n81_), .Y(mai_mai_n1349_));
  NO2        m1300(.A(mai_mai_n933_), .B(mai_mai_n71_), .Y(mai_mai_n1350_));
  NA2        m1301(.A(mai_mai_n1350_), .B(mai_mai_n1349_), .Y(mai_mai_n1351_));
  NO2        m1302(.A(mai_mai_n980_), .B(x6), .Y(mai_mai_n1352_));
  NA3        m1303(.A(mai_mai_n1352_), .B(mai_mai_n597_), .C(mai_mai_n416_), .Y(mai_mai_n1353_));
  AN4        m1304(.A(mai_mai_n1353_), .B(mai_mai_n1351_), .C(mai_mai_n1348_), .D(mai_mai_n1346_), .Y(mai_mai_n1354_));
  NA4        m1305(.A(mai_mai_n1354_), .B(mai_mai_n1345_), .C(mai_mai_n1339_), .D(mai_mai_n1333_), .Y(mai_mai_n1355_));
  NA2        m1306(.A(mai_mai_n165_), .B(mai_mai_n739_), .Y(mai_mai_n1356_));
  NO2        m1307(.A(mai_mai_n650_), .B(x2), .Y(mai_mai_n1357_));
  OAI210     m1308(.A0(mai_mai_n68_), .A1(mai_mai_n53_), .B0(mai_mai_n145_), .Y(mai_mai_n1358_));
  OAI210     m1309(.A0(mai_mai_n1357_), .A1(mai_mai_n85_), .B0(mai_mai_n1358_), .Y(mai_mai_n1359_));
  AOI210     m1310(.A0(mai_mai_n1359_), .A1(mai_mai_n1356_), .B0(mai_mai_n322_), .Y(mai_mai_n1360_));
  NO3        m1311(.A(mai_mai_n1312_), .B(mai_mai_n268_), .C(mai_mai_n249_), .Y(mai_mai_n1361_));
  NA3        m1312(.A(mai_mai_n57_), .B(x1), .C(x0), .Y(mai_mai_n1362_));
  NA3        m1313(.A(mai_mai_n71_), .B(x5), .C(x2), .Y(mai_mai_n1363_));
  NA4        m1314(.A(x7), .B(x3), .C(mai_mai_n53_), .D(x0), .Y(mai_mai_n1364_));
  OAI220     m1315(.A0(mai_mai_n1364_), .A1(x6), .B0(mai_mai_n1363_), .B1(mai_mai_n1362_), .Y(mai_mai_n1365_));
  NO2        m1316(.A(mai_mai_n1365_), .B(mai_mai_n1361_), .Y(mai_mai_n1366_));
  NAi21      m1317(.An(mai_mai_n116_), .B(mai_mai_n749_), .Y(mai_mai_n1367_));
  NA4        m1318(.A(mai_mai_n1367_), .B(mai_mai_n320_), .C(mai_mai_n290_), .D(mai_mai_n627_), .Y(mai_mai_n1368_));
  OAI220     m1319(.A0(mai_mai_n325_), .A1(x7), .B0(mai_mai_n132_), .B1(mai_mai_n71_), .Y(mai_mai_n1369_));
  NA3        m1320(.A(mai_mai_n1369_), .B(mai_mai_n792_), .C(mai_mai_n1099_), .Y(mai_mai_n1370_));
  NA2        m1321(.A(mai_mai_n82_), .B(mai_mai_n50_), .Y(mai_mai_n1371_));
  AO210      m1322(.A0(mai_mai_n1371_), .A1(mai_mai_n315_), .B0(mai_mai_n157_), .Y(mai_mai_n1372_));
  NA4        m1323(.A(mai_mai_n1372_), .B(mai_mai_n1370_), .C(mai_mai_n1368_), .D(mai_mai_n1366_), .Y(mai_mai_n1373_));
  OAI210     m1324(.A0(mai_mai_n1373_), .A1(mai_mai_n1360_), .B0(mai_mai_n56_), .Y(mai_mai_n1374_));
  AOI210     m1325(.A0(mai_mai_n691_), .A1(x4), .B0(mai_mai_n959_), .Y(mai_mai_n1375_));
  OAI220     m1326(.A0(mai_mai_n1375_), .A1(mai_mai_n301_), .B0(mai_mai_n1026_), .B1(mai_mai_n947_), .Y(mai_mai_n1376_));
  NA2        m1327(.A(mai_mai_n835_), .B(mai_mai_n409_), .Y(mai_mai_n1377_));
  OAI210     m1328(.A0(mai_mai_n1349_), .A1(mai_mai_n1341_), .B0(mai_mai_n291_), .Y(mai_mai_n1378_));
  OAI210     m1329(.A0(mai_mai_n1377_), .A1(mai_mai_n847_), .B0(mai_mai_n1378_), .Y(mai_mai_n1379_));
  OAI210     m1330(.A0(mai_mai_n1379_), .A1(mai_mai_n1376_), .B0(x6), .Y(mai_mai_n1380_));
  NO2        m1331(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n1381_));
  NO2        m1332(.A(x7), .B(x5), .Y(mai_mai_n1382_));
  AOI220     m1333(.A0(mai_mai_n856_), .A1(mai_mai_n1381_), .B0(mai_mai_n539_), .B1(mai_mai_n1382_), .Y(mai_mai_n1383_));
  NA2        m1334(.A(mai_mai_n764_), .B(mai_mai_n291_), .Y(mai_mai_n1384_));
  NA3        m1335(.A(mai_mai_n619_), .B(mai_mai_n293_), .C(mai_mai_n244_), .Y(mai_mai_n1385_));
  NA3        m1336(.A(mai_mai_n1385_), .B(mai_mai_n1384_), .C(mai_mai_n1383_), .Y(mai_mai_n1386_));
  NA2        m1337(.A(mai_mai_n1386_), .B(mai_mai_n427_), .Y(mai_mai_n1387_));
  AOI210     m1338(.A0(mai_mai_n381_), .A1(mai_mai_n342_), .B0(mai_mai_n55_), .Y(mai_mai_n1388_));
  NA4        m1339(.A(mai_mai_n1388_), .B(mai_mai_n1387_), .C(mai_mai_n1380_), .D(mai_mai_n1374_), .Y(mai_mai_n1389_));
  AO220      m1340(.A0(mai_mai_n1389_), .A1(mai_mai_n1355_), .B0(mai_mai_n1324_), .B1(mai_mai_n1318_), .Y(mai16));
  NO2        m1341(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n1391_));
  NA2        m1342(.A(mai_mai_n664_), .B(mai_mai_n536_), .Y(mai_mai_n1392_));
  NA3        m1343(.A(mai_mai_n233_), .B(mai_mai_n434_), .C(mai_mai_n959_), .Y(mai_mai_n1393_));
  NA2        m1344(.A(mai_mai_n135_), .B(mai_mai_n209_), .Y(mai_mai_n1394_));
  AOI210     m1345(.A0(mai_mai_n1393_), .A1(mai_mai_n1392_), .B0(mai_mai_n1394_), .Y(mai_mai_n1395_));
  NO3        m1346(.A(x8), .B(x6), .C(mai_mai_n50_), .Y(mai_mai_n1396_));
  NO2        m1347(.A(mai_mai_n737_), .B(mai_mai_n187_), .Y(mai_mai_n1397_));
  OAI210     m1348(.A0(mai_mai_n1396_), .A1(mai_mai_n241_), .B0(mai_mai_n1397_), .Y(mai_mai_n1398_));
  NO2        m1349(.A(mai_mai_n161_), .B(x5), .Y(mai_mai_n1399_));
  NA2        m1350(.A(mai_mai_n1399_), .B(mai_mai_n1357_), .Y(mai_mai_n1400_));
  NA3        m1351(.A(mai_mai_n582_), .B(mai_mai_n538_), .C(mai_mai_n478_), .Y(mai_mai_n1401_));
  NA3        m1352(.A(mai_mai_n1401_), .B(mai_mai_n1400_), .C(mai_mai_n1398_), .Y(mai_mai_n1402_));
  OAI210     m1353(.A0(mai_mai_n1402_), .A1(mai_mai_n1395_), .B0(mai_mai_n1391_), .Y(mai_mai_n1403_));
  NO2        m1354(.A(mai_mai_n322_), .B(x7), .Y(mai_mai_n1404_));
  NA2        m1355(.A(mai_mai_n1078_), .B(mai_mai_n200_), .Y(mai_mai_n1405_));
  NA2        m1356(.A(mai_mai_n55_), .B(mai_mai_n108_), .Y(mai_mai_n1406_));
  NA2        m1357(.A(mai_mai_n1406_), .B(mai_mai_n685_), .Y(mai_mai_n1407_));
  NA2        m1358(.A(mai_mai_n380_), .B(mai_mai_n1082_), .Y(mai_mai_n1408_));
  OA220      m1359(.A0(mai_mai_n1408_), .A1(mai_mai_n1407_), .B0(mai_mai_n1405_), .B1(mai_mai_n635_), .Y(mai_mai_n1409_));
  NO2        m1360(.A(mai_mai_n1409_), .B(mai_mai_n654_), .Y(mai_mai_n1410_));
  INV        m1361(.A(mai_mai_n1022_), .Y(mai_mai_n1411_));
  NO2        m1362(.A(mai_mai_n1411_), .B(mai_mai_n62_), .Y(mai_mai_n1412_));
  AOI220     m1363(.A0(mai_mai_n1412_), .A1(mai_mai_n272_), .B0(mai_mai_n1257_), .B1(mai_mai_n128_), .Y(mai_mai_n1413_));
  AOI220     m1364(.A0(mai_mai_n640_), .A1(mai_mai_n365_), .B0(mai_mai_n627_), .B1(mai_mai_n88_), .Y(mai_mai_n1414_));
  NA3        m1365(.A(mai_mai_n465_), .B(mai_mai_n589_), .C(mai_mai_n194_), .Y(mai_mai_n1415_));
  OAI220     m1366(.A0(mai_mai_n1415_), .A1(mai_mai_n1414_), .B0(mai_mai_n1413_), .B1(mai_mai_n311_), .Y(mai_mai_n1416_));
  NO2        m1367(.A(mai_mai_n1416_), .B(mai_mai_n1410_), .Y(mai_mai_n1417_));
  NO3        m1368(.A(x6), .B(x4), .C(x3), .Y(mai_mai_n1418_));
  NA2        m1369(.A(mai_mai_n1418_), .B(mai_mai_n535_), .Y(mai_mai_n1419_));
  NA4        m1370(.A(mai_mai_n709_), .B(mai_mai_n187_), .C(mai_mai_n58_), .D(x6), .Y(mai_mai_n1420_));
  AOI210     m1371(.A0(mai_mai_n1420_), .A1(mai_mai_n1419_), .B0(mai_mai_n54_), .Y(mai_mai_n1421_));
  NO2        m1372(.A(mai_mai_n725_), .B(x3), .Y(mai_mai_n1422_));
  AOI210     m1373(.A0(mai_mai_n663_), .A1(mai_mai_n148_), .B0(mai_mai_n1064_), .Y(mai_mai_n1423_));
  OA210      m1374(.A0(mai_mai_n1422_), .A1(mai_mai_n427_), .B0(mai_mai_n1423_), .Y(mai_mai_n1424_));
  NO3        m1375(.A(mai_mai_n500_), .B(mai_mai_n222_), .C(mai_mai_n75_), .Y(mai_mai_n1425_));
  NO2        m1376(.A(mai_mai_n764_), .B(mai_mai_n512_), .Y(mai_mai_n1426_));
  NO3        m1377(.A(mai_mai_n1426_), .B(mai_mai_n262_), .C(mai_mai_n156_), .Y(mai_mai_n1427_));
  NO4        m1378(.A(mai_mai_n1427_), .B(mai_mai_n1425_), .C(mai_mai_n1424_), .D(mai_mai_n1421_), .Y(mai_mai_n1428_));
  NA2        m1379(.A(mai_mai_n410_), .B(mai_mai_n959_), .Y(mai_mai_n1429_));
  NA4        m1380(.A(mai_mai_n484_), .B(mai_mai_n373_), .C(mai_mai_n224_), .D(x6), .Y(mai_mai_n1430_));
  OAI210     m1381(.A0(mai_mai_n725_), .A1(mai_mai_n1429_), .B0(mai_mai_n1430_), .Y(mai_mai_n1431_));
  NA2        m1382(.A(mai_mai_n910_), .B(mai_mai_n1301_), .Y(mai_mai_n1432_));
  NA2        m1383(.A(mai_mai_n734_), .B(x7), .Y(mai_mai_n1433_));
  OAI210     m1384(.A0(mai_mai_n1433_), .A1(mai_mai_n391_), .B0(mai_mai_n1432_), .Y(mai_mai_n1434_));
  NA2        m1385(.A(mai_mai_n277_), .B(x2), .Y(mai_mai_n1435_));
  NO3        m1386(.A(mai_mai_n1435_), .B(mai_mai_n597_), .C(mai_mai_n72_), .Y(mai_mai_n1436_));
  OA210      m1387(.A0(mai_mai_n1256_), .A1(mai_mai_n58_), .B0(mai_mai_n781_), .Y(mai_mai_n1437_));
  AOI210     m1388(.A0(mai_mai_n582_), .A1(mai_mai_n50_), .B0(mai_mai_n592_), .Y(mai_mai_n1438_));
  OAI210     m1389(.A0(mai_mai_n929_), .A1(mai_mai_n946_), .B0(mai_mai_n386_), .Y(mai_mai_n1439_));
  OAI220     m1390(.A0(mai_mai_n1439_), .A1(mai_mai_n1438_), .B0(mai_mai_n1437_), .B1(mai_mai_n192_), .Y(mai_mai_n1440_));
  NO4        m1391(.A(mai_mai_n1440_), .B(mai_mai_n1436_), .C(mai_mai_n1434_), .D(mai_mai_n1431_), .Y(mai_mai_n1441_));
  OA220      m1392(.A0(mai_mai_n1441_), .A1(mai_mai_n447_), .B0(mai_mai_n1428_), .B1(mai_mai_n207_), .Y(mai_mai_n1442_));
  NO2        m1393(.A(mai_mai_n924_), .B(mai_mai_n55_), .Y(mai_mai_n1443_));
  NA2        m1394(.A(mai_mai_n421_), .B(mai_mai_n806_), .Y(mai_mai_n1444_));
  NO2        m1395(.A(mai_mai_n1444_), .B(mai_mai_n1443_), .Y(mai_mai_n1445_));
  NO3        m1396(.A(mai_mai_n960_), .B(mai_mai_n335_), .C(x8), .Y(mai_mai_n1446_));
  OAI210     m1397(.A0(mai_mai_n1446_), .A1(mai_mai_n1445_), .B0(x6), .Y(mai_mai_n1447_));
  NO2        m1398(.A(mai_mai_n1094_), .B(mai_mai_n1056_), .Y(mai_mai_n1448_));
  NA2        m1399(.A(mai_mai_n192_), .B(x7), .Y(mai_mai_n1449_));
  OAI220     m1400(.A0(mai_mai_n1449_), .A1(mai_mai_n1448_), .B0(mai_mai_n766_), .B1(mai_mai_n87_), .Y(mai_mai_n1450_));
  NA2        m1401(.A(mai_mai_n1450_), .B(mai_mai_n929_), .Y(mai_mai_n1451_));
  NA2        m1402(.A(mai_mai_n876_), .B(mai_mai_n71_), .Y(mai_mai_n1452_));
  INV        m1403(.A(mai_mai_n1011_), .Y(mai_mai_n1453_));
  AOI210     m1404(.A0(mai_mai_n500_), .A1(mai_mai_n57_), .B0(mai_mai_n635_), .Y(mai_mai_n1454_));
  NA3        m1405(.A(mai_mai_n230_), .B(mai_mai_n76_), .C(mai_mai_n71_), .Y(mai_mai_n1455_));
  OAI210     m1406(.A0(mai_mai_n920_), .A1(mai_mai_n233_), .B0(mai_mai_n1455_), .Y(mai_mai_n1456_));
  AOI210     m1407(.A0(mai_mai_n1454_), .A1(mai_mai_n1453_), .B0(mai_mai_n1456_), .Y(mai_mai_n1457_));
  NA3        m1408(.A(mai_mai_n1457_), .B(mai_mai_n1451_), .C(mai_mai_n1447_), .Y(mai_mai_n1458_));
  NO2        m1409(.A(mai_mai_n641_), .B(x6), .Y(mai_mai_n1459_));
  OAI210     m1410(.A0(mai_mai_n386_), .A1(mai_mai_n84_), .B0(mai_mai_n384_), .Y(mai_mai_n1460_));
  OA210      m1411(.A0(mai_mai_n1460_), .A1(mai_mai_n1459_), .B0(mai_mai_n133_), .Y(mai_mai_n1461_));
  NO3        m1412(.A(mai_mai_n449_), .B(mai_mai_n389_), .C(x7), .Y(mai_mai_n1462_));
  NO3        m1413(.A(mai_mai_n161_), .B(mai_mai_n75_), .C(x2), .Y(mai_mai_n1463_));
  NO3        m1414(.A(mai_mai_n1463_), .B(mai_mai_n1462_), .C(mai_mai_n1461_), .Y(mai_mai_n1464_));
  NO2        m1415(.A(mai_mai_n233_), .B(x1), .Y(mai_mai_n1465_));
  OAI210     m1416(.A0(mai_mai_n1465_), .A1(mai_mai_n454_), .B0(mai_mai_n512_), .Y(mai_mai_n1466_));
  NO2        m1417(.A(mai_mai_n57_), .B(mai_mai_n108_), .Y(mai_mai_n1467_));
  NA2        m1418(.A(mai_mai_n1087_), .B(mai_mai_n1467_), .Y(mai_mai_n1468_));
  AOI210     m1419(.A0(mai_mai_n1468_), .A1(mai_mai_n1466_), .B0(mai_mai_n56_), .Y(mai_mai_n1469_));
  AOI220     m1420(.A0(mai_mai_n766_), .A1(mai_mai_n777_), .B0(mai_mai_n515_), .B1(mai_mai_n281_), .Y(mai_mai_n1470_));
  NO2        m1421(.A(mai_mai_n1470_), .B(mai_mai_n1301_), .Y(mai_mai_n1471_));
  NO3        m1422(.A(mai_mai_n535_), .B(mai_mai_n174_), .C(mai_mai_n1056_), .Y(mai_mai_n1472_));
  NA2        m1423(.A(mai_mai_n946_), .B(x4), .Y(mai_mai_n1473_));
  OAI220     m1424(.A0(mai_mai_n1473_), .A1(mai_mai_n690_), .B0(mai_mai_n648_), .B1(mai_mai_n613_), .Y(mai_mai_n1474_));
  NO4        m1425(.A(mai_mai_n1474_), .B(mai_mai_n1472_), .C(mai_mai_n1471_), .D(mai_mai_n1469_), .Y(mai_mai_n1475_));
  OAI210     m1426(.A0(mai_mai_n1464_), .A1(x5), .B0(mai_mai_n1475_), .Y(mai_mai_n1476_));
  AOI220     m1427(.A0(mai_mai_n1476_), .A1(mai_mai_n99_), .B0(mai_mai_n1458_), .B1(mai_mai_n342_), .Y(mai_mai_n1477_));
  NA4        m1428(.A(mai_mai_n1477_), .B(mai_mai_n1442_), .C(mai_mai_n1417_), .D(mai_mai_n1403_), .Y(mai17));
  NO4        m1429(.A(mai_mai_n604_), .B(mai_mai_n703_), .C(mai_mai_n102_), .D(mai_mai_n101_), .Y(mai_mai_n1479_));
  NO2        m1430(.A(mai_mai_n126_), .B(mai_mai_n1164_), .Y(mai_mai_n1480_));
  AOI220     m1431(.A0(mai_mai_n1480_), .A1(mai_mai_n719_), .B0(mai_mai_n1479_), .B1(mai_mai_n506_), .Y(mai_mai_n1481_));
  NA2        m1432(.A(mai_mai_n165_), .B(mai_mai_n78_), .Y(mai_mai_n1482_));
  NOi21      m1433(.An(mai_mai_n384_), .B(mai_mai_n84_), .Y(mai_mai_n1483_));
  OAI210     m1434(.A0(mai_mai_n627_), .A1(mai_mai_n55_), .B0(mai_mai_n1483_), .Y(mai_mai_n1484_));
  NA2        m1435(.A(mai_mai_n1217_), .B(mai_mai_n1017_), .Y(mai_mai_n1485_));
  NA4        m1436(.A(mai_mai_n1485_), .B(mai_mai_n1484_), .C(mai_mai_n737_), .D(mai_mai_n57_), .Y(mai_mai_n1486_));
  OAI210     m1437(.A0(mai_mai_n709_), .A1(x8), .B0(mai_mai_n1301_), .Y(mai_mai_n1487_));
  NA3        m1438(.A(mai_mai_n1487_), .B(mai_mai_n1243_), .C(mai_mai_n403_), .Y(mai_mai_n1488_));
  NA3        m1439(.A(mai_mai_n397_), .B(mai_mai_n272_), .C(mai_mai_n588_), .Y(mai_mai_n1489_));
  OA210      m1440(.A0(mai_mai_n1312_), .A1(mai_mai_n1157_), .B0(mai_mai_n757_), .Y(mai_mai_n1490_));
  NA4        m1441(.A(mai_mai_n1490_), .B(mai_mai_n1489_), .C(mai_mai_n1488_), .D(mai_mai_n1486_), .Y(mai_mai_n1491_));
  NA3        m1442(.A(mai_mai_n164_), .B(mai_mai_n633_), .C(mai_mai_n1056_), .Y(mai_mai_n1492_));
  AOI210     m1443(.A0(mai_mai_n1084_), .A1(mai_mai_n307_), .B0(mai_mai_n59_), .Y(mai_mai_n1493_));
  NA2        m1444(.A(mai_mai_n1493_), .B(mai_mai_n1492_), .Y(mai_mai_n1494_));
  AOI210     m1445(.A0(mai_mai_n1491_), .A1(x1), .B0(mai_mai_n1494_), .Y(mai_mai_n1495_));
  NO2        m1446(.A(mai_mai_n985_), .B(mai_mai_n500_), .Y(mai_mai_n1496_));
  OAI210     m1447(.A0(mai_mai_n1496_), .A1(mai_mai_n1068_), .B0(mai_mai_n610_), .Y(mai_mai_n1497_));
  NO3        m1448(.A(mai_mai_n635_), .B(mai_mai_n557_), .C(mai_mai_n526_), .Y(mai_mai_n1498_));
  OAI210     m1449(.A0(mai_mai_n1498_), .A1(mai_mai_n909_), .B0(mai_mai_n1422_), .Y(mai_mai_n1499_));
  AOI210     m1450(.A0(mai_mai_n1499_), .A1(mai_mai_n1497_), .B0(x8), .Y(mai_mai_n1500_));
  NA3        m1451(.A(mai_mai_n635_), .B(mai_mai_n274_), .C(mai_mai_n123_), .Y(mai_mai_n1501_));
  NO2        m1452(.A(mai_mai_n145_), .B(mai_mai_n144_), .Y(mai_mai_n1502_));
  NO3        m1453(.A(mai_mai_n904_), .B(mai_mai_n777_), .C(mai_mai_n703_), .Y(mai_mai_n1503_));
  AOI210     m1454(.A0(mai_mai_n1503_), .A1(mai_mai_n1502_), .B0(x0), .Y(mai_mai_n1504_));
  OAI210     m1455(.A0(mai_mai_n1501_), .A1(mai_mai_n251_), .B0(mai_mai_n1504_), .Y(mai_mai_n1505_));
  NO2        m1456(.A(mai_mai_n1505_), .B(mai_mai_n1500_), .Y(mai_mai_n1506_));
  OAI220     m1457(.A0(mai_mai_n1506_), .A1(mai_mai_n1495_), .B0(mai_mai_n1482_), .B1(mai_mai_n1481_), .Y(mai18));
  AOI210     m1458(.A0(x8), .A1(x0), .B0(x5), .Y(mai_mai_n1508_));
  NOi31      m1459(.An(mai_mai_n307_), .B(mai_mai_n1508_), .C(mai_mai_n1054_), .Y(mai_mai_n1509_));
  NA2        m1460(.A(mai_mai_n604_), .B(mai_mai_n59_), .Y(mai_mai_n1510_));
  AOI210     m1461(.A0(mai_mai_n1405_), .A1(mai_mai_n353_), .B0(mai_mai_n1510_), .Y(mai_mai_n1511_));
  NO2        m1462(.A(mai_mai_n620_), .B(mai_mai_n778_), .Y(mai_mai_n1512_));
  NO4        m1463(.A(mai_mai_n258_), .B(mai_mai_n816_), .C(mai_mai_n155_), .D(mai_mai_n70_), .Y(mai_mai_n1513_));
  NO4        m1464(.A(mai_mai_n1513_), .B(mai_mai_n1512_), .C(mai_mai_n1511_), .D(mai_mai_n1509_), .Y(mai_mai_n1514_));
  NA3        m1465(.A(mai_mai_n521_), .B(mai_mai_n218_), .C(x0), .Y(mai_mai_n1515_));
  NAi21      m1466(.An(mai_mai_n390_), .B(mai_mai_n1515_), .Y(mai_mai_n1516_));
  NO2        m1467(.A(mai_mai_n894_), .B(x5), .Y(mai_mai_n1517_));
  AOI210     m1468(.A0(mai_mai_n1142_), .A1(x5), .B0(mai_mai_n1517_), .Y(mai_mai_n1518_));
  OA220      m1469(.A0(mai_mai_n521_), .A1(mai_mai_n335_), .B0(mai_mai_n403_), .B1(x5), .Y(mai_mai_n1519_));
  OAI220     m1470(.A0(mai_mai_n1519_), .A1(mai_mai_n295_), .B0(mai_mai_n1518_), .B1(mai_mai_n216_), .Y(mai_mai_n1520_));
  AOI210     m1471(.A0(mai_mai_n1516_), .A1(mai_mai_n293_), .B0(mai_mai_n1520_), .Y(mai_mai_n1521_));
  AOI210     m1472(.A0(mai_mai_n1521_), .A1(mai_mai_n1514_), .B0(x6), .Y(mai_mai_n1522_));
  NA3        m1473(.A(mai_mai_n525_), .B(mai_mai_n424_), .C(x2), .Y(mai_mai_n1523_));
  NA3        m1474(.A(mai_mai_n1054_), .B(mai_mai_n51_), .C(mai_mai_n57_), .Y(mai_mai_n1524_));
  AOI210     m1475(.A0(mai_mai_n1524_), .A1(mai_mai_n1523_), .B0(mai_mai_n792_), .Y(mai_mai_n1525_));
  AOI210     m1476(.A0(mai_mai_n428_), .A1(mai_mai_n140_), .B0(mai_mai_n790_), .Y(mai_mai_n1526_));
  NA2        m1477(.A(mai_mai_n272_), .B(x6), .Y(mai_mai_n1527_));
  OAI210     m1478(.A0(mai_mai_n180_), .A1(mai_mai_n110_), .B0(mai_mai_n1148_), .Y(mai_mai_n1528_));
  OAI220     m1479(.A0(mai_mai_n1528_), .A1(mai_mai_n1527_), .B0(mai_mai_n1526_), .B1(mai_mai_n749_), .Y(mai_mai_n1529_));
  OAI210     m1480(.A0(mai_mai_n1529_), .A1(mai_mai_n1525_), .B0(mai_mai_n53_), .Y(mai_mai_n1530_));
  NO2        m1481(.A(mai_mai_n689_), .B(mai_mai_n265_), .Y(mai_mai_n1531_));
  NO2        m1482(.A(mai_mai_n268_), .B(x3), .Y(mai_mai_n1532_));
  NO3        m1483(.A(mai_mai_n438_), .B(mai_mai_n604_), .C(mai_mai_n840_), .Y(mai_mai_n1533_));
  OAI210     m1484(.A0(mai_mai_n1533_), .A1(mai_mai_n1531_), .B0(mai_mai_n1532_), .Y(mai_mai_n1534_));
  AOI210     m1485(.A0(mai_mai_n1151_), .A1(mai_mai_n619_), .B0(x4), .Y(mai_mai_n1535_));
  OAI210     m1486(.A0(mai_mai_n557_), .A1(mai_mai_n604_), .B0(mai_mai_n59_), .Y(mai_mai_n1536_));
  OAI210     m1487(.A0(mai_mai_n627_), .A1(mai_mai_n650_), .B0(mai_mai_n1536_), .Y(mai_mai_n1537_));
  AO220      m1488(.A0(mai_mai_n1260_), .A1(mai_mai_n737_), .B0(mai_mai_n558_), .B1(mai_mai_n358_), .Y(mai_mai_n1538_));
  AOI220     m1489(.A0(mai_mai_n1538_), .A1(x1), .B0(mai_mai_n1537_), .B1(mai_mai_n162_), .Y(mai_mai_n1539_));
  NA4        m1490(.A(mai_mai_n1539_), .B(mai_mai_n1535_), .C(mai_mai_n1534_), .D(mai_mai_n1530_), .Y(mai_mai_n1540_));
  NO3        m1491(.A(mai_mai_n1075_), .B(mai_mai_n133_), .C(mai_mai_n132_), .Y(mai_mai_n1541_));
  OAI210     m1492(.A0(mai_mai_n1541_), .A1(mai_mai_n655_), .B0(mai_mai_n108_), .Y(mai_mai_n1542_));
  AOI210     m1493(.A0(mai_mai_n1542_), .A1(mai_mai_n563_), .B0(mai_mai_n792_), .Y(mai_mai_n1543_));
  NA3        m1494(.A(mai_mai_n1209_), .B(mai_mai_n192_), .C(mai_mai_n143_), .Y(mai_mai_n1544_));
  NA3        m1495(.A(mai_mai_n1078_), .B(mai_mai_n780_), .C(mai_mai_n346_), .Y(mai_mai_n1545_));
  NA2        m1496(.A(mai_mai_n172_), .B(mai_mai_n777_), .Y(mai_mai_n1546_));
  OAI210     m1497(.A0(mai_mai_n1546_), .A1(mai_mai_n1315_), .B0(mai_mai_n1545_), .Y(mai_mai_n1547_));
  AOI210     m1498(.A0(mai_mai_n1544_), .A1(mai_mai_n179_), .B0(mai_mai_n1547_), .Y(mai_mai_n1548_));
  OAI210     m1499(.A0(mai_mai_n1548_), .A1(mai_mai_n544_), .B0(x4), .Y(mai_mai_n1549_));
  OAI220     m1500(.A0(mai_mai_n1549_), .A1(mai_mai_n1543_), .B0(mai_mai_n1540_), .B1(mai_mai_n1522_), .Y(mai_mai_n1550_));
  NO2        m1501(.A(mai_mai_n147_), .B(mai_mai_n124_), .Y(mai_mai_n1551_));
  NO2        m1502(.A(mai_mai_n192_), .B(mai_mai_n806_), .Y(mai_mai_n1552_));
  AOI210     m1503(.A0(mai_mai_n605_), .A1(mai_mai_n512_), .B0(mai_mai_n1552_), .Y(mai_mai_n1553_));
  NO2        m1504(.A(mai_mai_n1553_), .B(x6), .Y(mai_mai_n1554_));
  NO2        m1505(.A(mai_mai_n389_), .B(mai_mai_n257_), .Y(mai_mai_n1555_));
  NO2        m1506(.A(mai_mai_n133_), .B(mai_mai_n739_), .Y(mai_mai_n1556_));
  NO2        m1507(.A(mai_mai_n960_), .B(mai_mai_n588_), .Y(mai_mai_n1557_));
  AO220      m1508(.A0(mai_mai_n1557_), .A1(mai_mai_n1556_), .B0(mai_mai_n1555_), .B1(mai_mai_n126_), .Y(mai_mai_n1558_));
  NO3        m1509(.A(mai_mai_n1558_), .B(mai_mai_n1554_), .C(mai_mai_n1551_), .Y(mai_mai_n1559_));
  NA2        m1510(.A(mai_mai_n1075_), .B(x3), .Y(mai_mai_n1560_));
  NA2        m1511(.A(mai_mai_n1352_), .B(mai_mai_n135_), .Y(mai_mai_n1561_));
  OAI220     m1512(.A0(mai_mai_n1561_), .A1(mai_mai_n1560_), .B0(mai_mai_n1559_), .B1(x3), .Y(mai_mai_n1562_));
  NO3        m1513(.A(mai_mai_n1007_), .B(mai_mai_n689_), .C(mai_mai_n330_), .Y(mai_mai_n1563_));
  AO210      m1514(.A0(mai_mai_n1036_), .A1(mai_mai_n300_), .B0(mai_mai_n1563_), .Y(mai_mai_n1564_));
  AOI220     m1515(.A0(mai_mai_n1564_), .A1(x8), .B0(mai_mai_n1352_), .B1(mai_mai_n439_), .Y(mai_mai_n1565_));
  NA2        m1516(.A(mai_mai_n753_), .B(mai_mai_n321_), .Y(mai_mai_n1566_));
  NO4        m1517(.A(mai_mai_n371_), .B(mai_mai_n205_), .C(mai_mai_n341_), .D(x2), .Y(mai_mai_n1567_));
  NA2        m1518(.A(mai_mai_n1406_), .B(mai_mai_n110_), .Y(mai_mai_n1568_));
  NO3        m1519(.A(mai_mai_n1211_), .B(mai_mai_n1000_), .C(mai_mai_n1148_), .Y(mai_mai_n1569_));
  AOI210     m1520(.A0(mai_mai_n1569_), .A1(mai_mai_n1568_), .B0(mai_mai_n1567_), .Y(mai_mai_n1570_));
  OA220      m1521(.A0(mai_mai_n1570_), .A1(mai_mai_n960_), .B0(mai_mai_n1566_), .B1(mai_mai_n572_), .Y(mai_mai_n1571_));
  OAI210     m1522(.A0(mai_mai_n1565_), .A1(mai_mai_n413_), .B0(mai_mai_n1571_), .Y(mai_mai_n1572_));
  AOI210     m1523(.A0(mai_mai_n1562_), .A1(mai_mai_n140_), .B0(mai_mai_n1572_), .Y(mai_mai_n1573_));
  NA2        m1524(.A(mai_mai_n1573_), .B(mai_mai_n1550_), .Y(mai19));
  NO2        m1525(.A(mai_mai_n1452_), .B(mai_mai_n261_), .Y(mai_mai_n1575_));
  NA2        m1526(.A(mai_mai_n650_), .B(x3), .Y(mai_mai_n1576_));
  OAI210     m1527(.A0(mai_mai_n155_), .A1(mai_mai_n109_), .B0(mai_mai_n81_), .Y(mai_mai_n1577_));
  NA3        m1528(.A(mai_mai_n1577_), .B(mai_mai_n1576_), .C(mai_mai_n244_), .Y(mai_mai_n1578_));
  NO2        m1529(.A(mai_mai_n1310_), .B(mai_mai_n172_), .Y(mai_mai_n1579_));
  AOI210     m1530(.A0(mai_mai_n1479_), .A1(mai_mai_n356_), .B0(mai_mai_n1579_), .Y(mai_mai_n1580_));
  AOI210     m1531(.A0(mai_mai_n1580_), .A1(mai_mai_n1578_), .B0(mai_mai_n56_), .Y(mai_mai_n1581_));
  NO2        m1532(.A(mai_mai_n865_), .B(mai_mai_n1224_), .Y(mai_mai_n1582_));
  OAI210     m1533(.A0(mai_mai_n1581_), .A1(mai_mai_n1575_), .B0(mai_mai_n1582_), .Y(mai_mai_n1583_));
  NOi21      m1534(.An(mai_mai_n614_), .B(mai_mai_n654_), .Y(mai_mai_n1584_));
  AOI210     m1535(.A0(mai_mai_n356_), .A1(x6), .B0(mai_mai_n123_), .Y(mai_mai_n1585_));
  NO3        m1536(.A(mai_mai_n1585_), .B(mai_mai_n762_), .C(mai_mai_n128_), .Y(mai_mai_n1586_));
  NA2        m1537(.A(mai_mai_n1204_), .B(mai_mai_n124_), .Y(mai_mai_n1587_));
  NO4        m1538(.A(mai_mai_n1587_), .B(mai_mai_n1007_), .C(mai_mai_n894_), .D(mai_mai_n77_), .Y(mai_mai_n1588_));
  NO3        m1539(.A(mai_mai_n1588_), .B(mai_mai_n1586_), .C(mai_mai_n1033_), .Y(mai_mai_n1589_));
  NO2        m1540(.A(mai_mai_n544_), .B(mai_mai_n623_), .Y(mai_mai_n1590_));
  NA2        m1541(.A(mai_mai_n1256_), .B(mai_mai_n50_), .Y(mai_mai_n1591_));
  NO3        m1542(.A(mai_mai_n519_), .B(mai_mai_n309_), .C(mai_mai_n64_), .Y(mai_mai_n1592_));
  AOI220     m1543(.A0(mai_mai_n1592_), .A1(mai_mai_n1591_), .B0(mai_mai_n1590_), .B1(mai_mai_n780_), .Y(mai_mai_n1593_));
  OAI210     m1544(.A0(mai_mai_n1589_), .A1(mai_mai_n57_), .B0(mai_mai_n1593_), .Y(mai_mai_n1594_));
  AOI210     m1545(.A0(mai_mai_n1594_), .A1(mai_mai_n777_), .B0(mai_mai_n1584_), .Y(mai_mai_n1595_));
  AOI210     m1546(.A0(mai_mai_n826_), .A1(mai_mai_n739_), .B0(mai_mai_n767_), .Y(mai_mai_n1596_));
  NO2        m1547(.A(mai_mai_n1596_), .B(x4), .Y(mai_mai_n1597_));
  NA3        m1548(.A(mai_mai_n737_), .B(mai_mai_n260_), .C(x7), .Y(mai_mai_n1598_));
  AOI220     m1549(.A0(mai_mai_n1404_), .A1(mai_mai_n792_), .B0(mai_mai_n703_), .B1(mai_mai_n1164_), .Y(mai_mai_n1599_));
  AOI210     m1550(.A0(mai_mai_n1599_), .A1(mai_mai_n1598_), .B0(mai_mai_n504_), .Y(mai_mai_n1600_));
  OAI210     m1551(.A0(mai_mai_n1600_), .A1(mai_mai_n1597_), .B0(mai_mai_n816_), .Y(mai_mai_n1601_));
  NO2        m1552(.A(mai_mai_n749_), .B(mai_mai_n325_), .Y(mai_mai_n1602_));
  NO2        m1553(.A(mai_mai_n155_), .B(mai_mai_n1032_), .Y(mai_mai_n1603_));
  AOI220     m1554(.A0(mai_mai_n1603_), .A1(mai_mai_n1272_), .B0(mai_mai_n1602_), .B1(mai_mai_n479_), .Y(mai_mai_n1604_));
  AO210      m1555(.A0(mai_mai_n1604_), .A1(mai_mai_n1601_), .B0(x1), .Y(mai_mai_n1605_));
  NA2        m1556(.A(mai_mai_n635_), .B(mai_mai_n1056_), .Y(mai_mai_n1606_));
  NA2        m1557(.A(mai_mai_n148_), .B(mai_mai_n111_), .Y(mai_mai_n1607_));
  NOi21      m1558(.An(x1), .B(x6), .Y(mai_mai_n1608_));
  NA2        m1559(.A(mai_mai_n1608_), .B(mai_mai_n84_), .Y(mai_mai_n1609_));
  NA3        m1560(.A(mai_mai_n1609_), .B(mai_mai_n1607_), .C(mai_mai_n1606_), .Y(mai_mai_n1610_));
  AOI220     m1561(.A0(mai_mai_n1610_), .A1(x3), .B0(mai_mai_n1212_), .B1(mai_mai_n385_), .Y(mai_mai_n1611_));
  NA3        m1562(.A(mai_mai_n1217_), .B(mai_mai_n801_), .C(mai_mai_n606_), .Y(mai_mai_n1612_));
  AOI220     m1563(.A0(mai_mai_n1260_), .A1(mai_mai_n123_), .B0(mai_mai_n924_), .B1(mai_mai_n818_), .Y(mai_mai_n1613_));
  AOI210     m1564(.A0(mai_mai_n1613_), .A1(mai_mai_n1612_), .B0(mai_mai_n325_), .Y(mai_mai_n1614_));
  NA2        m1565(.A(mai_mai_n946_), .B(mai_mai_n50_), .Y(mai_mai_n1615_));
  NA3        m1566(.A(mai_mai_n1204_), .B(mai_mai_n386_), .C(mai_mai_n110_), .Y(mai_mai_n1616_));
  AOI210     m1567(.A0(mai_mai_n1616_), .A1(mai_mai_n1615_), .B0(mai_mai_n970_), .Y(mai_mai_n1617_));
  NO3        m1568(.A(mai_mai_n621_), .B(mai_mai_n518_), .C(mai_mai_n1230_), .Y(mai_mai_n1618_));
  NO3        m1569(.A(mai_mai_n1618_), .B(mai_mai_n1617_), .C(mai_mai_n1614_), .Y(mai_mai_n1619_));
  OAI210     m1570(.A0(mai_mai_n1611_), .A1(mai_mai_n852_), .B0(mai_mai_n1619_), .Y(mai_mai_n1620_));
  NO2        m1571(.A(mai_mai_n557_), .B(mai_mai_n68_), .Y(mai_mai_n1621_));
  OAI220     m1572(.A0(mai_mai_n1621_), .A1(mai_mai_n1576_), .B0(mai_mai_n308_), .B1(mai_mai_n902_), .Y(mai_mai_n1622_));
  AOI220     m1573(.A0(mai_mai_n1622_), .A1(mai_mai_n56_), .B0(mai_mai_n1357_), .B1(mai_mai_n734_), .Y(mai_mai_n1623_));
  NO2        m1574(.A(mai_mai_n54_), .B(mai_mai_n71_), .Y(mai_mai_n1624_));
  AO220      m1575(.A0(mai_mai_n1624_), .A1(mai_mai_n1007_), .B0(mai_mai_n818_), .B1(mai_mai_n959_), .Y(mai_mai_n1625_));
  NA2        m1576(.A(mai_mai_n1188_), .B(mai_mai_n363_), .Y(mai_mai_n1626_));
  NA2        m1577(.A(mai_mai_n500_), .B(mai_mai_n734_), .Y(mai_mai_n1627_));
  OAI210     m1578(.A0(mai_mai_n1627_), .A1(mai_mai_n2667_), .B0(mai_mai_n1626_), .Y(mai_mai_n1628_));
  AOI210     m1579(.A0(mai_mai_n1625_), .A1(x2), .B0(mai_mai_n1628_), .Y(mai_mai_n1629_));
  OAI220     m1580(.A0(mai_mai_n1629_), .A1(mai_mai_n155_), .B0(mai_mai_n1623_), .B1(mai_mai_n54_), .Y(mai_mai_n1630_));
  OAI210     m1581(.A0(mai_mai_n1630_), .A1(mai_mai_n1620_), .B0(x8), .Y(mai_mai_n1631_));
  NA4        m1582(.A(mai_mai_n1631_), .B(mai_mai_n1605_), .C(mai_mai_n1595_), .D(mai_mai_n1583_), .Y(mai20));
  NA4        m1583(.A(mai_mai_n396_), .B(mai_mai_n281_), .C(mai_mai_n384_), .D(mai_mai_n62_), .Y(mai_mai_n1633_));
  NA2        m1584(.A(mai_mai_n479_), .B(mai_mai_n417_), .Y(mai_mai_n1634_));
  AOI210     m1585(.A0(mai_mai_n1634_), .A1(mai_mai_n1633_), .B0(mai_mai_n87_), .Y(mai_mai_n1635_));
  AOI210     m1586(.A0(mai_mai_n1060_), .A1(mai_mai_n62_), .B0(mai_mai_n1590_), .Y(mai_mai_n1636_));
  AOI210     m1587(.A0(mai_mai_n994_), .A1(mai_mai_n352_), .B0(mai_mai_n1195_), .Y(mai_mai_n1637_));
  OAI210     m1588(.A0(mai_mai_n1636_), .A1(mai_mai_n685_), .B0(mai_mai_n1637_), .Y(mai_mai_n1638_));
  OAI210     m1589(.A0(mai_mai_n1638_), .A1(mai_mai_n1635_), .B0(mai_mai_n1113_), .Y(mai_mai_n1639_));
  NAi21      m1590(.An(mai_mai_n553_), .B(mai_mai_n405_), .Y(mai_mai_n1640_));
  NA3        m1591(.A(mai_mai_n1640_), .B(mai_mai_n992_), .C(mai_mai_n959_), .Y(mai_mai_n1641_));
  NA3        m1592(.A(mai_mai_n1112_), .B(mai_mai_n281_), .C(mai_mai_n587_), .Y(mai_mai_n1642_));
  AOI210     m1593(.A0(mai_mai_n1642_), .A1(mai_mai_n1641_), .B0(mai_mai_n1301_), .Y(mai_mai_n1643_));
  NO2        m1594(.A(mai_mai_n753_), .B(mai_mai_n980_), .Y(mai_mai_n1644_));
  NOi31      m1595(.An(mai_mai_n1644_), .B(mai_mai_n1180_), .C(mai_mai_n531_), .Y(mai_mai_n1645_));
  OAI210     m1596(.A0(mai_mai_n1645_), .A1(mai_mai_n1643_), .B0(mai_mai_n330_), .Y(mai_mai_n1646_));
  NA2        m1597(.A(mai_mai_n321_), .B(mai_mai_n93_), .Y(mai_mai_n1647_));
  NA2        m1598(.A(mai_mai_n331_), .B(mai_mai_n108_), .Y(mai_mai_n1648_));
  NA2        m1599(.A(mai_mai_n427_), .B(mai_mai_n52_), .Y(mai_mai_n1649_));
  OAI220     m1600(.A0(mai_mai_n1649_), .A1(mai_mai_n1648_), .B0(mai_mai_n1647_), .B1(mai_mai_n276_), .Y(mai_mai_n1650_));
  NA2        m1601(.A(mai_mai_n1650_), .B(mai_mai_n224_), .Y(mai_mai_n1651_));
  NO2        m1602(.A(mai_mai_n669_), .B(mai_mai_n610_), .Y(mai_mai_n1652_));
  NA2        m1603(.A(mai_mai_n960_), .B(mai_mai_n50_), .Y(mai_mai_n1653_));
  NO3        m1604(.A(mai_mai_n1653_), .B(mai_mai_n369_), .C(mai_mai_n232_), .Y(mai_mai_n1654_));
  NA4        m1605(.A(mai_mai_n342_), .B(mai_mai_n241_), .C(mai_mai_n806_), .D(mai_mai_n64_), .Y(mai_mai_n1655_));
  OAI220     m1606(.A0(mai_mai_n1655_), .A1(mai_mai_n679_), .B0(mai_mai_n1473_), .B1(mai_mai_n1045_), .Y(mai_mai_n1656_));
  AOI210     m1607(.A0(mai_mai_n1654_), .A1(mai_mai_n1652_), .B0(mai_mai_n1656_), .Y(mai_mai_n1657_));
  NA4        m1608(.A(mai_mai_n1657_), .B(mai_mai_n1651_), .C(mai_mai_n1646_), .D(mai_mai_n1639_), .Y(mai21));
  OAI210     m1609(.A0(mai_mai_n410_), .A1(mai_mai_n54_), .B0(x7), .Y(mai_mai_n1659_));
  OAI220     m1610(.A0(mai_mai_n1659_), .A1(mai_mai_n1290_), .B0(mai_mai_n1061_), .B1(mai_mai_n96_), .Y(mai_mai_n1660_));
  NA2        m1611(.A(mai_mai_n1660_), .B(mai_mai_n78_), .Y(mai_mai_n1661_));
  NA2        m1612(.A(mai_mai_n293_), .B(mai_mai_n863_), .Y(mai_mai_n1662_));
  AOI220     m1613(.A0(mai_mai_n1662_), .A1(mai_mai_n311_), .B0(mai_mai_n572_), .B1(mai_mai_n463_), .Y(mai_mai_n1663_));
  NA2        m1614(.A(mai_mai_n946_), .B(mai_mai_n275_), .Y(mai_mai_n1664_));
  NA2        m1615(.A(mai_mai_n539_), .B(mai_mai_n464_), .Y(mai_mai_n1665_));
  NA4        m1616(.A(mai_mai_n1665_), .B(mai_mai_n1664_), .C(mai_mai_n1384_), .D(mai_mai_n56_), .Y(mai_mai_n1666_));
  NO2        m1617(.A(mai_mai_n780_), .B(mai_mai_n438_), .Y(mai_mai_n1667_));
  NO3        m1618(.A(mai_mai_n1667_), .B(mai_mai_n726_), .C(mai_mai_n253_), .Y(mai_mai_n1668_));
  NOi31      m1619(.An(mai_mai_n195_), .B(mai_mai_n635_), .C(mai_mai_n1099_), .Y(mai_mai_n1669_));
  NO4        m1620(.A(mai_mai_n1669_), .B(mai_mai_n1668_), .C(mai_mai_n1666_), .D(mai_mai_n1663_), .Y(mai_mai_n1670_));
  NO3        m1621(.A(mai_mai_n438_), .B(mai_mai_n279_), .C(mai_mai_n52_), .Y(mai_mai_n1671_));
  OA210      m1622(.A0(mai_mai_n1671_), .A1(mai_mai_n891_), .B0(x3), .Y(mai_mai_n1672_));
  OAI210     m1623(.A0(mai_mai_n791_), .A1(mai_mai_n592_), .B0(mai_mai_n344_), .Y(mai_mai_n1673_));
  NO2        m1624(.A(mai_mai_n70_), .B(x2), .Y(mai_mai_n1674_));
  OAI210     m1625(.A0(mai_mai_n179_), .A1(x0), .B0(mai_mai_n1674_), .Y(mai_mai_n1675_));
  NA2        m1626(.A(mai_mai_n1675_), .B(mai_mai_n1673_), .Y(mai_mai_n1676_));
  OAI210     m1627(.A0(mai_mai_n1676_), .A1(mai_mai_n1672_), .B0(x8), .Y(mai_mai_n1677_));
  NO3        m1628(.A(mai_mai_n778_), .B(mai_mai_n624_), .C(mai_mai_n588_), .Y(mai_mai_n1678_));
  NA2        m1629(.A(mai_mai_n55_), .B(mai_mai_n50_), .Y(mai_mai_n1679_));
  MUX2       m1630(.S(mai_mai_n604_), .A(mai_mai_n1679_), .B(mai_mai_n107_), .Y(mai_mai_n1680_));
  AOI210     m1631(.A0(mai_mai_n1362_), .A1(mai_mai_n242_), .B0(mai_mai_n1680_), .Y(mai_mai_n1681_));
  OAI210     m1632(.A0(mai_mai_n646_), .A1(mai_mai_n587_), .B0(x4), .Y(mai_mai_n1682_));
  NO3        m1633(.A(mai_mai_n1682_), .B(mai_mai_n1681_), .C(mai_mai_n1678_), .Y(mai_mai_n1683_));
  AO220      m1634(.A0(mai_mai_n1683_), .A1(mai_mai_n1677_), .B0(mai_mai_n1670_), .B1(mai_mai_n1661_), .Y(mai_mai_n1684_));
  AO220      m1635(.A0(mai_mai_n636_), .A1(mai_mai_n325_), .B0(mai_mai_n593_), .B1(x8), .Y(mai_mai_n1685_));
  NO2        m1636(.A(mai_mai_n865_), .B(x0), .Y(mai_mai_n1686_));
  NO3        m1637(.A(mai_mai_n1686_), .B(mai_mai_n549_), .C(mai_mai_n88_), .Y(mai_mai_n1687_));
  NO2        m1638(.A(mai_mai_n161_), .B(x2), .Y(mai_mai_n1688_));
  NO3        m1639(.A(mai_mai_n382_), .B(mai_mai_n258_), .C(mai_mai_n187_), .Y(mai_mai_n1689_));
  AOI210     m1640(.A0(mai_mai_n1688_), .A1(mai_mai_n68_), .B0(mai_mai_n1689_), .Y(mai_mai_n1690_));
  OAI210     m1641(.A0(mai_mai_n1687_), .A1(mai_mai_n403_), .B0(mai_mai_n1690_), .Y(mai_mai_n1691_));
  AOI220     m1642(.A0(mai_mai_n1691_), .A1(x5), .B0(mai_mai_n1685_), .B1(mai_mai_n753_), .Y(mai_mai_n1692_));
  AOI210     m1643(.A0(mai_mai_n1692_), .A1(mai_mai_n1684_), .B0(mai_mai_n71_), .Y(mai_mai_n1693_));
  NO2        m1644(.A(mai_mai_n914_), .B(mai_mai_n170_), .Y(mai_mai_n1694_));
  NOi41      m1645(.An(mai_mai_n1435_), .B(mai_mai_n1508_), .C(mai_mai_n1163_), .D(mai_mai_n856_), .Y(mai_mai_n1695_));
  NA2        m1646(.A(mai_mai_n1695_), .B(mai_mai_n1694_), .Y(mai_mai_n1696_));
  NO2        m1647(.A(mai_mai_n78_), .B(x4), .Y(mai_mai_n1697_));
  OAI210     m1648(.A0(mai_mai_n291_), .A1(mai_mai_n159_), .B0(mai_mai_n1697_), .Y(mai_mai_n1698_));
  OAI210     m1649(.A0(mai_mai_n412_), .A1(mai_mai_n428_), .B0(mai_mai_n232_), .Y(mai_mai_n1699_));
  NO2        m1650(.A(mai_mai_n260_), .B(mai_mai_n50_), .Y(mai_mai_n1700_));
  NO2        m1651(.A(mai_mai_n1700_), .B(mai_mai_n57_), .Y(mai_mai_n1701_));
  NA2        m1652(.A(mai_mai_n1701_), .B(mai_mai_n1699_), .Y(mai_mai_n1702_));
  AOI210     m1653(.A0(mai_mai_n1698_), .A1(mai_mai_n1696_), .B0(mai_mai_n1702_), .Y(mai_mai_n1703_));
  NA2        m1654(.A(mai_mai_n764_), .B(mai_mai_n553_), .Y(mai_mai_n1704_));
  AO210      m1655(.A0(mai_mai_n1704_), .A1(mai_mai_n970_), .B0(mai_mai_n50_), .Y(mai_mai_n1705_));
  NO2        m1656(.A(mai_mai_n1640_), .B(mai_mai_n1224_), .Y(mai_mai_n1706_));
  AOI220     m1657(.A0(mai_mai_n1706_), .A1(mai_mai_n1173_), .B0(mai_mai_n1329_), .B1(mai_mai_n1054_), .Y(mai_mai_n1707_));
  AOI210     m1658(.A0(mai_mai_n1707_), .A1(mai_mai_n1705_), .B0(mai_mai_n110_), .Y(mai_mai_n1708_));
  NA2        m1659(.A(mai_mai_n300_), .B(mai_mai_n108_), .Y(mai_mai_n1709_));
  NA2        m1660(.A(mai_mai_n901_), .B(mai_mai_n55_), .Y(mai_mai_n1710_));
  NO2        m1661(.A(mai_mai_n1710_), .B(mai_mai_n1709_), .Y(mai_mai_n1711_));
  NO2        m1662(.A(mai_mai_n674_), .B(mai_mai_n1064_), .Y(mai_mai_n1712_));
  NO4        m1663(.A(mai_mai_n1712_), .B(mai_mai_n1711_), .C(mai_mai_n1708_), .D(mai_mai_n1703_), .Y(mai_mai_n1713_));
  NO2        m1664(.A(mai_mai_n1713_), .B(x6), .Y(mai_mai_n1714_));
  AOI210     m1665(.A0(mai_mai_n613_), .A1(mai_mai_n1064_), .B0(mai_mai_n1508_), .Y(mai_mai_n1715_));
  OAI210     m1666(.A0(mai_mai_n1715_), .A1(mai_mai_n692_), .B0(mai_mai_n56_), .Y(mai_mai_n1716_));
  NO2        m1667(.A(mai_mai_n755_), .B(mai_mai_n54_), .Y(mai_mai_n1717_));
  NO2        m1668(.A(mai_mai_n870_), .B(x5), .Y(mai_mai_n1718_));
  NO3        m1669(.A(mai_mai_n1718_), .B(mai_mai_n1717_), .C(mai_mai_n953_), .Y(mai_mai_n1719_));
  AOI210     m1670(.A0(mai_mai_n1719_), .A1(mai_mai_n1716_), .B0(mai_mai_n50_), .Y(mai_mai_n1720_));
  NA2        m1671(.A(mai_mai_n161_), .B(mai_mai_n108_), .Y(mai_mai_n1721_));
  OA220      m1672(.A0(mai_mai_n1721_), .A1(mai_mai_n442_), .B0(mai_mai_n469_), .B1(mai_mai_n753_), .Y(mai_mai_n1722_));
  NA3        m1673(.A(mai_mai_n55_), .B(x2), .C(x0), .Y(mai_mai_n1723_));
  AOI220     m1674(.A0(mai_mai_n1723_), .A1(mai_mai_n172_), .B0(mai_mai_n870_), .B1(mai_mai_n157_), .Y(mai_mai_n1724_));
  NO2        m1675(.A(mai_mai_n685_), .B(mai_mai_n260_), .Y(mai_mai_n1725_));
  NO3        m1676(.A(mai_mai_n248_), .B(mai_mai_n230_), .C(mai_mai_n363_), .Y(mai_mai_n1726_));
  NO3        m1677(.A(mai_mai_n1726_), .B(mai_mai_n1725_), .C(mai_mai_n1724_), .Y(mai_mai_n1727_));
  OAI220     m1678(.A0(mai_mai_n1727_), .A1(mai_mai_n56_), .B0(mai_mai_n1722_), .B1(mai_mai_n701_), .Y(mai_mai_n1728_));
  OAI210     m1679(.A0(mai_mai_n1728_), .A1(mai_mai_n1720_), .B0(mai_mai_n116_), .Y(mai_mai_n1729_));
  NO2        m1680(.A(mai_mai_n618_), .B(mai_mai_n306_), .Y(mai_mai_n1730_));
  AOI210     m1681(.A0(mai_mai_n611_), .A1(x5), .B0(mai_mai_n1730_), .Y(mai_mai_n1731_));
  NO2        m1682(.A(mai_mai_n1731_), .B(mai_mai_n110_), .Y(mai_mai_n1732_));
  NA2        m1683(.A(mai_mai_n709_), .B(mai_mai_n81_), .Y(mai_mai_n1733_));
  NA3        m1684(.A(mai_mai_n1733_), .B(mai_mai_n435_), .C(mai_mai_n57_), .Y(mai_mai_n1734_));
  OAI210     m1685(.A0(mai_mai_n1710_), .A1(mai_mai_n1709_), .B0(mai_mai_n1734_), .Y(mai_mai_n1735_));
  OAI210     m1686(.A0(mai_mai_n1735_), .A1(mai_mai_n1732_), .B0(x1), .Y(mai_mai_n1736_));
  NO4        m1687(.A(mai_mai_n421_), .B(mai_mai_n78_), .C(mai_mai_n149_), .D(x3), .Y(mai_mai_n1737_));
  NO2        m1688(.A(mai_mai_n331_), .B(mai_mai_n112_), .Y(mai_mai_n1738_));
  OAI210     m1689(.A0(mai_mai_n1737_), .A1(mai_mai_n1302_), .B0(mai_mai_n1738_), .Y(mai_mai_n1739_));
  NO2        m1690(.A(mai_mai_n60_), .B(mai_mai_n108_), .Y(mai_mai_n1740_));
  NO4        m1691(.A(mai_mai_n1709_), .B(mai_mai_n968_), .C(mai_mai_n669_), .D(mai_mai_n50_), .Y(mai_mai_n1741_));
  AOI210     m1692(.A0(mai_mai_n1740_), .A1(mai_mai_n1552_), .B0(mai_mai_n1741_), .Y(mai_mai_n1742_));
  NA4        m1693(.A(mai_mai_n1742_), .B(mai_mai_n1739_), .C(mai_mai_n1736_), .D(mai_mai_n1729_), .Y(mai_mai_n1743_));
  NO3        m1694(.A(mai_mai_n1743_), .B(mai_mai_n1714_), .C(mai_mai_n1693_), .Y(mai22));
  AOI210     m1695(.A0(mai_mai_n525_), .A1(mai_mai_n71_), .B0(mai_mai_n472_), .Y(mai_mai_n1745_));
  NO3        m1696(.A(mai_mai_n1200_), .B(mai_mai_n557_), .C(mai_mai_n703_), .Y(mai_mai_n1746_));
  AOI210     m1697(.A0(x5), .A1(x2), .B0(x8), .Y(mai_mai_n1747_));
  NA2        m1698(.A(mai_mai_n1747_), .B(mai_mai_n59_), .Y(mai_mai_n1748_));
  OAI220     m1699(.A0(mai_mai_n1748_), .A1(mai_mai_n1746_), .B0(mai_mai_n1745_), .B1(mai_mai_n403_), .Y(mai_mai_n1749_));
  NA2        m1700(.A(mai_mai_n587_), .B(mai_mai_n87_), .Y(mai_mai_n1750_));
  NA2        m1701(.A(mai_mai_n276_), .B(mai_mai_n77_), .Y(mai_mai_n1751_));
  OA220      m1702(.A0(mai_mai_n1751_), .A1(mai_mai_n1750_), .B0(mai_mai_n849_), .B1(mai_mai_n1017_), .Y(mai_mai_n1752_));
  NO4        m1703(.A(mai_mai_n389_), .B(mai_mai_n222_), .C(mai_mai_n71_), .D(x3), .Y(mai_mai_n1753_));
  NO3        m1704(.A(mai_mai_n1253_), .B(mai_mai_n87_), .C(x0), .Y(mai_mai_n1754_));
  OAI210     m1705(.A0(mai_mai_n403_), .A1(mai_mai_n207_), .B0(x4), .Y(mai_mai_n1755_));
  NO2        m1706(.A(mai_mai_n1755_), .B(mai_mai_n1753_), .Y(mai_mai_n1756_));
  OAI210     m1707(.A0(mai_mai_n1752_), .A1(mai_mai_n200_), .B0(mai_mai_n1756_), .Y(mai_mai_n1757_));
  AOI210     m1708(.A0(mai_mai_n1749_), .A1(mai_mai_n53_), .B0(mai_mai_n1757_), .Y(mai_mai_n1758_));
  NA2        m1709(.A(mai_mai_n304_), .B(mai_mai_n309_), .Y(mai_mai_n1759_));
  NA3        m1710(.A(mai_mai_n1759_), .B(mai_mai_n224_), .C(mai_mai_n308_), .Y(mai_mai_n1760_));
  NA2        m1711(.A(mai_mai_n582_), .B(mai_mai_n247_), .Y(mai_mai_n1761_));
  NO3        m1712(.A(mai_mai_n500_), .B(mai_mai_n268_), .C(mai_mai_n216_), .Y(mai_mai_n1762_));
  NAi31      m1713(.An(mai_mai_n1762_), .B(mai_mai_n1761_), .C(mai_mai_n1760_), .Y(mai_mai_n1763_));
  NO2        m1714(.A(mai_mai_n469_), .B(mai_mai_n262_), .Y(mai_mai_n1764_));
  NO2        m1715(.A(mai_mai_n1253_), .B(x3), .Y(mai_mai_n1765_));
  AOI210     m1716(.A0(mai_mai_n1765_), .A1(mai_mai_n352_), .B0(mai_mai_n1764_), .Y(mai_mai_n1766_));
  OAI210     m1717(.A0(mai_mai_n1094_), .A1(mai_mai_n189_), .B0(mai_mai_n56_), .Y(mai_mai_n1767_));
  NA3        m1718(.A(mai_mai_n55_), .B(mai_mai_n71_), .C(x0), .Y(mai_mai_n1768_));
  OAI220     m1719(.A0(mai_mai_n1768_), .A1(mai_mai_n1064_), .B0(mai_mai_n369_), .B1(mai_mai_n215_), .Y(mai_mai_n1769_));
  NO2        m1720(.A(mai_mai_n1769_), .B(mai_mai_n1767_), .Y(mai_mai_n1770_));
  OAI210     m1721(.A0(mai_mai_n1766_), .A1(mai_mai_n260_), .B0(mai_mai_n1770_), .Y(mai_mai_n1771_));
  AOI210     m1722(.A0(mai_mai_n1763_), .A1(mai_mai_n108_), .B0(mai_mai_n1771_), .Y(mai_mai_n1772_));
  AOI210     m1723(.A0(mai_mai_n957_), .A1(mai_mai_n779_), .B0(mai_mai_n874_), .Y(mai_mai_n1773_));
  OAI210     m1724(.A0(mai_mai_n808_), .A1(mai_mai_n161_), .B0(mai_mai_n943_), .Y(mai_mai_n1774_));
  OAI210     m1725(.A0(mai_mai_n1774_), .A1(mai_mai_n1773_), .B0(mai_mai_n617_), .Y(mai_mai_n1775_));
  OA210      m1726(.A0(mai_mai_n1772_), .A1(mai_mai_n1758_), .B0(mai_mai_n1775_), .Y(mai_mai_n1776_));
  OAI210     m1727(.A0(mai_mai_n1182_), .A1(mai_mai_n708_), .B0(mai_mai_n696_), .Y(mai_mai_n1777_));
  NO2        m1728(.A(mai_mai_n357_), .B(x0), .Y(mai_mai_n1778_));
  NA3        m1729(.A(mai_mai_n1778_), .B(mai_mai_n352_), .C(mai_mai_n56_), .Y(mai_mai_n1779_));
  AOI210     m1730(.A0(mai_mai_n1779_), .A1(mai_mai_n1777_), .B0(mai_mai_n403_), .Y(mai_mai_n1780_));
  NO3        m1731(.A(mai_mai_n172_), .B(mai_mai_n161_), .C(mai_mai_n62_), .Y(mai_mai_n1781_));
  OAI210     m1732(.A0(mai_mai_n1781_), .A1(mai_mai_n423_), .B0(mai_mai_n110_), .Y(mai_mai_n1782_));
  NA2        m1733(.A(mai_mai_n143_), .B(mai_mai_n792_), .Y(mai_mai_n1783_));
  NA2        m1734(.A(mai_mai_n421_), .B(x3), .Y(mai_mai_n1784_));
  NAi31      m1735(.An(mai_mai_n1784_), .B(mai_mai_n1783_), .C(mai_mai_n1568_), .Y(mai_mai_n1785_));
  NO3        m1736(.A(mai_mai_n865_), .B(mai_mai_n468_), .C(mai_mai_n110_), .Y(mai_mai_n1786_));
  NO2        m1737(.A(mai_mai_n1096_), .B(mai_mai_n144_), .Y(mai_mai_n1787_));
  NO3        m1738(.A(mai_mai_n904_), .B(mai_mai_n417_), .C(mai_mai_n305_), .Y(mai_mai_n1788_));
  AOI220     m1739(.A0(mai_mai_n1788_), .A1(mai_mai_n1787_), .B0(mai_mai_n1786_), .B1(mai_mai_n1778_), .Y(mai_mai_n1789_));
  NA3        m1740(.A(mai_mai_n417_), .B(mai_mai_n93_), .C(mai_mai_n81_), .Y(mai_mai_n1790_));
  AOI210     m1741(.A0(mai_mai_n613_), .A1(mai_mai_n460_), .B0(mai_mai_n498_), .Y(mai_mai_n1791_));
  NA2        m1742(.A(mai_mai_n1184_), .B(x3), .Y(mai_mai_n1792_));
  OAI210     m1743(.A0(mai_mai_n1792_), .A1(mai_mai_n1791_), .B0(mai_mai_n1790_), .Y(mai_mai_n1793_));
  NA3        m1744(.A(mai_mai_n56_), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n1794_));
  NOi21      m1745(.An(mai_mai_n83_), .B(mai_mai_n737_), .Y(mai_mai_n1795_));
  NA3        m1746(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n1796_));
  NA3        m1747(.A(mai_mai_n1796_), .B(mai_mai_n1000_), .C(mai_mai_n269_), .Y(mai_mai_n1797_));
  OAI220     m1748(.A0(mai_mai_n1797_), .A1(mai_mai_n1795_), .B0(mai_mai_n1067_), .B1(mai_mai_n1794_), .Y(mai_mai_n1798_));
  AOI220     m1749(.A0(mai_mai_n1798_), .A1(mai_mai_n1078_), .B0(mai_mai_n1793_), .B1(mai_mai_n352_), .Y(mai_mai_n1799_));
  NA4        m1750(.A(mai_mai_n1799_), .B(mai_mai_n1789_), .C(mai_mai_n1785_), .D(mai_mai_n1782_), .Y(mai_mai_n1800_));
  AOI210     m1751(.A0(mai_mai_n1800_), .A1(x7), .B0(mai_mai_n1780_), .Y(mai_mai_n1801_));
  OAI210     m1752(.A0(mai_mai_n1776_), .A1(x7), .B0(mai_mai_n1801_), .Y(mai23));
  OR2        m1753(.A(mai_mai_n519_), .B(mai_mai_n224_), .Y(mai_mai_n1803_));
  AOI220     m1754(.A0(mai_mai_n1803_), .A1(mai_mai_n1644_), .B0(mai_mai_n619_), .B1(mai_mai_n296_), .Y(mai_mai_n1804_));
  NO3        m1755(.A(mai_mai_n849_), .B(mai_mai_n596_), .C(mai_mai_n491_), .Y(mai_mai_n1805_));
  NO3        m1756(.A(mai_mai_n961_), .B(mai_mai_n150_), .C(mai_mai_n117_), .Y(mai_mai_n1806_));
  AOI210     m1757(.A0(mai_mai_n1806_), .A1(mai_mai_n1039_), .B0(mai_mai_n1805_), .Y(mai_mai_n1807_));
  OAI210     m1758(.A0(mai_mai_n1804_), .A1(mai_mai_n155_), .B0(mai_mai_n1807_), .Y(mai_mai_n1808_));
  NA2        m1759(.A(mai_mai_n1808_), .B(mai_mai_n55_), .Y(mai_mai_n1809_));
  NO2        m1760(.A(mai_mai_n968_), .B(mai_mai_n517_), .Y(mai_mai_n1810_));
  AO220      m1761(.A0(mai_mai_n1286_), .A1(mai_mai_n183_), .B0(mai_mai_n1007_), .B1(mai_mai_n753_), .Y(mai_mai_n1811_));
  OAI210     m1762(.A0(mai_mai_n1811_), .A1(mai_mai_n1810_), .B0(mai_mai_n593_), .Y(mai_mai_n1812_));
  NA2        m1763(.A(mai_mai_n180_), .B(mai_mai_n170_), .Y(mai_mai_n1813_));
  NA2        m1764(.A(mai_mai_n409_), .B(mai_mai_n162_), .Y(mai_mai_n1814_));
  AOI210     m1765(.A0(mai_mai_n1814_), .A1(mai_mai_n1813_), .B0(mai_mai_n239_), .Y(mai_mai_n1815_));
  NA3        m1766(.A(mai_mai_n874_), .B(mai_mai_n428_), .C(mai_mai_n260_), .Y(mai_mai_n1816_));
  AOI210     m1767(.A0(mai_mai_n1816_), .A1(mai_mai_n502_), .B0(mai_mai_n386_), .Y(mai_mai_n1817_));
  OAI210     m1768(.A0(mai_mai_n1817_), .A1(mai_mai_n1815_), .B0(mai_mai_n300_), .Y(mai_mai_n1818_));
  NA3        m1769(.A(mai_mai_n57_), .B(x4), .C(x3), .Y(mai_mai_n1819_));
  NO3        m1770(.A(mai_mai_n1819_), .B(mai_mai_n750_), .C(mai_mai_n143_), .Y(mai_mai_n1820_));
  INV        m1771(.A(mai_mai_n1820_), .Y(mai_mai_n1821_));
  NA4        m1772(.A(mai_mai_n1821_), .B(mai_mai_n1818_), .C(mai_mai_n1812_), .D(mai_mai_n1809_), .Y(mai24));
  NO2        m1773(.A(mai_mai_n244_), .B(x1), .Y(mai_mai_n1823_));
  NA2        m1774(.A(mai_mai_n342_), .B(mai_mai_n495_), .Y(mai_mai_n1824_));
  BUFFER     m1775(.A(mai_mai_n1823_), .Y(mai_mai_n1825_));
  NO3        m1776(.A(mai_mai_n544_), .B(mai_mai_n688_), .C(mai_mai_n157_), .Y(mai_mai_n1826_));
  AOI210     m1777(.A0(mai_mai_n1825_), .A1(mai_mai_n93_), .B0(mai_mai_n1826_), .Y(mai_mai_n1827_));
  NA2        m1778(.A(mai_mai_n102_), .B(x8), .Y(mai_mai_n1828_));
  AN2        m1779(.A(mai_mai_n1274_), .B(mai_mai_n330_), .Y(mai_mai_n1829_));
  NA2        m1780(.A(mai_mai_n460_), .B(x8), .Y(mai_mai_n1830_));
  NA2        m1781(.A(mai_mai_n670_), .B(mai_mai_n126_), .Y(mai_mai_n1831_));
  OAI220     m1782(.A0(mai_mai_n1831_), .A1(mai_mai_n1444_), .B0(mai_mai_n1830_), .B1(mai_mai_n847_), .Y(mai_mai_n1832_));
  AOI220     m1783(.A0(mai_mai_n1832_), .A1(mai_mai_n1700_), .B0(mai_mai_n1829_), .B1(mai_mai_n1039_), .Y(mai_mai_n1833_));
  OAI210     m1784(.A0(mai_mai_n1828_), .A1(mai_mai_n1827_), .B0(mai_mai_n1833_), .Y(mai25));
  NA2        m1785(.A(mai_mai_n331_), .B(mai_mai_n59_), .Y(mai_mai_n1835_));
  NO2        m1786(.A(mai_mai_n1835_), .B(mai_mai_n322_), .Y(mai_mai_n1836_));
  OAI210     m1787(.A0(mai_mai_n1836_), .A1(mai_mai_n1189_), .B0(mai_mai_n116_), .Y(mai_mai_n1837_));
  NA2        m1788(.A(mai_mai_n1602_), .B(mai_mai_n1190_), .Y(mai_mai_n1838_));
  AOI210     m1789(.A0(mai_mai_n1838_), .A1(mai_mai_n1837_), .B0(mai_mai_n683_), .Y(mai_mai_n1839_));
  NO3        m1790(.A(mai_mai_n1051_), .B(mai_mai_n145_), .C(mai_mai_n78_), .Y(mai_mai_n1840_));
  OAI210     m1791(.A0(mai_mai_n200_), .A1(mai_mai_n276_), .B0(mai_mai_n332_), .Y(mai_mai_n1841_));
  OAI210     m1792(.A0(mai_mai_n1841_), .A1(mai_mai_n1840_), .B0(mai_mai_n1188_), .Y(mai_mai_n1842_));
  NO2        m1793(.A(mai_mai_n1396_), .B(mai_mai_n453_), .Y(mai_mai_n1843_));
  NO3        m1794(.A(mai_mai_n1843_), .B(mai_mai_n535_), .C(mai_mai_n99_), .Y(mai_mai_n1844_));
  NA2        m1795(.A(mai_mai_n512_), .B(mai_mai_n55_), .Y(mai_mai_n1845_));
  OAI220     m1796(.A0(mai_mai_n1845_), .A1(mai_mai_n244_), .B0(mai_mai_n590_), .B1(mai_mai_n276_), .Y(mai_mai_n1846_));
  OAI210     m1797(.A0(mai_mai_n1846_), .A1(mai_mai_n1844_), .B0(mai_mai_n640_), .Y(mai_mai_n1847_));
  NA2        m1798(.A(mai_mai_n1764_), .B(mai_mai_n1142_), .Y(mai_mai_n1848_));
  NA3        m1799(.A(mai_mai_n1848_), .B(mai_mai_n1847_), .C(mai_mai_n1842_), .Y(mai_mai_n1849_));
  AO210      m1800(.A0(mai_mai_n1849_), .A1(mai_mai_n108_), .B0(mai_mai_n1839_), .Y(mai26));
  NA2        m1801(.A(mai_mai_n777_), .B(mai_mai_n50_), .Y(mai_mai_n1851_));
  OAI220     m1802(.A0(mai_mai_n306_), .A1(mai_mai_n253_), .B0(mai_mai_n1851_), .B1(x7), .Y(mai_mai_n1852_));
  AOI220     m1803(.A0(mai_mai_n1852_), .A1(mai_mai_n93_), .B0(mai_mai_n1302_), .B1(mai_mai_n1148_), .Y(mai_mai_n1853_));
  NA2        m1804(.A(mai_mai_n628_), .B(mai_mai_n582_), .Y(mai_mai_n1854_));
  OAI210     m1805(.A0(mai_mai_n636_), .A1(mai_mai_n628_), .B0(mai_mai_n753_), .Y(mai_mai_n1855_));
  AOI210     m1806(.A0(mai_mai_n1854_), .A1(mai_mai_n1211_), .B0(mai_mai_n1855_), .Y(mai_mai_n1856_));
  NA2        m1807(.A(mai_mai_n1787_), .B(mai_mai_n1467_), .Y(mai_mai_n1857_));
  NO2        m1808(.A(mai_mai_n1096_), .B(mai_mai_n75_), .Y(mai_mai_n1858_));
  NA2        m1809(.A(mai_mai_n816_), .B(mai_mai_n179_), .Y(mai_mai_n1859_));
  NO2        m1810(.A(mai_mai_n1859_), .B(mai_mai_n540_), .Y(mai_mai_n1860_));
  AOI210     m1811(.A0(mai_mai_n1858_), .A1(mai_mai_n589_), .B0(mai_mai_n1860_), .Y(mai_mai_n1861_));
  OAI220     m1812(.A0(mai_mai_n1861_), .A1(mai_mai_n108_), .B0(mai_mai_n1857_), .B1(mai_mai_n53_), .Y(mai_mai_n1862_));
  NA2        m1813(.A(mai_mai_n605_), .B(mai_mai_n512_), .Y(mai_mai_n1863_));
  NO2        m1814(.A(mai_mai_n136_), .B(mai_mai_n133_), .Y(mai_mai_n1864_));
  NA2        m1815(.A(mai_mai_n1864_), .B(mai_mai_n123_), .Y(mai_mai_n1865_));
  NA2        m1816(.A(mai_mai_n753_), .B(x3), .Y(mai_mai_n1866_));
  AOI210     m1817(.A0(mai_mai_n1865_), .A1(mai_mai_n1863_), .B0(mai_mai_n1866_), .Y(mai_mai_n1867_));
  NO2        m1818(.A(mai_mai_n1017_), .B(x3), .Y(mai_mai_n1868_));
  AOI210     m1819(.A0(mai_mai_n451_), .A1(mai_mai_n108_), .B0(mai_mai_n1868_), .Y(mai_mai_n1869_));
  NA3        m1820(.A(mai_mai_n573_), .B(mai_mai_n51_), .C(mai_mai_n56_), .Y(mai_mai_n1870_));
  AOI210     m1821(.A0(mai_mai_n1652_), .A1(mai_mai_n1068_), .B0(x0), .Y(mai_mai_n1871_));
  OAI210     m1822(.A0(mai_mai_n1870_), .A1(mai_mai_n1869_), .B0(mai_mai_n1871_), .Y(mai_mai_n1872_));
  NO4        m1823(.A(mai_mai_n1872_), .B(mai_mai_n1867_), .C(mai_mai_n1862_), .D(mai_mai_n1856_), .Y(mai_mai_n1873_));
  AOI210     m1824(.A0(x8), .A1(x6), .B0(x5), .Y(mai_mai_n1874_));
  AO220      m1825(.A0(mai_mai_n1874_), .A1(mai_mai_n146_), .B0(mai_mai_n596_), .B1(mai_mai_n143_), .Y(mai_mai_n1875_));
  NA2        m1826(.A(mai_mai_n1875_), .B(mai_mai_n452_), .Y(mai_mai_n1876_));
  NO2        m1827(.A(mai_mai_n763_), .B(mai_mai_n146_), .Y(mai_mai_n1877_));
  NA3        m1828(.A(mai_mai_n1877_), .B(mai_mai_n1674_), .C(mai_mai_n137_), .Y(mai_mai_n1878_));
  NO2        m1829(.A(mai_mai_n403_), .B(mai_mai_n1382_), .Y(mai_mai_n1879_));
  OAI210     m1830(.A0(mai_mai_n1879_), .A1(mai_mai_n1349_), .B0(mai_mai_n451_), .Y(mai_mai_n1880_));
  NA3        m1831(.A(mai_mai_n377_), .B(mai_mai_n863_), .C(mai_mai_n257_), .Y(mai_mai_n1881_));
  NA4        m1832(.A(mai_mai_n1881_), .B(mai_mai_n1880_), .C(mai_mai_n1878_), .D(mai_mai_n1876_), .Y(mai_mai_n1882_));
  AOI210     m1833(.A0(mai_mai_n226_), .A1(x2), .B0(mai_mai_n496_), .Y(mai_mai_n1883_));
  NO2        m1834(.A(mai_mai_n1883_), .B(mai_mai_n117_), .Y(mai_mai_n1884_));
  NA3        m1835(.A(mai_mai_n818_), .B(mai_mai_n1017_), .C(x7), .Y(mai_mai_n1885_));
  AOI210     m1836(.A0(mai_mai_n346_), .A1(mai_mai_n218_), .B0(mai_mai_n1885_), .Y(mai_mai_n1886_));
  OAI220     m1837(.A0(mai_mai_n907_), .A1(mai_mai_n306_), .B0(mai_mai_n646_), .B1(mai_mai_n688_), .Y(mai_mai_n1887_));
  NO3        m1838(.A(mai_mai_n1887_), .B(mai_mai_n1886_), .C(mai_mai_n1884_), .Y(mai_mai_n1888_));
  NA3        m1839(.A(mai_mai_n670_), .B(mai_mai_n194_), .C(mai_mai_n959_), .Y(mai_mai_n1889_));
  NA2        m1840(.A(mai_mai_n1889_), .B(mai_mai_n646_), .Y(mai_mai_n1890_));
  NA2        m1841(.A(mai_mai_n143_), .B(mai_mai_n135_), .Y(mai_mai_n1891_));
  OAI210     m1842(.A0(mai_mai_n1891_), .A1(mai_mai_n1430_), .B0(x0), .Y(mai_mai_n1892_));
  AOI210     m1843(.A0(mai_mai_n1890_), .A1(mai_mai_n1418_), .B0(mai_mai_n1892_), .Y(mai_mai_n1893_));
  OAI210     m1844(.A0(mai_mai_n1888_), .A1(mai_mai_n53_), .B0(mai_mai_n1893_), .Y(mai_mai_n1894_));
  AOI210     m1845(.A0(mai_mai_n1882_), .A1(x4), .B0(mai_mai_n1894_), .Y(mai_mai_n1895_));
  OA220      m1846(.A0(mai_mai_n1895_), .A1(mai_mai_n1873_), .B0(mai_mai_n1853_), .B1(mai_mai_n109_), .Y(mai27));
  NA2        m1847(.A(mai_mai_n1152_), .B(mai_mai_n451_), .Y(mai_mai_n1897_));
  NO2        m1848(.A(mai_mai_n1897_), .B(mai_mai_n301_), .Y(mai_mai_n1898_));
  NA2        m1849(.A(mai_mai_n924_), .B(mai_mai_n818_), .Y(mai_mai_n1899_));
  NA3        m1850(.A(mai_mai_n824_), .B(mai_mai_n366_), .C(mai_mai_n1032_), .Y(mai_mai_n1900_));
  AOI210     m1851(.A0(mai_mai_n1900_), .A1(mai_mai_n1899_), .B0(mai_mai_n218_), .Y(mai_mai_n1901_));
  OAI210     m1852(.A0(mai_mai_n1901_), .A1(mai_mai_n1898_), .B0(mai_mai_n704_), .Y(mai_mai_n1902_));
  XO2        m1853(.A(x8), .B(x4), .Y(mai_mai_n1903_));
  NO3        m1854(.A(mai_mai_n1903_), .B(mai_mai_n451_), .C(mai_mai_n172_), .Y(mai_mai_n1904_));
  OA210      m1855(.A0(mai_mai_n1904_), .A1(mai_mai_n1257_), .B0(mai_mai_n279_), .Y(mai_mai_n1905_));
  NO2        m1856(.A(mai_mai_n398_), .B(mai_mai_n166_), .Y(mai_mai_n1906_));
  OAI210     m1857(.A0(mai_mai_n1906_), .A1(mai_mai_n1905_), .B0(mai_mai_n1130_), .Y(mai_mai_n1907_));
  AOI210     m1858(.A0(mai_mai_n636_), .A1(mai_mai_n56_), .B0(mai_mai_n1858_), .Y(mai_mai_n1908_));
  OAI220     m1859(.A0(mai_mai_n1908_), .A1(mai_mai_n1256_), .B0(mai_mai_n1209_), .B1(mai_mai_n209_), .Y(mai_mai_n1909_));
  NO2        m1860(.A(mai_mai_n701_), .B(mai_mai_n145_), .Y(mai_mai_n1910_));
  NO2        m1861(.A(mai_mai_n1194_), .B(mai_mai_n260_), .Y(mai_mai_n1911_));
  AOI220     m1862(.A0(mai_mai_n1911_), .A1(mai_mai_n1910_), .B0(mai_mai_n1909_), .B1(mai_mai_n539_), .Y(mai_mai_n1912_));
  NA3        m1863(.A(mai_mai_n1912_), .B(mai_mai_n1907_), .C(mai_mai_n1902_), .Y(mai28));
  NO3        m1864(.A(mai_mai_n1903_), .B(mai_mai_n1391_), .C(mai_mai_n148_), .Y(mai_mai_n1914_));
  OAI210     m1865(.A0(mai_mai_n1914_), .A1(mai_mai_n1276_), .B0(mai_mai_n588_), .Y(mai_mai_n1915_));
  NA3        m1866(.A(mai_mai_n1190_), .B(mai_mai_n901_), .C(x7), .Y(mai_mai_n1916_));
  NA3        m1867(.A(mai_mai_n498_), .B(mai_mai_n78_), .C(mai_mai_n610_), .Y(mai_mai_n1917_));
  NA3        m1868(.A(mai_mai_n1917_), .B(mai_mai_n1916_), .C(mai_mai_n1915_), .Y(mai_mai_n1918_));
  NA2        m1869(.A(mai_mai_n1253_), .B(mai_mai_n449_), .Y(mai_mai_n1919_));
  NA3        m1870(.A(mai_mai_n1919_), .B(mai_mai_n1407_), .C(mai_mai_n416_), .Y(mai_mai_n1920_));
  NO2        m1871(.A(mai_mai_n309_), .B(x4), .Y(mai_mai_n1921_));
  AOI220     m1872(.A0(mai_mai_n1921_), .A1(mai_mai_n1868_), .B0(mai_mai_n1131_), .B1(mai_mai_n678_), .Y(mai_mai_n1922_));
  NA2        m1873(.A(mai_mai_n1922_), .B(mai_mai_n1920_), .Y(mai_mai_n1923_));
  NO2        m1874(.A(mai_mai_n1253_), .B(mai_mai_n1230_), .Y(mai_mai_n1924_));
  NO4        m1875(.A(x6), .B(mai_mai_n56_), .C(x2), .D(x0), .Y(mai_mai_n1925_));
  OAI210     m1876(.A0(mai_mai_n1925_), .A1(mai_mai_n1924_), .B0(mai_mai_n1054_), .Y(mai_mai_n1926_));
  NA2        m1877(.A(mai_mai_n1184_), .B(mai_mai_n108_), .Y(mai_mai_n1927_));
  NA2        m1878(.A(mai_mai_n1092_), .B(mai_mai_n107_), .Y(mai_mai_n1928_));
  OAI210     m1879(.A0(mai_mai_n1928_), .A1(mai_mai_n1927_), .B0(mai_mai_n1926_), .Y(mai_mai_n1929_));
  OAI210     m1880(.A0(mai_mai_n1929_), .A1(mai_mai_n1923_), .B0(x7), .Y(mai_mai_n1930_));
  NO2        m1881(.A(mai_mai_n389_), .B(x7), .Y(mai_mai_n1931_));
  NO3        m1882(.A(mai_mai_n403_), .B(mai_mai_n274_), .C(mai_mai_n124_), .Y(mai_mai_n1932_));
  OAI210     m1883(.A0(mai_mai_n874_), .A1(mai_mai_n262_), .B0(mai_mai_n81_), .Y(mai_mai_n1933_));
  OAI220     m1884(.A0(mai_mai_n1933_), .A1(mai_mai_n1932_), .B0(mai_mai_n1931_), .B1(mai_mai_n111_), .Y(mai_mai_n1934_));
  NA2        m1885(.A(mai_mai_n1796_), .B(mai_mai_n658_), .Y(mai_mai_n1935_));
  NO2        m1886(.A(mai_mai_n1845_), .B(mai_mai_n77_), .Y(mai_mai_n1936_));
  AOI220     m1887(.A0(mai_mai_n1936_), .A1(mai_mai_n1935_), .B0(mai_mai_n480_), .B1(mai_mai_n50_), .Y(mai_mai_n1937_));
  AOI210     m1888(.A0(mai_mai_n1937_), .A1(mai_mai_n1934_), .B0(mai_mai_n59_), .Y(mai_mai_n1938_));
  AOI220     m1889(.A0(mai_mai_n1396_), .A1(mai_mai_n676_), .B0(mai_mai_n415_), .B1(mai_mai_n460_), .Y(mai_mai_n1939_));
  OAI210     m1890(.A0(mai_mai_n1939_), .A1(mai_mai_n145_), .B0(x1), .Y(mai_mai_n1940_));
  NO2        m1891(.A(mai_mai_n1940_), .B(mai_mai_n1938_), .Y(mai_mai_n1941_));
  AOI210     m1892(.A0(mai_mai_n1587_), .A1(mai_mai_n403_), .B0(mai_mai_n668_), .Y(mai_mai_n1942_));
  NO2        m1893(.A(mai_mai_n403_), .B(x5), .Y(mai_mai_n1943_));
  NO2        m1894(.A(mai_mai_n1943_), .B(mai_mai_n230_), .Y(mai_mai_n1944_));
  NO2        m1895(.A(mai_mai_n1944_), .B(mai_mai_n1942_), .Y(mai_mai_n1945_));
  NOi21      m1896(.An(mai_mai_n709_), .B(mai_mai_n1007_), .Y(mai_mai_n1946_));
  NA3        m1897(.A(mai_mai_n1946_), .B(mai_mai_n1092_), .C(mai_mai_n874_), .Y(mai_mai_n1947_));
  OAI210     m1898(.A0(mai_mai_n1363_), .A1(mai_mai_n1679_), .B0(mai_mai_n1947_), .Y(mai_mai_n1948_));
  OAI210     m1899(.A0(mai_mai_n1948_), .A1(mai_mai_n1945_), .B0(mai_mai_n1130_), .Y(mai_mai_n1949_));
  OAI210     m1900(.A0(mai_mai_n449_), .A1(mai_mai_n51_), .B0(mai_mai_n1026_), .Y(mai_mai_n1950_));
  AOI220     m1901(.A0(mai_mai_n1950_), .A1(mai_mai_n464_), .B0(mai_mai_n449_), .B1(mai_mai_n390_), .Y(mai_mai_n1951_));
  NO2        m1902(.A(mai_mai_n1951_), .B(mai_mai_n155_), .Y(mai_mai_n1952_));
  OAI220     m1903(.A0(mai_mai_n689_), .A1(mai_mai_n265_), .B0(mai_mai_n685_), .B1(x6), .Y(mai_mai_n1953_));
  NO2        m1904(.A(mai_mai_n304_), .B(x4), .Y(mai_mai_n1954_));
  AOI220     m1905(.A0(mai_mai_n1954_), .A1(mai_mai_n366_), .B0(mai_mai_n1953_), .B1(x4), .Y(mai_mai_n1955_));
  NO3        m1906(.A(mai_mai_n1955_), .B(mai_mai_n325_), .C(x5), .Y(mai_mai_n1956_));
  NO2        m1907(.A(mai_mai_n709_), .B(mai_mai_n57_), .Y(mai_mai_n1957_));
  OAI210     m1908(.A0(mai_mai_n1957_), .A1(mai_mai_n1910_), .B0(mai_mai_n451_), .Y(mai_mai_n1958_));
  AOI220     m1909(.A0(mai_mai_n666_), .A1(mai_mai_n739_), .B0(mai_mai_n496_), .B1(mai_mai_n240_), .Y(mai_mai_n1959_));
  AOI210     m1910(.A0(mai_mai_n1959_), .A1(mai_mai_n1958_), .B0(mai_mai_n260_), .Y(mai_mai_n1960_));
  NO4        m1911(.A(mai_mai_n1960_), .B(mai_mai_n1956_), .C(x1), .D(mai_mai_n1952_), .Y(mai_mai_n1961_));
  AOI220     m1912(.A0(mai_mai_n1961_), .A1(mai_mai_n1949_), .B0(mai_mai_n1941_), .B1(mai_mai_n1930_), .Y(mai_mai_n1962_));
  AOI210     m1913(.A0(mai_mai_n1918_), .A1(x3), .B0(mai_mai_n1962_), .Y(mai29));
  OAI210     m1914(.A0(mai_mai_n558_), .A1(mai_mai_n266_), .B0(mai_mai_n734_), .Y(mai_mai_n1964_));
  NA2        m1915(.A(mai_mai_n755_), .B(mai_mai_n1054_), .Y(mai_mai_n1965_));
  AO210      m1916(.A0(mai_mai_n1165_), .A1(mai_mai_n1174_), .B0(mai_mai_n1965_), .Y(mai_mai_n1966_));
  AOI210     m1917(.A0(mai_mai_n184_), .A1(mai_mai_n168_), .B0(mai_mai_n709_), .Y(mai_mai_n1967_));
  AOI210     m1918(.A0(mai_mai_n1422_), .A1(mai_mai_n78_), .B0(mai_mai_n1967_), .Y(mai_mai_n1968_));
  NA3        m1919(.A(mai_mai_n1968_), .B(mai_mai_n1966_), .C(mai_mai_n1964_), .Y(mai_mai_n1969_));
  NO3        m1920(.A(mai_mai_n668_), .B(mai_mai_n1148_), .C(mai_mai_n50_), .Y(mai_mai_n1970_));
  NO3        m1921(.A(mai_mai_n1970_), .B(mai_mai_n1252_), .C(mai_mai_n558_), .Y(mai_mai_n1971_));
  NO2        m1922(.A(mai_mai_n447_), .B(mai_mai_n58_), .Y(mai_mai_n1972_));
  AOI220     m1923(.A0(mai_mai_n1972_), .A1(mai_mai_n1211_), .B0(mai_mai_n673_), .B1(mai_mai_n1381_), .Y(mai_mai_n1973_));
  OAI210     m1924(.A0(mai_mai_n1971_), .A1(mai_mai_n544_), .B0(mai_mai_n1973_), .Y(mai_mai_n1974_));
  AOI210     m1925(.A0(mai_mai_n1969_), .A1(x6), .B0(mai_mai_n1974_), .Y(mai_mai_n1975_));
  OAI210     m1926(.A0(x8), .A1(x4), .B0(x5), .Y(mai_mai_n1976_));
  NA2        m1927(.A(mai_mai_n1976_), .B(mai_mai_n112_), .Y(mai_mai_n1977_));
  NA2        m1928(.A(mai_mai_n304_), .B(mai_mai_n148_), .Y(mai_mai_n1978_));
  NA4        m1929(.A(mai_mai_n1978_), .B(mai_mai_n1977_), .C(mai_mai_n667_), .D(mai_mai_n64_), .Y(mai_mai_n1979_));
  AOI210     m1930(.A0(mai_mai_n1321_), .A1(mai_mai_n274_), .B0(mai_mai_n1730_), .Y(mai_mai_n1980_));
  AOI210     m1931(.A0(mai_mai_n1980_), .A1(mai_mai_n1979_), .B0(mai_mai_n894_), .Y(mai_mai_n1981_));
  NA4        m1932(.A(mai_mai_n668_), .B(mai_mai_n309_), .C(mai_mai_n184_), .D(mai_mai_n168_), .Y(mai_mai_n1982_));
  NA3        m1933(.A(mai_mai_n634_), .B(mai_mai_n297_), .C(mai_mai_n806_), .Y(mai_mai_n1983_));
  AOI210     m1934(.A0(mai_mai_n1983_), .A1(mai_mai_n1982_), .B0(mai_mai_n1211_), .Y(mai_mai_n1984_));
  OAI210     m1935(.A0(mai_mai_n901_), .A1(x8), .B0(x7), .Y(mai_mai_n1985_));
  NO2        m1936(.A(mai_mai_n1985_), .B(mai_mai_n129_), .Y(mai_mai_n1986_));
  OA210      m1937(.A0(mai_mai_n874_), .A1(mai_mai_n276_), .B0(mai_mai_n1976_), .Y(mai_mai_n1987_));
  OAI220     m1938(.A0(mai_mai_n1987_), .A1(mai_mai_n590_), .B0(mai_mai_n1510_), .B1(mai_mai_n398_), .Y(mai_mai_n1988_));
  NO4        m1939(.A(mai_mai_n1988_), .B(mai_mai_n1986_), .C(mai_mai_n1984_), .D(mai_mai_n1981_), .Y(mai_mai_n1989_));
  OAI210     m1940(.A0(mai_mai_n1975_), .A1(x2), .B0(mai_mai_n1989_), .Y(mai_mai_n1990_));
  NA3        m1941(.A(x6), .B(mai_mai_n50_), .C(x2), .Y(mai_mai_n1991_));
  OAI210     m1942(.A0(mai_mai_n1230_), .A1(mai_mai_n356_), .B0(mai_mai_n1991_), .Y(mai_mai_n1992_));
  NO3        m1943(.A(mai_mai_n449_), .B(x3), .C(x0), .Y(mai_mai_n1993_));
  AO220      m1944(.A0(mai_mai_n1993_), .A1(x5), .B0(mai_mai_n1925_), .B1(mai_mai_n81_), .Y(mai_mai_n1994_));
  AOI210     m1945(.A0(mai_mai_n1992_), .A1(mai_mai_n346_), .B0(mai_mai_n1994_), .Y(mai_mai_n1995_));
  NO3        m1946(.A(mai_mai_n702_), .B(mai_mai_n367_), .C(mai_mai_n144_), .Y(mai_mai_n1996_));
  AOI210     m1947(.A0(mai_mai_n733_), .A1(mai_mai_n617_), .B0(mai_mai_n1996_), .Y(mai_mai_n1997_));
  OAI210     m1948(.A0(mai_mai_n1995_), .A1(x7), .B0(mai_mai_n1997_), .Y(mai_mai_n1998_));
  AOI210     m1949(.A0(mai_mai_n1102_), .A1(mai_mai_n403_), .B0(mai_mai_n1406_), .Y(mai_mai_n1999_));
  NO2        m1950(.A(mai_mai_n148_), .B(x2), .Y(mai_mai_n2000_));
  OA210      m1951(.A0(mai_mai_n2000_), .A1(mai_mai_n632_), .B0(mai_mai_n668_), .Y(mai_mai_n2001_));
  OAI210     m1952(.A0(mai_mai_n2001_), .A1(mai_mai_n1999_), .B0(mai_mai_n68_), .Y(mai_mai_n2002_));
  NO2        m1953(.A(mai_mai_n200_), .B(mai_mai_n85_), .Y(mai_mai_n2003_));
  OAI210     m1954(.A0(mai_mai_n2003_), .A1(mai_mai_n793_), .B0(mai_mai_n1108_), .Y(mai_mai_n2004_));
  NA3        m1955(.A(mai_mai_n1943_), .B(mai_mai_n233_), .C(mai_mai_n83_), .Y(mai_mai_n2005_));
  NA3        m1956(.A(mai_mai_n2005_), .B(mai_mai_n2004_), .C(mai_mai_n2002_), .Y(mai_mai_n2006_));
  AOI210     m1957(.A0(mai_mai_n1998_), .A1(x8), .B0(mai_mai_n2006_), .Y(mai_mai_n2007_));
  OAI210     m1958(.A0(mai_mai_n447_), .A1(mai_mai_n249_), .B0(mai_mai_n970_), .Y(mai_mai_n2008_));
  OAI210     m1959(.A0(mai_mai_n2008_), .A1(mai_mai_n1131_), .B0(mai_mai_n678_), .Y(mai_mai_n2009_));
  NO3        m1960(.A(mai_mai_n1030_), .B(mai_mai_n357_), .C(mai_mai_n149_), .Y(mai_mai_n2010_));
  NA3        m1961(.A(mai_mai_n2010_), .B(mai_mai_n1301_), .C(mai_mai_n50_), .Y(mai_mai_n2011_));
  NO2        m1962(.A(mai_mai_n137_), .B(mai_mai_n93_), .Y(mai_mai_n2012_));
  AOI220     m1963(.A0(mai_mai_n2012_), .A1(mai_mai_n591_), .B0(mai_mai_n1924_), .B1(mai_mai_n363_), .Y(mai_mai_n2013_));
  NOi31      m1964(.An(mai_mai_n1132_), .B(mai_mai_n1874_), .C(mai_mai_n627_), .Y(mai_mai_n2014_));
  NA2        m1965(.A(mai_mai_n174_), .B(x4), .Y(mai_mai_n2015_));
  NO3        m1966(.A(mai_mai_n1483_), .B(mai_mai_n244_), .C(mai_mai_n71_), .Y(mai_mai_n2016_));
  AOI210     m1967(.A0(mai_mai_n2016_), .A1(mai_mai_n2015_), .B0(mai_mai_n2014_), .Y(mai_mai_n2017_));
  NA4        m1968(.A(mai_mai_n2017_), .B(mai_mai_n2013_), .C(mai_mai_n2011_), .D(mai_mai_n2009_), .Y(mai_mai_n2018_));
  NO4        m1969(.A(mai_mai_n1230_), .B(mai_mai_n172_), .C(mai_mai_n55_), .D(mai_mai_n71_), .Y(mai_mai_n2019_));
  NO4        m1970(.A(mai_mai_n1204_), .B(mai_mai_n504_), .C(mai_mai_n1381_), .D(mai_mai_n108_), .Y(mai_mai_n2020_));
  OAI210     m1971(.A0(mai_mai_n2020_), .A1(mai_mai_n2019_), .B0(mai_mai_n110_), .Y(mai_mai_n2021_));
  AOI210     m1972(.A0(mai_mai_n308_), .A1(x4), .B0(mai_mai_n194_), .Y(mai_mai_n2022_));
  OAI210     m1973(.A0(mai_mai_n2022_), .A1(mai_mai_n1972_), .B0(mai_mai_n728_), .Y(mai_mai_n2023_));
  OR3        m1974(.A(mai_mai_n1751_), .B(mai_mai_n1433_), .C(mai_mai_n1094_), .Y(mai_mai_n2024_));
  NA2        m1975(.A(mai_mai_n1925_), .B(mai_mai_n813_), .Y(mai_mai_n2025_));
  OA220      m1976(.A0(mai_mai_n2025_), .A1(mai_mai_n249_), .B0(mai_mai_n583_), .B1(mai_mai_n1794_), .Y(mai_mai_n2026_));
  NA4        m1977(.A(mai_mai_n2026_), .B(mai_mai_n2024_), .C(mai_mai_n2023_), .D(mai_mai_n2021_), .Y(mai_mai_n2027_));
  AOI210     m1978(.A0(mai_mai_n2018_), .A1(mai_mai_n293_), .B0(mai_mai_n2027_), .Y(mai_mai_n2028_));
  OAI210     m1979(.A0(mai_mai_n2007_), .A1(x1), .B0(mai_mai_n2028_), .Y(mai_mai_n2029_));
  AO210      m1980(.A0(mai_mai_n1990_), .A1(x1), .B0(mai_mai_n2029_), .Y(mai30));
  NO3        m1981(.A(mai_mai_n1778_), .B(mai_mai_n579_), .C(mai_mai_n99_), .Y(mai_mai_n2031_));
  NO3        m1982(.A(mai_mai_n1146_), .B(mai_mai_n140_), .C(mai_mai_n386_), .Y(mai_mai_n2032_));
  AOI210     m1983(.A0(mai_mai_n728_), .A1(mai_mai_n257_), .B0(mai_mai_n2032_), .Y(mai_mai_n2033_));
  AOI210     m1984(.A0(mai_mai_n2033_), .A1(mai_mai_n2031_), .B0(mai_mai_n56_), .Y(mai_mai_n2034_));
  NA2        m1985(.A(mai_mai_n818_), .B(mai_mai_n344_), .Y(mai_mai_n2035_));
  NA2        m1986(.A(mai_mai_n2035_), .B(mai_mai_n1364_), .Y(mai_mai_n2036_));
  OAI210     m1987(.A0(mai_mai_n2036_), .A1(mai_mai_n2034_), .B0(mai_mai_n110_), .Y(mai_mai_n2037_));
  OAI210     m1988(.A0(mai_mai_n1007_), .A1(mai_mai_n573_), .B0(mai_mai_n678_), .Y(mai_mai_n2038_));
  AOI220     m1989(.A0(mai_mai_n452_), .A1(mai_mai_n946_), .B0(mai_mai_n330_), .B1(mai_mai_n460_), .Y(mai_mai_n2039_));
  AOI210     m1990(.A0(mai_mai_n2039_), .A1(mai_mai_n2038_), .B0(mai_mai_n260_), .Y(mai_mai_n2040_));
  NO3        m1991(.A(mai_mai_n282_), .B(mai_mai_n125_), .C(x0), .Y(mai_mai_n2041_));
  AOI210     m1992(.A0(mai_mai_n506_), .A1(x6), .B0(mai_mai_n2041_), .Y(mai_mai_n2042_));
  AOI220     m1993(.A0(mai_mai_n1142_), .A1(mai_mai_n427_), .B0(mai_mai_n766_), .B1(mai_mai_n92_), .Y(mai_mai_n2043_));
  OAI220     m1994(.A0(mai_mai_n2043_), .A1(mai_mai_n249_), .B0(mai_mai_n2042_), .B1(mai_mai_n54_), .Y(mai_mai_n2044_));
  NA3        m1995(.A(mai_mai_n326_), .B(mai_mai_n165_), .C(mai_mai_n71_), .Y(mai_mai_n2045_));
  AO210      m1996(.A0(mai_mai_n572_), .A1(mai_mai_n520_), .B0(x5), .Y(mai_mai_n2046_));
  AOI210     m1997(.A0(mai_mai_n2045_), .A1(mai_mai_n725_), .B0(mai_mai_n2046_), .Y(mai_mai_n2047_));
  AOI210     m1998(.A0(mai_mai_n1608_), .A1(mai_mai_n50_), .B0(mai_mai_n460_), .Y(mai_mai_n2048_));
  NA2        m1999(.A(mai_mai_n199_), .B(x2), .Y(mai_mai_n2049_));
  OA220      m2000(.A0(mai_mai_n2049_), .A1(mai_mai_n2048_), .B0(mai_mai_n277_), .B1(x6), .Y(mai_mai_n2050_));
  OAI210     m2001(.A0(x7), .A1(x6), .B0(x1), .Y(mai_mai_n2051_));
  NA3        m2002(.A(mai_mai_n57_), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n2052_));
  AOI220     m2003(.A0(mai_mai_n2052_), .A1(mai_mai_n1371_), .B0(mai_mai_n2051_), .B1(mai_mai_n1819_), .Y(mai_mai_n2053_));
  NO3        m2004(.A(mai_mai_n1367_), .B(mai_mai_n346_), .C(mai_mai_n1032_), .Y(mai_mai_n2054_));
  NO2        m2005(.A(mai_mai_n518_), .B(mai_mai_n867_), .Y(mai_mai_n2055_));
  NOi21      m2006(.An(mai_mai_n2055_), .B(mai_mai_n852_), .Y(mai_mai_n2056_));
  NO3        m2007(.A(mai_mai_n1301_), .B(mai_mai_n235_), .C(mai_mai_n650_), .Y(mai_mai_n2057_));
  NO4        m2008(.A(mai_mai_n2057_), .B(mai_mai_n2056_), .C(mai_mai_n2054_), .D(mai_mai_n2053_), .Y(mai_mai_n2058_));
  OAI210     m2009(.A0(mai_mai_n2050_), .A1(mai_mai_n762_), .B0(mai_mai_n2058_), .Y(mai_mai_n2059_));
  NO4        m2010(.A(mai_mai_n2059_), .B(mai_mai_n2047_), .C(mai_mai_n2044_), .D(mai_mai_n2040_), .Y(mai_mai_n2060_));
  AOI210     m2011(.A0(mai_mai_n2060_), .A1(mai_mai_n2037_), .B0(x8), .Y(mai_mai_n2061_));
  NO3        m2012(.A(mai_mai_n494_), .B(mai_mai_n790_), .C(mai_mai_n53_), .Y(mai_mai_n2062_));
  OAI220     m2013(.A0(mai_mai_n1794_), .A1(mai_mai_n346_), .B0(mai_mai_n486_), .B1(mai_mai_n587_), .Y(mai_mai_n2063_));
  OAI210     m2014(.A0(mai_mai_n2063_), .A1(mai_mai_n2062_), .B0(x6), .Y(mai_mai_n2064_));
  OAI210     m2015(.A0(mai_mai_n1047_), .A1(mai_mai_n539_), .B0(mai_mai_n818_), .Y(mai_mai_n2065_));
  OAI210     m2016(.A0(mai_mai_n1740_), .A1(mai_mai_n333_), .B0(mai_mai_n128_), .Y(mai_mai_n2066_));
  AOI210     m2017(.A0(mai_mai_n382_), .A1(mai_mai_n232_), .B0(mai_mai_n72_), .Y(mai_mai_n2067_));
  AOI210     m2018(.A0(mai_mai_n1007_), .A1(mai_mai_n753_), .B0(mai_mai_n2067_), .Y(mai_mai_n2068_));
  NA4        m2019(.A(mai_mai_n2068_), .B(mai_mai_n2066_), .C(mai_mai_n2065_), .D(mai_mai_n2064_), .Y(mai_mai_n2069_));
  NA2        m2020(.A(mai_mai_n1099_), .B(mai_mai_n59_), .Y(mai_mai_n2070_));
  AOI210     m2021(.A0(mai_mai_n929_), .A1(mai_mai_n495_), .B0(mai_mai_n684_), .Y(mai_mai_n2071_));
  OAI220     m2022(.A0(mai_mai_n2071_), .A1(mai_mai_n308_), .B0(mai_mai_n2070_), .B1(mai_mai_n485_), .Y(mai_mai_n2072_));
  AOI210     m2023(.A0(mai_mai_n2069_), .A1(x8), .B0(mai_mai_n2072_), .Y(mai_mai_n2073_));
  NO2        m2024(.A(mai_mai_n2073_), .B(mai_mai_n57_), .Y(mai_mai_n2074_));
  NA2        m2025(.A(mai_mai_n438_), .B(mai_mai_n852_), .Y(mai_mai_n2075_));
  NO2        m2026(.A(mai_mai_n928_), .B(mai_mai_n664_), .Y(mai_mai_n2076_));
  AOI210     m2027(.A0(mai_mai_n2076_), .A1(mai_mai_n2075_), .B0(mai_mai_n449_), .Y(mai_mai_n2077_));
  NO3        m2028(.A(mai_mai_n640_), .B(mai_mai_n412_), .C(mai_mai_n1146_), .Y(mai_mai_n2078_));
  NO3        m2029(.A(mai_mai_n2078_), .B(mai_mai_n1256_), .C(mai_mai_n1381_), .Y(mai_mai_n2079_));
  AOI210     m2030(.A0(mai_mai_n305_), .A1(x1), .B0(mai_mai_n149_), .Y(mai_mai_n2080_));
  NO2        m2031(.A(mai_mai_n311_), .B(x5), .Y(mai_mai_n2081_));
  NO2        m2032(.A(mai_mai_n2081_), .B(mai_mai_n860_), .Y(mai_mai_n2082_));
  OAI220     m2033(.A0(mai_mai_n2082_), .A1(mai_mai_n1065_), .B0(mai_mai_n2080_), .B1(mai_mai_n209_), .Y(mai_mai_n2083_));
  NO3        m2034(.A(mai_mai_n2083_), .B(mai_mai_n2079_), .C(mai_mai_n2077_), .Y(mai_mai_n2084_));
  NA2        m2035(.A(mai_mai_n968_), .B(mai_mai_n82_), .Y(mai_mai_n2085_));
  AO210      m2036(.A0(mai_mai_n2085_), .A1(mai_mai_n1609_), .B0(x3), .Y(mai_mai_n2086_));
  NO2        m2037(.A(mai_mai_n221_), .B(mai_mai_n56_), .Y(mai_mai_n2087_));
  NO2        m2038(.A(mai_mai_n357_), .B(mai_mai_n235_), .Y(mai_mai_n2088_));
  AOI220     m2039(.A0(mai_mai_n2088_), .A1(x2), .B0(mai_mai_n2087_), .B1(mai_mai_n1624_), .Y(mai_mai_n2089_));
  AOI210     m2040(.A0(mai_mai_n2089_), .A1(mai_mai_n2086_), .B0(mai_mai_n265_), .Y(mai_mai_n2090_));
  NO2        m2041(.A(mai_mai_n305_), .B(mai_mai_n124_), .Y(mai_mai_n2091_));
  NO3        m2042(.A(mai_mai_n823_), .B(mai_mai_n703_), .C(mai_mai_n168_), .Y(mai_mai_n2092_));
  OAI210     m2043(.A0(mai_mai_n2092_), .A1(mai_mai_n2091_), .B0(mai_mai_n156_), .Y(mai_mai_n2093_));
  NA3        m2044(.A(x5), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n2094_));
  AOI210     m2045(.A0(mai_mai_n2094_), .A1(mai_mai_n1309_), .B0(mai_mai_n540_), .Y(mai_mai_n2095_));
  AOI210     m2046(.A0(mai_mai_n1329_), .A1(x2), .B0(mai_mai_n2095_), .Y(mai_mai_n2096_));
  AOI210     m2047(.A0(mai_mai_n2096_), .A1(mai_mai_n2093_), .B0(mai_mai_n50_), .Y(mai_mai_n2097_));
  NA3        m2048(.A(mai_mai_n1480_), .B(mai_mai_n1140_), .C(mai_mai_n478_), .Y(mai_mai_n2098_));
  AOI210     m2049(.A0(mai_mai_n2098_), .A1(mai_mai_n2085_), .B0(mai_mai_n613_), .Y(mai_mai_n2099_));
  AOI210     m2050(.A0(mai_mai_n1032_), .A1(x1), .B0(mai_mai_n1321_), .Y(mai_mai_n2100_));
  OAI220     m2051(.A0(mai_mai_n309_), .A1(x4), .B0(mai_mai_n51_), .B1(x6), .Y(mai_mai_n2101_));
  NO2        m2052(.A(mai_mai_n123_), .B(mai_mai_n112_), .Y(mai_mai_n2102_));
  AOI220     m2053(.A0(mai_mai_n2102_), .A1(mai_mai_n2101_), .B0(mai_mai_n1167_), .B1(mai_mai_n627_), .Y(mai_mai_n2103_));
  OAI210     m2054(.A0(mai_mai_n2100_), .A1(mai_mai_n489_), .B0(mai_mai_n2103_), .Y(mai_mai_n2104_));
  NO4        m2055(.A(mai_mai_n2104_), .B(mai_mai_n2099_), .C(mai_mai_n2097_), .D(mai_mai_n2090_), .Y(mai_mai_n2105_));
  OAI210     m2056(.A0(mai_mai_n2084_), .A1(mai_mai_n137_), .B0(mai_mai_n2105_), .Y(mai_mai_n2106_));
  NO3        m2057(.A(mai_mai_n2106_), .B(mai_mai_n2074_), .C(mai_mai_n2061_), .Y(mai31));
  NA2        m2058(.A(mai_mai_n992_), .B(mai_mai_n358_), .Y(mai_mai_n2108_));
  NO2        m2059(.A(mai_mai_n453_), .B(mai_mai_n678_), .Y(mai_mai_n2109_));
  AOI210     m2060(.A0(mai_mai_n2109_), .A1(mai_mai_n2108_), .B0(mai_mai_n58_), .Y(mai_mai_n2110_));
  NO2        m2061(.A(mai_mai_n792_), .B(mai_mai_n56_), .Y(mai_mai_n2111_));
  AOI220     m2062(.A0(mai_mai_n2111_), .A1(x2), .B0(mai_mai_n91_), .B1(x0), .Y(mai_mai_n2112_));
  NA3        m2063(.A(mai_mai_n2112_), .B(mai_mai_n2025_), .C(mai_mai_n1854_), .Y(mai_mai_n2113_));
  OAI210     m2064(.A0(mai_mai_n2113_), .A1(mai_mai_n2110_), .B0(mai_mai_n53_), .Y(mai_mai_n2114_));
  NO2        m2065(.A(mai_mai_n435_), .B(mai_mai_n678_), .Y(mai_mai_n2115_));
  NO3        m2066(.A(mai_mai_n1954_), .B(mai_mai_n1925_), .C(mai_mai_n895_), .Y(mai_mai_n2116_));
  OA220      m2067(.A0(mai_mai_n2116_), .A1(mai_mai_n478_), .B0(mai_mai_n2115_), .B1(mai_mai_n1473_), .Y(mai_mai_n2117_));
  AOI210     m2068(.A0(mai_mai_n2117_), .A1(mai_mai_n2114_), .B0(mai_mai_n108_), .Y(mai_mai_n2118_));
  NO2        m2069(.A(mai_mai_n500_), .B(mai_mai_n75_), .Y(mai_mai_n2119_));
  NA2        m2070(.A(mai_mai_n449_), .B(mai_mai_n57_), .Y(mai_mai_n2120_));
  AOI210     m2071(.A0(mai_mai_n308_), .A1(mai_mai_n86_), .B0(mai_mai_n2120_), .Y(mai_mai_n2121_));
  OAI210     m2072(.A0(mai_mai_n2121_), .A1(mai_mai_n2119_), .B0(mai_mai_n777_), .Y(mai_mai_n2122_));
  NO4        m2073(.A(mai_mai_n1163_), .B(mai_mai_n367_), .C(mai_mai_n1608_), .D(mai_mai_n67_), .Y(mai_mai_n2123_));
  AOI210     m2074(.A0(mai_mai_n1647_), .A1(mai_mai_n1356_), .B0(mai_mai_n447_), .Y(mai_mai_n2124_));
  OAI220     m2075(.A0(mai_mai_n1310_), .A1(mai_mai_n960_), .B0(mai_mai_n779_), .B1(mai_mai_n117_), .Y(mai_mai_n2125_));
  NO3        m2076(.A(mai_mai_n2125_), .B(mai_mai_n2124_), .C(mai_mai_n2123_), .Y(mai_mai_n2126_));
  AOI210     m2077(.A0(mai_mai_n2126_), .A1(mai_mai_n2122_), .B0(x5), .Y(mai_mai_n2127_));
  AOI220     m2078(.A0(mai_mai_n451_), .A1(mai_mai_n627_), .B0(mai_mai_n573_), .B1(mai_mai_n63_), .Y(mai_mai_n2128_));
  AOI210     m2079(.A0(mai_mai_n2128_), .A1(mai_mai_n583_), .B0(mai_mai_n1230_), .Y(mai_mai_n2129_));
  AOI220     m2080(.A0(mai_mai_n969_), .A1(mai_mai_n739_), .B0(mai_mai_n1146_), .B1(mai_mai_n122_), .Y(mai_mai_n2130_));
  OAI220     m2081(.A0(mai_mai_n2130_), .A1(mai_mai_n389_), .B0(mai_mai_n485_), .B1(mai_mai_n778_), .Y(mai_mai_n2131_));
  NO4        m2082(.A(mai_mai_n2131_), .B(mai_mai_n2129_), .C(mai_mai_n2127_), .D(mai_mai_n2118_), .Y(mai_mai_n2132_));
  NA2        m2083(.A(mai_mai_n495_), .B(mai_mai_n59_), .Y(mai_mai_n2133_));
  AOI210     m2084(.A0(mai_mai_n544_), .A1(mai_mai_n2133_), .B0(mai_mai_n143_), .Y(mai_mai_n2134_));
  OAI210     m2085(.A0(mai_mai_n104_), .A1(mai_mai_n276_), .B0(mai_mai_n2070_), .Y(mai_mai_n2135_));
  OAI210     m2086(.A0(mai_mai_n2135_), .A1(mai_mai_n2134_), .B0(x7), .Y(mai_mai_n2136_));
  NA2        m2087(.A(mai_mai_n1096_), .B(mai_mai_n92_), .Y(mai_mai_n2137_));
  AOI210     m2088(.A0(mai_mai_n907_), .A1(mai_mai_n112_), .B0(mai_mai_n2137_), .Y(mai_mai_n2138_));
  NA2        m2089(.A(mai_mai_n1555_), .B(x6), .Y(mai_mai_n2139_));
  AOI210     m2090(.A0(mai_mai_n2139_), .A1(mai_mai_n292_), .B0(mai_mai_n108_), .Y(mai_mai_n2140_));
  NA2        m2091(.A(mai_mai_n1190_), .B(mai_mai_n321_), .Y(mai_mai_n2141_));
  AOI210     m2092(.A0(mai_mai_n2141_), .A1(mai_mai_n646_), .B0(mai_mai_n53_), .Y(mai_mai_n2142_));
  NO3        m2093(.A(mai_mai_n2142_), .B(mai_mai_n2140_), .C(mai_mai_n2138_), .Y(mai_mai_n2143_));
  AOI210     m2094(.A0(mai_mai_n2143_), .A1(mai_mai_n2136_), .B0(mai_mai_n688_), .Y(mai_mai_n2144_));
  NOi21      m2095(.An(mai_mai_n1768_), .B(mai_mai_n1069_), .Y(mai_mai_n2145_));
  OAI220     m2096(.A0(mai_mai_n2145_), .A1(mai_mai_n1927_), .B0(mai_mai_n930_), .B1(mai_mai_n2133_), .Y(mai_mai_n2146_));
  NA2        m2097(.A(mai_mai_n2146_), .B(x3), .Y(mai_mai_n2147_));
  AOI220     m2098(.A0(mai_mai_n1391_), .A1(x8), .B0(mai_mai_n60_), .B1(x1), .Y(mai_mai_n2148_));
  NO3        m2099(.A(mai_mai_n2148_), .B(mai_mai_n1120_), .C(x6), .Y(mai_mai_n2149_));
  AOI220     m2100(.A0(mai_mai_n617_), .A1(mai_mai_n412_), .B0(mai_mai_n495_), .B1(mai_mai_n78_), .Y(mai_mai_n2150_));
  NA2        m2101(.A(mai_mai_n118_), .B(mai_mai_n531_), .Y(mai_mai_n2151_));
  OAI220     m2102(.A0(mai_mai_n2151_), .A1(mai_mai_n1927_), .B0(mai_mai_n2150_), .B1(x4), .Y(mai_mai_n2152_));
  NO2        m2103(.A(mai_mai_n2152_), .B(mai_mai_n2149_), .Y(mai_mai_n2153_));
  AOI210     m2104(.A0(mai_mai_n2153_), .A1(mai_mai_n2147_), .B0(mai_mai_n187_), .Y(mai_mai_n2154_));
  NO4        m2105(.A(mai_mai_n618_), .B(mai_mai_n591_), .C(mai_mai_n704_), .D(mai_mai_n703_), .Y(mai_mai_n2155_));
  OAI210     m2106(.A0(mai_mai_n2155_), .A1(mai_mai_n1087_), .B0(x3), .Y(mai_mai_n2156_));
  NO4        m2107(.A(mai_mai_n809_), .B(mai_mai_n1230_), .C(mai_mai_n777_), .D(x5), .Y(mai_mai_n2157_));
  NO3        m2108(.A(x6), .B(mai_mai_n56_), .C(x1), .Y(mai_mai_n2158_));
  NA2        m2109(.A(mai_mai_n2158_), .B(mai_mai_n288_), .Y(mai_mai_n2159_));
  OAI210     m2110(.A0(mai_mai_n1897_), .A1(mai_mai_n382_), .B0(mai_mai_n2159_), .Y(mai_mai_n2160_));
  NA4        m2111(.A(mai_mai_n640_), .B(mai_mai_n180_), .C(x6), .D(mai_mai_n108_), .Y(mai_mai_n2161_));
  NO2        m2112(.A(mai_mai_n861_), .B(mai_mai_n253_), .Y(mai_mai_n2162_));
  NOi41      m2113(.An(mai_mai_n2161_), .B(mai_mai_n2162_), .C(mai_mai_n2160_), .D(mai_mai_n2157_), .Y(mai_mai_n2163_));
  AOI210     m2114(.A0(mai_mai_n2163_), .A1(mai_mai_n2156_), .B0(mai_mai_n535_), .Y(mai_mai_n2164_));
  OAI210     m2115(.A0(mai_mai_n617_), .A1(mai_mai_n472_), .B0(mai_mai_n946_), .Y(mai_mai_n2165_));
  NO3        m2116(.A(mai_mai_n377_), .B(mai_mai_n77_), .C(mai_mai_n53_), .Y(mai_mai_n2166_));
  NO3        m2117(.A(mai_mai_n464_), .B(mai_mai_n352_), .C(mai_mai_n50_), .Y(mai_mai_n2167_));
  OAI210     m2118(.A0(mai_mai_n2167_), .A1(mai_mai_n2166_), .B0(mai_mai_n1164_), .Y(mai_mai_n2168_));
  AOI210     m2119(.A0(mai_mai_n2168_), .A1(mai_mai_n2165_), .B0(mai_mai_n396_), .Y(mai_mai_n2169_));
  NO2        m2120(.A(mai_mai_n218_), .B(mai_mai_n540_), .Y(mai_mai_n2170_));
  OAI210     m2121(.A0(mai_mai_n140_), .A1(x2), .B0(mai_mai_n2170_), .Y(mai_mai_n2171_));
  NO2        m2122(.A(mai_mai_n2171_), .B(mai_mai_n64_), .Y(mai_mai_n2172_));
  NA2        m2123(.A(mai_mai_n123_), .B(mai_mai_n57_), .Y(mai_mai_n2173_));
  AOI220     m2124(.A0(mai_mai_n1587_), .A1(mai_mai_n914_), .B0(mai_mai_n275_), .B1(x4), .Y(mai_mai_n2174_));
  AOI220     m2125(.A0(mai_mai_n1640_), .A1(mai_mai_n619_), .B0(mai_mai_n726_), .B1(mai_mai_n777_), .Y(mai_mai_n2175_));
  OAI220     m2126(.A0(mai_mai_n2175_), .A1(mai_mai_n2173_), .B0(mai_mai_n2174_), .B1(mai_mai_n192_), .Y(mai_mai_n2176_));
  OR3        m2127(.A(mai_mai_n2176_), .B(mai_mai_n2172_), .C(mai_mai_n2169_), .Y(mai_mai_n2177_));
  NO4        m2128(.A(mai_mai_n2177_), .B(mai_mai_n2164_), .C(mai_mai_n2154_), .D(mai_mai_n2144_), .Y(mai_mai_n2178_));
  OAI210     m2129(.A0(mai_mai_n2132_), .A1(x3), .B0(mai_mai_n2178_), .Y(mai32));
  OAI210     m2130(.A0(mai_mai_n566_), .A1(mai_mai_n53_), .B0(mai_mai_n417_), .Y(mai_mai_n2180_));
  NA2        m2131(.A(mai_mai_n515_), .B(x2), .Y(mai_mai_n2181_));
  AOI210     m2132(.A0(mai_mai_n2181_), .A1(mai_mai_n2180_), .B0(mai_mai_n57_), .Y(mai_mai_n2182_));
  OAI210     m2133(.A0(mai_mai_n2182_), .A1(mai_mai_n793_), .B0(mai_mai_n56_), .Y(mai_mai_n2183_));
  OAI210     m2134(.A0(mai_mai_n1710_), .A1(mai_mai_n1452_), .B0(mai_mai_n1482_), .Y(mai_mai_n2184_));
  AOI210     m2135(.A0(mai_mai_n2111_), .A1(mai_mai_n279_), .B0(mai_mai_n2184_), .Y(mai_mai_n2185_));
  AOI210     m2136(.A0(mai_mai_n2185_), .A1(mai_mai_n2183_), .B0(mai_mai_n50_), .Y(mai_mai_n2186_));
  NA3        m2137(.A(mai_mai_n1556_), .B(mai_mai_n807_), .C(mai_mai_n291_), .Y(mai_mai_n2187_));
  NA2        m2138(.A(mai_mai_n750_), .B(mai_mai_n548_), .Y(mai_mai_n2188_));
  OAI220     m2139(.A0(mai_mai_n1064_), .A1(mai_mai_n233_), .B0(mai_mai_n685_), .B1(mai_mai_n209_), .Y(mai_mai_n2189_));
  NO3        m2140(.A(mai_mai_n378_), .B(mai_mai_n576_), .C(mai_mai_n813_), .Y(mai_mai_n2190_));
  NO2        m2141(.A(mai_mai_n1367_), .B(mai_mai_n587_), .Y(mai_mai_n2191_));
  NO4        m2142(.A(mai_mai_n2191_), .B(mai_mai_n2190_), .C(mai_mai_n2189_), .D(mai_mai_n2188_), .Y(mai_mai_n2192_));
  AOI210     m2143(.A0(mai_mai_n2192_), .A1(mai_mai_n2187_), .B0(mai_mai_n144_), .Y(mai_mai_n2193_));
  OAI220     m2144(.A0(mai_mai_n405_), .A1(x7), .B0(mai_mai_n304_), .B1(mai_mai_n297_), .Y(mai_mai_n2194_));
  NA2        m2145(.A(mai_mai_n2194_), .B(mai_mai_n968_), .Y(mai_mai_n2195_));
  NO2        m2146(.A(mai_mai_n553_), .B(mai_mai_n867_), .Y(mai_mai_n2196_));
  AOI220     m2147(.A0(mai_mai_n2196_), .A1(mai_mai_n1877_), .B0(mai_mai_n532_), .B1(mai_mai_n133_), .Y(mai_mai_n2197_));
  AOI210     m2148(.A0(mai_mai_n2197_), .A1(mai_mai_n2195_), .B0(mai_mai_n110_), .Y(mai_mai_n2198_));
  NA3        m2149(.A(mai_mai_n1320_), .B(mai_mai_n1148_), .C(mai_mai_n117_), .Y(mai_mai_n2199_));
  NA2        m2150(.A(mai_mai_n1357_), .B(mai_mai_n704_), .Y(mai_mai_n2200_));
  AOI210     m2151(.A0(mai_mai_n2200_), .A1(mai_mai_n2199_), .B0(mai_mai_n56_), .Y(mai_mai_n2201_));
  NA2        m2152(.A(mai_mai_n968_), .B(mai_mai_n57_), .Y(mai_mai_n2202_));
  NOi21      m2153(.An(mai_mai_n2202_), .B(mai_mai_n133_), .Y(mai_mai_n2203_));
  NA2        m2154(.A(mai_mai_n1022_), .B(mai_mai_n253_), .Y(mai_mai_n2204_));
  NO3        m2155(.A(mai_mai_n2204_), .B(mai_mai_n2203_), .C(mai_mai_n59_), .Y(mai_mai_n2205_));
  OR4        m2156(.A(mai_mai_n2205_), .B(mai_mai_n2201_), .C(mai_mai_n2198_), .D(mai_mai_n2193_), .Y(mai_mai_n2206_));
  OAI210     m2157(.A0(mai_mai_n2206_), .A1(mai_mai_n2186_), .B0(mai_mai_n108_), .Y(mai_mai_n2207_));
  NO3        m2158(.A(mai_mai_n1230_), .B(mai_mai_n146_), .C(mai_mai_n126_), .Y(mai_mai_n2208_));
  NO2        m2159(.A(mai_mai_n384_), .B(mai_mai_n55_), .Y(mai_mai_n2209_));
  NA2        m2160(.A(mai_mai_n2209_), .B(mai_mai_n116_), .Y(mai_mai_n2210_));
  OAI210     m2161(.A0(mai_mai_n636_), .A1(mai_mai_n593_), .B0(mai_mai_n818_), .Y(mai_mai_n2211_));
  NA2        m2162(.A(mai_mai_n2211_), .B(mai_mai_n2210_), .Y(mai_mai_n2212_));
  OAI210     m2163(.A0(mai_mai_n2212_), .A1(mai_mai_n2208_), .B0(x3), .Y(mai_mai_n2213_));
  OAI210     m2164(.A0(mai_mai_n901_), .A1(mai_mai_n274_), .B0(mai_mai_n50_), .Y(mai_mai_n2214_));
  AOI210     m2165(.A0(mai_mai_n62_), .A1(mai_mai_n110_), .B0(mai_mai_n2214_), .Y(mai_mai_n2215_));
  OAI210     m2166(.A0(mai_mai_n2215_), .A1(mai_mai_n1858_), .B0(mai_mai_n703_), .Y(mai_mai_n2216_));
  NO3        m2167(.A(mai_mai_n306_), .B(mai_mai_n174_), .C(mai_mai_n124_), .Y(mai_mai_n2217_));
  NO3        m2168(.A(mai_mai_n807_), .B(mai_mai_n365_), .C(mai_mai_n144_), .Y(mai_mai_n2218_));
  OAI210     m2169(.A0(mai_mai_n2218_), .A1(mai_mai_n2217_), .B0(mai_mai_n59_), .Y(mai_mai_n2219_));
  NA2        m2170(.A(mai_mai_n1152_), .B(mai_mai_n71_), .Y(mai_mai_n2220_));
  NO2        m2171(.A(mai_mai_n1931_), .B(mai_mai_n593_), .Y(mai_mai_n2221_));
  AOI210     m2172(.A0(mai_mai_n2221_), .A1(mai_mai_n1859_), .B0(mai_mai_n2220_), .Y(mai_mai_n2222_));
  NO2        m2173(.A(mai_mai_n276_), .B(mai_mai_n57_), .Y(mai_mai_n2223_));
  NO2        m2174(.A(mai_mai_n2223_), .B(mai_mai_n1014_), .Y(mai_mai_n2224_));
  NOi31      m2175(.An(mai_mai_n728_), .B(mai_mai_n2224_), .C(mai_mai_n282_), .Y(mai_mai_n2225_));
  NO3        m2176(.A(mai_mai_n1312_), .B(mai_mai_n218_), .C(mai_mai_n260_), .Y(mai_mai_n2226_));
  NO4        m2177(.A(mai_mai_n2226_), .B(mai_mai_n2225_), .C(mai_mai_n2222_), .D(x1), .Y(mai_mai_n2227_));
  NA4        m2178(.A(mai_mai_n2227_), .B(mai_mai_n2219_), .C(mai_mai_n2216_), .D(mai_mai_n2213_), .Y(mai_mai_n2228_));
  AO210      m2179(.A0(mai_mai_n1102_), .A1(mai_mai_n400_), .B0(mai_mai_n1017_), .Y(mai_mai_n2229_));
  NA3        m2180(.A(mai_mai_n1903_), .B(mai_mai_n557_), .C(mai_mai_n276_), .Y(mai_mai_n2230_));
  AOI210     m2181(.A0(mai_mai_n2230_), .A1(mai_mai_n2229_), .B0(mai_mai_n306_), .Y(mai_mai_n2231_));
  NA4        m2182(.A(mai_mai_n1265_), .B(mai_mai_n529_), .C(mai_mai_n389_), .D(mai_mai_n233_), .Y(mai_mai_n2232_));
  NO3        m2183(.A(mai_mai_n1433_), .B(mai_mai_n1017_), .C(x2), .Y(mai_mai_n2233_));
  NO2        m2184(.A(mai_mai_n1835_), .B(mai_mai_n64_), .Y(mai_mai_n2234_));
  NO3        m2185(.A(mai_mai_n2234_), .B(mai_mai_n2233_), .C(mai_mai_n53_), .Y(mai_mai_n2235_));
  NO3        m2186(.A(mai_mai_n468_), .B(mai_mai_n1096_), .C(mai_mai_n123_), .Y(mai_mai_n2236_));
  OAI220     m2187(.A0(mai_mai_n688_), .A1(mai_mai_n174_), .B0(mai_mai_n357_), .B1(mai_mai_n144_), .Y(mai_mai_n2237_));
  OAI210     m2188(.A0(mai_mai_n2237_), .A1(mai_mai_n2236_), .B0(mai_mai_n68_), .Y(mai_mai_n2238_));
  NO2        m2189(.A(mai_mai_n1976_), .B(mai_mai_n369_), .Y(mai_mai_n2239_));
  OAI210     m2190(.A0(mai_mai_n1864_), .A1(mai_mai_n611_), .B0(mai_mai_n2239_), .Y(mai_mai_n2240_));
  NA4        m2191(.A(mai_mai_n2240_), .B(mai_mai_n2238_), .C(mai_mai_n2235_), .D(mai_mai_n2232_), .Y(mai_mai_n2241_));
  OAI210     m2192(.A0(mai_mai_n2241_), .A1(mai_mai_n2231_), .B0(mai_mai_n2228_), .Y(mai_mai_n2242_));
  NO3        m2193(.A(mai_mai_n1217_), .B(mai_mai_n107_), .C(mai_mai_n71_), .Y(mai_mai_n2243_));
  NO2        m2194(.A(mai_mai_n566_), .B(mai_mai_n373_), .Y(mai_mai_n2244_));
  OAI210     m2195(.A0(mai_mai_n2243_), .A1(mai_mai_n1412_), .B0(mai_mai_n2244_), .Y(mai_mai_n2245_));
  NO3        m2196(.A(x8), .B(mai_mai_n71_), .C(x2), .Y(mai_mai_n2246_));
  OAI220     m2197(.A0(mai_mai_n2246_), .A1(mai_mai_n627_), .B0(mai_mai_n1422_), .B1(mai_mai_n91_), .Y(mai_mai_n2247_));
  AOI220     m2198(.A0(mai_mai_n558_), .A1(mai_mai_n818_), .B0(mai_mai_n678_), .B1(mai_mai_n258_), .Y(mai_mai_n2248_));
  AOI210     m2199(.A0(mai_mai_n2248_), .A1(mai_mai_n2247_), .B0(mai_mai_n268_), .Y(mai_mai_n2249_));
  NA2        m2200(.A(mai_mai_n1022_), .B(mai_mai_n1146_), .Y(mai_mai_n2250_));
  AOI210     m2201(.A0(mai_mai_n674_), .A1(mai_mai_n688_), .B0(mai_mai_n2250_), .Y(mai_mai_n2251_));
  AOI210     m2202(.A0(mai_mai_n591_), .A1(mai_mai_n627_), .B0(mai_mai_n694_), .Y(mai_mai_n2252_));
  NO2        m2203(.A(mai_mai_n2252_), .B(mai_mai_n1819_), .Y(mai_mai_n2253_));
  NO2        m2204(.A(mai_mai_n454_), .B(mai_mai_n435_), .Y(mai_mai_n2254_));
  NOi31      m2205(.An(mai_mai_n1502_), .B(mai_mai_n2254_), .C(mai_mai_n591_), .Y(mai_mai_n2255_));
  NO4        m2206(.A(mai_mai_n2255_), .B(mai_mai_n2253_), .C(mai_mai_n2251_), .D(mai_mai_n2249_), .Y(mai_mai_n2256_));
  NA4        m2207(.A(mai_mai_n2256_), .B(mai_mai_n2245_), .C(mai_mai_n2242_), .D(mai_mai_n2207_), .Y(mai33));
  OAI210     m2208(.A0(mai_mai_n814_), .A1(x1), .B0(mai_mai_n203_), .Y(mai_mai_n2258_));
  OAI210     m2209(.A0(mai_mai_n2081_), .A1(mai_mai_n179_), .B0(mai_mai_n331_), .Y(mai_mai_n2259_));
  OAI220     m2210(.A0(mai_mai_n1082_), .A1(mai_mai_n813_), .B0(mai_mai_n1674_), .B1(mai_mai_n356_), .Y(mai_mai_n2260_));
  NA3        m2211(.A(mai_mai_n2260_), .B(mai_mai_n2259_), .C(mai_mai_n639_), .Y(mai_mai_n2261_));
  AOI210     m2212(.A0(mai_mai_n2258_), .A1(x5), .B0(mai_mai_n2261_), .Y(mai_mai_n2262_));
  NA2        m2213(.A(mai_mai_n232_), .B(mai_mai_n76_), .Y(mai_mai_n2263_));
  NA4        m2214(.A(mai_mai_n1747_), .B(mai_mai_n567_), .C(mai_mai_n249_), .D(x4), .Y(mai_mai_n2264_));
  AOI210     m2215(.A0(mai_mai_n2264_), .A1(mai_mai_n2263_), .B0(mai_mai_n356_), .Y(mai_mai_n2265_));
  OAI210     m2216(.A0(mai_mai_n438_), .A1(mai_mai_n272_), .B0(mai_mai_n53_), .Y(mai_mai_n2266_));
  AOI210     m2217(.A0(mai_mai_n2266_), .A1(mai_mai_n440_), .B0(mai_mai_n64_), .Y(mai_mai_n2267_));
  NA2        m2218(.A(mai_mai_n1662_), .B(mai_mai_n71_), .Y(mai_mai_n2268_));
  NO3        m2219(.A(mai_mai_n2268_), .B(mai_mai_n2267_), .C(mai_mai_n2265_), .Y(mai_mai_n2269_));
  OAI210     m2220(.A0(mai_mai_n2262_), .A1(x4), .B0(mai_mai_n2269_), .Y(mai_mai_n2270_));
  INV        m2221(.A(mai_mai_n242_), .Y(mai_mai_n2271_));
  NA2        m2222(.A(mai_mai_n187_), .B(x4), .Y(mai_mai_n2272_));
  NA2        m2223(.A(mai_mai_n311_), .B(mai_mai_n288_), .Y(mai_mai_n2273_));
  NO2        m2224(.A(mai_mai_n968_), .B(mai_mai_n230_), .Y(mai_mai_n2274_));
  NA2        m2225(.A(mai_mai_n641_), .B(x7), .Y(mai_mai_n2275_));
  OAI220     m2226(.A0(mai_mai_n2275_), .A1(mai_mai_n2274_), .B0(mai_mai_n2273_), .B1(mai_mai_n2272_), .Y(mai_mai_n2276_));
  AOI210     m2227(.A0(mai_mai_n2271_), .A1(mai_mai_n1030_), .B0(mai_mai_n2276_), .Y(mai_mai_n2277_));
  NA2        m2228(.A(mai_mai_n214_), .B(mai_mai_n959_), .Y(mai_mai_n2278_));
  AOI210     m2229(.A0(mai_mai_n2278_), .A1(mai_mai_n2202_), .B0(mai_mai_n216_), .Y(mai_mai_n2279_));
  OAI210     m2230(.A0(mai_mai_n867_), .A1(mai_mai_n51_), .B0(x6), .Y(mai_mai_n2280_));
  NA3        m2231(.A(mai_mai_n924_), .B(mai_mai_n734_), .C(mai_mai_n55_), .Y(mai_mai_n2281_));
  OAI210     m2232(.A0(mai_mai_n621_), .A1(mai_mai_n506_), .B0(mai_mai_n2281_), .Y(mai_mai_n2282_));
  NO3        m2233(.A(mai_mai_n2282_), .B(mai_mai_n2280_), .C(mai_mai_n2279_), .Y(mai_mai_n2283_));
  OAI210     m2234(.A0(mai_mai_n2277_), .A1(mai_mai_n50_), .B0(mai_mai_n2283_), .Y(mai_mai_n2284_));
  NA3        m2235(.A(mai_mai_n2284_), .B(mai_mai_n2270_), .C(mai_mai_n59_), .Y(mai_mai_n2285_));
  NA2        m2236(.A(mai_mai_n536_), .B(mai_mai_n109_), .Y(mai_mai_n2286_));
  NO3        m2237(.A(mai_mai_n1568_), .B(mai_mai_n377_), .C(x4), .Y(mai_mai_n2287_));
  AOI210     m2238(.A0(mai_mai_n2287_), .A1(mai_mai_n2286_), .B0(mai_mai_n441_), .Y(mai_mai_n2288_));
  NA2        m2239(.A(mai_mai_n816_), .B(mai_mai_n108_), .Y(mai_mai_n2289_));
  NA2        m2240(.A(mai_mai_n2289_), .B(mai_mai_n463_), .Y(mai_mai_n2290_));
  NO2        m2241(.A(mai_mai_n709_), .B(mai_mai_n378_), .Y(mai_mai_n2291_));
  NA2        m2242(.A(mai_mai_n502_), .B(mai_mai_n53_), .Y(mai_mai_n2292_));
  AOI210     m2243(.A0(mai_mai_n2291_), .A1(mai_mai_n2290_), .B0(mai_mai_n2292_), .Y(mai_mai_n2293_));
  OAI210     m2244(.A0(mai_mai_n2288_), .A1(mai_mai_n59_), .B0(mai_mai_n2293_), .Y(mai_mai_n2294_));
  AOI220     m2245(.A0(mai_mai_n688_), .A1(mai_mai_n239_), .B0(mai_mai_n389_), .B1(mai_mai_n233_), .Y(mai_mai_n2295_));
  NA2        m2246(.A(mai_mai_n735_), .B(mai_mai_n980_), .Y(mai_mai_n2296_));
  OAI210     m2247(.A0(mai_mai_n2296_), .A1(mai_mai_n2295_), .B0(mai_mai_n305_), .Y(mai_mai_n2297_));
  AOI210     m2248(.A0(mai_mai_n2111_), .A1(mai_mai_n217_), .B0(mai_mai_n53_), .Y(mai_mai_n2298_));
  NO2        m2249(.A(mai_mai_n144_), .B(mai_mai_n341_), .Y(mai_mai_n2299_));
  AOI220     m2250(.A0(mai_mai_n2299_), .A1(mai_mai_n1000_), .B0(mai_mai_n673_), .B1(mai_mai_n356_), .Y(mai_mai_n2300_));
  NA2        m2251(.A(mai_mai_n449_), .B(mai_mai_n500_), .Y(mai_mai_n2301_));
  NO3        m2252(.A(mai_mai_n2301_), .B(mai_mai_n1036_), .C(mai_mai_n184_), .Y(mai_mai_n2302_));
  AOI210     m2253(.A0(mai_mai_n1795_), .A1(mai_mai_n1190_), .B0(mai_mai_n2302_), .Y(mai_mai_n2303_));
  NA4        m2254(.A(mai_mai_n2303_), .B(mai_mai_n2300_), .C(mai_mai_n2298_), .D(mai_mai_n2297_), .Y(mai_mai_n2304_));
  NA3        m2255(.A(mai_mai_n2304_), .B(mai_mai_n2294_), .C(mai_mai_n57_), .Y(mai_mai_n2305_));
  NAi21      m2256(.An(mai_mai_n1192_), .B(mai_mai_n491_), .Y(mai_mai_n2306_));
  NA4        m2257(.A(mai_mai_n641_), .B(mai_mai_n1301_), .C(mai_mai_n472_), .D(mai_mai_n50_), .Y(mai_mai_n2307_));
  OAI210     m2258(.A0(mai_mai_n2299_), .A1(mai_mai_n2055_), .B0(x2), .Y(mai_mai_n2308_));
  NA4        m2259(.A(mai_mai_n288_), .B(mai_mai_n157_), .C(mai_mai_n277_), .D(mai_mai_n123_), .Y(mai_mai_n2309_));
  NA3        m2260(.A(mai_mai_n2309_), .B(mai_mai_n2308_), .C(mai_mai_n2307_), .Y(mai_mai_n2310_));
  AO220      m2261(.A0(mai_mai_n2310_), .A1(x0), .B0(mai_mai_n2306_), .B1(mai_mai_n141_), .Y(mai_mai_n2311_));
  NA3        m2262(.A(mai_mai_n777_), .B(mai_mai_n356_), .C(mai_mai_n60_), .Y(mai_mai_n2312_));
  NO2        m2263(.A(mai_mai_n2246_), .B(mai_mai_n416_), .Y(mai_mai_n2313_));
  NA2        m2264(.A(mai_mai_n640_), .B(mai_mai_n518_), .Y(mai_mai_n2314_));
  OAI220     m2265(.A0(mai_mai_n2314_), .A1(mai_mai_n2313_), .B0(mai_mai_n2312_), .B1(mai_mai_n71_), .Y(mai_mai_n2315_));
  OAI210     m2266(.A0(mai_mai_n1532_), .A1(mai_mai_n352_), .B0(mai_mai_n111_), .Y(mai_mai_n2316_));
  AOI210     m2267(.A0(mai_mai_n591_), .A1(mai_mai_n468_), .B0(mai_mai_n141_), .Y(mai_mai_n2317_));
  OAI210     m2268(.A0(mai_mai_n2317_), .A1(mai_mai_n389_), .B0(mai_mai_n2316_), .Y(mai_mai_n2318_));
  OAI210     m2269(.A0(mai_mai_n2318_), .A1(mai_mai_n2315_), .B0(mai_mai_n102_), .Y(mai_mai_n2319_));
  NA3        m2270(.A(mai_mai_n1209_), .B(mai_mai_n134_), .C(mai_mai_n384_), .Y(mai_mai_n2320_));
  NA2        m2271(.A(mai_mai_n2320_), .B(mai_mai_n1823_), .Y(mai_mai_n2321_));
  NA2        m2272(.A(mai_mai_n1189_), .B(mai_mai_n712_), .Y(mai_mai_n2322_));
  NA2        m2273(.A(mai_mai_n1357_), .B(mai_mai_n1170_), .Y(mai_mai_n2323_));
  NA4        m2274(.A(mai_mai_n2323_), .B(mai_mai_n2322_), .C(mai_mai_n2321_), .D(mai_mai_n2319_), .Y(mai_mai_n2324_));
  AOI210     m2275(.A0(mai_mai_n2311_), .A1(x7), .B0(mai_mai_n2324_), .Y(mai_mai_n2325_));
  NA3        m2276(.A(mai_mai_n2325_), .B(mai_mai_n2305_), .C(mai_mai_n2285_), .Y(mai34));
  NA2        m2277(.A(mai_mai_n435_), .B(x4), .Y(mai_mai_n2327_));
  NO2        m2278(.A(mai_mai_n1954_), .B(mai_mai_n860_), .Y(mai_mai_n2328_));
  AOI210     m2279(.A0(mai_mai_n2328_), .A1(mai_mai_n2327_), .B0(mai_mai_n322_), .Y(mai_mai_n2329_));
  NA2        m2280(.A(mai_mai_n288_), .B(mai_mai_n124_), .Y(mai_mai_n2330_));
  NO2        m2281(.A(mai_mai_n978_), .B(mai_mai_n2330_), .Y(mai_mai_n2331_));
  AOI210     m2282(.A0(mai_mai_n2035_), .A1(mai_mai_n544_), .B0(mai_mai_n143_), .Y(mai_mai_n2332_));
  NA2        m2283(.A(mai_mai_n1954_), .B(x0), .Y(mai_mai_n2333_));
  OAI210     m2284(.A0(mai_mai_n1830_), .A1(mai_mai_n982_), .B0(mai_mai_n2333_), .Y(mai_mai_n2334_));
  NO4        m2285(.A(mai_mai_n2334_), .B(mai_mai_n2332_), .C(mai_mai_n2331_), .D(mai_mai_n2329_), .Y(mai_mai_n2335_));
  NO2        m2286(.A(mai_mai_n2335_), .B(mai_mai_n478_), .Y(mai_mai_n2336_));
  NA2        m2287(.A(mai_mai_n737_), .B(x8), .Y(mai_mai_n2337_));
  AO210      m2288(.A0(mai_mai_n2337_), .A1(mai_mai_n488_), .B0(mai_mai_n663_), .Y(mai_mai_n2338_));
  NA2        m2289(.A(mai_mai_n673_), .B(mai_mai_n632_), .Y(mai_mai_n2339_));
  AOI210     m2290(.A0(mai_mai_n2339_), .A1(mai_mai_n2338_), .B0(mai_mai_n268_), .Y(mai_mai_n2340_));
  OAI210     m2291(.A0(mai_mai_n123_), .A1(mai_mai_n1056_), .B0(mai_mai_n1467_), .Y(mai_mai_n2341_));
  OAI210     m2292(.A0(mai_mai_n1608_), .A1(mai_mai_n58_), .B0(mai_mai_n2341_), .Y(mai_mai_n2342_));
  NA3        m2293(.A(mai_mai_n2342_), .B(mai_mai_n342_), .C(x8), .Y(mai_mai_n2343_));
  NO3        m2294(.A(mai_mai_n999_), .B(mai_mai_n709_), .C(mai_mai_n459_), .Y(mai_mai_n2344_));
  AOI210     m2295(.A0(mai_mai_n1590_), .A1(mai_mai_n330_), .B0(mai_mai_n2344_), .Y(mai_mai_n2345_));
  NA2        m2296(.A(mai_mai_n667_), .B(mai_mai_n322_), .Y(mai_mai_n2346_));
  NA2        m2297(.A(mai_mai_n137_), .B(x0), .Y(mai_mai_n2347_));
  NAi31      m2298(.An(mai_mai_n2347_), .B(mai_mai_n2346_), .C(mai_mai_n801_), .Y(mai_mai_n2348_));
  NA3        m2299(.A(mai_mai_n1603_), .B(mai_mai_n1399_), .C(mai_mai_n50_), .Y(mai_mai_n2349_));
  NA4        m2300(.A(mai_mai_n2349_), .B(mai_mai_n2348_), .C(mai_mai_n2345_), .D(mai_mai_n2343_), .Y(mai_mai_n2350_));
  NA2        m2301(.A(mai_mai_n1112_), .B(mai_mai_n753_), .Y(mai_mai_n2351_));
  NA3        m2302(.A(mai_mai_n1148_), .B(mai_mai_n168_), .C(mai_mai_n1099_), .Y(mai_mai_n2352_));
  AOI210     m2303(.A0(mai_mai_n2352_), .A1(mai_mai_n2351_), .B0(mai_mai_n763_), .Y(mai_mai_n2353_));
  AOI210     m2304(.A0(mai_mai_n1778_), .A1(mai_mai_n133_), .B0(mai_mai_n2353_), .Y(mai_mai_n2354_));
  AOI210     m2305(.A0(mai_mai_n558_), .A1(mai_mai_n818_), .B0(mai_mai_n257_), .Y(mai_mai_n2355_));
  OAI220     m2306(.A0(mai_mai_n2355_), .A1(mai_mai_n59_), .B0(mai_mai_n1123_), .B1(mai_mai_n55_), .Y(mai_mai_n2356_));
  NA3        m2307(.A(mai_mai_n2356_), .B(mai_mai_n737_), .C(mai_mai_n56_), .Y(mai_mai_n2357_));
  OAI210     m2308(.A0(mai_mai_n2354_), .A1(mai_mai_n144_), .B0(mai_mai_n2357_), .Y(mai_mai_n2358_));
  NO4        m2309(.A(mai_mai_n2358_), .B(mai_mai_n2350_), .C(mai_mai_n2340_), .D(mai_mai_n2336_), .Y(mai_mai_n2359_));
  NO2        m2310(.A(mai_mai_n312_), .B(mai_mai_n959_), .Y(mai_mai_n2360_));
  NO3        m2311(.A(mai_mai_n2360_), .B(mai_mai_n447_), .C(mai_mai_n330_), .Y(mai_mai_n2361_));
  NA2        m2312(.A(mai_mai_n787_), .B(mai_mai_n161_), .Y(mai_mai_n2362_));
  NO3        m2313(.A(mai_mai_n2223_), .B(mai_mai_n305_), .C(mai_mai_n1099_), .Y(mai_mai_n2363_));
  OAI220     m2314(.A0(mai_mai_n2363_), .A1(mai_mai_n1560_), .B0(mai_mai_n2362_), .B1(mai_mai_n1174_), .Y(mai_mai_n2364_));
  OAI210     m2315(.A0(mai_mai_n2364_), .A1(mai_mai_n2361_), .B0(x2), .Y(mai_mai_n2365_));
  OAI210     m2316(.A0(mai_mai_n870_), .A1(mai_mai_n373_), .B0(mai_mai_n2365_), .Y(mai_mai_n2366_));
  NA2        m2317(.A(mai_mai_n315_), .B(x4), .Y(mai_mai_n2367_));
  OAI220     m2318(.A0(mai_mai_n749_), .A1(mai_mai_n55_), .B0(mai_mai_n281_), .B1(mai_mai_n107_), .Y(mai_mai_n2368_));
  NO4        m2319(.A(mai_mai_n451_), .B(mai_mai_n77_), .C(x7), .D(x3), .Y(mai_mai_n2369_));
  NO2        m2320(.A(mai_mai_n1112_), .B(mai_mai_n289_), .Y(mai_mai_n2370_));
  NO4        m2321(.A(mai_mai_n2370_), .B(mai_mai_n2369_), .C(mai_mai_n2368_), .D(mai_mai_n2367_), .Y(mai_mai_n2371_));
  NA2        m2322(.A(mai_mai_n1244_), .B(mai_mai_n1054_), .Y(mai_mai_n2372_));
  NA4        m2323(.A(mai_mai_n737_), .B(mai_mai_n180_), .C(mai_mai_n57_), .D(mai_mai_n108_), .Y(mai_mai_n2373_));
  NA3        m2324(.A(mai_mai_n1396_), .B(mai_mai_n260_), .C(x7), .Y(mai_mai_n2374_));
  NA3        m2325(.A(mai_mai_n2374_), .B(mai_mai_n2373_), .C(mai_mai_n2372_), .Y(mai_mai_n2375_));
  OAI210     m2326(.A0(mai_mai_n2375_), .A1(mai_mai_n2371_), .B0(mai_mai_n165_), .Y(mai_mai_n2376_));
  NA3        m2327(.A(mai_mai_n865_), .B(mai_mai_n87_), .C(x0), .Y(mai_mai_n2377_));
  NA4        m2328(.A(mai_mai_n2377_), .B(mai_mai_n1152_), .C(mai_mai_n298_), .D(mai_mai_n589_), .Y(mai_mai_n2378_));
  NA2        m2329(.A(mai_mai_n1156_), .B(mai_mai_n678_), .Y(mai_mai_n2379_));
  OAI210     m2330(.A0(mai_mai_n2379_), .A1(mai_mai_n269_), .B0(mai_mai_n2161_), .Y(mai_mai_n2380_));
  AOI220     m2331(.A0(mai_mai_n2380_), .A1(x7), .B0(mai_mai_n1021_), .B1(mai_mai_n664_), .Y(mai_mai_n2381_));
  OAI210     m2332(.A0(mai_mai_n2048_), .A1(mai_mai_n265_), .B0(mai_mai_n741_), .Y(mai_mai_n2382_));
  AOI220     m2333(.A0(mai_mai_n412_), .A1(x8), .B0(mai_mai_n92_), .B1(x2), .Y(mai_mai_n2383_));
  AOI210     m2334(.A0(mai_mai_n273_), .A1(mai_mai_n53_), .B0(mai_mai_n655_), .Y(mai_mai_n2384_));
  OAI220     m2335(.A0(mai_mai_n2384_), .A1(mai_mai_n97_), .B0(mai_mai_n2383_), .B1(mai_mai_n1343_), .Y(mai_mai_n2385_));
  AOI220     m2336(.A0(mai_mai_n2385_), .A1(mai_mai_n1321_), .B0(mai_mai_n2382_), .B1(mai_mai_n1517_), .Y(mai_mai_n2386_));
  NA4        m2337(.A(mai_mai_n2386_), .B(mai_mai_n2381_), .C(mai_mai_n2378_), .D(mai_mai_n2376_), .Y(mai_mai_n2387_));
  AOI210     m2338(.A0(mai_mai_n2366_), .A1(mai_mai_n818_), .B0(mai_mai_n2387_), .Y(mai_mai_n2388_));
  OAI210     m2339(.A0(mai_mai_n2359_), .A1(x2), .B0(mai_mai_n2388_), .Y(mai35));
  AOI220     m2340(.A0(mai_mai_n640_), .A1(mai_mai_n55_), .B0(mai_mai_n777_), .B1(mai_mai_n1224_), .Y(mai_mai_n2390_));
  NO2        m2341(.A(mai_mai_n2390_), .B(mai_mai_n71_), .Y(mai_mai_n2391_));
  NO3        m2342(.A(mai_mai_n514_), .B(mai_mai_n468_), .C(mai_mai_n341_), .Y(mai_mai_n2392_));
  OAI210     m2343(.A0(mai_mai_n2392_), .A1(mai_mai_n2391_), .B0(x2), .Y(mai_mai_n2393_));
  AOI210     m2344(.A0(mai_mai_n218_), .A1(x0), .B0(mai_mai_n275_), .Y(mai_mai_n2394_));
  OAI220     m2345(.A0(mai_mai_n2394_), .A1(mai_mai_n669_), .B0(mai_mai_n200_), .B1(x4), .Y(mai_mai_n2395_));
  NA2        m2346(.A(mai_mai_n2395_), .B(mai_mai_n141_), .Y(mai_mai_n2396_));
  NO2        m2347(.A(mai_mai_n1723_), .B(mai_mai_n688_), .Y(mai_mai_n2397_));
  OAI210     m2348(.A0(mai_mai_n2312_), .A1(x6), .B0(mai_mai_n752_), .Y(mai_mai_n2398_));
  NO2        m2349(.A(mai_mai_n2398_), .B(mai_mai_n2397_), .Y(mai_mai_n2399_));
  NA3        m2350(.A(mai_mai_n2399_), .B(mai_mai_n2396_), .C(mai_mai_n2393_), .Y(mai_mai_n2400_));
  NAi21      m2351(.An(mai_mai_n1688_), .B(mai_mai_n1297_), .Y(mai_mai_n2401_));
  NA2        m2352(.A(mai_mai_n216_), .B(mai_mai_n576_), .Y(mai_mai_n2402_));
  NO2        m2353(.A(mai_mai_n435_), .B(mai_mai_n428_), .Y(mai_mai_n2403_));
  AOI220     m2354(.A0(mai_mai_n2403_), .A1(mai_mai_n2402_), .B0(mai_mai_n2401_), .B1(mai_mai_n56_), .Y(mai_mai_n2404_));
  NA2        m2355(.A(mai_mai_n766_), .B(mai_mai_n701_), .Y(mai_mai_n2405_));
  NO3        m2356(.A(mai_mai_n683_), .B(mai_mai_n55_), .C(x6), .Y(mai_mai_n2406_));
  OAI210     m2357(.A0(mai_mai_n2406_), .A1(mai_mai_n712_), .B0(mai_mai_n221_), .Y(mai_mai_n2407_));
  NA2        m2358(.A(mai_mai_n1329_), .B(mai_mai_n63_), .Y(mai_mai_n2408_));
  OAI210     m2359(.A0(mai_mai_n1078_), .A1(x6), .B0(mai_mai_n473_), .Y(mai_mai_n2409_));
  NA3        m2360(.A(mai_mai_n2409_), .B(mai_mai_n2408_), .C(mai_mai_n2407_), .Y(mai_mai_n2410_));
  NA3        m2361(.A(mai_mai_n1273_), .B(mai_mai_n755_), .C(x3), .Y(mai_mai_n2411_));
  NO3        m2362(.A(mai_mai_n2411_), .B(mai_mai_n685_), .C(mai_mai_n209_), .Y(mai_mai_n2412_));
  AOI210     m2363(.A0(mai_mai_n2410_), .A1(mai_mai_n50_), .B0(mai_mai_n2412_), .Y(mai_mai_n2413_));
  OAI210     m2364(.A0(mai_mai_n2405_), .A1(mai_mai_n2404_), .B0(mai_mai_n2413_), .Y(mai_mai_n2414_));
  AOI210     m2365(.A0(mai_mai_n2400_), .A1(mai_mai_n57_), .B0(mai_mai_n2414_), .Y(mai_mai_n2415_));
  NA2        m2366(.A(mai_mai_n968_), .B(mai_mai_n63_), .Y(mai_mai_n2416_));
  NO3        m2367(.A(mai_mai_n1078_), .B(mai_mai_n566_), .C(mai_mai_n124_), .Y(mai_mai_n2417_));
  OAI210     m2368(.A0(mai_mai_n158_), .A1(mai_mai_n67_), .B0(mai_mai_n2417_), .Y(mai_mai_n2418_));
  AOI210     m2369(.A0(mai_mai_n2418_), .A1(mai_mai_n2416_), .B0(mai_mai_n50_), .Y(mai_mai_n2419_));
  NA3        m2370(.A(mai_mai_n468_), .B(mai_mai_n876_), .C(mai_mai_n104_), .Y(mai_mai_n2420_));
  OAI210     m2371(.A0(mai_mai_n968_), .A1(mai_mai_n258_), .B0(mai_mai_n756_), .Y(mai_mai_n2421_));
  OAI210     m2372(.A0(mai_mai_n258_), .A1(mai_mai_n588_), .B0(mai_mai_n2158_), .Y(mai_mai_n2422_));
  NA3        m2373(.A(mai_mai_n2422_), .B(mai_mai_n2421_), .C(mai_mai_n2420_), .Y(mai_mai_n2423_));
  OAI210     m2374(.A0(mai_mai_n2423_), .A1(mai_mai_n2419_), .B0(mai_mai_n59_), .Y(mai_mai_n2424_));
  AOI210     m2375(.A0(mai_mai_n865_), .A1(mai_mai_n535_), .B0(mai_mai_n1903_), .Y(mai_mai_n2425_));
  AOI210     m2376(.A0(mai_mai_n566_), .A1(mai_mai_n610_), .B0(mai_mai_n2425_), .Y(mai_mai_n2426_));
  NO4        m2377(.A(mai_mai_n960_), .B(mai_mai_n566_), .C(mai_mai_n365_), .D(mai_mai_n410_), .Y(mai_mai_n2427_));
  XN2        m2378(.A(x4), .B(x3), .Y(mai_mai_n2428_));
  NO3        m2379(.A(mai_mai_n2428_), .B(mai_mai_n668_), .C(mai_mai_n311_), .Y(mai_mai_n2429_));
  NO3        m2380(.A(mai_mai_n2429_), .B(mai_mai_n2427_), .C(mai_mai_n1463_), .Y(mai_mai_n2430_));
  OAI210     m2381(.A0(mai_mai_n2426_), .A1(x3), .B0(mai_mai_n2430_), .Y(mai_mai_n2431_));
  NO3        m2382(.A(mai_mai_n749_), .B(mai_mai_n867_), .C(mai_mai_n276_), .Y(mai_mai_n2432_));
  OAI210     m2383(.A0(mai_mai_n2432_), .A1(mai_mai_n1463_), .B0(mai_mai_n50_), .Y(mai_mai_n2433_));
  NA3        m2384(.A(mai_mai_n1086_), .B(mai_mai_n816_), .C(mai_mai_n257_), .Y(mai_mai_n2434_));
  NA2        m2385(.A(mai_mai_n2434_), .B(mai_mai_n2433_), .Y(mai_mai_n2435_));
  AOI210     m2386(.A0(mai_mai_n2431_), .A1(mai_mai_n591_), .B0(mai_mai_n2435_), .Y(mai_mai_n2436_));
  AOI210     m2387(.A0(mai_mai_n1433_), .A1(mai_mai_n645_), .B0(mai_mai_n685_), .Y(mai_mai_n2437_));
  NO2        m2388(.A(mai_mai_n876_), .B(mai_mai_n56_), .Y(mai_mai_n2438_));
  OAI210     m2389(.A0(mai_mai_n1957_), .A1(mai_mai_n610_), .B0(mai_mai_n2246_), .Y(mai_mai_n2439_));
  OAI210     m2390(.A0(mai_mai_n2337_), .A1(mai_mai_n2438_), .B0(mai_mai_n2439_), .Y(mai_mai_n2440_));
  OAI210     m2391(.A0(mai_mai_n2440_), .A1(mai_mai_n2437_), .B0(mai_mai_n92_), .Y(mai_mai_n2441_));
  NO2        m2392(.A(mai_mai_n858_), .B(mai_mai_n665_), .Y(mai_mai_n2442_));
  NO2        m2393(.A(mai_mai_n289_), .B(x6), .Y(mai_mai_n2443_));
  OAI210     m2394(.A0(mai_mai_n2442_), .A1(mai_mai_n1786_), .B0(mai_mai_n2443_), .Y(mai_mai_n2444_));
  NA4        m2395(.A(mai_mai_n2444_), .B(mai_mai_n2441_), .C(mai_mai_n2436_), .D(mai_mai_n2424_), .Y(mai_mai_n2445_));
  NA4        m2396(.A(mai_mai_n618_), .B(mai_mai_n688_), .C(mai_mai_n434_), .D(x6), .Y(mai_mai_n2446_));
  AOI210     m2397(.A0(mai_mai_n2446_), .A1(mai_mai_n429_), .B0(x1), .Y(mai_mai_n2447_));
  NO2        m2398(.A(mai_mai_n735_), .B(mai_mai_n685_), .Y(mai_mai_n2448_));
  OAI210     m2399(.A0(mai_mai_n468_), .A1(mai_mai_n169_), .B0(mai_mai_n799_), .Y(mai_mai_n2449_));
  AOI210     m2400(.A0(mai_mai_n2449_), .A1(mai_mai_n1026_), .B0(mai_mai_n53_), .Y(mai_mai_n2450_));
  NO3        m2401(.A(mai_mai_n2450_), .B(mai_mai_n2448_), .C(mai_mai_n2447_), .Y(mai_mai_n2451_));
  NA3        m2402(.A(mai_mai_n1435_), .B(mai_mai_n1274_), .C(mai_mai_n822_), .Y(mai_mai_n2452_));
  AOI220     m2403(.A0(mai_mai_n1946_), .A1(mai_mai_n141_), .B0(mai_mai_n421_), .B1(mai_mai_n128_), .Y(mai_mai_n2453_));
  AOI210     m2404(.A0(mai_mai_n2453_), .A1(mai_mai_n2452_), .B0(mai_mai_n1510_), .Y(mai_mai_n2454_));
  NO2        m2405(.A(mai_mai_n640_), .B(x3), .Y(mai_mai_n2455_));
  NO3        m2406(.A(mai_mai_n696_), .B(mai_mai_n1608_), .C(x2), .Y(mai_mai_n2456_));
  AOI220     m2407(.A0(mai_mai_n2456_), .A1(mai_mai_n2455_), .B0(mai_mai_n1919_), .B1(mai_mai_n773_), .Y(mai_mai_n2457_));
  NA3        m2408(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n2458_));
  OAI220     m2409(.A0(mai_mai_n2458_), .A1(mai_mai_n199_), .B0(mai_mai_n683_), .B1(mai_mai_n531_), .Y(mai_mai_n2459_));
  OAI220     m2410(.A0(mai_mai_n1310_), .A1(x8), .B0(mai_mai_n377_), .B1(mai_mai_n355_), .Y(mai_mai_n2460_));
  AOI220     m2411(.A0(mai_mai_n2460_), .A1(mai_mai_n421_), .B0(mai_mai_n2459_), .B1(mai_mai_n923_), .Y(mai_mai_n2461_));
  OAI210     m2412(.A0(mai_mai_n2457_), .A1(mai_mai_n1165_), .B0(mai_mai_n2461_), .Y(mai_mai_n2462_));
  NO2        m2413(.A(mai_mai_n2462_), .B(mai_mai_n2454_), .Y(mai_mai_n2463_));
  OAI210     m2414(.A0(mai_mai_n2451_), .A1(mai_mai_n315_), .B0(mai_mai_n2463_), .Y(mai_mai_n2464_));
  AOI210     m2415(.A0(mai_mai_n2445_), .A1(x5), .B0(mai_mai_n2464_), .Y(mai_mai_n2465_));
  OAI210     m2416(.A0(mai_mai_n2415_), .A1(x5), .B0(mai_mai_n2465_), .Y(mai36));
  NO2        m2417(.A(mai_mai_n867_), .B(mai_mai_n304_), .Y(mai_mai_n2467_));
  NO3        m2418(.A(mai_mai_n123_), .B(mai_mai_n1056_), .C(mai_mai_n55_), .Y(mai_mai_n2468_));
  NO3        m2419(.A(mai_mai_n2468_), .B(mai_mai_n1976_), .C(mai_mai_n1078_), .Y(mai_mai_n2469_));
  OAI210     m2420(.A0(mai_mai_n2469_), .A1(mai_mai_n2467_), .B0(mai_mai_n110_), .Y(mai_mai_n2470_));
  OR4        m2421(.A(mai_mai_n961_), .B(mai_mai_n809_), .C(mai_mai_n380_), .D(mai_mai_n495_), .Y(mai_mai_n2471_));
  INV        m2422(.A(mai_mai_n1011_), .Y(mai_mai_n2472_));
  OAI210     m2423(.A0(mai_mai_n2209_), .A1(mai_mai_n2472_), .B0(mai_mai_n281_), .Y(mai_mai_n2473_));
  NA3        m2424(.A(mai_mai_n449_), .B(mai_mai_n230_), .C(mai_mai_n122_), .Y(mai_mai_n2474_));
  NA4        m2425(.A(mai_mai_n2474_), .B(mai_mai_n2473_), .C(mai_mai_n2471_), .D(mai_mai_n2470_), .Y(mai_mai_n2475_));
  NO2        m2426(.A(mai_mai_n1000_), .B(x8), .Y(mai_mai_n2476_));
  NO3        m2427(.A(mai_mai_n2476_), .B(mai_mai_n996_), .C(mai_mai_n540_), .Y(mai_mai_n2477_));
  AOI220     m2428(.A0(mai_mai_n305_), .A1(x1), .B0(mai_mai_n140_), .B1(x6), .Y(mai_mai_n2478_));
  AOI210     m2429(.A0(mai_mai_n1099_), .A1(x6), .B0(mai_mai_n425_), .Y(mai_mai_n2479_));
  OAI220     m2430(.A0(mai_mai_n2479_), .A1(mai_mai_n364_), .B0(mai_mai_n2478_), .B1(mai_mai_n469_), .Y(mai_mai_n2480_));
  OAI210     m2431(.A0(mai_mai_n2480_), .A1(mai_mai_n2477_), .B0(mai_mai_n468_), .Y(mai_mai_n2481_));
  NA2        m2432(.A(mai_mai_n673_), .B(mai_mai_n495_), .Y(mai_mai_n2482_));
  AOI210     m2433(.A0(mai_mai_n2482_), .A1(mai_mai_n652_), .B0(mai_mai_n269_), .Y(mai_mai_n2483_));
  NO3        m2434(.A(mai_mai_n1874_), .B(mai_mai_n1607_), .C(mai_mai_n277_), .Y(mai_mai_n2484_));
  NO2        m2435(.A(mai_mai_n2416_), .B(mai_mai_n232_), .Y(mai_mai_n2485_));
  NO4        m2436(.A(mai_mai_n2485_), .B(mai_mai_n2484_), .C(mai_mai_n2483_), .D(mai_mai_n423_), .Y(mai_mai_n2486_));
  OAI210     m2437(.A0(mai_mai_n641_), .A1(mai_mai_n808_), .B0(mai_mai_n986_), .Y(mai_mai_n2487_));
  OAI220     m2438(.A0(mai_mai_n1653_), .A1(mai_mai_n1648_), .B0(mai_mai_n986_), .B1(mai_mai_n1099_), .Y(mai_mai_n2488_));
  AOI220     m2439(.A0(mai_mai_n2488_), .A1(mai_mai_n121_), .B0(mai_mai_n2487_), .B1(mai_mai_n632_), .Y(mai_mai_n2489_));
  NA3        m2440(.A(mai_mai_n2489_), .B(mai_mai_n2486_), .C(mai_mai_n2481_), .Y(mai_mai_n2490_));
  AOI210     m2441(.A0(mai_mai_n2475_), .A1(mai_mai_n342_), .B0(mai_mai_n2490_), .Y(mai_mai_n2491_));
  OAI210     m2442(.A0(mai_mai_n596_), .A1(mai_mai_n519_), .B0(mai_mai_n169_), .Y(mai_mai_n2492_));
  OAI210     m2443(.A0(mai_mai_n1991_), .A1(mai_mai_n70_), .B0(mai_mai_n2492_), .Y(mai_mai_n2493_));
  OAI210     m2444(.A0(mai_mai_n498_), .A1(mai_mai_n241_), .B0(mai_mai_n258_), .Y(mai_mai_n2494_));
  NO2        m2445(.A(mai_mai_n2000_), .B(mai_mai_n176_), .Y(mai_mai_n2495_));
  NA2        m2446(.A(mai_mai_n1211_), .B(mai_mai_n55_), .Y(mai_mai_n2496_));
  OAI210     m2447(.A0(mai_mai_n2496_), .A1(mai_mai_n2495_), .B0(mai_mai_n2494_), .Y(mai_mai_n2497_));
  OAI210     m2448(.A0(mai_mai_n2497_), .A1(mai_mai_n2493_), .B0(mai_mai_n901_), .Y(mai_mai_n2498_));
  AOI210     m2449(.A0(mai_mai_n107_), .A1(mai_mai_n110_), .B0(mai_mai_n344_), .Y(mai_mai_n2499_));
  NA2        m2450(.A(mai_mai_n673_), .B(mai_mai_n1608_), .Y(mai_mai_n2500_));
  OAI220     m2451(.A0(mai_mai_n2500_), .A1(mai_mai_n2499_), .B0(mai_mai_n752_), .B1(mai_mai_n1256_), .Y(mai_mai_n2501_));
  NO2        m2452(.A(mai_mai_n1399_), .B(mai_mai_n582_), .Y(mai_mai_n2502_));
  NO3        m2453(.A(mai_mai_n2502_), .B(mai_mai_n1794_), .C(mai_mai_n696_), .Y(mai_mai_n2503_));
  NO2        m2454(.A(mai_mai_n2503_), .B(mai_mai_n2501_), .Y(mai_mai_n2504_));
  AOI210     m2455(.A0(mai_mai_n2504_), .A1(mai_mai_n2498_), .B0(x7), .Y(mai_mai_n2505_));
  AOI210     m2456(.A0(mai_mai_n591_), .A1(mai_mai_n627_), .B0(mai_mai_n1190_), .Y(mai_mai_n2506_));
  NA3        m2457(.A(mai_mai_n2506_), .B(mai_mai_n999_), .C(mai_mai_n894_), .Y(mai_mai_n2507_));
  NA2        m2458(.A(mai_mai_n2507_), .B(mai_mai_n506_), .Y(mai_mai_n2508_));
  AOI220     m2459(.A0(mai_mai_n1747_), .A1(mai_mai_n261_), .B0(mai_mai_n1054_), .B1(mai_mai_n128_), .Y(mai_mai_n2509_));
  NO2        m2460(.A(mai_mai_n2509_), .B(mai_mai_n449_), .Y(mai_mai_n2510_));
  NO2        m2461(.A(mai_mai_n410_), .B(mai_mai_n230_), .Y(mai_mai_n2511_));
  NO3        m2462(.A(mai_mai_n2511_), .B(mai_mai_n1278_), .C(mai_mai_n59_), .Y(mai_mai_n2512_));
  AOI210     m2463(.A0(mai_mai_n1228_), .A1(mai_mai_n411_), .B0(x6), .Y(mai_mai_n2513_));
  NA3        m2464(.A(mai_mai_n1679_), .B(mai_mai_n281_), .C(mai_mai_n273_), .Y(mai_mai_n2514_));
  NA2        m2465(.A(mai_mai_n2514_), .B(mai_mai_n1634_), .Y(mai_mai_n2515_));
  NO4        m2466(.A(mai_mai_n2515_), .B(mai_mai_n2513_), .C(mai_mai_n2512_), .D(mai_mai_n2510_), .Y(mai_mai_n2516_));
  AOI210     m2467(.A0(mai_mai_n2516_), .A1(mai_mai_n2508_), .B0(mai_mai_n459_), .Y(mai_mai_n2517_));
  NO3        m2468(.A(mai_mai_n2428_), .B(mai_mai_n907_), .C(mai_mai_n505_), .Y(mai_mai_n2518_));
  AOI210     m2469(.A0(mai_mai_n1276_), .A1(mai_mai_n272_), .B0(mai_mai_n2518_), .Y(mai_mai_n2519_));
  OAI210     m2470(.A0(mai_mai_n874_), .A1(mai_mai_n276_), .B0(mai_mai_n400_), .Y(mai_mai_n2520_));
  NA2        m2471(.A(mai_mai_n1211_), .B(mai_mai_n174_), .Y(mai_mai_n2521_));
  NO2        m2472(.A(mai_mai_n617_), .B(mai_mai_n110_), .Y(mai_mai_n2522_));
  AO210      m2473(.A0(mai_mai_n2522_), .A1(mai_mai_n2521_), .B0(mai_mai_n1764_), .Y(mai_mai_n2523_));
  NO2        m2474(.A(mai_mai_n464_), .B(mai_mai_n422_), .Y(mai_mai_n2524_));
  AOI220     m2475(.A0(mai_mai_n2524_), .A1(mai_mai_n2523_), .B0(mai_mai_n2520_), .B1(mai_mai_n296_), .Y(mai_mai_n2525_));
  OAI210     m2476(.A0(mai_mai_n2519_), .A1(x1), .B0(mai_mai_n2525_), .Y(mai_mai_n2526_));
  NO3        m2477(.A(mai_mai_n2526_), .B(mai_mai_n2517_), .C(mai_mai_n2505_), .Y(mai_mai_n2527_));
  OAI210     m2478(.A0(mai_mai_n2491_), .A1(mai_mai_n57_), .B0(mai_mai_n2527_), .Y(mai37));
  NA3        m2479(.A(mai_mai_n1075_), .B(mai_mai_n143_), .C(x3), .Y(mai_mai_n2529_));
  NA3        m2480(.A(mai_mai_n787_), .B(mai_mai_n161_), .C(mai_mai_n50_), .Y(mai_mai_n2530_));
  AOI210     m2481(.A0(mai_mai_n2530_), .A1(mai_mai_n2529_), .B0(mai_mai_n689_), .Y(mai_mai_n2531_));
  NO3        m2482(.A(mai_mai_n1075_), .B(mai_mai_n380_), .C(mai_mai_n513_), .Y(mai_mai_n2532_));
  OAI210     m2483(.A0(mai_mai_n2532_), .A1(mai_mai_n2531_), .B0(mai_mai_n56_), .Y(mai_mai_n2533_));
  NA2        m2484(.A(mai_mai_n605_), .B(mai_mai_n753_), .Y(mai_mai_n2534_));
  AOI210     m2485(.A0(mai_mai_n2534_), .A1(mai_mai_n1055_), .B0(x3), .Y(mai_mai_n2535_));
  AOI220     m2486(.A0(mai_mai_n605_), .A1(mai_mai_n753_), .B0(mai_mai_n468_), .B1(mai_mai_n1054_), .Y(mai_mai_n2536_));
  NO2        m2487(.A(mai_mai_n668_), .B(mai_mai_n183_), .Y(mai_mai_n2537_));
  OAI220     m2488(.A0(mai_mai_n2537_), .A1(mai_mai_n843_), .B0(mai_mai_n2536_), .B1(mai_mai_n110_), .Y(mai_mai_n2538_));
  OAI210     m2489(.A0(mai_mai_n2538_), .A1(mai_mai_n2535_), .B0(mai_mai_n71_), .Y(mai_mai_n2539_));
  NA2        m2490(.A(mai_mai_n1192_), .B(mai_mai_n1078_), .Y(mai_mai_n2540_));
  OAI210     m2491(.A0(mai_mai_n1213_), .A1(mai_mai_n193_), .B0(mai_mai_n460_), .Y(mai_mai_n2541_));
  NA4        m2492(.A(mai_mai_n2541_), .B(mai_mai_n2540_), .C(mai_mai_n2539_), .D(mai_mai_n2533_), .Y(mai_mai_n2542_));
  NA2        m2493(.A(mai_mai_n428_), .B(mai_mai_n140_), .Y(mai_mai_n2543_));
  NO2        m2494(.A(mai_mai_n1710_), .B(mai_mai_n109_), .Y(mai_mai_n2544_));
  AOI210     m2495(.A0(mai_mai_n1978_), .A1(mai_mai_n868_), .B0(mai_mai_n2544_), .Y(mai_mai_n2545_));
  OAI220     m2496(.A0(mai_mai_n2545_), .A1(mai_mai_n51_), .B0(mai_mai_n1609_), .B1(mai_mai_n2543_), .Y(mai_mai_n2546_));
  AOI210     m2497(.A0(mai_mai_n2542_), .A1(mai_mai_n68_), .B0(mai_mai_n2546_), .Y(mai_mai_n2547_));
  OAI210     m2498(.A0(mai_mai_n273_), .A1(mai_mai_n1103_), .B0(mai_mai_n489_), .Y(mai_mai_n2548_));
  NA3        m2499(.A(mai_mai_n2548_), .B(mai_mai_n269_), .C(mai_mai_n1056_), .Y(mai_mai_n2549_));
  OAI210     m2500(.A0(mai_mai_n233_), .A1(mai_mai_n221_), .B0(mai_mai_n1723_), .Y(mai_mai_n2550_));
  NA2        m2501(.A(mai_mai_n350_), .B(mai_mai_n275_), .Y(mai_mai_n2551_));
  NA3        m2502(.A(mai_mai_n406_), .B(mai_mai_n822_), .C(mai_mai_n110_), .Y(mai_mai_n2552_));
  NO2        m2503(.A(mai_mai_n532_), .B(mai_mai_n56_), .Y(mai_mai_n2553_));
  NA3        m2504(.A(mai_mai_n2553_), .B(mai_mai_n2552_), .C(mai_mai_n2551_), .Y(mai_mai_n2554_));
  AOI210     m2505(.A0(mai_mai_n2550_), .A1(mai_mai_n513_), .B0(mai_mai_n2554_), .Y(mai_mai_n2555_));
  NO2        m2506(.A(mai_mai_n1183_), .B(mai_mai_n276_), .Y(mai_mai_n2556_));
  OAI210     m2507(.A0(mai_mai_n296_), .A1(mai_mai_n267_), .B0(mai_mai_n2556_), .Y(mai_mai_n2557_));
  OAI210     m2508(.A0(mai_mai_n670_), .A1(mai_mai_n141_), .B0(x3), .Y(mai_mai_n2558_));
  AOI210     m2509(.A0(mai_mai_n670_), .A1(mai_mai_n369_), .B0(mai_mai_n2558_), .Y(mai_mai_n2559_));
  AOI210     m2510(.A0(mai_mai_n1608_), .A1(mai_mai_n50_), .B0(mai_mai_n350_), .Y(mai_mai_n2560_));
  OAI210     m2511(.A0(mai_mai_n2560_), .A1(mai_mai_n405_), .B0(mai_mai_n56_), .Y(mai_mai_n2561_));
  NO2        m2512(.A(mai_mai_n2561_), .B(mai_mai_n2559_), .Y(mai_mai_n2562_));
  AOI220     m2513(.A0(mai_mai_n2562_), .A1(mai_mai_n2557_), .B0(mai_mai_n2555_), .B1(mai_mai_n2549_), .Y(mai_mai_n2563_));
  OAI210     m2514(.A0(mai_mai_n2563_), .A1(mai_mai_n1762_), .B0(mai_mai_n102_), .Y(mai_mai_n2564_));
  NA2        m2515(.A(mai_mai_n696_), .B(mai_mai_n1197_), .Y(mai_mai_n2565_));
  NOi21      m2516(.An(mai_mai_n1363_), .B(mai_mai_n111_), .Y(mai_mai_n2566_));
  AOI210     m2517(.A0(mai_mai_n2566_), .A1(mai_mai_n2565_), .B0(mai_mai_n438_), .Y(mai_mai_n2567_));
  NO2        m2518(.A(mai_mai_n2220_), .B(mai_mai_n55_), .Y(mai_mai_n2568_));
  OAI210     m2519(.A0(mai_mai_n2568_), .A1(mai_mai_n2567_), .B0(mai_mai_n1823_), .Y(mai_mai_n2569_));
  AOI210     m2520(.A0(mai_mai_n357_), .A1(mai_mai_n143_), .B0(mai_mai_n144_), .Y(mai_mai_n2570_));
  NA2        m2521(.A(mai_mai_n2570_), .B(mai_mai_n350_), .Y(mai_mai_n2571_));
  AOI210     m2522(.A0(mai_mai_n618_), .A1(mai_mai_n438_), .B0(mai_mai_n1286_), .Y(mai_mai_n2572_));
  NO3        m2523(.A(mai_mai_n2572_), .B(mai_mai_n269_), .C(mai_mai_n63_), .Y(mai_mai_n2573_));
  OAI220     m2524(.A0(mai_mai_n2337_), .A1(mai_mai_n486_), .B0(mai_mai_n2094_), .B1(mai_mai_n389_), .Y(mai_mai_n2574_));
  OAI210     m2525(.A0(mai_mai_n2574_), .A1(mai_mai_n2573_), .B0(mai_mai_n53_), .Y(mai_mai_n2575_));
  NO4        m2526(.A(mai_mai_n2347_), .B(mai_mai_n939_), .C(mai_mai_n439_), .D(mai_mai_n224_), .Y(mai_mai_n2576_));
  NO4        m2527(.A(mai_mai_n737_), .B(mai_mai_n606_), .C(mai_mai_n447_), .D(mai_mai_n1064_), .Y(mai_mai_n2577_));
  NO3        m2528(.A(mai_mai_n2577_), .B(mai_mai_n2576_), .C(mai_mai_n1070_), .Y(mai_mai_n2578_));
  NA4        m2529(.A(mai_mai_n2578_), .B(mai_mai_n2575_), .C(mai_mai_n2571_), .D(mai_mai_n2569_), .Y(mai_mai_n2579_));
  NO3        m2530(.A(mai_mai_n253_), .B(mai_mai_n356_), .C(mai_mai_n84_), .Y(mai_mai_n2580_));
  NO2        m2531(.A(mai_mai_n279_), .B(mai_mai_n777_), .Y(mai_mai_n2581_));
  NO3        m2532(.A(mai_mai_n2581_), .B(mai_mai_n1211_), .C(mai_mai_n1230_), .Y(mai_mai_n2582_));
  OAI220     m2533(.A0(mai_mai_n2582_), .A1(mai_mai_n2580_), .B0(mai_mai_n468_), .B1(mai_mai_n85_), .Y(mai_mai_n2583_));
  OR2        m2534(.A(mai_mai_n945_), .B(mai_mai_n755_), .Y(mai_mai_n2584_));
  NA2        m2535(.A(mai_mai_n1224_), .B(mai_mai_n55_), .Y(mai_mai_n2585_));
  NOi21      m2536(.An(mai_mai_n2585_), .B(mai_mai_n390_), .Y(mai_mai_n2586_));
  AOI210     m2537(.A0(mai_mai_n2586_), .A1(mai_mai_n2584_), .B0(x1), .Y(mai_mai_n2587_));
  NA2        m2538(.A(mai_mai_n268_), .B(mai_mai_n84_), .Y(mai_mai_n2588_));
  AOI210     m2539(.A0(mai_mai_n1560_), .A1(mai_mai_n405_), .B0(mai_mai_n2588_), .Y(mai_mai_n2589_));
  NA2        m2540(.A(mai_mai_n1112_), .B(mai_mai_n62_), .Y(mai_mai_n2590_));
  NA2        m2541(.A(mai_mai_n1156_), .B(mai_mai_n176_), .Y(mai_mai_n2591_));
  OAI210     m2542(.A0(mai_mai_n2590_), .A1(mai_mai_n314_), .B0(mai_mai_n2591_), .Y(mai_mai_n2592_));
  NO3        m2543(.A(mai_mai_n2592_), .B(mai_mai_n2589_), .C(mai_mai_n2587_), .Y(mai_mai_n2593_));
  OAI210     m2544(.A0(mai_mai_n2593_), .A1(x6), .B0(mai_mai_n2583_), .Y(mai_mai_n2594_));
  AOI220     m2545(.A0(mai_mai_n2594_), .A1(mai_mai_n1467_), .B0(mai_mai_n2579_), .B1(mai_mai_n57_), .Y(mai_mai_n2595_));
  NA3        m2546(.A(mai_mai_n2595_), .B(mai_mai_n2564_), .C(mai_mai_n2547_), .Y(mai38));
  AOI210     m2547(.A0(mai_mai_n1665_), .A1(mai_mai_n189_), .B0(mai_mai_n980_), .Y(mai_mai_n2597_));
  AOI210     m2548(.A0(mai_mai_n1228_), .A1(mai_mai_n581_), .B0(mai_mai_n1096_), .Y(mai_mai_n2598_));
  AOI210     m2549(.A0(mai_mai_n2585_), .A1(mai_mai_n1851_), .B0(mai_mai_n232_), .Y(mai_mai_n2599_));
  NO3        m2550(.A(mai_mai_n2599_), .B(mai_mai_n2598_), .C(mai_mai_n2597_), .Y(mai_mai_n2600_));
  NO2        m2551(.A(mai_mai_n2600_), .B(x6), .Y(mai_mai_n2601_));
  NA4        m2552(.A(mai_mai_n382_), .B(mai_mai_n260_), .C(mai_mai_n192_), .D(x8), .Y(mai_mai_n2602_));
  NA2        m2553(.A(mai_mai_n404_), .B(mai_mai_n108_), .Y(mai_mai_n2603_));
  AOI210     m2554(.A0(mai_mai_n2603_), .A1(mai_mai_n2602_), .B0(mai_mai_n144_), .Y(mai_mai_n2604_));
  AOI210     m2555(.A0(mai_mai_n439_), .A1(mai_mai_n409_), .B0(mai_mai_n1733_), .Y(mai_mai_n2605_));
  NO2        m2556(.A(mai_mai_n816_), .B(mai_mai_n92_), .Y(mai_mai_n2606_));
  OAI210     m2557(.A0(mai_mai_n1030_), .A1(mai_mai_n149_), .B0(mai_mai_n363_), .Y(mai_mai_n2607_));
  OAI220     m2558(.A0(mai_mai_n2607_), .A1(mai_mai_n2606_), .B0(mai_mai_n2605_), .B1(mai_mai_n192_), .Y(mai_mai_n2608_));
  OAI210     m2559(.A0(mai_mai_n2608_), .A1(mai_mai_n2604_), .B0(x6), .Y(mai_mai_n2609_));
  NO2        m2560(.A(mai_mai_n250_), .B(mai_mai_n777_), .Y(mai_mai_n2610_));
  NO3        m2561(.A(mai_mai_n2610_), .B(mai_mai_n1688_), .C(mai_mai_n260_), .Y(mai_mai_n2611_));
  NO3        m2562(.A(x3), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n2612_));
  OAI210     m2563(.A0(mai_mai_n525_), .A1(x2), .B0(mai_mai_n2612_), .Y(mai_mai_n2613_));
  NA3        m2564(.A(mai_mai_n438_), .B(mai_mai_n428_), .C(mai_mai_n295_), .Y(mai_mai_n2614_));
  NA2        m2565(.A(mai_mai_n2614_), .B(mai_mai_n2613_), .Y(mai_mai_n2615_));
  OAI210     m2566(.A0(mai_mai_n2615_), .A1(mai_mai_n2611_), .B0(mai_mai_n818_), .Y(mai_mai_n2616_));
  NO2        m2567(.A(mai_mai_n606_), .B(mai_mai_n277_), .Y(mai_mai_n2617_));
  AN3        m2568(.A(mai_mai_n823_), .B(mai_mai_n787_), .C(x0), .Y(mai_mai_n2618_));
  OAI210     m2569(.A0(mai_mai_n2618_), .A1(mai_mai_n2617_), .B0(mai_mai_n331_), .Y(mai_mai_n2619_));
  OAI220     m2570(.A0(mai_mai_n606_), .A1(mai_mai_n277_), .B0(mai_mai_n822_), .B1(mai_mai_n93_), .Y(mai_mai_n2620_));
  OAI210     m2571(.A0(mai_mai_n688_), .A1(x0), .B0(mai_mai_n51_), .Y(mai_mai_n2621_));
  AOI210     m2572(.A0(mai_mai_n587_), .A1(x4), .B0(mai_mai_n231_), .Y(mai_mai_n2622_));
  AOI220     m2573(.A0(mai_mai_n2622_), .A1(mai_mai_n2621_), .B0(mai_mai_n2620_), .B1(mai_mai_n406_), .Y(mai_mai_n2623_));
  NA4        m2574(.A(mai_mai_n2623_), .B(mai_mai_n2619_), .C(mai_mai_n2616_), .D(mai_mai_n2609_), .Y(mai_mai_n2624_));
  OAI210     m2575(.A0(mai_mai_n2624_), .A1(mai_mai_n2601_), .B0(x7), .Y(mai_mai_n2625_));
  AOI210     m2576(.A0(mai_mai_n378_), .A1(x1), .B0(mai_mai_n1236_), .Y(mai_mai_n2626_));
  NO2        m2577(.A(mai_mai_n2626_), .B(mai_mai_n51_), .Y(mai_mai_n2627_));
  AOI210     m2578(.A0(mai_mai_n92_), .A1(mai_mai_n71_), .B0(mai_mai_n2246_), .Y(mai_mai_n2628_));
  NA2        m2579(.A(mai_mai_n389_), .B(x3), .Y(mai_mai_n2629_));
  NO2        m2580(.A(mai_mai_n1754_), .B(mai_mai_n532_), .Y(mai_mai_n2630_));
  OAI210     m2581(.A0(mai_mai_n2629_), .A1(mai_mai_n2628_), .B0(mai_mai_n2630_), .Y(mai_mai_n2631_));
  OAI210     m2582(.A0(mai_mai_n2631_), .A1(mai_mai_n2627_), .B0(x4), .Y(mai_mai_n2632_));
  NO2        m2583(.A(mai_mai_n1765_), .B(mai_mai_n462_), .Y(mai_mai_n2633_));
  NO3        m2584(.A(mai_mai_n2633_), .B(mai_mai_n405_), .C(mai_mai_n121_), .Y(mai_mai_n2634_));
  AOI210     m2585(.A0(mai_mai_n1064_), .A1(mai_mai_n244_), .B0(mai_mai_n398_), .Y(mai_mai_n2635_));
  AO210      m2586(.A0(mai_mai_n1302_), .A1(x6), .B0(mai_mai_n2635_), .Y(mai_mai_n2636_));
  NO2        m2587(.A(mai_mai_n1418_), .B(mai_mai_n141_), .Y(mai_mai_n2637_));
  NA2        m2588(.A(mai_mai_n1954_), .B(mai_mai_n325_), .Y(mai_mai_n2638_));
  OAI220     m2589(.A0(mai_mai_n2638_), .A1(mai_mai_n1083_), .B0(mai_mai_n2637_), .B1(mai_mai_n1835_), .Y(mai_mai_n2639_));
  NO3        m2590(.A(mai_mai_n2639_), .B(mai_mai_n2636_), .C(mai_mai_n2634_), .Y(mai_mai_n2640_));
  AOI210     m2591(.A0(mai_mai_n2640_), .A1(mai_mai_n2632_), .B0(mai_mai_n108_), .Y(mai_mai_n2641_));
  NA3        m2592(.A(mai_mai_n1946_), .B(mai_mai_n606_), .C(mai_mai_n165_), .Y(mai_mai_n2642_));
  AOI210     m2593(.A0(mai_mai_n2642_), .A1(mai_mai_n1429_), .B0(mai_mai_n233_), .Y(mai_mai_n2643_));
  AOI210     m2594(.A0(mai_mai_n506_), .A1(mai_mai_n495_), .B0(mai_mai_n684_), .Y(mai_mai_n2644_));
  OAI220     m2595(.A0(mai_mai_n2644_), .A1(mai_mai_n469_), .B0(mai_mai_n200_), .B1(mai_mai_n119_), .Y(mai_mai_n2645_));
  OAI210     m2596(.A0(mai_mai_n2645_), .A1(mai_mai_n2643_), .B0(x0), .Y(mai_mai_n2646_));
  NA3        m2597(.A(mai_mai_n409_), .B(mai_mai_n822_), .C(mai_mai_n277_), .Y(mai_mai_n2647_));
  AOI210     m2598(.A0(mai_mai_n2647_), .A1(mai_mai_n720_), .B0(mai_mai_n2204_), .Y(mai_mai_n2648_));
  NA2        m2599(.A(mai_mai_n1132_), .B(mai_mai_n959_), .Y(mai_mai_n2649_));
  NA4        m2600(.A(mai_mai_n683_), .B(mai_mai_n606_), .C(mai_mai_n180_), .D(x3), .Y(mai_mai_n2650_));
  AOI210     m2601(.A0(mai_mai_n2650_), .A1(mai_mai_n2649_), .B0(mai_mai_n500_), .Y(mai_mai_n2651_));
  NO4        m2602(.A(mai_mai_n1411_), .B(mai_mai_n521_), .C(mai_mai_n1230_), .D(mai_mai_n777_), .Y(mai_mai_n2652_));
  NO2        m2603(.A(mai_mai_n1784_), .B(mai_mai_n2289_), .Y(mai_mai_n2653_));
  NO4        m2604(.A(mai_mai_n2653_), .B(mai_mai_n2652_), .C(mai_mai_n2651_), .D(mai_mai_n2648_), .Y(mai_mai_n2654_));
  NA2        m2605(.A(mai_mai_n2654_), .B(mai_mai_n2646_), .Y(mai_mai_n2655_));
  OAI210     m2606(.A0(mai_mai_n2655_), .A1(mai_mai_n2641_), .B0(mai_mai_n57_), .Y(mai_mai_n2656_));
  AOI210     m2607(.A0(mai_mai_n1824_), .A1(mai_mai_n277_), .B0(mai_mai_n685_), .Y(mai_mai_n2657_));
  OAI210     m2608(.A0(mai_mai_n1761_), .A1(mai_mai_n216_), .B0(mai_mai_n497_), .Y(mai_mai_n2658_));
  OAI210     m2609(.A0(mai_mai_n2658_), .A1(mai_mai_n2657_), .B0(mai_mai_n634_), .Y(mai_mai_n2659_));
  NO2        m2610(.A(mai_mai_n1768_), .B(mai_mai_n277_), .Y(mai_mai_n2660_));
  NA2        m2611(.A(mai_mai_n1868_), .B(mai_mai_n358_), .Y(mai_mai_n2661_));
  OAI220     m2612(.A0(mai_mai_n2661_), .A1(mai_mai_n641_), .B0(mai_mai_n695_), .B1(mai_mai_n151_), .Y(mai_mai_n2662_));
  AOI210     m2613(.A0(mai_mai_n2660_), .A1(mai_mai_n1000_), .B0(mai_mai_n2662_), .Y(mai_mai_n2663_));
  NA4        m2614(.A(mai_mai_n2663_), .B(mai_mai_n2659_), .C(mai_mai_n2656_), .D(mai_mai_n2625_), .Y(mai39));
  INV        m2615(.A(mai_mai_n1608_), .Y(mai_mai_n2667_));
  INV        u0000(.A(x3), .Y(men_men_n50_));
  NA2        u0001(.A(men_men_n50_), .B(x2), .Y(men_men_n51_));
  NA2        u0002(.A(x7), .B(x0), .Y(men_men_n52_));
  INV        u0003(.A(x1), .Y(men_men_n53_));
  NA2        u0004(.A(x5), .B(men_men_n53_), .Y(men_men_n54_));
  INV        u0005(.A(x8), .Y(men_men_n55_));
  INV        u0006(.A(x4), .Y(men_men_n56_));
  INV        u0007(.A(x7), .Y(men_men_n57_));
  NA2        u0008(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0009(.A(x0), .Y(men_men_n59_));
  NA2        u0010(.A(x4), .B(men_men_n59_), .Y(men_men_n60_));
  NA4        u0011(.A(men_men_n60_), .B(men_men_n58_), .C(men_men_n55_), .D(x6), .Y(men_men_n61_));
  NA2        u0012(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n62_));
  NO2        u0013(.A(men_men_n55_), .B(x6), .Y(men_men_n63_));
  NA2        u0014(.A(men_men_n57_), .B(x4), .Y(men_men_n64_));
  NA3        u0015(.A(men_men_n64_), .B(men_men_n63_), .C(men_men_n62_), .Y(men_men_n65_));
  AOI210     u0016(.A0(men_men_n65_), .A1(men_men_n61_), .B0(men_men_n54_), .Y(men_men_n66_));
  NO2        u0017(.A(x8), .B(men_men_n57_), .Y(men_men_n67_));
  NO2        u0018(.A(x7), .B(men_men_n59_), .Y(men_men_n68_));
  NO2        u0019(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi21      u0020(.An(x5), .B(x1), .Y(men_men_n70_));
  INV        u0021(.A(x6), .Y(men_men_n71_));
  NA2        u0022(.A(men_men_n71_), .B(x4), .Y(men_men_n72_));
  NO3        u0023(.A(men_men_n72_), .B(men_men_n70_), .C(men_men_n69_), .Y(men_men_n73_));
  OAI210     u0024(.A0(men_men_n73_), .A1(men_men_n66_), .B0(men_men_n52_), .Y(men_men_n74_));
  NA2        u0025(.A(x7), .B(x4), .Y(men_men_n75_));
  NO2        u0026(.A(men_men_n75_), .B(x1), .Y(men_men_n76_));
  NO2        u0027(.A(men_men_n71_), .B(x5), .Y(men_men_n77_));
  NO2        u0028(.A(x8), .B(men_men_n59_), .Y(men_men_n78_));
  NA3        u0029(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n76_), .Y(men_men_n79_));
  AOI210     u0030(.A0(men_men_n79_), .A1(men_men_n74_), .B0(men_men_n51_), .Y(men_men_n80_));
  NA2        u0031(.A(x5), .B(x3), .Y(men_men_n81_));
  NO2        u0032(.A(x6), .B(x0), .Y(men_men_n82_));
  NO2        u0033(.A(men_men_n82_), .B(x4), .Y(men_men_n83_));
  NO2        u0034(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u0035(.A(men_men_n71_), .B(men_men_n59_), .Y(men_men_n85_));
  NO2        u0036(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n86_));
  NA2        u0037(.A(x8), .B(x1), .Y(men_men_n87_));
  NO2        u0038(.A(men_men_n87_), .B(x7), .Y(men_men_n88_));
  INV        u0039(.A(men_men_n88_), .Y(men_men_n89_));
  OR3        u0040(.A(men_men_n89_), .B(men_men_n86_), .C(men_men_n83_), .Y(men_men_n90_));
  NO3        u0041(.A(x8), .B(men_men_n57_), .C(x6), .Y(men_men_n91_));
  NO2        u0042(.A(x1), .B(men_men_n59_), .Y(men_men_n92_));
  NO2        u0043(.A(men_men_n56_), .B(x2), .Y(men_men_n93_));
  NA3        u0044(.A(men_men_n93_), .B(men_men_n92_), .C(men_men_n91_), .Y(men_men_n94_));
  AOI210     u0045(.A0(men_men_n94_), .A1(men_men_n90_), .B0(men_men_n81_), .Y(men_men_n95_));
  XO2        u0046(.A(x7), .B(x1), .Y(men_men_n96_));
  INV        u0047(.A(men_men_n96_), .Y(men_men_n97_));
  NO2        u0048(.A(men_men_n97_), .B(x6), .Y(men_men_n98_));
  NO2        u0049(.A(men_men_n50_), .B(x0), .Y(men_men_n99_));
  NA2        u0050(.A(men_men_n99_), .B(men_men_n55_), .Y(men_men_n100_));
  NO2        u0051(.A(x6), .B(x5), .Y(men_men_n101_));
  NO2        u0052(.A(men_men_n57_), .B(x5), .Y(men_men_n102_));
  NO2        u0053(.A(men_men_n102_), .B(men_men_n101_), .Y(men_men_n103_));
  NA2        u0054(.A(x6), .B(x1), .Y(men_men_n104_));
  NA2        u0055(.A(men_men_n104_), .B(men_men_n84_), .Y(men_men_n105_));
  NO4        u0056(.A(men_men_n105_), .B(men_men_n103_), .C(men_men_n100_), .D(men_men_n98_), .Y(men_men_n106_));
  NA2        u0057(.A(x3), .B(x0), .Y(men_men_n107_));
  INV        u0058(.A(x5), .Y(men_men_n108_));
  NA2        u0059(.A(men_men_n71_), .B(men_men_n108_), .Y(men_men_n109_));
  INV        u0060(.A(x2), .Y(men_men_n110_));
  NO2        u0061(.A(men_men_n56_), .B(men_men_n110_), .Y(men_men_n111_));
  NA2        u0062(.A(men_men_n57_), .B(men_men_n108_), .Y(men_men_n112_));
  NA3        u0063(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n109_), .Y(men_men_n113_));
  NO3        u0064(.A(men_men_n113_), .B(men_men_n107_), .C(men_men_n53_), .Y(men_men_n114_));
  NO4        u0065(.A(men_men_n114_), .B(men_men_n106_), .C(men_men_n95_), .D(men_men_n80_), .Y(men00));
  NO2        u0066(.A(x7), .B(x6), .Y(men_men_n116_));
  INV        u0067(.A(men_men_n116_), .Y(men_men_n117_));
  NO2        u0068(.A(men_men_n55_), .B(men_men_n53_), .Y(men_men_n118_));
  NA2        u0069(.A(men_men_n118_), .B(men_men_n56_), .Y(men_men_n119_));
  XN2        u0070(.A(x6), .B(x1), .Y(men_men_n120_));
  INV        u0071(.A(men_men_n120_), .Y(men_men_n121_));
  NO2        u0072(.A(x6), .B(x4), .Y(men_men_n122_));
  NA2        u0073(.A(x6), .B(x4), .Y(men_men_n123_));
  NAi21      u0074(.An(men_men_n122_), .B(men_men_n123_), .Y(men_men_n124_));
  XN2        u0075(.A(x7), .B(x6), .Y(men_men_n125_));
  NO2        u0076(.A(x3), .B(men_men_n110_), .Y(men_men_n126_));
  NA2        u0077(.A(men_men_n126_), .B(men_men_n108_), .Y(men_men_n127_));
  NA2        u0078(.A(x3), .B(men_men_n110_), .Y(men_men_n128_));
  NO2        u0079(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n129_));
  NA2        u0080(.A(men_men_n129_), .B(men_men_n56_), .Y(men_men_n130_));
  NA2        u0081(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n131_));
  NA2        u0082(.A(men_men_n131_), .B(x2), .Y(men_men_n132_));
  NA2        u0083(.A(x8), .B(x3), .Y(men_men_n133_));
  NA2        u0084(.A(men_men_n133_), .B(men_men_n75_), .Y(men_men_n134_));
  OAI220     u0085(.A0(men_men_n134_), .A1(men_men_n132_), .B0(men_men_n130_), .B1(men_men_n128_), .Y(men_men_n135_));
  NO2        u0086(.A(x5), .B(x0), .Y(men_men_n136_));
  NO2        u0087(.A(x6), .B(x1), .Y(men_men_n137_));
  NA3        u0088(.A(men_men_n137_), .B(men_men_n136_), .C(men_men_n135_), .Y(men_men_n138_));
  NA2        u0089(.A(x8), .B(men_men_n108_), .Y(men_men_n139_));
  NA2        u0090(.A(x4), .B(men_men_n50_), .Y(men_men_n140_));
  NO3        u0091(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n104_), .Y(men_men_n141_));
  NAi21      u0092(.An(x7), .B(x2), .Y(men_men_n142_));
  NO2        u0093(.A(men_men_n142_), .B(x0), .Y(men_men_n143_));
  XO2        u0094(.A(x8), .B(x7), .Y(men_men_n144_));
  NA2        u0095(.A(men_men_n144_), .B(men_men_n110_), .Y(men_men_n145_));
  NA2        u0096(.A(x6), .B(x5), .Y(men_men_n146_));
  NO2        u0097(.A(men_men_n56_), .B(x0), .Y(men_men_n147_));
  NO2        u0098(.A(men_men_n50_), .B(x1), .Y(men_men_n148_));
  NA2        u0099(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n149_));
  NO3        u0100(.A(men_men_n149_), .B(men_men_n146_), .C(men_men_n145_), .Y(men_men_n150_));
  AOI210     u0101(.A0(men_men_n143_), .A1(men_men_n141_), .B0(men_men_n150_), .Y(men_men_n151_));
  NA2        u0102(.A(men_men_n151_), .B(men_men_n138_), .Y(men01));
  NA2        u0103(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n153_));
  NO2        u0104(.A(x2), .B(x1), .Y(men_men_n154_));
  NA2        u0105(.A(x2), .B(x1), .Y(men_men_n155_));
  NOi21      u0106(.An(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  NA2        u0107(.A(men_men_n108_), .B(men_men_n53_), .Y(men_men_n157_));
  NO2        u0108(.A(men_men_n157_), .B(x8), .Y(men_men_n158_));
  NAi21      u0109(.An(x8), .B(x1), .Y(men_men_n159_));
  NO2        u0110(.A(men_men_n159_), .B(x3), .Y(men_men_n160_));
  OAI210     u0111(.A0(men_men_n160_), .A1(men_men_n158_), .B0(men_men_n156_), .Y(men_men_n161_));
  NO2        u0112(.A(x5), .B(men_men_n50_), .Y(men_men_n162_));
  NO2        u0113(.A(men_men_n110_), .B(x1), .Y(men_men_n163_));
  NA2        u0114(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  AOI210     u0115(.A0(men_men_n164_), .A1(men_men_n161_), .B0(men_men_n153_), .Y(men_men_n165_));
  NAi21      u0116(.An(x7), .B(x0), .Y(men_men_n166_));
  NO2        u0117(.A(men_men_n55_), .B(x2), .Y(men_men_n167_));
  NO2        u0118(.A(men_men_n81_), .B(x1), .Y(men_men_n168_));
  NA2        u0119(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NA2        u0120(.A(x5), .B(men_men_n50_), .Y(men_men_n170_));
  NO2        u0121(.A(men_men_n170_), .B(men_men_n159_), .Y(men_men_n171_));
  NA2        u0122(.A(x8), .B(x5), .Y(men_men_n172_));
  NO2        u0123(.A(men_men_n172_), .B(men_men_n51_), .Y(men_men_n173_));
  NO3        u0124(.A(x3), .B(men_men_n110_), .C(men_men_n53_), .Y(men_men_n174_));
  NO3        u0125(.A(men_men_n174_), .B(men_men_n173_), .C(men_men_n171_), .Y(men_men_n175_));
  AOI210     u0126(.A0(men_men_n175_), .A1(men_men_n169_), .B0(men_men_n166_), .Y(men_men_n176_));
  NO2        u0127(.A(men_men_n57_), .B(x3), .Y(men_men_n177_));
  NO2        u0128(.A(men_men_n55_), .B(x0), .Y(men_men_n178_));
  NA3        u0129(.A(men_men_n108_), .B(men_men_n110_), .C(x1), .Y(men_men_n179_));
  NO2        u0130(.A(men_men_n179_), .B(men_men_n178_), .Y(men_men_n180_));
  NO2        u0131(.A(men_men_n87_), .B(men_men_n50_), .Y(men_men_n181_));
  NA2        u0132(.A(men_men_n108_), .B(x0), .Y(men_men_n182_));
  NO2        u0133(.A(men_men_n182_), .B(x2), .Y(men_men_n183_));
  AOI220     u0134(.A0(men_men_n183_), .A1(men_men_n181_), .B0(men_men_n180_), .B1(men_men_n177_), .Y(men_men_n184_));
  NA2        u0135(.A(x7), .B(men_men_n110_), .Y(men_men_n185_));
  NA2        u0136(.A(men_men_n162_), .B(x8), .Y(men_men_n186_));
  NA4        u0137(.A(x5), .B(x3), .C(x1), .D(x0), .Y(men_men_n187_));
  AO210      u0138(.A0(men_men_n187_), .A1(men_men_n186_), .B0(men_men_n185_), .Y(men_men_n188_));
  NO2        u0139(.A(men_men_n155_), .B(men_men_n50_), .Y(men_men_n189_));
  NAi21      u0140(.An(x1), .B(x2), .Y(men_men_n190_));
  NO2        u0141(.A(men_men_n170_), .B(men_men_n190_), .Y(men_men_n191_));
  NA2        u0142(.A(x8), .B(x7), .Y(men_men_n192_));
  NO2        u0143(.A(men_men_n192_), .B(x0), .Y(men_men_n193_));
  OAI210     u0144(.A0(men_men_n191_), .A1(men_men_n189_), .B0(men_men_n193_), .Y(men_men_n194_));
  NA3        u0145(.A(men_men_n194_), .B(men_men_n188_), .C(men_men_n184_), .Y(men_men_n195_));
  NO3        u0146(.A(men_men_n195_), .B(men_men_n176_), .C(men_men_n165_), .Y(men_men_n196_));
  NA2        u0147(.A(x3), .B(x1), .Y(men_men_n197_));
  NA2        u0148(.A(men_men_n50_), .B(men_men_n110_), .Y(men_men_n198_));
  NO2        u0149(.A(men_men_n198_), .B(men_men_n70_), .Y(men_men_n199_));
  OAI210     u0150(.A0(men_men_n199_), .A1(men_men_n191_), .B0(men_men_n67_), .Y(men_men_n200_));
  NA2        u0151(.A(men_men_n129_), .B(men_men_n110_), .Y(men_men_n201_));
  OAI210     u0152(.A0(men_men_n201_), .A1(men_men_n197_), .B0(men_men_n200_), .Y(men_men_n202_));
  XO2        u0153(.A(x5), .B(x3), .Y(men_men_n203_));
  NA2        u0154(.A(men_men_n203_), .B(x8), .Y(men_men_n204_));
  NA2        u0155(.A(x8), .B(men_men_n59_), .Y(men_men_n205_));
  NA2        u0156(.A(men_men_n205_), .B(men_men_n133_), .Y(men_men_n206_));
  NA2        u0157(.A(x7), .B(men_men_n71_), .Y(men_men_n207_));
  NO2        u0158(.A(men_men_n190_), .B(men_men_n207_), .Y(men_men_n208_));
  OA210      u0159(.A0(men_men_n206_), .A1(men_men_n203_), .B0(men_men_n208_), .Y(men_men_n209_));
  AOI220     u0160(.A0(men_men_n209_), .A1(men_men_n204_), .B0(men_men_n202_), .B1(x0), .Y(men_men_n210_));
  OAI210     u0161(.A0(men_men_n196_), .A1(men_men_n71_), .B0(men_men_n210_), .Y(men_men_n211_));
  NO2        u0162(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n212_));
  NA4        u0163(.A(men_men_n55_), .B(x5), .C(x3), .D(x2), .Y(men_men_n213_));
  NA2        u0164(.A(x8), .B(men_men_n50_), .Y(men_men_n214_));
  NA2        u0165(.A(men_men_n214_), .B(x2), .Y(men_men_n215_));
  NA2        u0166(.A(men_men_n55_), .B(x3), .Y(men_men_n216_));
  NA3        u0167(.A(men_men_n215_), .B(men_men_n203_), .C(men_men_n82_), .Y(men_men_n217_));
  AOI210     u0168(.A0(men_men_n217_), .A1(men_men_n213_), .B0(men_men_n53_), .Y(men_men_n218_));
  NO2        u0169(.A(men_men_n110_), .B(men_men_n59_), .Y(men_men_n219_));
  NA2        u0170(.A(x5), .B(x1), .Y(men_men_n220_));
  NO2        u0171(.A(men_men_n220_), .B(x6), .Y(men_men_n221_));
  NO2        u0172(.A(x3), .B(x1), .Y(men_men_n222_));
  AOI210     u0173(.A0(men_men_n222_), .A1(men_men_n77_), .B0(men_men_n221_), .Y(men_men_n223_));
  NO2        u0174(.A(men_men_n81_), .B(men_men_n55_), .Y(men_men_n224_));
  NO2        u0175(.A(men_men_n104_), .B(men_men_n50_), .Y(men_men_n225_));
  NO2        u0176(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  OAI210     u0177(.A0(men_men_n223_), .A1(x8), .B0(men_men_n226_), .Y(men_men_n227_));
  NO2        u0178(.A(men_men_n55_), .B(x5), .Y(men_men_n228_));
  NA2        u0179(.A(men_men_n228_), .B(men_men_n71_), .Y(men_men_n229_));
  NAi21      u0180(.An(x2), .B(x5), .Y(men_men_n230_));
  NA2        u0181(.A(x8), .B(x6), .Y(men_men_n231_));
  OAI210     u0182(.A0(men_men_n231_), .A1(men_men_n230_), .B0(men_men_n229_), .Y(men_men_n232_));
  NA2        u0183(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n233_));
  NO2        u0184(.A(men_men_n233_), .B(men_men_n59_), .Y(men_men_n234_));
  AO220      u0185(.A0(men_men_n234_), .A1(men_men_n232_), .B0(men_men_n227_), .B1(men_men_n219_), .Y(men_men_n235_));
  OAI210     u0186(.A0(men_men_n235_), .A1(men_men_n218_), .B0(men_men_n212_), .Y(men_men_n236_));
  NA2        u0187(.A(men_men_n71_), .B(men_men_n56_), .Y(men_men_n237_));
  NO2        u0188(.A(men_men_n237_), .B(x7), .Y(men_men_n238_));
  NO2        u0189(.A(men_men_n108_), .B(men_men_n53_), .Y(men_men_n239_));
  NA2        u0190(.A(men_men_n239_), .B(men_men_n110_), .Y(men_men_n240_));
  AOI210     u0191(.A0(men_men_n240_), .A1(men_men_n164_), .B0(men_men_n59_), .Y(men_men_n241_));
  NA2        u0192(.A(x3), .B(men_men_n59_), .Y(men_men_n242_));
  NO2        u0193(.A(men_men_n179_), .B(men_men_n242_), .Y(men_men_n243_));
  OA210      u0194(.A0(men_men_n243_), .A1(men_men_n241_), .B0(x8), .Y(men_men_n244_));
  NO2        u0195(.A(x1), .B(x0), .Y(men_men_n245_));
  NA2        u0196(.A(men_men_n245_), .B(men_men_n110_), .Y(men_men_n246_));
  NA2        u0197(.A(men_men_n108_), .B(men_men_n50_), .Y(men_men_n247_));
  XN2        u0198(.A(x3), .B(x2), .Y(men_men_n248_));
  NA2        u0199(.A(men_men_n248_), .B(men_men_n156_), .Y(men_men_n249_));
  NO2        u0200(.A(men_men_n108_), .B(x0), .Y(men_men_n250_));
  NA2        u0201(.A(x8), .B(men_men_n53_), .Y(men_men_n251_));
  NA2        u0202(.A(men_men_n251_), .B(men_men_n250_), .Y(men_men_n252_));
  OAI220     u0203(.A0(men_men_n252_), .A1(men_men_n249_), .B0(men_men_n247_), .B1(men_men_n246_), .Y(men_men_n253_));
  OAI210     u0204(.A0(men_men_n253_), .A1(men_men_n244_), .B0(men_men_n238_), .Y(men_men_n254_));
  NO2        u0205(.A(x7), .B(x1), .Y(men_men_n255_));
  NOi21      u0206(.An(x8), .B(x3), .Y(men_men_n256_));
  NA2        u0207(.A(men_men_n256_), .B(men_men_n59_), .Y(men_men_n257_));
  NA2        u0208(.A(x5), .B(x0), .Y(men_men_n258_));
  NAi21      u0209(.An(men_men_n136_), .B(men_men_n258_), .Y(men_men_n259_));
  NA2        u0210(.A(men_men_n71_), .B(men_men_n50_), .Y(men_men_n260_));
  OAI210     u0211(.A0(men_men_n260_), .A1(men_men_n259_), .B0(men_men_n257_), .Y(men_men_n261_));
  NA3        u0212(.A(men_men_n261_), .B(men_men_n139_), .C(men_men_n255_), .Y(men_men_n262_));
  NA2        u0213(.A(x8), .B(men_men_n57_), .Y(men_men_n263_));
  NO2        u0214(.A(men_men_n263_), .B(x5), .Y(men_men_n264_));
  NO2        u0215(.A(men_men_n148_), .B(men_men_n71_), .Y(men_men_n265_));
  NA2        u0216(.A(x1), .B(x0), .Y(men_men_n266_));
  NA2        u0217(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n267_));
  NA4        u0218(.A(men_men_n267_), .B(men_men_n266_), .C(men_men_n265_), .D(men_men_n264_), .Y(men_men_n268_));
  NA3        u0219(.A(men_men_n268_), .B(men_men_n262_), .C(men_men_n187_), .Y(men_men_n269_));
  NO2        u0220(.A(men_men_n108_), .B(x3), .Y(men_men_n270_));
  NO2        u0221(.A(men_men_n110_), .B(x0), .Y(men_men_n271_));
  NA2        u0222(.A(men_men_n271_), .B(men_men_n270_), .Y(men_men_n272_));
  NO2        u0223(.A(men_men_n55_), .B(x7), .Y(men_men_n273_));
  NA2        u0224(.A(men_men_n273_), .B(men_men_n137_), .Y(men_men_n274_));
  NO3        u0225(.A(x8), .B(men_men_n50_), .C(x0), .Y(men_men_n275_));
  NAi21      u0226(.An(x8), .B(x0), .Y(men_men_n276_));
  NAi21      u0227(.An(x1), .B(x3), .Y(men_men_n277_));
  NO2        u0228(.A(men_men_n277_), .B(men_men_n276_), .Y(men_men_n278_));
  NO2        u0229(.A(x2), .B(men_men_n53_), .Y(men_men_n279_));
  AOI210     u0230(.A0(men_men_n279_), .A1(men_men_n275_), .B0(men_men_n278_), .Y(men_men_n280_));
  NOi21      u0231(.An(x5), .B(x6), .Y(men_men_n281_));
  NO2        u0232(.A(men_men_n57_), .B(x4), .Y(men_men_n282_));
  NA2        u0233(.A(men_men_n282_), .B(men_men_n281_), .Y(men_men_n283_));
  OAI220     u0234(.A0(men_men_n283_), .A1(men_men_n280_), .B0(men_men_n274_), .B1(men_men_n272_), .Y(men_men_n284_));
  AOI210     u0235(.A0(men_men_n269_), .A1(men_men_n111_), .B0(men_men_n284_), .Y(men_men_n285_));
  NA3        u0236(.A(men_men_n285_), .B(men_men_n254_), .C(men_men_n236_), .Y(men_men_n286_));
  AOI210     u0237(.A0(men_men_n211_), .A1(men_men_n56_), .B0(men_men_n286_), .Y(men02));
  NO2        u0238(.A(x8), .B(men_men_n108_), .Y(men_men_n288_));
  XN2        u0239(.A(x7), .B(x3), .Y(men_men_n289_));
  INV        u0240(.A(men_men_n289_), .Y(men_men_n290_));
  NO2        u0241(.A(x2), .B(x0), .Y(men_men_n291_));
  NA2        u0242(.A(men_men_n291_), .B(men_men_n71_), .Y(men_men_n292_));
  NO2        u0243(.A(men_men_n57_), .B(x1), .Y(men_men_n293_));
  NO3        u0244(.A(men_men_n293_), .B(men_men_n292_), .C(men_men_n290_), .Y(men_men_n294_));
  NA2        u0245(.A(men_men_n53_), .B(x0), .Y(men_men_n295_));
  NO2        u0246(.A(men_men_n277_), .B(x6), .Y(men_men_n296_));
  XO2        u0247(.A(x7), .B(x0), .Y(men_men_n297_));
  NO2        u0248(.A(men_men_n297_), .B(men_men_n291_), .Y(men_men_n298_));
  NA2        u0249(.A(men_men_n298_), .B(men_men_n296_), .Y(men_men_n299_));
  AN2        u0250(.A(x7), .B(x2), .Y(men_men_n300_));
  NA2        u0251(.A(men_men_n300_), .B(men_men_n50_), .Y(men_men_n301_));
  OAI210     u0252(.A0(men_men_n301_), .A1(men_men_n295_), .B0(men_men_n299_), .Y(men_men_n302_));
  OAI210     u0253(.A0(men_men_n302_), .A1(men_men_n294_), .B0(men_men_n288_), .Y(men_men_n303_));
  NAi21      u0254(.An(x8), .B(x6), .Y(men_men_n304_));
  NO2        u0255(.A(men_men_n108_), .B(men_men_n59_), .Y(men_men_n305_));
  NA2        u0256(.A(x7), .B(x3), .Y(men_men_n306_));
  NO2        u0257(.A(men_men_n306_), .B(x2), .Y(men_men_n307_));
  NA2        u0258(.A(x2), .B(x0), .Y(men_men_n308_));
  NA2        u0259(.A(men_men_n110_), .B(men_men_n59_), .Y(men_men_n309_));
  NA2        u0260(.A(men_men_n309_), .B(men_men_n308_), .Y(men_men_n310_));
  NAi21      u0261(.An(x7), .B(x1), .Y(men_men_n311_));
  NO2        u0262(.A(men_men_n311_), .B(x3), .Y(men_men_n312_));
  AOI220     u0263(.A0(men_men_n312_), .A1(men_men_n310_), .B0(men_men_n307_), .B1(men_men_n305_), .Y(men_men_n313_));
  NA2        u0264(.A(men_men_n279_), .B(men_men_n50_), .Y(men_men_n314_));
  NA3        u0265(.A(x7), .B(men_men_n108_), .C(x0), .Y(men_men_n315_));
  NA2        u0266(.A(men_men_n271_), .B(men_men_n53_), .Y(men_men_n316_));
  NA2        u0267(.A(men_men_n162_), .B(men_men_n57_), .Y(men_men_n317_));
  OA220      u0268(.A0(men_men_n317_), .A1(men_men_n316_), .B0(men_men_n315_), .B1(men_men_n314_), .Y(men_men_n318_));
  AOI210     u0269(.A0(men_men_n318_), .A1(men_men_n313_), .B0(men_men_n304_), .Y(men_men_n319_));
  INV        u0270(.A(men_men_n297_), .Y(men_men_n320_));
  NO2        u0271(.A(x7), .B(men_men_n71_), .Y(men_men_n321_));
  NA2        u0272(.A(men_men_n108_), .B(x3), .Y(men_men_n322_));
  NO2        u0273(.A(men_men_n322_), .B(men_men_n321_), .Y(men_men_n323_));
  NA2        u0274(.A(men_men_n323_), .B(men_men_n320_), .Y(men_men_n324_));
  NA2        u0275(.A(men_men_n50_), .B(x0), .Y(men_men_n325_));
  NO2        u0276(.A(men_men_n325_), .B(x7), .Y(men_men_n326_));
  NA2        u0277(.A(men_men_n167_), .B(x1), .Y(men_men_n327_));
  NO2        u0278(.A(men_men_n324_), .B(men_men_n327_), .Y(men_men_n328_));
  NO2        u0279(.A(men_men_n57_), .B(men_men_n50_), .Y(men_men_n329_));
  NO2        u0280(.A(men_men_n55_), .B(men_men_n110_), .Y(men_men_n330_));
  NA3        u0281(.A(men_men_n330_), .B(men_men_n329_), .C(men_men_n59_), .Y(men_men_n331_));
  NO2        u0282(.A(men_men_n157_), .B(x6), .Y(men_men_n332_));
  NO2        u0283(.A(men_men_n104_), .B(men_men_n108_), .Y(men_men_n333_));
  NA2        u0284(.A(men_men_n57_), .B(men_men_n110_), .Y(men_men_n334_));
  NO2        u0285(.A(men_men_n334_), .B(men_men_n267_), .Y(men_men_n335_));
  OAI210     u0286(.A0(men_men_n333_), .A1(men_men_n332_), .B0(men_men_n335_), .Y(men_men_n336_));
  OAI210     u0287(.A0(men_men_n331_), .A1(men_men_n104_), .B0(men_men_n336_), .Y(men_men_n337_));
  NO3        u0288(.A(men_men_n337_), .B(men_men_n328_), .C(men_men_n319_), .Y(men_men_n338_));
  AOI210     u0289(.A0(men_men_n338_), .A1(men_men_n303_), .B0(x4), .Y(men_men_n339_));
  NA2        u0290(.A(x8), .B(men_men_n71_), .Y(men_men_n340_));
  NO2        u0291(.A(x3), .B(men_men_n59_), .Y(men_men_n341_));
  NA3        u0292(.A(men_men_n341_), .B(men_men_n108_), .C(men_men_n53_), .Y(men_men_n342_));
  NO2        u0293(.A(x3), .B(x0), .Y(men_men_n343_));
  NAi21      u0294(.An(men_men_n343_), .B(men_men_n107_), .Y(men_men_n344_));
  NA2        u0295(.A(x5), .B(x2), .Y(men_men_n345_));
  NO2        u0296(.A(men_men_n345_), .B(men_men_n222_), .Y(men_men_n346_));
  AOI210     u0297(.A0(men_men_n346_), .A1(men_men_n344_), .B0(men_men_n243_), .Y(men_men_n347_));
  AO210      u0298(.A0(men_men_n347_), .A1(men_men_n342_), .B0(men_men_n340_), .Y(men_men_n348_));
  NO2        u0299(.A(men_men_n110_), .B(men_men_n53_), .Y(men_men_n349_));
  NA2        u0300(.A(men_men_n349_), .B(x3), .Y(men_men_n350_));
  NO2        u0301(.A(men_men_n55_), .B(x1), .Y(men_men_n351_));
  NA2        u0302(.A(men_men_n351_), .B(men_men_n110_), .Y(men_men_n352_));
  OAI210     u0303(.A0(men_men_n352_), .A1(men_men_n170_), .B0(men_men_n350_), .Y(men_men_n353_));
  NAi32      u0304(.An(x3), .Bn(x0), .C(x2), .Y(men_men_n354_));
  NO2        u0305(.A(men_men_n50_), .B(x2), .Y(men_men_n355_));
  NAi21      u0306(.An(x6), .B(x5), .Y(men_men_n356_));
  NO2        u0307(.A(x2), .B(men_men_n59_), .Y(men_men_n357_));
  NO4        u0308(.A(men_men_n357_), .B(men_men_n356_), .C(men_men_n159_), .D(men_men_n355_), .Y(men_men_n358_));
  AOI220     u0309(.A0(men_men_n358_), .A1(men_men_n354_), .B0(men_men_n353_), .B1(men_men_n85_), .Y(men_men_n359_));
  AOI210     u0310(.A0(men_men_n359_), .A1(men_men_n348_), .B0(men_men_n75_), .Y(men_men_n360_));
  NA2        u0311(.A(men_men_n351_), .B(men_men_n56_), .Y(men_men_n361_));
  NO2        u0312(.A(men_men_n108_), .B(men_men_n50_), .Y(men_men_n362_));
  NO2        u0313(.A(men_men_n291_), .B(men_men_n219_), .Y(men_men_n363_));
  XO2        u0314(.A(x7), .B(x2), .Y(men_men_n364_));
  INV        u0315(.A(men_men_n364_), .Y(men_men_n365_));
  XO2        u0316(.A(x6), .B(x2), .Y(men_men_n366_));
  NA4        u0317(.A(men_men_n366_), .B(men_men_n365_), .C(men_men_n363_), .D(men_men_n362_), .Y(men_men_n367_));
  NAi21      u0318(.An(x0), .B(x6), .Y(men_men_n368_));
  AOI210     u0319(.A0(men_men_n368_), .A1(men_men_n142_), .B0(men_men_n271_), .Y(men_men_n369_));
  XN2        u0320(.A(x7), .B(x5), .Y(men_men_n370_));
  NA2        u0321(.A(men_men_n370_), .B(men_men_n71_), .Y(men_men_n371_));
  NA2        u0322(.A(x7), .B(x5), .Y(men_men_n372_));
  AOI210     u0323(.A0(men_men_n372_), .A1(x6), .B0(men_men_n354_), .Y(men_men_n373_));
  AOI220     u0324(.A0(men_men_n373_), .A1(men_men_n371_), .B0(men_men_n369_), .B1(men_men_n323_), .Y(men_men_n374_));
  AOI210     u0325(.A0(men_men_n374_), .A1(men_men_n367_), .B0(men_men_n361_), .Y(men_men_n375_));
  NO2        u0326(.A(x8), .B(x6), .Y(men_men_n376_));
  NAi21      u0327(.An(men_men_n376_), .B(men_men_n231_), .Y(men_men_n377_));
  AOI210     u0328(.A0(men_men_n377_), .A1(men_men_n92_), .B0(x3), .Y(men_men_n378_));
  NA2        u0329(.A(men_men_n108_), .B(x2), .Y(men_men_n379_));
  NO2        u0330(.A(men_men_n379_), .B(men_men_n64_), .Y(men_men_n380_));
  NA2        u0331(.A(x1), .B(men_men_n59_), .Y(men_men_n381_));
  NO2        u0332(.A(men_men_n381_), .B(men_men_n231_), .Y(men_men_n382_));
  OAI210     u0333(.A0(men_men_n382_), .A1(men_men_n50_), .B0(men_men_n380_), .Y(men_men_n383_));
  NA2        u0334(.A(x4), .B(x2), .Y(men_men_n384_));
  NO2        u0335(.A(men_men_n384_), .B(men_men_n108_), .Y(men_men_n385_));
  NAi21      u0336(.An(x1), .B(x6), .Y(men_men_n386_));
  NA2        u0337(.A(men_men_n343_), .B(men_men_n273_), .Y(men_men_n387_));
  OAI220     u0338(.A0(men_men_n387_), .A1(men_men_n386_), .B0(men_men_n107_), .B1(men_men_n53_), .Y(men_men_n388_));
  NA2        u0339(.A(x8), .B(x2), .Y(men_men_n389_));
  NO2        u0340(.A(men_men_n389_), .B(men_men_n50_), .Y(men_men_n390_));
  INV        u0341(.A(men_men_n221_), .Y(men_men_n391_));
  NA2        u0342(.A(men_men_n388_), .B(men_men_n385_), .Y(men_men_n392_));
  OAI210     u0343(.A0(men_men_n383_), .A1(men_men_n378_), .B0(men_men_n392_), .Y(men_men_n393_));
  NO4        u0344(.A(men_men_n393_), .B(men_men_n375_), .C(men_men_n360_), .D(men_men_n339_), .Y(men03));
  NAi21      u0345(.An(x2), .B(x0), .Y(men_men_n395_));
  NO3        u0346(.A(x8), .B(x6), .C(x4), .Y(men_men_n396_));
  INV        u0347(.A(men_men_n396_), .Y(men_men_n397_));
  NO2        u0348(.A(men_men_n397_), .B(men_men_n395_), .Y(men_men_n398_));
  NA2        u0349(.A(men_men_n111_), .B(men_men_n59_), .Y(men_men_n399_));
  NO2        u0350(.A(men_men_n399_), .B(men_men_n55_), .Y(men_men_n400_));
  OAI210     u0351(.A0(men_men_n400_), .A1(men_men_n398_), .B0(men_men_n162_), .Y(men_men_n401_));
  NA2        u0352(.A(x3), .B(x2), .Y(men_men_n402_));
  NO2        u0353(.A(men_men_n159_), .B(x0), .Y(men_men_n403_));
  NA2        u0354(.A(x8), .B(x0), .Y(men_men_n404_));
  NO2        u0355(.A(men_men_n404_), .B(x6), .Y(men_men_n405_));
  AOI210     u0356(.A0(men_men_n405_), .A1(x5), .B0(men_men_n403_), .Y(men_men_n406_));
  NO2        u0357(.A(men_men_n406_), .B(men_men_n402_), .Y(men_men_n407_));
  NO2        u0358(.A(x5), .B(men_men_n59_), .Y(men_men_n408_));
  NO2        u0359(.A(x3), .B(x2), .Y(men_men_n409_));
  NA2        u0360(.A(men_men_n409_), .B(men_men_n408_), .Y(men_men_n410_));
  NO2        u0361(.A(men_men_n53_), .B(x0), .Y(men_men_n411_));
  NA2        u0362(.A(men_men_n411_), .B(x5), .Y(men_men_n412_));
  AOI210     u0363(.A0(men_men_n412_), .A1(men_men_n410_), .B0(men_men_n304_), .Y(men_men_n413_));
  NA2        u0364(.A(men_men_n257_), .B(men_men_n172_), .Y(men_men_n414_));
  NO2        u0365(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n415_));
  NO2        u0366(.A(men_men_n71_), .B(x0), .Y(men_men_n416_));
  NO4        u0367(.A(men_men_n416_), .B(men_men_n415_), .C(x2), .D(men_men_n53_), .Y(men_men_n417_));
  AO210      u0368(.A0(men_men_n417_), .A1(men_men_n414_), .B0(men_men_n413_), .Y(men_men_n418_));
  OAI210     u0369(.A0(men_men_n418_), .A1(men_men_n407_), .B0(x4), .Y(men_men_n419_));
  NO2        u0370(.A(x4), .B(men_men_n53_), .Y(men_men_n420_));
  NA2        u0371(.A(men_men_n420_), .B(men_men_n59_), .Y(men_men_n421_));
  NO3        u0372(.A(men_men_n421_), .B(men_men_n231_), .C(x5), .Y(men_men_n422_));
  NA2        u0373(.A(x7), .B(men_men_n108_), .Y(men_men_n423_));
  NO3        u0374(.A(x5), .B(men_men_n53_), .C(x0), .Y(men_men_n424_));
  INV        u0375(.A(men_men_n424_), .Y(men_men_n425_));
  NO2        u0376(.A(x6), .B(men_men_n56_), .Y(men_men_n426_));
  NO2        u0377(.A(x8), .B(men_men_n50_), .Y(men_men_n427_));
  NA2        u0378(.A(men_men_n427_), .B(men_men_n426_), .Y(men_men_n428_));
  OAI210     u0379(.A0(men_men_n428_), .A1(men_men_n425_), .B0(men_men_n423_), .Y(men_men_n429_));
  AOI210     u0380(.A0(men_men_n422_), .A1(x2), .B0(men_men_n429_), .Y(men_men_n430_));
  AOI220     u0381(.A0(men_men_n430_), .A1(men_men_n419_), .B0(men_men_n401_), .B1(x7), .Y(men_men_n431_));
  NA2        u0382(.A(x7), .B(men_men_n53_), .Y(men_men_n432_));
  NO2        u0383(.A(men_men_n256_), .B(men_men_n110_), .Y(men_men_n433_));
  NO2        u0384(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n434_));
  NO3        u0385(.A(men_men_n434_), .B(men_men_n433_), .C(men_men_n146_), .Y(men_men_n435_));
  AOI210     u0386(.A0(men_men_n206_), .A1(men_men_n101_), .B0(men_men_n435_), .Y(men_men_n436_));
  NO2        u0387(.A(x5), .B(x2), .Y(men_men_n437_));
  NO2        u0388(.A(x8), .B(x3), .Y(men_men_n438_));
  NA2        u0389(.A(men_men_n438_), .B(men_men_n437_), .Y(men_men_n439_));
  NO2        u0390(.A(men_men_n439_), .B(x6), .Y(men_men_n440_));
  NA2        u0391(.A(men_men_n205_), .B(x2), .Y(men_men_n441_));
  NO3        u0392(.A(men_men_n438_), .B(men_men_n344_), .C(men_men_n356_), .Y(men_men_n442_));
  AOI210     u0393(.A0(men_men_n442_), .A1(men_men_n441_), .B0(men_men_n440_), .Y(men_men_n443_));
  OAI210     u0394(.A0(men_men_n436_), .A1(men_men_n291_), .B0(men_men_n443_), .Y(men_men_n444_));
  NA2        u0395(.A(men_men_n444_), .B(x4), .Y(men_men_n445_));
  NA2        u0396(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n446_));
  NO2        u0397(.A(men_men_n446_), .B(x5), .Y(men_men_n447_));
  NAi21      u0398(.An(x4), .B(x6), .Y(men_men_n448_));
  NO2        u0399(.A(men_men_n448_), .B(men_men_n51_), .Y(men_men_n449_));
  NO2        u0400(.A(men_men_n55_), .B(men_men_n71_), .Y(men_men_n450_));
  NO2        u0401(.A(men_men_n50_), .B(men_men_n110_), .Y(men_men_n451_));
  NO2        u0402(.A(men_men_n231_), .B(x0), .Y(men_men_n452_));
  NO2        u0403(.A(men_men_n356_), .B(x8), .Y(men_men_n453_));
  OAI210     u0404(.A0(men_men_n453_), .A1(men_men_n452_), .B0(men_men_n451_), .Y(men_men_n454_));
  OAI210     u0405(.A0(men_men_n410_), .A1(men_men_n450_), .B0(men_men_n454_), .Y(men_men_n455_));
  AOI220     u0406(.A0(men_men_n455_), .A1(men_men_n56_), .B0(men_men_n449_), .B1(men_men_n447_), .Y(men_men_n456_));
  AOI210     u0407(.A0(men_men_n456_), .A1(men_men_n445_), .B0(men_men_n432_), .Y(men_men_n457_));
  NA2        u0408(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n458_));
  NO2        u0409(.A(men_men_n71_), .B(men_men_n56_), .Y(men_men_n459_));
  NA2        u0410(.A(men_men_n355_), .B(men_men_n59_), .Y(men_men_n460_));
  OAI220     u0411(.A0(men_men_n460_), .A1(men_men_n55_), .B0(men_men_n198_), .B1(men_men_n276_), .Y(men_men_n461_));
  NA2        u0412(.A(men_men_n461_), .B(men_men_n459_), .Y(men_men_n462_));
  NO3        u0413(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n463_));
  NA2        u0414(.A(men_men_n434_), .B(x5), .Y(men_men_n464_));
  NO2        u0415(.A(x8), .B(x5), .Y(men_men_n465_));
  NAi21      u0416(.An(men_men_n465_), .B(men_men_n172_), .Y(men_men_n466_));
  OAI210     u0417(.A0(men_men_n466_), .A1(men_men_n309_), .B0(men_men_n464_), .Y(men_men_n467_));
  NA2        u0418(.A(men_men_n363_), .B(men_men_n77_), .Y(men_men_n468_));
  NOi21      u0419(.An(x3), .B(x4), .Y(men_men_n469_));
  NA2        u0420(.A(men_men_n55_), .B(men_men_n110_), .Y(men_men_n470_));
  NA2        u0421(.A(men_men_n470_), .B(men_men_n469_), .Y(men_men_n471_));
  NO2        u0422(.A(men_men_n51_), .B(x6), .Y(men_men_n472_));
  NO2        u0423(.A(men_men_n146_), .B(men_men_n55_), .Y(men_men_n473_));
  NO3        u0424(.A(men_men_n56_), .B(x2), .C(x0), .Y(men_men_n474_));
  AOI220     u0425(.A0(men_men_n474_), .A1(men_men_n473_), .B0(men_men_n472_), .B1(men_men_n447_), .Y(men_men_n475_));
  OAI210     u0426(.A0(men_men_n471_), .A1(men_men_n468_), .B0(men_men_n475_), .Y(men_men_n476_));
  AOI210     u0427(.A0(men_men_n467_), .A1(men_men_n463_), .B0(men_men_n476_), .Y(men_men_n477_));
  AOI210     u0428(.A0(men_men_n477_), .A1(men_men_n462_), .B0(men_men_n458_), .Y(men_men_n478_));
  NA2        u0429(.A(x7), .B(x1), .Y(men_men_n479_));
  NO3        u0430(.A(x5), .B(x4), .C(x2), .Y(men_men_n480_));
  AN2        u0431(.A(men_men_n480_), .B(men_men_n376_), .Y(men_men_n481_));
  NO2        u0432(.A(men_men_n481_), .B(men_men_n385_), .Y(men_men_n482_));
  NA2        u0433(.A(men_men_n376_), .B(men_men_n343_), .Y(men_men_n483_));
  NO2        u0434(.A(men_men_n483_), .B(men_men_n482_), .Y(men_men_n484_));
  NO2        u0435(.A(x4), .B(men_men_n110_), .Y(men_men_n485_));
  NA2        u0436(.A(men_men_n485_), .B(x6), .Y(men_men_n486_));
  NA3        u0437(.A(men_men_n108_), .B(x4), .C(men_men_n110_), .Y(men_men_n487_));
  AOI210     u0438(.A0(men_men_n487_), .A1(men_men_n486_), .B0(men_men_n100_), .Y(men_men_n488_));
  NA2        u0439(.A(men_men_n469_), .B(men_men_n71_), .Y(men_men_n489_));
  NA2        u0440(.A(men_men_n167_), .B(men_men_n59_), .Y(men_men_n490_));
  NO2        u0441(.A(men_men_n490_), .B(men_men_n489_), .Y(men_men_n491_));
  NA2        u0442(.A(men_men_n451_), .B(x4), .Y(men_men_n492_));
  NO3        u0443(.A(men_men_n492_), .B(men_men_n376_), .C(men_men_n416_), .Y(men_men_n493_));
  NO4        u0444(.A(men_men_n493_), .B(men_men_n491_), .C(men_men_n488_), .D(men_men_n484_), .Y(men_men_n494_));
  NA2        u0445(.A(x5), .B(x4), .Y(men_men_n495_));
  NO2        u0446(.A(men_men_n71_), .B(men_men_n53_), .Y(men_men_n496_));
  NO3        u0447(.A(x8), .B(x3), .C(x2), .Y(men_men_n497_));
  NA3        u0448(.A(men_men_n497_), .B(men_men_n496_), .C(men_men_n59_), .Y(men_men_n498_));
  NO3        u0449(.A(x6), .B(x5), .C(x2), .Y(men_men_n499_));
  NA3        u0450(.A(men_men_n499_), .B(men_men_n293_), .C(men_men_n78_), .Y(men_men_n500_));
  OAI210     u0451(.A0(men_men_n498_), .A1(men_men_n495_), .B0(men_men_n500_), .Y(men_men_n501_));
  NA2        u0452(.A(men_men_n71_), .B(x2), .Y(men_men_n502_));
  NO3        u0453(.A(x4), .B(x3), .C(men_men_n59_), .Y(men_men_n503_));
  NA2        u0454(.A(men_men_n503_), .B(men_men_n228_), .Y(men_men_n504_));
  NO3        u0455(.A(men_men_n504_), .B(men_men_n502_), .C(men_men_n96_), .Y(men_men_n505_));
  XO2        u0456(.A(x4), .B(x0), .Y(men_men_n506_));
  NA2        u0457(.A(men_men_n267_), .B(x5), .Y(men_men_n507_));
  NO2        u0458(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n508_));
  NO2        u0459(.A(men_men_n508_), .B(men_men_n63_), .Y(men_men_n509_));
  NO4        u0460(.A(men_men_n509_), .B(men_men_n507_), .C(men_men_n506_), .D(men_men_n155_), .Y(men_men_n510_));
  NO3        u0461(.A(men_men_n510_), .B(men_men_n505_), .C(men_men_n501_), .Y(men_men_n511_));
  OAI210     u0462(.A0(men_men_n494_), .A1(men_men_n479_), .B0(men_men_n511_), .Y(men_men_n512_));
  NO4        u0463(.A(men_men_n512_), .B(men_men_n478_), .C(men_men_n457_), .D(men_men_n431_), .Y(men04));
  NO2        u0464(.A(x7), .B(x2), .Y(men_men_n514_));
  NO2        u0465(.A(x3), .B(men_men_n53_), .Y(men_men_n515_));
  NO2        u0466(.A(men_men_n515_), .B(men_men_n148_), .Y(men_men_n516_));
  XN2        u0467(.A(x8), .B(x1), .Y(men_men_n517_));
  NO2        u0468(.A(men_men_n517_), .B(men_men_n146_), .Y(men_men_n518_));
  NA2        u0469(.A(men_men_n518_), .B(men_men_n516_), .Y(men_men_n519_));
  NA2        u0470(.A(x6), .B(x3), .Y(men_men_n520_));
  NO2        u0471(.A(men_men_n520_), .B(x5), .Y(men_men_n521_));
  NA2        u0472(.A(men_men_n71_), .B(x1), .Y(men_men_n522_));
  NO2        u0473(.A(men_men_n465_), .B(men_men_n256_), .Y(men_men_n523_));
  NO3        u0474(.A(men_men_n523_), .B(men_men_n438_), .C(men_men_n522_), .Y(men_men_n524_));
  AOI210     u0475(.A0(men_men_n521_), .A1(men_men_n351_), .B0(men_men_n524_), .Y(men_men_n525_));
  AOI210     u0476(.A0(men_men_n525_), .A1(men_men_n519_), .B0(x0), .Y(men_men_n526_));
  NOi21      u0477(.An(men_men_n172_), .B(men_men_n465_), .Y(men_men_n527_));
  NA2        u0478(.A(men_men_n109_), .B(x1), .Y(men_men_n528_));
  NO3        u0479(.A(men_men_n528_), .B(men_men_n527_), .C(men_men_n325_), .Y(men_men_n529_));
  OAI210     u0480(.A0(men_men_n529_), .A1(men_men_n526_), .B0(men_men_n514_), .Y(men_men_n530_));
  NA2        u0481(.A(men_men_n133_), .B(men_men_n242_), .Y(men_men_n531_));
  OR4        u0482(.A(men_men_n531_), .B(men_men_n377_), .C(men_men_n82_), .D(men_men_n54_), .Y(men_men_n532_));
  OR2        u0483(.A(x6), .B(x0), .Y(men_men_n533_));
  NO3        u0484(.A(men_men_n533_), .B(x3), .C(x1), .Y(men_men_n534_));
  AOI220     u0485(.A0(men_men_n534_), .A1(men_men_n108_), .B0(men_men_n281_), .B1(men_men_n275_), .Y(men_men_n535_));
  AOI210     u0486(.A0(men_men_n535_), .A1(men_men_n532_), .B0(men_men_n185_), .Y(men_men_n536_));
  NA2        u0487(.A(x7), .B(x2), .Y(men_men_n537_));
  INV        u0488(.A(men_men_n133_), .Y(men_men_n538_));
  OAI210     u0489(.A0(men_men_n171_), .A1(men_men_n538_), .B0(men_men_n82_), .Y(men_men_n539_));
  NO2        u0490(.A(men_men_n322_), .B(men_men_n55_), .Y(men_men_n540_));
  NO3        u0491(.A(x3), .B(x1), .C(x0), .Y(men_men_n541_));
  OR2        u0492(.A(x6), .B(x1), .Y(men_men_n542_));
  NA2        u0493(.A(men_men_n542_), .B(x0), .Y(men_men_n543_));
  AOI220     u0494(.A0(men_men_n543_), .A1(men_men_n540_), .B0(men_men_n541_), .B1(men_men_n473_), .Y(men_men_n544_));
  AOI210     u0495(.A0(men_men_n544_), .A1(men_men_n539_), .B0(men_men_n537_), .Y(men_men_n545_));
  NA2        u0496(.A(men_men_n71_), .B(x0), .Y(men_men_n546_));
  NOi31      u0497(.An(men_men_n346_), .B(men_men_n546_), .C(men_men_n263_), .Y(men_men_n547_));
  NO4        u0498(.A(men_men_n547_), .B(men_men_n545_), .C(men_men_n536_), .D(men_men_n56_), .Y(men_men_n548_));
  NA2        u0499(.A(men_men_n548_), .B(men_men_n530_), .Y(men_men_n549_));
  NA3        u0500(.A(x8), .B(x7), .C(x0), .Y(men_men_n550_));
  INV        u0501(.A(men_men_n550_), .Y(men_men_n551_));
  NA2        u0502(.A(men_men_n434_), .B(men_men_n57_), .Y(men_men_n552_));
  NO2        u0503(.A(x8), .B(x0), .Y(men_men_n553_));
  NA2        u0504(.A(men_men_n553_), .B(men_men_n365_), .Y(men_men_n554_));
  AOI210     u0505(.A0(men_men_n554_), .A1(men_men_n552_), .B0(men_men_n277_), .Y(men_men_n555_));
  NA2        u0506(.A(men_men_n555_), .B(men_men_n281_), .Y(men_men_n556_));
  NO2        u0507(.A(men_men_n71_), .B(men_men_n110_), .Y(men_men_n557_));
  NO2        u0508(.A(men_men_n372_), .B(x8), .Y(men_men_n558_));
  NO2        u0509(.A(men_men_n558_), .B(men_men_n264_), .Y(men_men_n559_));
  NO3        u0510(.A(men_men_n559_), .B(men_men_n381_), .C(men_men_n270_), .Y(men_men_n560_));
  NO2        u0511(.A(men_men_n290_), .B(x8), .Y(men_men_n561_));
  OAI210     u0512(.A0(men_men_n465_), .A1(men_men_n329_), .B0(men_men_n245_), .Y(men_men_n562_));
  NA2        u0513(.A(men_men_n351_), .B(men_men_n177_), .Y(men_men_n563_));
  OAI220     u0514(.A0(men_men_n563_), .A1(men_men_n59_), .B0(men_men_n562_), .B1(men_men_n561_), .Y(men_men_n564_));
  OAI210     u0515(.A0(men_men_n564_), .A1(men_men_n560_), .B0(men_men_n557_), .Y(men_men_n565_));
  NO2        u0516(.A(x8), .B(x2), .Y(men_men_n566_));
  NO2        u0517(.A(men_men_n222_), .B(men_men_n57_), .Y(men_men_n567_));
  NA3        u0518(.A(men_men_n567_), .B(men_men_n566_), .C(men_men_n344_), .Y(men_men_n568_));
  NO2        u0519(.A(men_men_n246_), .B(men_men_n133_), .Y(men_men_n569_));
  AOI210     u0520(.A0(men_men_n326_), .A1(men_men_n163_), .B0(men_men_n569_), .Y(men_men_n570_));
  AOI210     u0521(.A0(men_men_n570_), .A1(men_men_n568_), .B0(men_men_n109_), .Y(men_men_n571_));
  NA2        u0522(.A(men_men_n341_), .B(x2), .Y(men_men_n572_));
  NO2        u0523(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n573_));
  NA2        u0524(.A(men_men_n573_), .B(men_men_n63_), .Y(men_men_n574_));
  AOI210     u0525(.A0(men_men_n572_), .A1(men_men_n460_), .B0(men_men_n574_), .Y(men_men_n575_));
  NA2        u0526(.A(men_men_n110_), .B(men_men_n53_), .Y(men_men_n576_));
  NO2        u0527(.A(men_men_n576_), .B(x8), .Y(men_men_n577_));
  NA2        u0528(.A(x7), .B(men_men_n50_), .Y(men_men_n578_));
  NO2        u0529(.A(men_men_n182_), .B(men_men_n578_), .Y(men_men_n579_));
  AN2        u0530(.A(men_men_n579_), .B(men_men_n577_), .Y(men_men_n580_));
  NA2        u0531(.A(men_men_n408_), .B(men_men_n148_), .Y(men_men_n581_));
  NO2        u0532(.A(men_men_n71_), .B(x2), .Y(men_men_n582_));
  NA2        u0533(.A(men_men_n582_), .B(men_men_n273_), .Y(men_men_n583_));
  OAI210     u0534(.A0(men_men_n583_), .A1(men_men_n581_), .B0(men_men_n56_), .Y(men_men_n584_));
  NO4        u0535(.A(men_men_n584_), .B(men_men_n580_), .C(men_men_n575_), .D(men_men_n571_), .Y(men_men_n585_));
  NA3        u0536(.A(men_men_n585_), .B(men_men_n565_), .C(men_men_n556_), .Y(men_men_n586_));
  NA2        u0537(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n587_));
  NOi21      u0538(.An(x2), .B(x7), .Y(men_men_n588_));
  NO2        u0539(.A(x6), .B(x3), .Y(men_men_n589_));
  NA2        u0540(.A(men_men_n589_), .B(men_men_n588_), .Y(men_men_n590_));
  NO2        u0541(.A(x6), .B(men_men_n59_), .Y(men_men_n591_));
  NO3        u0542(.A(men_men_n57_), .B(x2), .C(x1), .Y(men_men_n592_));
  NO3        u0543(.A(men_men_n57_), .B(x2), .C(x0), .Y(men_men_n593_));
  AOI220     u0544(.A0(men_men_n593_), .A1(men_men_n225_), .B0(men_men_n592_), .B1(men_men_n591_), .Y(men_men_n594_));
  OAI210     u0545(.A0(men_men_n590_), .A1(men_men_n587_), .B0(men_men_n594_), .Y(men_men_n595_));
  NO2        u0546(.A(men_men_n101_), .B(men_men_n53_), .Y(men_men_n596_));
  NA2        u0547(.A(men_men_n220_), .B(men_men_n57_), .Y(men_men_n597_));
  OAI210     u0548(.A0(men_men_n596_), .A1(men_men_n453_), .B0(men_men_n597_), .Y(men_men_n598_));
  NO3        u0549(.A(men_men_n598_), .B(men_men_n492_), .C(men_men_n59_), .Y(men_men_n599_));
  AO210      u0550(.A0(men_men_n595_), .A1(men_men_n465_), .B0(men_men_n599_), .Y(men_men_n600_));
  AOI210     u0551(.A0(men_men_n586_), .A1(men_men_n549_), .B0(men_men_n600_), .Y(men05));
  AOI210     u0552(.A0(men_men_n162_), .A1(men_men_n55_), .B0(men_men_n508_), .Y(men_men_n602_));
  OR2        u0553(.A(men_men_n602_), .B(men_men_n57_), .Y(men_men_n603_));
  NO2        u0554(.A(x7), .B(men_men_n108_), .Y(men_men_n604_));
  NO2        u0555(.A(x8), .B(men_men_n56_), .Y(men_men_n605_));
  NA2        u0556(.A(x5), .B(men_men_n56_), .Y(men_men_n606_));
  NO2        u0557(.A(men_men_n606_), .B(men_men_n578_), .Y(men_men_n607_));
  AOI210     u0558(.A0(men_men_n605_), .A1(men_men_n604_), .B0(men_men_n607_), .Y(men_men_n608_));
  AOI210     u0559(.A0(men_men_n608_), .A1(men_men_n603_), .B0(men_men_n110_), .Y(men_men_n609_));
  NO2        u0560(.A(x7), .B(x4), .Y(men_men_n610_));
  NO2        u0561(.A(men_men_n64_), .B(men_men_n55_), .Y(men_men_n611_));
  NO2        u0562(.A(men_men_n198_), .B(x5), .Y(men_men_n612_));
  NA2        u0563(.A(men_men_n108_), .B(men_men_n110_), .Y(men_men_n613_));
  NO2        u0564(.A(men_men_n613_), .B(men_men_n216_), .Y(men_men_n614_));
  AN2        u0565(.A(men_men_n614_), .B(men_men_n610_), .Y(men_men_n615_));
  OAI210     u0566(.A0(men_men_n615_), .A1(men_men_n609_), .B0(men_men_n496_), .Y(men_men_n616_));
  NO2        u0567(.A(x6), .B(men_men_n50_), .Y(men_men_n617_));
  NA2        u0568(.A(men_men_n55_), .B(x4), .Y(men_men_n618_));
  NO2        u0569(.A(men_men_n108_), .B(men_men_n110_), .Y(men_men_n619_));
  NA2        u0570(.A(men_men_n619_), .B(x7), .Y(men_men_n620_));
  NA2        u0571(.A(men_men_n437_), .B(men_men_n255_), .Y(men_men_n621_));
  AOI210     u0572(.A0(men_men_n621_), .A1(men_men_n620_), .B0(men_men_n618_), .Y(men_men_n622_));
  NA2        u0573(.A(men_men_n108_), .B(x4), .Y(men_men_n623_));
  XO2        u0574(.A(x7), .B(x5), .Y(men_men_n624_));
  NO2        u0575(.A(men_men_n624_), .B(men_men_n53_), .Y(men_men_n625_));
  NA3        u0576(.A(men_men_n625_), .B(men_men_n623_), .C(men_men_n330_), .Y(men_men_n626_));
  NO2        u0577(.A(men_men_n108_), .B(x2), .Y(men_men_n627_));
  NO2        u0578(.A(men_men_n75_), .B(men_men_n55_), .Y(men_men_n628_));
  NA2        u0579(.A(men_men_n628_), .B(men_men_n627_), .Y(men_men_n629_));
  NA2        u0580(.A(men_men_n629_), .B(men_men_n626_), .Y(men_men_n630_));
  OAI210     u0581(.A0(men_men_n630_), .A1(men_men_n622_), .B0(men_men_n617_), .Y(men_men_n631_));
  NO2        u0582(.A(men_men_n71_), .B(men_men_n50_), .Y(men_men_n632_));
  NO2        u0583(.A(men_men_n192_), .B(x4), .Y(men_men_n633_));
  NO2        u0584(.A(x5), .B(men_men_n56_), .Y(men_men_n634_));
  XO2        u0585(.A(x5), .B(x2), .Y(men_men_n635_));
  NO3        u0586(.A(x8), .B(x7), .C(men_men_n110_), .Y(men_men_n636_));
  AO220      u0587(.A0(men_men_n636_), .A1(men_men_n634_), .B0(men_men_n635_), .B1(men_men_n633_), .Y(men_men_n637_));
  NA3        u0588(.A(men_men_n637_), .B(men_men_n632_), .C(men_men_n53_), .Y(men_men_n638_));
  NA2        u0589(.A(men_men_n270_), .B(men_men_n588_), .Y(men_men_n639_));
  NOi21      u0590(.An(x4), .B(x1), .Y(men_men_n640_));
  NA2        u0591(.A(men_men_n640_), .B(men_men_n63_), .Y(men_men_n641_));
  NA2        u0592(.A(x4), .B(x1), .Y(men_men_n642_));
  NO2        u0593(.A(men_men_n642_), .B(men_men_n50_), .Y(men_men_n643_));
  AOI210     u0594(.A0(men_men_n643_), .A1(men_men_n619_), .B0(men_men_n59_), .Y(men_men_n644_));
  OA210      u0595(.A0(men_men_n641_), .A1(men_men_n639_), .B0(men_men_n644_), .Y(men_men_n645_));
  NA4        u0596(.A(men_men_n645_), .B(men_men_n638_), .C(men_men_n631_), .D(men_men_n616_), .Y(men_men_n646_));
  NA2        u0597(.A(men_men_n632_), .B(men_men_n56_), .Y(men_men_n647_));
  NA2        u0598(.A(men_men_n566_), .B(men_men_n604_), .Y(men_men_n648_));
  NO2        u0599(.A(men_men_n648_), .B(men_men_n647_), .Y(men_men_n649_));
  NA2        u0600(.A(men_men_n273_), .B(men_men_n122_), .Y(men_men_n650_));
  OAI210     u0601(.A0(men_men_n650_), .A1(men_men_n164_), .B0(men_men_n59_), .Y(men_men_n651_));
  NA2        u0602(.A(men_men_n57_), .B(x6), .Y(men_men_n652_));
  AOI210     u0603(.A0(men_men_n652_), .A1(x3), .B0(men_men_n91_), .Y(men_men_n653_));
  NA2        u0604(.A(men_men_n634_), .B(men_men_n154_), .Y(men_men_n654_));
  NO3        u0605(.A(men_men_n654_), .B(men_men_n653_), .C(men_men_n427_), .Y(men_men_n655_));
  NA2        u0606(.A(men_men_n282_), .B(men_men_n71_), .Y(men_men_n656_));
  NO2        u0607(.A(men_men_n389_), .B(x3), .Y(men_men_n657_));
  NO2        u0608(.A(men_men_n427_), .B(men_men_n633_), .Y(men_men_n658_));
  NO2        u0609(.A(men_men_n469_), .B(men_men_n108_), .Y(men_men_n659_));
  NO2        u0610(.A(men_men_n576_), .B(x6), .Y(men_men_n660_));
  NA2        u0611(.A(men_men_n660_), .B(men_men_n659_), .Y(men_men_n661_));
  NO2        u0612(.A(men_men_n661_), .B(men_men_n658_), .Y(men_men_n662_));
  NO4        u0613(.A(men_men_n662_), .B(men_men_n655_), .C(men_men_n651_), .D(men_men_n649_), .Y(men_men_n663_));
  NA2        u0614(.A(men_men_n57_), .B(x5), .Y(men_men_n664_));
  NO2        u0615(.A(men_men_n664_), .B(x1), .Y(men_men_n665_));
  NA2        u0616(.A(x8), .B(men_men_n56_), .Y(men_men_n666_));
  NO2        u0617(.A(men_men_n666_), .B(men_men_n128_), .Y(men_men_n667_));
  NA2        u0618(.A(x8), .B(x4), .Y(men_men_n668_));
  NO2        u0619(.A(x8), .B(x4), .Y(men_men_n669_));
  NAi21      u0620(.An(men_men_n669_), .B(men_men_n668_), .Y(men_men_n670_));
  NAi21      u0621(.An(men_men_n566_), .B(men_men_n389_), .Y(men_men_n671_));
  NO4        u0622(.A(men_men_n671_), .B(men_men_n670_), .C(men_men_n427_), .D(men_men_n71_), .Y(men_men_n672_));
  OAI210     u0623(.A0(men_men_n672_), .A1(men_men_n667_), .B0(men_men_n665_), .Y(men_men_n673_));
  NO3        u0624(.A(x8), .B(men_men_n108_), .C(x4), .Y(men_men_n674_));
  INV        u0625(.A(men_men_n674_), .Y(men_men_n675_));
  NO2        u0626(.A(men_men_n675_), .B(men_men_n110_), .Y(men_men_n676_));
  NO2        u0627(.A(x5), .B(x4), .Y(men_men_n677_));
  NA3        u0628(.A(men_men_n677_), .B(men_men_n63_), .C(men_men_n110_), .Y(men_men_n678_));
  NO2        u0629(.A(x6), .B(men_men_n110_), .Y(men_men_n679_));
  NA2        u0630(.A(men_men_n666_), .B(men_men_n679_), .Y(men_men_n680_));
  OAI210     u0631(.A0(men_men_n680_), .A1(men_men_n527_), .B0(men_men_n678_), .Y(men_men_n681_));
  OAI210     u0632(.A0(men_men_n681_), .A1(men_men_n676_), .B0(men_men_n312_), .Y(men_men_n682_));
  NA3        u0633(.A(men_men_n682_), .B(men_men_n673_), .C(men_men_n663_), .Y(men_men_n683_));
  OR2        u0634(.A(x4), .B(x1), .Y(men_men_n684_));
  NO2        u0635(.A(men_men_n684_), .B(x3), .Y(men_men_n685_));
  NA2        u0636(.A(men_men_n55_), .B(x2), .Y(men_men_n686_));
  NO3        u0637(.A(men_men_n370_), .B(men_men_n686_), .C(x6), .Y(men_men_n687_));
  AOI220     u0638(.A0(men_men_n687_), .A1(men_men_n685_), .B0(men_men_n683_), .B1(men_men_n646_), .Y(men06));
  NA2        u0639(.A(men_men_n56_), .B(x3), .Y(men_men_n689_));
  NA2        u0640(.A(x6), .B(men_men_n110_), .Y(men_men_n690_));
  NA2        u0641(.A(men_men_n690_), .B(men_men_n55_), .Y(men_men_n691_));
  NA2        u0642(.A(x5), .B(men_men_n59_), .Y(men_men_n692_));
  NO2        u0643(.A(men_men_n692_), .B(men_men_n118_), .Y(men_men_n693_));
  NA3        u0644(.A(men_men_n693_), .B(men_men_n691_), .C(men_men_n502_), .Y(men_men_n694_));
  NO2        u0645(.A(men_men_n389_), .B(x0), .Y(men_men_n695_));
  NA2        u0646(.A(men_men_n340_), .B(x2), .Y(men_men_n696_));
  NOi21      u0647(.An(x6), .B(x8), .Y(men_men_n697_));
  NO2        u0648(.A(men_men_n697_), .B(x2), .Y(men_men_n698_));
  NO3        u0649(.A(men_men_n698_), .B(men_men_n70_), .C(men_men_n59_), .Y(men_men_n699_));
  AOI220     u0650(.A0(men_men_n699_), .A1(men_men_n696_), .B0(men_men_n695_), .B1(men_men_n332_), .Y(men_men_n700_));
  AOI210     u0651(.A0(men_men_n700_), .A1(men_men_n694_), .B0(men_men_n689_), .Y(men_men_n701_));
  NA2        u0652(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n702_));
  NA2        u0653(.A(men_men_n368_), .B(men_men_n356_), .Y(men_men_n703_));
  NO2        u0654(.A(men_men_n71_), .B(men_men_n108_), .Y(men_men_n704_));
  NO2        u0655(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n705_));
  NO4        u0656(.A(men_men_n705_), .B(men_men_n686_), .C(men_men_n704_), .D(men_men_n496_), .Y(men_men_n706_));
  AOI220     u0657(.A0(men_men_n706_), .A1(men_men_n703_), .B0(men_men_n424_), .B1(men_men_n63_), .Y(men_men_n707_));
  NO2        u0658(.A(men_men_n707_), .B(men_men_n702_), .Y(men_men_n708_));
  NO2        u0659(.A(men_men_n54_), .B(x0), .Y(men_men_n709_));
  NA2        u0660(.A(x4), .B(x3), .Y(men_men_n710_));
  NO2        u0661(.A(men_men_n104_), .B(men_men_n56_), .Y(men_men_n711_));
  INV        u0662(.A(men_men_n385_), .Y(men_men_n712_));
  NO2        u0663(.A(men_men_n411_), .B(x8), .Y(men_men_n713_));
  NO2        u0664(.A(men_men_n257_), .B(men_men_n522_), .Y(men_men_n714_));
  AOI210     u0665(.A0(men_men_n713_), .A1(men_men_n265_), .B0(men_men_n714_), .Y(men_men_n715_));
  NO2        u0666(.A(x5), .B(x3), .Y(men_men_n716_));
  NA3        u0667(.A(men_men_n553_), .B(men_men_n716_), .C(x1), .Y(men_men_n717_));
  NA2        u0668(.A(men_men_n605_), .B(men_men_n557_), .Y(men_men_n718_));
  OA220      u0669(.A0(men_men_n718_), .A1(men_men_n581_), .B0(men_men_n717_), .B1(men_men_n502_), .Y(men_men_n719_));
  OAI210     u0670(.A0(men_men_n715_), .A1(men_men_n712_), .B0(men_men_n719_), .Y(men_men_n720_));
  OR3        u0671(.A(men_men_n720_), .B(men_men_n708_), .C(men_men_n701_), .Y(men_men_n721_));
  NA2        u0672(.A(x7), .B(men_men_n56_), .Y(men_men_n722_));
  NO2        u0673(.A(men_men_n619_), .B(men_men_n59_), .Y(men_men_n723_));
  NA2        u0674(.A(men_men_n723_), .B(men_men_n632_), .Y(men_men_n724_));
  NO2        u0675(.A(men_men_n170_), .B(x6), .Y(men_men_n725_));
  NA2        u0676(.A(men_men_n725_), .B(men_men_n291_), .Y(men_men_n726_));
  AOI210     u0677(.A0(men_men_n726_), .A1(men_men_n724_), .B0(men_men_n722_), .Y(men_men_n727_));
  AN2        u0678(.A(men_men_n474_), .B(men_men_n323_), .Y(men_men_n728_));
  OAI210     u0679(.A0(men_men_n728_), .A1(men_men_n727_), .B0(men_men_n351_), .Y(men_men_n729_));
  NO2        u0680(.A(men_men_n308_), .B(men_men_n108_), .Y(men_men_n730_));
  NO2        u0681(.A(men_men_n56_), .B(x3), .Y(men_men_n731_));
  NA2        u0682(.A(men_men_n731_), .B(men_men_n71_), .Y(men_men_n732_));
  NO2        u0683(.A(men_men_n732_), .B(men_men_n251_), .Y(men_men_n733_));
  NO2        u0684(.A(men_men_n71_), .B(x3), .Y(men_men_n734_));
  NA3        u0685(.A(men_men_n734_), .B(men_men_n573_), .C(men_men_n56_), .Y(men_men_n735_));
  NO2        u0686(.A(men_men_n57_), .B(x6), .Y(men_men_n736_));
  NA3        u0687(.A(men_men_n605_), .B(men_men_n329_), .C(men_men_n71_), .Y(men_men_n737_));
  NA2        u0688(.A(men_men_n737_), .B(men_men_n735_), .Y(men_men_n738_));
  OR3        u0689(.A(men_men_n738_), .B(men_men_n733_), .C(men_men_n643_), .Y(men_men_n739_));
  NA2        u0690(.A(men_men_n739_), .B(men_men_n730_), .Y(men_men_n740_));
  NA2        u0691(.A(men_men_n709_), .B(men_men_n632_), .Y(men_men_n741_));
  NA4        u0692(.A(men_men_n266_), .B(men_men_n589_), .C(men_men_n220_), .D(men_men_n258_), .Y(men_men_n742_));
  NA2        u0693(.A(men_men_n485_), .B(men_men_n67_), .Y(men_men_n743_));
  AOI210     u0694(.A0(men_men_n742_), .A1(men_men_n741_), .B0(men_men_n743_), .Y(men_men_n744_));
  NA2        u0695(.A(x7), .B(x6), .Y(men_men_n745_));
  NA3        u0696(.A(x2), .B(x1), .C(x0), .Y(men_men_n746_));
  NO3        u0697(.A(men_men_n746_), .B(men_men_n745_), .C(men_men_n602_), .Y(men_men_n747_));
  NA2        u0698(.A(men_men_n497_), .B(men_men_n147_), .Y(men_men_n748_));
  NO2        u0699(.A(x5), .B(x1), .Y(men_men_n749_));
  NA2        u0700(.A(men_men_n749_), .B(men_men_n736_), .Y(men_men_n750_));
  NA2        u0701(.A(x4), .B(x0), .Y(men_men_n751_));
  NO3        u0702(.A(men_men_n57_), .B(x6), .C(x2), .Y(men_men_n752_));
  NA2        u0703(.A(men_men_n752_), .B(men_men_n224_), .Y(men_men_n753_));
  OAI220     u0704(.A0(men_men_n753_), .A1(men_men_n751_), .B0(men_men_n750_), .B1(men_men_n748_), .Y(men_men_n754_));
  NO3        u0705(.A(men_men_n754_), .B(men_men_n747_), .C(men_men_n744_), .Y(men_men_n755_));
  NA3        u0706(.A(men_men_n755_), .B(men_men_n740_), .C(men_men_n729_), .Y(men_men_n756_));
  AOI210     u0707(.A0(men_men_n721_), .A1(men_men_n57_), .B0(men_men_n756_), .Y(men07));
  NA2        u0708(.A(men_men_n108_), .B(men_men_n59_), .Y(men_men_n758_));
  NOi21      u0709(.An(men_men_n745_), .B(men_men_n116_), .Y(men_men_n759_));
  NO4        u0710(.A(men_men_n759_), .B(men_men_n632_), .C(men_men_n251_), .D(men_men_n758_), .Y(men_men_n760_));
  NO3        u0711(.A(men_men_n57_), .B(x5), .C(x1), .Y(men_men_n761_));
  NA2        u0712(.A(men_men_n761_), .B(men_men_n376_), .Y(men_men_n762_));
  NO2        u0713(.A(men_men_n57_), .B(men_men_n71_), .Y(men_men_n763_));
  NO2        u0714(.A(men_men_n153_), .B(men_men_n109_), .Y(men_men_n764_));
  AOI210     u0715(.A0(men_men_n763_), .A1(men_men_n92_), .B0(men_men_n764_), .Y(men_men_n765_));
  OAI220     u0716(.A0(men_men_n765_), .A1(men_men_n133_), .B0(men_men_n762_), .B1(men_men_n325_), .Y(men_men_n766_));
  OAI210     u0717(.A0(men_men_n766_), .A1(men_men_n760_), .B0(x2), .Y(men_men_n767_));
  NAi21      u0718(.An(men_men_n154_), .B(men_men_n155_), .Y(men_men_n768_));
  NA3        u0719(.A(men_men_n768_), .B(men_men_n91_), .C(x3), .Y(men_men_n769_));
  NO3        u0720(.A(men_men_n55_), .B(x3), .C(x1), .Y(men_men_n770_));
  NO2        u0721(.A(men_men_n515_), .B(x2), .Y(men_men_n771_));
  AOI210     u0722(.A0(men_men_n771_), .A1(men_men_n517_), .B0(men_men_n770_), .Y(men_men_n772_));
  OAI210     u0723(.A0(men_men_n772_), .A1(men_men_n652_), .B0(men_men_n769_), .Y(men_men_n773_));
  NO2        u0724(.A(x8), .B(men_men_n53_), .Y(men_men_n774_));
  NA2        u0725(.A(men_men_n774_), .B(men_men_n59_), .Y(men_men_n775_));
  NA2        u0726(.A(men_men_n357_), .B(men_men_n351_), .Y(men_men_n776_));
  NO2        u0727(.A(x7), .B(x3), .Y(men_men_n777_));
  NA2        u0728(.A(men_men_n777_), .B(men_men_n101_), .Y(men_men_n778_));
  AOI210     u0729(.A0(men_men_n776_), .A1(men_men_n775_), .B0(men_men_n778_), .Y(men_men_n779_));
  AOI210     u0730(.A0(men_men_n773_), .A1(men_men_n250_), .B0(men_men_n779_), .Y(men_men_n780_));
  AOI210     u0731(.A0(men_men_n780_), .A1(men_men_n767_), .B0(x4), .Y(men_men_n781_));
  NA3        u0732(.A(men_men_n749_), .B(men_men_n321_), .C(men_men_n55_), .Y(men_men_n782_));
  AOI210     u0733(.A0(men_men_n782_), .A1(men_men_n598_), .B0(men_men_n110_), .Y(men_men_n783_));
  XO2        u0734(.A(x5), .B(x1), .Y(men_men_n784_));
  NO4        u0735(.A(men_men_n784_), .B(men_men_n163_), .C(men_men_n207_), .D(men_men_n55_), .Y(men_men_n785_));
  OAI210     u0736(.A0(men_men_n785_), .A1(men_men_n783_), .B0(men_men_n415_), .Y(men_men_n786_));
  NO3        u0737(.A(men_men_n50_), .B(x2), .C(x0), .Y(men_men_n787_));
  NO2        u0738(.A(men_men_n311_), .B(men_men_n108_), .Y(men_men_n788_));
  NA2        u0739(.A(x6), .B(x0), .Y(men_men_n789_));
  NO2        u0740(.A(men_men_n686_), .B(men_men_n789_), .Y(men_men_n790_));
  NO2        u0741(.A(men_men_n784_), .B(men_men_n697_), .Y(men_men_n791_));
  OAI210     u0742(.A0(men_men_n749_), .A1(men_men_n63_), .B0(men_men_n57_), .Y(men_men_n792_));
  OAI210     u0743(.A0(men_men_n792_), .A1(men_men_n791_), .B0(men_men_n762_), .Y(men_men_n793_));
  AOI220     u0744(.A0(men_men_n793_), .A1(men_men_n787_), .B0(men_men_n790_), .B1(men_men_n788_), .Y(men_men_n794_));
  AOI210     u0745(.A0(men_men_n794_), .A1(men_men_n786_), .B0(men_men_n56_), .Y(men_men_n795_));
  NOi21      u0746(.An(men_men_n231_), .B(men_men_n376_), .Y(men_men_n796_));
  NO3        u0747(.A(men_men_n796_), .B(men_men_n240_), .C(men_men_n67_), .Y(men_men_n797_));
  NO2        u0748(.A(men_men_n190_), .B(men_men_n71_), .Y(men_men_n798_));
  NO2        u0749(.A(men_men_n311_), .B(x6), .Y(men_men_n799_));
  AO220      u0750(.A0(men_men_n799_), .A1(men_men_n330_), .B0(men_men_n798_), .B1(men_men_n558_), .Y(men_men_n800_));
  OAI210     u0751(.A0(men_men_n800_), .A1(men_men_n797_), .B0(men_men_n59_), .Y(men_men_n801_));
  NA2        u0752(.A(men_men_n92_), .B(men_men_n71_), .Y(men_men_n802_));
  NO2        u0753(.A(men_men_n802_), .B(men_men_n648_), .Y(men_men_n803_));
  NAi21      u0754(.An(x8), .B(x7), .Y(men_men_n804_));
  NA2        u0755(.A(men_men_n796_), .B(men_men_n804_), .Y(men_men_n805_));
  NA2        u0756(.A(men_men_n408_), .B(men_men_n110_), .Y(men_men_n806_));
  NO2        u0757(.A(men_men_n697_), .B(x1), .Y(men_men_n807_));
  NO3        u0758(.A(men_men_n807_), .B(men_men_n806_), .C(men_men_n573_), .Y(men_men_n808_));
  AOI210     u0759(.A0(men_men_n808_), .A1(men_men_n805_), .B0(men_men_n803_), .Y(men_men_n809_));
  AOI210     u0760(.A0(men_men_n809_), .A1(men_men_n801_), .B0(men_men_n140_), .Y(men_men_n810_));
  NO2        u0761(.A(x8), .B(x7), .Y(men_men_n811_));
  NO2        u0762(.A(men_men_n811_), .B(x3), .Y(men_men_n812_));
  NA3        u0763(.A(men_men_n812_), .B(men_men_n365_), .C(x1), .Y(men_men_n813_));
  NO2        u0764(.A(x8), .B(men_men_n110_), .Y(men_men_n814_));
  AOI220     u0765(.A0(men_men_n329_), .A1(men_men_n351_), .B0(men_men_n814_), .B1(men_men_n255_), .Y(men_men_n815_));
  NO2        u0766(.A(men_men_n71_), .B(x4), .Y(men_men_n816_));
  NA2        u0767(.A(men_men_n816_), .B(men_men_n305_), .Y(men_men_n817_));
  AOI210     u0768(.A0(men_men_n815_), .A1(men_men_n813_), .B0(men_men_n817_), .Y(men_men_n818_));
  NO4        u0769(.A(men_men_n818_), .B(men_men_n810_), .C(men_men_n795_), .D(men_men_n781_), .Y(men08));
  NA2        u0770(.A(men_men_n50_), .B(x1), .Y(men_men_n820_));
  XN2        u0771(.A(x5), .B(x4), .Y(men_men_n821_));
  INV        u0772(.A(men_men_n821_), .Y(men_men_n822_));
  AOI220     u0773(.A0(men_men_n822_), .A1(men_men_n357_), .B0(men_men_n136_), .B1(men_men_n56_), .Y(men_men_n823_));
  NO2        u0774(.A(men_men_n242_), .B(men_men_n108_), .Y(men_men_n824_));
  AOI210     u0775(.A0(men_men_n824_), .A1(men_men_n279_), .B0(men_men_n191_), .Y(men_men_n825_));
  OAI220     u0776(.A0(men_men_n825_), .A1(x4), .B0(men_men_n823_), .B1(men_men_n820_), .Y(men_men_n826_));
  NA2        u0777(.A(men_men_n826_), .B(men_men_n273_), .Y(men_men_n827_));
  AOI210     u0778(.A0(men_men_n272_), .A1(men_men_n806_), .B0(men_men_n618_), .Y(men_men_n828_));
  NA2        u0779(.A(men_men_n613_), .B(men_men_n170_), .Y(men_men_n829_));
  OAI220     u0780(.A0(men_men_n829_), .A1(men_men_n666_), .B0(men_men_n487_), .B1(men_men_n50_), .Y(men_men_n830_));
  AO210      u0781(.A0(men_men_n830_), .A1(men_men_n344_), .B0(men_men_n828_), .Y(men_men_n831_));
  NA2        u0782(.A(men_men_n279_), .B(men_men_n147_), .Y(men_men_n832_));
  NA2        u0783(.A(men_men_n140_), .B(x7), .Y(men_men_n833_));
  OR3        u0784(.A(men_men_n746_), .B(men_men_n469_), .C(men_men_n716_), .Y(men_men_n834_));
  OAI220     u0785(.A0(men_men_n834_), .A1(men_men_n833_), .B0(men_men_n832_), .B1(men_men_n204_), .Y(men_men_n835_));
  AOI210     u0786(.A0(men_men_n831_), .A1(men_men_n293_), .B0(men_men_n835_), .Y(men_men_n836_));
  AOI210     u0787(.A0(men_men_n836_), .A1(men_men_n827_), .B0(men_men_n71_), .Y(men_men_n837_));
  NO2        u0788(.A(men_men_n811_), .B(men_men_n110_), .Y(men_men_n838_));
  NA2        u0789(.A(men_men_n838_), .B(men_men_n192_), .Y(men_men_n839_));
  OAI210     u0790(.A0(men_men_n411_), .A1(men_men_n305_), .B0(men_men_n344_), .Y(men_men_n840_));
  NA2        u0791(.A(men_men_n437_), .B(men_men_n233_), .Y(men_men_n841_));
  NA2        u0792(.A(men_men_n713_), .B(men_men_n107_), .Y(men_men_n842_));
  OAI220     u0793(.A0(men_men_n842_), .A1(men_men_n841_), .B0(men_men_n840_), .B1(men_men_n839_), .Y(men_men_n843_));
  NA2        u0794(.A(men_men_n843_), .B(men_men_n289_), .Y(men_men_n844_));
  NA2        u0795(.A(men_men_n334_), .B(men_men_n53_), .Y(men_men_n845_));
  NO3        u0796(.A(men_men_n411_), .B(men_men_n133_), .C(men_men_n68_), .Y(men_men_n846_));
  NO2        u0797(.A(men_men_n705_), .B(men_men_n245_), .Y(men_men_n847_));
  NO3        u0798(.A(men_men_n567_), .B(men_men_n470_), .C(men_men_n99_), .Y(men_men_n848_));
  AO220      u0799(.A0(men_men_n848_), .A1(men_men_n847_), .B0(men_men_n846_), .B1(men_men_n845_), .Y(men_men_n849_));
  NA2        u0800(.A(x7), .B(men_men_n59_), .Y(men_men_n850_));
  NO3        u0801(.A(men_men_n314_), .B(men_men_n850_), .C(men_men_n288_), .Y(men_men_n851_));
  AOI210     u0802(.A0(men_men_n849_), .A1(x5), .B0(men_men_n851_), .Y(men_men_n852_));
  AOI210     u0803(.A0(men_men_n852_), .A1(men_men_n844_), .B0(men_men_n72_), .Y(men_men_n853_));
  NO2        u0804(.A(men_men_n70_), .B(x3), .Y(men_men_n854_));
  OAI210     u0805(.A0(men_men_n854_), .A1(men_men_n264_), .B0(men_men_n145_), .Y(men_men_n855_));
  MUX2       u0806(.S(x3), .A(men_men_n163_), .B(men_men_n768_), .Y(men_men_n856_));
  NA2        u0807(.A(men_men_n856_), .B(men_men_n558_), .Y(men_men_n857_));
  NO3        u0808(.A(x6), .B(x4), .C(x0), .Y(men_men_n858_));
  INV        u0809(.A(men_men_n858_), .Y(men_men_n859_));
  AOI210     u0810(.A0(men_men_n857_), .A1(men_men_n855_), .B0(men_men_n859_), .Y(men_men_n860_));
  NO3        u0811(.A(x5), .B(x3), .C(men_men_n110_), .Y(men_men_n861_));
  AOI220     u0812(.A0(men_men_n822_), .A1(men_men_n310_), .B0(men_men_n861_), .B1(men_men_n59_), .Y(men_men_n862_));
  OR2        u0813(.A(x8), .B(x1), .Y(men_men_n863_));
  NO3        u0814(.A(men_men_n863_), .B(men_men_n862_), .C(men_men_n731_), .Y(men_men_n864_));
  NAi21      u0815(.An(x4), .B(x1), .Y(men_men_n865_));
  NO2        u0816(.A(men_men_n865_), .B(x0), .Y(men_men_n866_));
  NA2        u0817(.A(men_men_n612_), .B(men_men_n866_), .Y(men_men_n867_));
  NA3        u0818(.A(men_men_n55_), .B(x1), .C(x0), .Y(men_men_n868_));
  OAI210     u0819(.A0(men_men_n868_), .A1(men_men_n712_), .B0(men_men_n867_), .Y(men_men_n869_));
  OAI210     u0820(.A0(men_men_n869_), .A1(men_men_n864_), .B0(men_men_n321_), .Y(men_men_n870_));
  AO210      u0821(.A0(men_men_n291_), .A1(men_men_n264_), .B0(men_men_n730_), .Y(men_men_n871_));
  NA2        u0822(.A(men_men_n108_), .B(men_men_n56_), .Y(men_men_n872_));
  NO2        u0823(.A(men_men_n872_), .B(men_men_n260_), .Y(men_men_n873_));
  NO2        u0824(.A(men_men_n57_), .B(x2), .Y(men_men_n874_));
  NO4        u0825(.A(men_men_n330_), .B(men_men_n874_), .C(men_men_n811_), .D(men_men_n295_), .Y(men_men_n875_));
  AOI220     u0826(.A0(men_men_n875_), .A1(men_men_n873_), .B0(men_men_n871_), .B1(men_men_n643_), .Y(men_men_n876_));
  NA2        u0827(.A(men_men_n876_), .B(men_men_n870_), .Y(men_men_n877_));
  NO4        u0828(.A(men_men_n877_), .B(men_men_n860_), .C(men_men_n853_), .D(men_men_n837_), .Y(men09));
  NO3        u0829(.A(men_men_n784_), .B(men_men_n120_), .C(men_men_n96_), .Y(men_men_n879_));
  AOI220     u0830(.A0(men_men_n300_), .A1(men_men_n70_), .B0(men_men_n588_), .B1(men_men_n542_), .Y(men_men_n880_));
  OAI210     u0831(.A0(men_men_n879_), .A1(x2), .B0(men_men_n880_), .Y(men_men_n881_));
  AOI210     u0832(.A0(men_men_n881_), .A1(men_men_n750_), .B0(men_men_n446_), .Y(men_men_n882_));
  NO2        u0833(.A(men_men_n587_), .B(men_men_n263_), .Y(men_men_n883_));
  NO2        u0834(.A(men_men_n749_), .B(men_men_n340_), .Y(men_men_n884_));
  NO3        u0835(.A(men_men_n604_), .B(men_men_n102_), .C(men_men_n110_), .Y(men_men_n885_));
  AO220      u0836(.A0(men_men_n885_), .A1(men_men_n884_), .B0(men_men_n883_), .B1(men_men_n619_), .Y(men_men_n886_));
  OAI210     u0837(.A0(men_men_n886_), .A1(men_men_n882_), .B0(x4), .Y(men_men_n887_));
  OAI220     u0838(.A0(men_men_n368_), .A1(men_men_n142_), .B0(men_men_n395_), .B1(men_men_n281_), .Y(men_men_n888_));
  NO2        u0839(.A(men_men_n190_), .B(men_men_n108_), .Y(men_men_n889_));
  AOI220     u0840(.A0(men_men_n889_), .A1(men_men_n125_), .B0(men_men_n888_), .B1(men_men_n625_), .Y(men_men_n890_));
  NO2        u0841(.A(men_men_n784_), .B(men_men_n96_), .Y(men_men_n891_));
  NAi21      u0842(.An(x0), .B(x2), .Y(men_men_n892_));
  NO2        u0843(.A(men_men_n304_), .B(men_men_n892_), .Y(men_men_n893_));
  OAI210     u0844(.A0(men_men_n479_), .A1(men_men_n276_), .B0(men_men_n190_), .Y(men_men_n894_));
  AOI210     u0845(.A0(men_men_n166_), .A1(men_men_n804_), .B0(men_men_n356_), .Y(men_men_n895_));
  AOI220     u0846(.A0(men_men_n895_), .A1(men_men_n894_), .B0(men_men_n893_), .B1(men_men_n891_), .Y(men_men_n896_));
  OAI210     u0847(.A0(men_men_n890_), .A1(men_men_n55_), .B0(men_men_n896_), .Y(men_men_n897_));
  NA2        u0848(.A(men_men_n897_), .B(men_men_n56_), .Y(men_men_n898_));
  NO2        u0849(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n899_));
  INV        u0850(.A(men_men_n125_), .Y(men_men_n900_));
  NA2        u0851(.A(men_men_n749_), .B(men_men_n55_), .Y(men_men_n901_));
  AOI210     u0852(.A0(x6), .A1(x1), .B0(x5), .Y(men_men_n902_));
  OAI210     u0853(.A0(men_men_n902_), .A1(men_men_n333_), .B0(x2), .Y(men_men_n903_));
  AOI210     u0854(.A0(men_men_n903_), .A1(men_men_n901_), .B0(men_men_n900_), .Y(men_men_n904_));
  NA2        u0855(.A(men_men_n557_), .B(men_men_n55_), .Y(men_men_n905_));
  NO4        u0856(.A(men_men_n57_), .B(x6), .C(x5), .D(x1), .Y(men_men_n906_));
  NO2        u0857(.A(men_men_n230_), .B(men_men_n386_), .Y(men_men_n907_));
  NO2        u0858(.A(men_men_n311_), .B(men_men_n146_), .Y(men_men_n908_));
  NO3        u0859(.A(men_men_n908_), .B(men_men_n907_), .C(men_men_n906_), .Y(men_men_n909_));
  OAI220     u0860(.A0(men_men_n909_), .A1(men_men_n55_), .B0(men_men_n905_), .B1(men_men_n458_), .Y(men_men_n910_));
  OAI210     u0861(.A0(men_men_n910_), .A1(men_men_n904_), .B0(men_men_n899_), .Y(men_men_n911_));
  NO2        u0862(.A(men_men_n404_), .B(men_men_n108_), .Y(men_men_n912_));
  NO2        u0863(.A(men_men_n334_), .B(men_men_n496_), .Y(men_men_n913_));
  AOI220     u0864(.A0(men_men_n913_), .A1(men_men_n912_), .B0(men_men_n208_), .B1(men_men_n228_), .Y(men_men_n914_));
  NA4        u0865(.A(men_men_n914_), .B(men_men_n911_), .C(men_men_n898_), .D(men_men_n887_), .Y(men_men_n915_));
  NA2        u0866(.A(men_men_n915_), .B(men_men_n50_), .Y(men_men_n916_));
  NO2        u0867(.A(men_men_n379_), .B(men_men_n159_), .Y(men_men_n917_));
  NO2        u0868(.A(men_men_n432_), .B(men_men_n814_), .Y(men_men_n918_));
  OAI210     u0869(.A0(men_men_n918_), .A1(men_men_n917_), .B0(x0), .Y(men_men_n919_));
  NO3        u0870(.A(x8), .B(x7), .C(x2), .Y(men_men_n920_));
  NO3        u0871(.A(men_men_n57_), .B(x5), .C(x2), .Y(men_men_n921_));
  OAI210     u0872(.A0(men_men_n921_), .A1(men_men_n920_), .B0(men_men_n517_), .Y(men_men_n922_));
  AOI210     u0873(.A0(men_men_n922_), .A1(men_men_n919_), .B0(x4), .Y(men_men_n923_));
  NO2        u0874(.A(men_men_n425_), .B(men_men_n145_), .Y(men_men_n924_));
  NO2        u0875(.A(men_men_n52_), .B(x2), .Y(men_men_n925_));
  NO2        u0876(.A(men_men_n108_), .B(men_men_n56_), .Y(men_men_n926_));
  NA2        u0877(.A(men_men_n926_), .B(x8), .Y(men_men_n927_));
  NA2        u0878(.A(men_men_n927_), .B(men_men_n901_), .Y(men_men_n928_));
  AO210      u0879(.A0(men_men_n928_), .A1(men_men_n925_), .B0(men_men_n924_), .Y(men_men_n929_));
  OAI210     u0880(.A0(men_men_n929_), .A1(men_men_n923_), .B0(men_men_n617_), .Y(men_men_n930_));
  NO2        u0881(.A(men_men_n259_), .B(men_men_n119_), .Y(men_men_n931_));
  OAI210     u0882(.A0(x4), .A1(x2), .B0(x0), .Y(men_men_n932_));
  NA3        u0883(.A(men_men_n606_), .B(men_men_n618_), .C(men_men_n345_), .Y(men_men_n933_));
  OAI210     u0884(.A0(men_men_n932_), .A1(men_men_n288_), .B0(men_men_n53_), .Y(men_men_n934_));
  AOI210     u0885(.A0(men_men_n933_), .A1(men_men_n932_), .B0(men_men_n934_), .Y(men_men_n935_));
  OAI210     u0886(.A0(men_men_n935_), .A1(men_men_n931_), .B0(men_men_n329_), .Y(men_men_n936_));
  AOI220     u0887(.A0(men_men_n668_), .A1(men_men_n349_), .B0(men_men_n351_), .B1(men_men_n93_), .Y(men_men_n937_));
  NA2        u0888(.A(men_men_n93_), .B(x5), .Y(men_men_n938_));
  OAI220     u0889(.A0(men_men_n938_), .A1(men_men_n863_), .B0(men_men_n937_), .B1(men_men_n322_), .Y(men_men_n939_));
  NA2        u0890(.A(men_men_n939_), .B(men_men_n68_), .Y(men_men_n940_));
  NA2        u0891(.A(men_men_n408_), .B(men_men_n768_), .Y(men_men_n941_));
  NA2        u0892(.A(men_men_n250_), .B(men_men_n163_), .Y(men_men_n942_));
  AO210      u0893(.A0(men_men_n942_), .A1(men_men_n941_), .B0(men_men_n130_), .Y(men_men_n943_));
  NO2        u0894(.A(men_men_n438_), .B(x2), .Y(men_men_n944_));
  NO2        u0895(.A(x7), .B(men_men_n53_), .Y(men_men_n945_));
  NA2        u0896(.A(men_men_n945_), .B(x5), .Y(men_men_n946_));
  NO2        u0897(.A(men_men_n946_), .B(men_men_n60_), .Y(men_men_n947_));
  AOI220     u0898(.A0(men_men_n947_), .A1(men_men_n944_), .B0(men_men_n669_), .B1(men_men_n243_), .Y(men_men_n948_));
  NA4        u0899(.A(men_men_n948_), .B(men_men_n943_), .C(men_men_n940_), .D(men_men_n936_), .Y(men_men_n949_));
  NO4        u0900(.A(men_men_n933_), .B(men_men_n634_), .C(men_men_n458_), .D(men_men_n50_), .Y(men_men_n950_));
  AOI220     u0901(.A0(men_men_n605_), .A1(men_men_n604_), .B0(men_men_n282_), .B1(x5), .Y(men_men_n951_));
  NO2        u0902(.A(men_men_n677_), .B(men_men_n190_), .Y(men_men_n952_));
  NA3        u0903(.A(men_men_n952_), .B(men_men_n670_), .C(x7), .Y(men_men_n953_));
  OAI210     u0904(.A0(men_men_n951_), .A1(men_men_n350_), .B0(men_men_n953_), .Y(men_men_n954_));
  OAI210     u0905(.A0(men_men_n954_), .A1(men_men_n950_), .B0(men_men_n82_), .Y(men_men_n955_));
  NA2        u0906(.A(men_men_n774_), .B(x2), .Y(men_men_n956_));
  NO2        u0907(.A(men_men_n956_), .B(men_men_n58_), .Y(men_men_n957_));
  NO2        u0908(.A(x5), .B(men_men_n53_), .Y(men_men_n958_));
  NAi21      u0909(.An(x1), .B(x4), .Y(men_men_n959_));
  NA2        u0910(.A(men_men_n959_), .B(men_men_n865_), .Y(men_men_n960_));
  NO3        u0911(.A(men_men_n960_), .B(men_men_n201_), .C(men_men_n958_), .Y(men_men_n961_));
  OAI210     u0912(.A0(men_men_n961_), .A1(men_men_n957_), .B0(men_men_n415_), .Y(men_men_n962_));
  NA3        u0913(.A(men_men_n398_), .B(men_men_n749_), .C(men_men_n57_), .Y(men_men_n963_));
  NA3        u0914(.A(men_men_n963_), .B(men_men_n962_), .C(men_men_n955_), .Y(men_men_n964_));
  AOI210     u0915(.A0(men_men_n949_), .A1(x6), .B0(men_men_n964_), .Y(men_men_n965_));
  NA3        u0916(.A(men_men_n965_), .B(men_men_n930_), .C(men_men_n916_), .Y(men10));
  NO2        u0917(.A(x4), .B(x1), .Y(men_men_n967_));
  NO2        u0918(.A(men_men_n967_), .B(men_men_n147_), .Y(men_men_n968_));
  NA3        u0919(.A(x5), .B(x4), .C(x0), .Y(men_men_n969_));
  OAI220     u0920(.A0(men_men_n969_), .A1(men_men_n277_), .B0(men_men_n705_), .B1(men_men_n247_), .Y(men_men_n970_));
  NA2        u0921(.A(men_men_n970_), .B(men_men_n968_), .Y(men_men_n971_));
  NO3        u0922(.A(men_men_n357_), .B(men_men_n322_), .C(men_men_n92_), .Y(men_men_n972_));
  NA3        u0923(.A(men_men_n972_), .B(men_men_n384_), .C(men_men_n62_), .Y(men_men_n973_));
  AOI210     u0924(.A0(men_men_n973_), .A1(men_men_n971_), .B0(men_men_n304_), .Y(men_men_n974_));
  NOi21      u0925(.An(men_men_n258_), .B(men_men_n136_), .Y(men_men_n975_));
  AOI210     u0926(.A0(men_men_n503_), .A1(men_men_n619_), .B0(men_men_n330_), .Y(men_men_n976_));
  NO2        u0927(.A(men_men_n899_), .B(men_men_n343_), .Y(men_men_n977_));
  NOi31      u0928(.An(men_men_n977_), .B(men_men_n976_), .C(men_men_n975_), .Y(men_men_n978_));
  NA2        u0929(.A(x4), .B(men_men_n110_), .Y(men_men_n979_));
  NO2        u0930(.A(men_men_n325_), .B(men_men_n979_), .Y(men_men_n980_));
  NA2        u0931(.A(men_men_n99_), .B(x5), .Y(men_men_n981_));
  NO3        u0932(.A(men_men_n981_), .B(men_men_n111_), .C(men_men_n55_), .Y(men_men_n982_));
  NO3        u0933(.A(men_men_n982_), .B(men_men_n980_), .C(men_men_n978_), .Y(men_men_n983_));
  NA2        u0934(.A(men_men_n958_), .B(men_men_n50_), .Y(men_men_n984_));
  NA2        u0935(.A(men_men_n605_), .B(men_men_n271_), .Y(men_men_n985_));
  NO2        u0936(.A(men_men_n985_), .B(men_men_n984_), .Y(men_men_n986_));
  OAI220     u0937(.A0(men_men_n927_), .A1(men_men_n107_), .B0(men_men_n872_), .B1(men_men_n446_), .Y(men_men_n987_));
  AOI210     u0938(.A0(men_men_n987_), .A1(men_men_n279_), .B0(men_men_n986_), .Y(men_men_n988_));
  OAI210     u0939(.A0(men_men_n983_), .A1(men_men_n386_), .B0(men_men_n988_), .Y(men_men_n989_));
  OAI210     u0940(.A0(men_men_n989_), .A1(men_men_n974_), .B0(x7), .Y(men_men_n990_));
  NA2        u0941(.A(men_men_n55_), .B(men_men_n71_), .Y(men_men_n991_));
  AOI210     u0942(.A0(men_men_n446_), .A1(men_men_n356_), .B0(men_men_n979_), .Y(men_men_n992_));
  NO3        u0943(.A(men_men_n448_), .B(men_men_n892_), .C(x5), .Y(men_men_n993_));
  OAI210     u0944(.A0(men_men_n993_), .A1(men_men_n992_), .B0(men_men_n991_), .Y(men_men_n994_));
  NO2        u0945(.A(men_men_n357_), .B(men_men_n139_), .Y(men_men_n995_));
  NA2        u0946(.A(men_men_n995_), .B(men_men_n426_), .Y(men_men_n996_));
  AOI210     u0947(.A0(men_men_n996_), .A1(men_men_n994_), .B0(x3), .Y(men_men_n997_));
  NO2        u0948(.A(x5), .B(men_men_n110_), .Y(men_men_n998_));
  NA2        u0949(.A(men_men_n237_), .B(men_men_n938_), .Y(men_men_n999_));
  NA3        u0950(.A(men_men_n465_), .B(men_men_n128_), .C(men_men_n426_), .Y(men_men_n1000_));
  OAI210     u0951(.A0(men_men_n448_), .A1(men_men_n213_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  AOI210     u0952(.A0(men_men_n999_), .A1(men_men_n256_), .B0(men_men_n1001_), .Y(men_men_n1002_));
  NO2        u0953(.A(men_men_n1002_), .B(men_men_n59_), .Y(men_men_n1003_));
  OAI210     u0954(.A0(men_men_n1003_), .A1(men_men_n997_), .B0(men_men_n945_), .Y(men_men_n1004_));
  NO2        u0955(.A(x4), .B(x3), .Y(men_men_n1005_));
  NO3        u0956(.A(men_men_n1005_), .B(men_men_n344_), .C(men_men_n87_), .Y(men_men_n1006_));
  OAI210     u0957(.A0(men_men_n1006_), .A1(men_men_n278_), .B0(men_men_n437_), .Y(men_men_n1007_));
  AOI210     u0958(.A0(men_men_n399_), .A1(men_men_n127_), .B0(men_men_n251_), .Y(men_men_n1008_));
  NA2        u0959(.A(men_men_n967_), .B(men_men_n55_), .Y(men_men_n1009_));
  NO2        u0960(.A(men_men_n1009_), .B(men_men_n981_), .Y(men_men_n1010_));
  NO2        u0961(.A(men_men_n527_), .B(men_men_n362_), .Y(men_men_n1011_));
  NO3        u0962(.A(x4), .B(men_men_n110_), .C(men_men_n59_), .Y(men_men_n1012_));
  NO2        u0963(.A(men_men_n438_), .B(x1), .Y(men_men_n1013_));
  NOi31      u0964(.An(men_men_n1012_), .B(men_men_n1013_), .C(men_men_n1011_), .Y(men_men_n1014_));
  NA2        u0965(.A(men_men_n55_), .B(x5), .Y(men_men_n1015_));
  NO4        u0966(.A(men_men_n968_), .B(men_men_n516_), .C(men_men_n1015_), .D(x2), .Y(men_men_n1016_));
  NO4        u0967(.A(men_men_n1016_), .B(men_men_n1014_), .C(men_men_n1010_), .D(men_men_n1008_), .Y(men_men_n1017_));
  AOI210     u0968(.A0(men_men_n1017_), .A1(men_men_n1007_), .B0(men_men_n207_), .Y(men_men_n1018_));
  NO2        u0969(.A(men_men_n666_), .B(men_men_n502_), .Y(men_men_n1019_));
  NO2        u0970(.A(x6), .B(x2), .Y(men_men_n1020_));
  NO3        u0971(.A(men_men_n1020_), .B(men_men_n697_), .C(men_men_n60_), .Y(men_men_n1021_));
  OAI210     u0972(.A0(men_men_n1021_), .A1(men_men_n1019_), .B0(men_men_n270_), .Y(men_men_n1022_));
  NO2        u0973(.A(men_men_n872_), .B(men_men_n446_), .Y(men_men_n1023_));
  NA3        u0974(.A(x4), .B(x3), .C(men_men_n110_), .Y(men_men_n1024_));
  NO3        u0975(.A(men_men_n1024_), .B(men_men_n703_), .C(men_men_n465_), .Y(men_men_n1025_));
  AOI210     u0976(.A0(men_men_n1023_), .A1(men_men_n472_), .B0(men_men_n1025_), .Y(men_men_n1026_));
  AOI210     u0977(.A0(men_men_n1026_), .A1(men_men_n1022_), .B0(men_men_n458_), .Y(men_men_n1027_));
  NO2        u0978(.A(men_men_n55_), .B(men_men_n56_), .Y(men_men_n1028_));
  OAI220     u0979(.A0(men_men_n822_), .A1(men_men_n460_), .B0(men_men_n751_), .B1(men_men_n127_), .Y(men_men_n1029_));
  NOi21      u0980(.An(men_men_n123_), .B(men_men_n122_), .Y(men_men_n1030_));
  NO3        u0981(.A(men_men_n345_), .B(men_men_n325_), .C(men_men_n1030_), .Y(men_men_n1031_));
  AOI220     u0982(.A0(men_men_n1031_), .A1(men_men_n255_), .B0(men_men_n1029_), .B1(men_men_n116_), .Y(men_men_n1032_));
  NO2        u0983(.A(men_men_n1032_), .B(men_men_n1028_), .Y(men_men_n1033_));
  NA2        u0984(.A(men_men_n520_), .B(men_men_n260_), .Y(men_men_n1034_));
  NO2        u0985(.A(men_men_n487_), .B(men_men_n587_), .Y(men_men_n1035_));
  NA3        u0986(.A(men_men_n1035_), .B(men_men_n1034_), .C(men_men_n55_), .Y(men_men_n1036_));
  NO2        u0987(.A(men_men_n182_), .B(men_men_n110_), .Y(men_men_n1037_));
  NA3        u0988(.A(men_men_n1037_), .B(men_men_n181_), .C(men_men_n122_), .Y(men_men_n1038_));
  NA2        u0989(.A(men_men_n1038_), .B(men_men_n1036_), .Y(men_men_n1039_));
  NO4        u0990(.A(men_men_n1039_), .B(men_men_n1033_), .C(men_men_n1027_), .D(men_men_n1018_), .Y(men_men_n1040_));
  NA3        u0991(.A(men_men_n1040_), .B(men_men_n1004_), .C(men_men_n990_), .Y(men11));
  NA2        u0992(.A(men_men_n377_), .B(men_men_n92_), .Y(men_men_n1042_));
  INV        u0993(.A(men_men_n893_), .Y(men_men_n1043_));
  OAI220     u0994(.A0(men_men_n1043_), .A1(men_men_n53_), .B0(men_men_n1042_), .B1(men_men_n366_), .Y(men_men_n1044_));
  NO2        u0995(.A(men_men_n768_), .B(x5), .Y(men_men_n1045_));
  NO2        u0996(.A(men_men_n167_), .B(men_men_n533_), .Y(men_men_n1046_));
  AOI220     u0997(.A0(men_men_n1046_), .A1(men_men_n1045_), .B0(men_men_n1044_), .B1(x5), .Y(men_men_n1047_));
  OAI220     u0998(.A0(men_men_n975_), .A1(men_men_n216_), .B0(men_men_n214_), .B1(men_men_n182_), .Y(men_men_n1048_));
  NO2        u0999(.A(men_men_n341_), .B(men_men_n427_), .Y(men_men_n1049_));
  AOI220     u1000(.A0(men_men_n1049_), .A1(men_men_n180_), .B0(men_men_n1048_), .B1(men_men_n163_), .Y(men_men_n1050_));
  NO2        u1001(.A(men_men_n1050_), .B(men_men_n448_), .Y(men_men_n1051_));
  NO2        u1002(.A(men_men_n251_), .B(x2), .Y(men_men_n1052_));
  OAI210     u1003(.A0(men_men_n917_), .A1(men_men_n1052_), .B0(men_men_n416_), .Y(men_men_n1053_));
  NO2        u1004(.A(men_men_n55_), .B(men_men_n108_), .Y(men_men_n1054_));
  NO2        u1005(.A(men_men_n71_), .B(x1), .Y(men_men_n1055_));
  NA2        u1006(.A(men_men_n1055_), .B(men_men_n78_), .Y(men_men_n1056_));
  OR2        u1007(.A(men_men_n1056_), .B(men_men_n613_), .Y(men_men_n1057_));
  AOI210     u1008(.A0(men_men_n1057_), .A1(men_men_n1053_), .B0(men_men_n710_), .Y(men_men_n1058_));
  NO2        u1009(.A(men_men_n305_), .B(men_men_n53_), .Y(men_men_n1059_));
  NO2        u1010(.A(men_men_n437_), .B(x3), .Y(men_men_n1060_));
  NA3        u1011(.A(men_men_n1060_), .B(men_men_n1059_), .C(men_men_n892_), .Y(men_men_n1061_));
  AOI210     u1012(.A0(men_men_n1061_), .A1(men_men_n942_), .B0(men_men_n397_), .Y(men_men_n1062_));
  NA2        u1013(.A(men_men_n110_), .B(x1), .Y(men_men_n1063_));
  NO2        u1014(.A(men_men_n619_), .B(men_men_n219_), .Y(men_men_n1064_));
  NA4        u1015(.A(men_men_n1064_), .B(men_men_n884_), .C(men_men_n469_), .D(men_men_n1063_), .Y(men_men_n1065_));
  NA3        u1016(.A(x6), .B(x5), .C(men_men_n110_), .Y(men_men_n1066_));
  NO2        u1017(.A(men_men_n1066_), .B(men_men_n277_), .Y(men_men_n1067_));
  NO2        u1018(.A(men_men_n448_), .B(x0), .Y(men_men_n1068_));
  NOi31      u1019(.An(men_men_n1068_), .B(men_men_n172_), .C(men_men_n51_), .Y(men_men_n1069_));
  AOI210     u1020(.A0(men_men_n1067_), .A1(men_men_n178_), .B0(men_men_n1069_), .Y(men_men_n1070_));
  NA2        u1021(.A(men_men_n1070_), .B(men_men_n1065_), .Y(men_men_n1071_));
  NO4        u1022(.A(men_men_n1071_), .B(men_men_n1062_), .C(men_men_n1058_), .D(men_men_n1051_), .Y(men_men_n1072_));
  OAI210     u1023(.A0(men_men_n1047_), .A1(men_men_n140_), .B0(men_men_n1072_), .Y(men_men_n1073_));
  NA2        u1024(.A(men_men_n863_), .B(men_men_n87_), .Y(men_men_n1074_));
  NO3        u1025(.A(men_men_n466_), .B(men_men_n774_), .C(men_men_n123_), .Y(men_men_n1075_));
  AOI210     u1026(.A0(men_men_n1074_), .A1(men_men_n101_), .B0(men_men_n1075_), .Y(men_men_n1076_));
  NO2        u1027(.A(x8), .B(x1), .Y(men_men_n1077_));
  NO3        u1028(.A(men_men_n1077_), .B(men_men_n689_), .C(men_men_n450_), .Y(men_men_n1078_));
  OAI210     u1029(.A0(men_men_n77_), .A1(men_men_n53_), .B0(men_men_n1078_), .Y(men_men_n1079_));
  OAI210     u1030(.A0(men_men_n1076_), .A1(x3), .B0(men_men_n1079_), .Y(men_men_n1080_));
  NO2        u1031(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n1081_));
  OAI210     u1032(.A0(men_men_n1081_), .A1(x2), .B0(men_men_n233_), .Y(men_men_n1082_));
  NO2        u1033(.A(men_men_n606_), .B(men_men_n231_), .Y(men_men_n1083_));
  NA2        u1034(.A(men_men_n1083_), .B(men_men_n1082_), .Y(men_men_n1084_));
  NO2        u1035(.A(men_men_n520_), .B(x4), .Y(men_men_n1085_));
  NO3        u1036(.A(men_men_n55_), .B(x6), .C(x1), .Y(men_men_n1086_));
  NA2        u1037(.A(men_men_n1085_), .B(men_men_n577_), .Y(men_men_n1087_));
  NA2        u1038(.A(men_men_n1087_), .B(men_men_n1084_), .Y(men_men_n1088_));
  AOI210     u1039(.A0(men_men_n1080_), .A1(x2), .B0(men_men_n1088_), .Y(men_men_n1089_));
  NO2        u1040(.A(men_men_n231_), .B(x2), .Y(men_men_n1090_));
  NA2        u1041(.A(men_men_n1090_), .B(men_men_n1005_), .Y(men_men_n1091_));
  NOi21      u1042(.An(men_men_n389_), .B(men_men_n566_), .Y(men_men_n1092_));
  NO3        u1043(.A(men_men_n1092_), .B(men_men_n605_), .C(men_men_n325_), .Y(men_men_n1093_));
  NA2        u1044(.A(x8), .B(men_men_n110_), .Y(men_men_n1094_));
  OAI220     u1045(.A0(men_men_n710_), .A1(men_men_n1094_), .B0(men_men_n325_), .B1(men_men_n384_), .Y(men_men_n1095_));
  OAI210     u1046(.A0(men_men_n1095_), .A1(men_men_n1093_), .B0(men_men_n71_), .Y(men_men_n1096_));
  NO2        u1047(.A(men_men_n108_), .B(x1), .Y(men_men_n1097_));
  NA2        u1048(.A(men_men_n1097_), .B(x7), .Y(men_men_n1098_));
  AOI210     u1049(.A0(men_men_n1096_), .A1(men_men_n1091_), .B0(men_men_n1098_), .Y(men_men_n1099_));
  NA2        u1050(.A(men_men_n84_), .B(men_men_n71_), .Y(men_men_n1100_));
  INV        u1051(.A(men_men_n248_), .Y(men_men_n1101_));
  NA2        u1052(.A(men_men_n1101_), .B(men_men_n147_), .Y(men_men_n1102_));
  OAI220     u1053(.A0(men_men_n1102_), .A1(men_men_n366_), .B0(men_men_n1100_), .B1(men_men_n325_), .Y(men_men_n1103_));
  NO2        u1054(.A(men_men_n157_), .B(men_men_n55_), .Y(men_men_n1104_));
  AOI210     u1055(.A0(men_men_n1104_), .A1(men_men_n1103_), .B0(men_men_n1099_), .Y(men_men_n1105_));
  OAI210     u1056(.A0(men_men_n1089_), .A1(men_men_n850_), .B0(men_men_n1105_), .Y(men_men_n1106_));
  AO210      u1057(.A0(men_men_n1073_), .A1(men_men_n57_), .B0(men_men_n1106_), .Y(men12));
  NA2        u1058(.A(men_men_n883_), .B(men_men_n247_), .Y(men_men_n1108_));
  NO2        u1059(.A(men_men_n623_), .B(x7), .Y(men_men_n1109_));
  NA2        u1060(.A(men_men_n1109_), .B(men_men_n278_), .Y(men_men_n1110_));
  NA2        u1061(.A(men_men_n702_), .B(men_men_n872_), .Y(men_men_n1111_));
  AOI210     u1062(.A0(men_men_n1110_), .A1(men_men_n1108_), .B0(men_men_n1111_), .Y(men_men_n1112_));
  NOi21      u1063(.An(men_men_n404_), .B(men_men_n553_), .Y(men_men_n1113_));
  NO2        u1064(.A(x7), .B(men_men_n50_), .Y(men_men_n1114_));
  NO2        u1065(.A(men_men_n606_), .B(men_men_n1114_), .Y(men_men_n1115_));
  NO3        u1066(.A(men_men_n865_), .B(men_men_n112_), .C(men_men_n99_), .Y(men_men_n1116_));
  AOI210     u1067(.A0(men_men_n1115_), .A1(men_men_n1013_), .B0(men_men_n1116_), .Y(men_men_n1117_));
  NA2        u1068(.A(men_men_n1054_), .B(men_men_n56_), .Y(men_men_n1118_));
  OAI220     u1069(.A0(men_men_n1118_), .A1(men_men_n578_), .B0(men_men_n1117_), .B1(men_men_n1113_), .Y(men_men_n1119_));
  OAI210     u1070(.A0(men_men_n1119_), .A1(men_men_n1112_), .B0(men_men_n582_), .Y(men_men_n1120_));
  NA2        u1071(.A(men_men_n87_), .B(x5), .Y(men_men_n1121_));
  OAI210     u1072(.A0(men_men_n1121_), .A1(men_men_n325_), .B0(men_men_n717_), .Y(men_men_n1122_));
  INV        u1073(.A(men_men_n1122_), .Y(men_men_n1123_));
  NA2        u1074(.A(men_men_n604_), .B(men_men_n53_), .Y(men_men_n1124_));
  NA2        u1075(.A(men_men_n288_), .B(men_men_n50_), .Y(men_men_n1125_));
  OAI220     u1076(.A0(men_men_n1125_), .A1(men_men_n311_), .B0(men_men_n1124_), .B1(men_men_n133_), .Y(men_men_n1126_));
  NA2        u1077(.A(men_men_n1126_), .B(men_men_n56_), .Y(men_men_n1127_));
  OAI210     u1078(.A0(men_men_n1123_), .A1(men_men_n64_), .B0(men_men_n1127_), .Y(men_men_n1128_));
  NO2        u1079(.A(men_men_n57_), .B(x0), .Y(men_men_n1129_));
  NO2        u1080(.A(men_men_n666_), .B(men_men_n322_), .Y(men_men_n1130_));
  NO2        u1081(.A(men_men_n751_), .B(x3), .Y(men_men_n1131_));
  NO2        u1082(.A(men_men_n664_), .B(x8), .Y(men_men_n1132_));
  AOI220     u1083(.A0(men_men_n1132_), .A1(men_men_n1131_), .B0(men_men_n1130_), .B1(men_men_n1129_), .Y(men_men_n1133_));
  AOI210     u1084(.A0(men_men_n689_), .A1(men_men_n247_), .B0(x7), .Y(men_men_n1134_));
  NO3        u1085(.A(men_men_n1134_), .B(men_men_n607_), .C(x8), .Y(men_men_n1135_));
  NA4        u1086(.A(men_men_n668_), .B(men_men_n660_), .C(men_men_n204_), .D(x0), .Y(men_men_n1136_));
  OAI220     u1087(.A0(men_men_n1136_), .A1(men_men_n1135_), .B0(men_men_n1133_), .B1(men_men_n576_), .Y(men_men_n1137_));
  AOI210     u1088(.A0(men_men_n1128_), .A1(men_men_n1020_), .B0(men_men_n1137_), .Y(men_men_n1138_));
  NO2        u1089(.A(men_men_n247_), .B(men_men_n55_), .Y(men_men_n1139_));
  NO2        u1090(.A(men_men_n255_), .B(x8), .Y(men_men_n1140_));
  NOi32      u1091(.An(men_men_n1140_), .Bn(men_men_n203_), .C(men_men_n567_), .Y(men_men_n1141_));
  NO2        u1092(.A(men_men_n88_), .B(men_men_n60_), .Y(men_men_n1142_));
  OAI210     u1093(.A0(men_men_n1141_), .A1(men_men_n1139_), .B0(men_men_n1142_), .Y(men_men_n1143_));
  NO2        u1094(.A(men_men_n945_), .B(men_men_n100_), .Y(men_men_n1144_));
  NO2        u1095(.A(men_men_n166_), .B(men_men_n53_), .Y(men_men_n1145_));
  AOI210     u1096(.A0(men_men_n341_), .A1(x8), .B0(men_men_n1145_), .Y(men_men_n1146_));
  AOI210     u1097(.A0(men_men_n216_), .A1(men_men_n96_), .B0(men_men_n1146_), .Y(men_men_n1147_));
  OAI210     u1098(.A0(men_men_n1147_), .A1(men_men_n1144_), .B0(men_men_n677_), .Y(men_men_n1148_));
  NO2        u1099(.A(x7), .B(x0), .Y(men_men_n1149_));
  NO3        u1100(.A(men_men_n157_), .B(men_men_n1149_), .C(men_men_n144_), .Y(men_men_n1150_));
  XN2        u1101(.A(x8), .B(x7), .Y(men_men_n1151_));
  NO3        u1102(.A(men_men_n1077_), .B(men_men_n258_), .C(men_men_n1151_), .Y(men_men_n1152_));
  OAI210     u1103(.A0(men_men_n1152_), .A1(men_men_n1150_), .B0(men_men_n731_), .Y(men_men_n1153_));
  NO2        u1104(.A(men_men_n267_), .B(men_men_n263_), .Y(men_men_n1154_));
  NO2        u1105(.A(men_men_n108_), .B(x4), .Y(men_men_n1155_));
  OAI210     u1106(.A0(men_men_n1154_), .A1(men_men_n278_), .B0(men_men_n1155_), .Y(men_men_n1156_));
  NA4        u1107(.A(men_men_n1156_), .B(men_men_n1153_), .C(men_men_n1148_), .D(men_men_n1143_), .Y(men_men_n1157_));
  NA2        u1108(.A(men_men_n1157_), .B(men_men_n557_), .Y(men_men_n1158_));
  NO2        u1109(.A(men_men_n55_), .B(x4), .Y(men_men_n1159_));
  NA2        u1110(.A(men_men_n1159_), .B(men_men_n162_), .Y(men_men_n1160_));
  NO2        u1111(.A(men_men_n670_), .B(men_men_n258_), .Y(men_men_n1161_));
  OAI210     u1112(.A0(men_men_n1161_), .A1(men_men_n1023_), .B0(men_men_n50_), .Y(men_men_n1162_));
  AOI210     u1113(.A0(men_men_n1162_), .A1(men_men_n1160_), .B0(men_men_n432_), .Y(men_men_n1163_));
  OAI220     u1114(.A0(men_men_n290_), .A1(men_men_n276_), .B0(men_men_n263_), .B1(men_men_n242_), .Y(men_men_n1164_));
  NA3        u1115(.A(men_men_n1164_), .B(men_men_n677_), .C(x1), .Y(men_men_n1165_));
  OAI210     u1116(.A0(x8), .A1(x0), .B0(x4), .Y(men_men_n1166_));
  NO2        u1117(.A(x7), .B(men_men_n56_), .Y(men_men_n1167_));
  NO2        u1118(.A(men_men_n68_), .B(men_men_n1167_), .Y(men_men_n1168_));
  NOi21      u1119(.An(men_men_n1166_), .B(men_men_n1168_), .Y(men_men_n1169_));
  NO2        u1120(.A(men_men_n668_), .B(men_men_n325_), .Y(men_men_n1170_));
  NO2        u1121(.A(men_men_n777_), .B(men_men_n220_), .Y(men_men_n1171_));
  OAI210     u1122(.A0(men_men_n1170_), .A1(men_men_n1169_), .B0(men_men_n1171_), .Y(men_men_n1172_));
  NO2        u1123(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n1173_));
  NO2        u1124(.A(men_men_n606_), .B(men_men_n446_), .Y(men_men_n1174_));
  OAI210     u1125(.A0(men_men_n1174_), .A1(men_men_n1173_), .B0(men_men_n255_), .Y(men_men_n1175_));
  NO2        u1126(.A(men_men_n820_), .B(men_men_n423_), .Y(men_men_n1176_));
  NA2        u1127(.A(men_men_n329_), .B(men_men_n59_), .Y(men_men_n1177_));
  NO2        u1128(.A(men_men_n1118_), .B(men_men_n1177_), .Y(men_men_n1178_));
  AOI210     u1129(.A0(men_men_n1176_), .A1(men_men_n178_), .B0(men_men_n1178_), .Y(men_men_n1179_));
  NA4        u1130(.A(men_men_n1179_), .B(men_men_n1175_), .C(men_men_n1172_), .D(men_men_n1165_), .Y(men_men_n1180_));
  OAI210     u1131(.A0(men_men_n1180_), .A1(men_men_n1163_), .B0(men_men_n679_), .Y(men_men_n1181_));
  NA4        u1132(.A(men_men_n1181_), .B(men_men_n1158_), .C(men_men_n1138_), .D(men_men_n1120_), .Y(men13));
  NO2        u1133(.A(men_men_n465_), .B(men_men_n351_), .Y(men_men_n1183_));
  NOi41      u1134(.An(men_men_n1183_), .B(men_men_n677_), .C(men_men_n292_), .D(men_men_n239_), .Y(men_men_n1184_));
  NO2        u1135(.A(men_men_n865_), .B(men_men_n182_), .Y(men_men_n1185_));
  NO2        u1136(.A(men_men_n156_), .B(men_men_n71_), .Y(men_men_n1186_));
  XN2        u1137(.A(x4), .B(x0), .Y(men_men_n1187_));
  NO3        u1138(.A(men_men_n1187_), .B(men_men_n111_), .C(men_men_n423_), .Y(men_men_n1188_));
  AO220      u1139(.A0(men_men_n1188_), .A1(men_men_n1186_), .B0(men_men_n1185_), .B1(men_men_n330_), .Y(men_men_n1189_));
  OAI210     u1140(.A0(men_men_n1189_), .A1(men_men_n1184_), .B0(x3), .Y(men_men_n1190_));
  NO2        u1141(.A(men_men_n865_), .B(x6), .Y(men_men_n1191_));
  NO2        u1142(.A(men_men_n1125_), .B(men_men_n395_), .Y(men_men_n1192_));
  NO3        u1143(.A(x8), .B(x5), .C(men_men_n110_), .Y(men_men_n1193_));
  NA2        u1144(.A(men_men_n1193_), .B(men_men_n643_), .Y(men_men_n1194_));
  NO2        u1145(.A(men_men_n606_), .B(men_men_n198_), .Y(men_men_n1195_));
  NA2        u1146(.A(men_men_n1195_), .B(men_men_n1086_), .Y(men_men_n1196_));
  NA2        u1147(.A(men_men_n450_), .B(men_men_n53_), .Y(men_men_n1197_));
  NO2        u1148(.A(men_men_n1197_), .B(men_men_n938_), .Y(men_men_n1198_));
  NA2        u1149(.A(men_men_n1118_), .B(men_men_n470_), .Y(men_men_n1199_));
  NA2        u1150(.A(men_men_n56_), .B(men_men_n110_), .Y(men_men_n1200_));
  NA2        u1151(.A(men_men_n1200_), .B(x1), .Y(men_men_n1201_));
  NO2        u1152(.A(men_men_n1201_), .B(men_men_n260_), .Y(men_men_n1202_));
  NO2        u1153(.A(men_men_n322_), .B(x6), .Y(men_men_n1203_));
  OAI210     u1154(.A0(men_men_n251_), .A1(men_men_n979_), .B0(men_men_n956_), .Y(men_men_n1204_));
  AOI220     u1155(.A0(men_men_n1204_), .A1(men_men_n1203_), .B0(men_men_n1202_), .B1(men_men_n1199_), .Y(men_men_n1205_));
  NAi41      u1156(.An(men_men_n1198_), .B(men_men_n1205_), .C(men_men_n1196_), .D(men_men_n1194_), .Y(men_men_n1206_));
  AOI220     u1157(.A0(men_men_n1206_), .A1(men_men_n68_), .B0(men_men_n1192_), .B1(men_men_n1191_), .Y(men_men_n1207_));
  NA2        u1158(.A(men_men_n71_), .B(x3), .Y(men_men_n1208_));
  NA2        u1159(.A(men_men_n1208_), .B(men_men_n901_), .Y(men_men_n1209_));
  OAI220     u1160(.A0(men_men_n304_), .A1(men_men_n820_), .B0(men_men_n87_), .B1(men_men_n77_), .Y(men_men_n1210_));
  AOI210     u1161(.A0(men_men_n1121_), .A1(men_men_n617_), .B0(men_men_n979_), .Y(men_men_n1211_));
  OA210      u1162(.A0(men_men_n1210_), .A1(men_men_n1209_), .B0(men_men_n1211_), .Y(men_men_n1212_));
  NA2        u1163(.A(men_men_n619_), .B(men_men_n55_), .Y(men_men_n1213_));
  NA2        u1164(.A(x6), .B(men_men_n50_), .Y(men_men_n1214_));
  NA2        u1165(.A(men_men_n1214_), .B(men_men_n542_), .Y(men_men_n1215_));
  NO2        u1166(.A(men_men_n159_), .B(men_men_n128_), .Y(men_men_n1216_));
  AOI210     u1167(.A0(men_men_n1215_), .A1(men_men_n433_), .B0(men_men_n1216_), .Y(men_men_n1217_));
  NO2        u1168(.A(men_men_n1217_), .B(men_men_n872_), .Y(men_men_n1218_));
  OAI210     u1169(.A0(men_men_n1218_), .A1(men_men_n1212_), .B0(men_men_n1149_), .Y(men_men_n1219_));
  NAi21      u1170(.An(men_men_n84_), .B(men_men_n384_), .Y(men_men_n1220_));
  NO2        u1171(.A(men_men_n1220_), .B(men_men_n71_), .Y(men_men_n1221_));
  AOI210     u1172(.A0(men_men_n162_), .A1(x4), .B0(men_men_n174_), .Y(men_men_n1222_));
  NO2        u1173(.A(men_men_n1222_), .B(x0), .Y(men_men_n1223_));
  NO2        u1174(.A(men_men_n170_), .B(men_men_n295_), .Y(men_men_n1224_));
  OAI210     u1175(.A0(men_men_n1224_), .A1(men_men_n1223_), .B0(men_men_n1221_), .Y(men_men_n1225_));
  NA3        u1176(.A(men_men_n1155_), .B(men_men_n189_), .C(men_men_n71_), .Y(men_men_n1226_));
  NO2        u1177(.A(x4), .B(x0), .Y(men_men_n1227_));
  NO3        u1178(.A(men_men_n998_), .B(men_men_n248_), .C(men_men_n542_), .Y(men_men_n1228_));
  OAI210     u1179(.A0(men_men_n1228_), .A1(men_men_n199_), .B0(men_men_n1227_), .Y(men_men_n1229_));
  NA3        u1180(.A(men_men_n1229_), .B(men_men_n1226_), .C(men_men_n1225_), .Y(men_men_n1230_));
  NA2        u1181(.A(men_men_n250_), .B(men_men_n731_), .Y(men_men_n1231_));
  NO2        u1182(.A(men_men_n1231_), .B(men_men_n522_), .Y(men_men_n1232_));
  NA2        u1183(.A(men_men_n56_), .B(x0), .Y(men_men_n1233_));
  NO3        u1184(.A(men_men_n1233_), .B(men_men_n496_), .C(men_men_n81_), .Y(men_men_n1234_));
  OAI210     u1185(.A0(men_men_n1234_), .A1(men_men_n1232_), .B0(x2), .Y(men_men_n1235_));
  NO2        u1186(.A(men_men_n325_), .B(men_men_n384_), .Y(men_men_n1236_));
  NO2        u1187(.A(men_men_n689_), .B(x0), .Y(men_men_n1237_));
  OAI210     u1188(.A0(men_men_n1237_), .A1(men_men_n1236_), .B0(men_men_n333_), .Y(men_men_n1238_));
  NO2        u1189(.A(men_men_n789_), .B(x1), .Y(men_men_n1239_));
  AOI220     u1190(.A0(men_men_n1239_), .A1(men_men_n612_), .B0(men_men_n480_), .B1(men_men_n296_), .Y(men_men_n1240_));
  NA2        u1191(.A(men_men_n502_), .B(men_men_n50_), .Y(men_men_n1241_));
  AOI220     u1192(.A0(men_men_n1241_), .A1(men_men_n1185_), .B0(men_men_n980_), .B1(men_men_n101_), .Y(men_men_n1242_));
  NA4        u1193(.A(men_men_n1242_), .B(men_men_n1240_), .C(men_men_n1238_), .D(men_men_n1235_), .Y(men_men_n1243_));
  AOI220     u1194(.A0(men_men_n1243_), .A1(men_men_n129_), .B0(men_men_n1230_), .B1(men_men_n67_), .Y(men_men_n1244_));
  NA4        u1195(.A(men_men_n1244_), .B(men_men_n1219_), .C(men_men_n1207_), .D(men_men_n1190_), .Y(men14));
  NO2        u1196(.A(men_men_n372_), .B(men_men_n71_), .Y(men_men_n1246_));
  NO3        u1197(.A(x7), .B(x6), .C(x0), .Y(men_men_n1247_));
  OAI210     u1198(.A0(men_men_n1247_), .A1(men_men_n1246_), .B0(x8), .Y(men_men_n1248_));
  NA2        u1199(.A(men_men_n1132_), .B(men_men_n85_), .Y(men_men_n1249_));
  AOI210     u1200(.A0(men_men_n1249_), .A1(men_men_n1248_), .B0(men_men_n155_), .Y(men_men_n1250_));
  AOI220     u1201(.A0(men_men_n376_), .A1(men_men_n850_), .B0(men_men_n450_), .B1(men_men_n423_), .Y(men_men_n1251_));
  NA2        u1202(.A(men_men_n279_), .B(men_men_n975_), .Y(men_men_n1252_));
  OAI220     u1203(.A0(men_men_n1252_), .A1(men_men_n1251_), .B0(men_men_n468_), .B1(men_men_n804_), .Y(men_men_n1253_));
  OA210      u1204(.A0(men_men_n1253_), .A1(men_men_n1250_), .B0(x4), .Y(men_men_n1254_));
  NO2        u1205(.A(men_men_n139_), .B(men_men_n610_), .Y(men_men_n1255_));
  NA2        u1206(.A(x6), .B(x2), .Y(men_men_n1256_));
  NO2        u1207(.A(men_men_n628_), .B(men_men_n1256_), .Y(men_men_n1257_));
  OA210      u1208(.A0(men_men_n1255_), .A1(men_men_n212_), .B0(men_men_n1257_), .Y(men_men_n1258_));
  NO4        u1209(.A(men_men_n606_), .B(men_men_n377_), .C(men_men_n300_), .D(men_men_n116_), .Y(men_men_n1259_));
  OAI210     u1210(.A0(men_men_n1259_), .A1(men_men_n1258_), .B0(men_men_n59_), .Y(men_men_n1260_));
  NA2        u1211(.A(x6), .B(men_men_n108_), .Y(men_men_n1261_));
  NO2        u1212(.A(men_men_n666_), .B(men_men_n1261_), .Y(men_men_n1262_));
  NA2        u1213(.A(men_men_n1262_), .B(men_men_n925_), .Y(men_men_n1263_));
  AOI210     u1214(.A0(men_men_n1132_), .A1(men_men_n1012_), .B0(x1), .Y(men_men_n1264_));
  NO2        u1215(.A(men_men_n537_), .B(x5), .Y(men_men_n1265_));
  NA3        u1216(.A(men_men_n1265_), .B(men_men_n122_), .C(x0), .Y(men_men_n1266_));
  NA4        u1217(.A(men_men_n696_), .B(men_men_n926_), .C(men_men_n304_), .D(men_men_n68_), .Y(men_men_n1267_));
  AN4        u1218(.A(men_men_n1267_), .B(men_men_n1266_), .C(men_men_n1264_), .D(men_men_n1263_), .Y(men_men_n1268_));
  NO2        u1219(.A(men_men_n703_), .B(men_men_n1094_), .Y(men_men_n1269_));
  NO2        u1220(.A(men_men_n77_), .B(men_men_n58_), .Y(men_men_n1270_));
  OAI210     u1221(.A0(men_men_n1269_), .A1(men_men_n447_), .B0(men_men_n1270_), .Y(men_men_n1271_));
  AO210      u1222(.A0(men_men_n1246_), .A1(men_men_n1012_), .B0(men_men_n53_), .Y(men_men_n1272_));
  AOI210     u1223(.A0(men_men_n764_), .A1(men_men_n814_), .B0(men_men_n1272_), .Y(men_men_n1273_));
  AOI220     u1224(.A0(men_men_n1273_), .A1(men_men_n1271_), .B0(men_men_n1268_), .B1(men_men_n1260_), .Y(men_men_n1274_));
  NO2        u1225(.A(men_men_n678_), .B(men_men_n166_), .Y(men_men_n1275_));
  NO3        u1226(.A(men_men_n1275_), .B(men_men_n1274_), .C(men_men_n1254_), .Y(men_men_n1276_));
  NO2        u1227(.A(men_men_n322_), .B(x2), .Y(men_men_n1277_));
  XN2        u1228(.A(x4), .B(x1), .Y(men_men_n1278_));
  NO2        u1229(.A(men_men_n1278_), .B(men_men_n304_), .Y(men_men_n1279_));
  NOi21      u1230(.An(men_men_n1279_), .B(men_men_n411_), .Y(men_men_n1280_));
  NO2        u1231(.A(men_men_n340_), .B(men_men_n60_), .Y(men_men_n1281_));
  OAI210     u1232(.A0(men_men_n1281_), .A1(men_men_n1280_), .B0(men_men_n1277_), .Y(men_men_n1282_));
  NA2        u1233(.A(men_men_n690_), .B(men_men_n56_), .Y(men_men_n1283_));
  OAI220     u1234(.A0(men_men_n1283_), .A1(men_men_n156_), .B0(men_men_n190_), .B1(men_men_n71_), .Y(men_men_n1284_));
  NO2        u1235(.A(men_men_n216_), .B(men_men_n258_), .Y(men_men_n1285_));
  AOI220     u1236(.A0(men_men_n136_), .A1(men_men_n56_), .B0(men_men_n93_), .B1(x5), .Y(men_men_n1286_));
  NA2        u1237(.A(men_men_n1086_), .B(men_men_n309_), .Y(men_men_n1287_));
  NA2        u1238(.A(men_men_n250_), .B(men_men_n355_), .Y(men_men_n1288_));
  NA2        u1239(.A(men_men_n642_), .B(men_men_n1030_), .Y(men_men_n1289_));
  OAI220     u1240(.A0(men_men_n1289_), .A1(men_men_n1288_), .B0(men_men_n1287_), .B1(men_men_n1286_), .Y(men_men_n1290_));
  AOI210     u1241(.A0(men_men_n1285_), .A1(men_men_n1284_), .B0(men_men_n1290_), .Y(men_men_n1291_));
  AOI210     u1242(.A0(men_men_n1291_), .A1(men_men_n1282_), .B0(x7), .Y(men_men_n1292_));
  NO2        u1243(.A(men_men_n495_), .B(x6), .Y(men_men_n1293_));
  AOI210     u1244(.A0(men_men_n816_), .A1(men_men_n958_), .B0(men_men_n1293_), .Y(men_men_n1294_));
  OAI220     u1245(.A0(men_men_n1294_), .A1(men_men_n55_), .B0(men_men_n495_), .B1(men_men_n104_), .Y(men_men_n1295_));
  NA2        u1246(.A(men_men_n1295_), .B(men_men_n357_), .Y(men_men_n1296_));
  NA3        u1247(.A(men_men_n613_), .B(men_men_n1063_), .C(men_men_n70_), .Y(men_men_n1297_));
  NO4        u1248(.A(men_men_n1297_), .B(men_men_n1233_), .C(men_men_n120_), .D(men_men_n55_), .Y(men_men_n1298_));
  NO3        u1249(.A(men_men_n1056_), .B(men_men_n822_), .C(men_men_n485_), .Y(men_men_n1299_));
  NO3        u1250(.A(men_men_n751_), .B(men_men_n502_), .C(men_men_n54_), .Y(men_men_n1300_));
  NO4        u1251(.A(men_men_n1300_), .B(men_men_n1299_), .C(men_men_n1298_), .D(men_men_n1035_), .Y(men_men_n1301_));
  AOI210     u1252(.A0(men_men_n1301_), .A1(men_men_n1296_), .B0(men_men_n306_), .Y(men_men_n1302_));
  NA2        u1253(.A(men_men_n899_), .B(men_men_n53_), .Y(men_men_n1303_));
  OAI210     u1254(.A0(men_men_n245_), .A1(men_men_n118_), .B0(x2), .Y(men_men_n1304_));
  NA2        u1255(.A(men_men_n368_), .B(men_men_n56_), .Y(men_men_n1305_));
  OA220      u1256(.A0(men_men_n1305_), .A1(men_men_n1304_), .B0(men_men_n1303_), .B1(men_men_n376_), .Y(men_men_n1306_));
  NA3        u1257(.A(men_men_n1035_), .B(men_men_n736_), .C(men_men_n55_), .Y(men_men_n1307_));
  NA2        u1258(.A(men_men_n56_), .B(x2), .Y(men_men_n1308_));
  NO2        u1259(.A(men_men_n1308_), .B(men_men_n197_), .Y(men_men_n1309_));
  NA4        u1260(.A(men_men_n1309_), .B(men_men_n368_), .C(men_men_n258_), .D(men_men_n67_), .Y(men_men_n1310_));
  NA3        u1261(.A(men_men_n1239_), .B(men_men_n619_), .C(men_men_n633_), .Y(men_men_n1311_));
  AN3        u1262(.A(men_men_n1311_), .B(men_men_n1310_), .C(men_men_n1307_), .Y(men_men_n1312_));
  OAI210     u1263(.A0(men_men_n1306_), .A1(men_men_n317_), .B0(men_men_n1312_), .Y(men_men_n1313_));
  NO3        u1264(.A(men_men_n1313_), .B(men_men_n1302_), .C(men_men_n1292_), .Y(men_men_n1314_));
  OAI210     u1265(.A0(men_men_n1276_), .A1(x3), .B0(men_men_n1314_), .Y(men15));
  NA2        u1266(.A(men_men_n588_), .B(men_men_n59_), .Y(men_men_n1316_));
  NAi41      u1267(.An(x2), .B(x7), .C(x6), .D(x0), .Y(men_men_n1317_));
  AOI210     u1268(.A0(men_men_n1317_), .A1(men_men_n1316_), .B0(men_men_n53_), .Y(men_men_n1318_));
  NA3        u1269(.A(men_men_n57_), .B(x6), .C(men_men_n110_), .Y(men_men_n1319_));
  NO2        u1270(.A(men_men_n1319_), .B(men_men_n295_), .Y(men_men_n1320_));
  OAI210     u1271(.A0(men_men_n1320_), .A1(men_men_n1318_), .B0(men_men_n1155_), .Y(men_men_n1321_));
  NA2        u1272(.A(men_men_n112_), .B(men_men_n110_), .Y(men_men_n1322_));
  NA4        u1273(.A(men_men_n1322_), .B(men_men_n640_), .C(men_men_n310_), .D(x6), .Y(men_men_n1323_));
  AOI210     u1274(.A0(men_men_n730_), .A1(men_men_n76_), .B0(x3), .Y(men_men_n1324_));
  NA3        u1275(.A(men_men_n1324_), .B(men_men_n1323_), .C(men_men_n1321_), .Y(men_men_n1325_));
  AOI210     u1276(.A0(men_men_n1068_), .A1(men_men_n592_), .B0(men_men_n50_), .Y(men_men_n1326_));
  NO2        u1277(.A(men_men_n295_), .B(men_men_n110_), .Y(men_men_n1327_));
  NO2        u1278(.A(men_men_n237_), .B(x5), .Y(men_men_n1328_));
  NA2        u1279(.A(men_men_n1328_), .B(men_men_n1327_), .Y(men_men_n1329_));
  NA3        u1280(.A(men_men_n1239_), .B(men_men_n627_), .C(men_men_n1167_), .Y(men_men_n1330_));
  NA4        u1281(.A(men_men_n1330_), .B(men_men_n1329_), .C(men_men_n1326_), .D(men_men_n1266_), .Y(men_men_n1331_));
  NA2        u1282(.A(men_men_n334_), .B(men_men_n343_), .Y(men_men_n1332_));
  AOI210     u1283(.A0(men_men_n1201_), .A1(men_men_n58_), .B0(men_men_n1332_), .Y(men_men_n1333_));
  NA4        u1284(.A(men_men_n1201_), .B(men_men_n702_), .C(men_men_n1129_), .D(men_men_n384_), .Y(men_men_n1334_));
  NA2        u1285(.A(men_men_n592_), .B(men_men_n469_), .Y(men_men_n1335_));
  NO2        u1286(.A(men_men_n751_), .B(men_men_n53_), .Y(men_men_n1336_));
  NO2        u1287(.A(men_men_n777_), .B(men_men_n300_), .Y(men_men_n1337_));
  NA2        u1288(.A(men_men_n1337_), .B(men_men_n1336_), .Y(men_men_n1338_));
  NA3        u1289(.A(men_men_n1338_), .B(men_men_n1335_), .C(men_men_n1334_), .Y(men_men_n1339_));
  OAI210     u1290(.A0(men_men_n1339_), .A1(men_men_n1333_), .B0(men_men_n77_), .Y(men_men_n1340_));
  NA2        u1291(.A(men_men_n370_), .B(men_men_n705_), .Y(men_men_n1341_));
  NA2        u1292(.A(men_men_n573_), .B(men_men_n56_), .Y(men_men_n1342_));
  NA3        u1293(.A(men_men_n1342_), .B(men_men_n343_), .C(men_men_n112_), .Y(men_men_n1343_));
  AOI210     u1294(.A0(men_men_n1343_), .A1(men_men_n1341_), .B0(men_men_n502_), .Y(men_men_n1344_));
  NO3        u1295(.A(men_men_n802_), .B(men_men_n624_), .C(men_men_n198_), .Y(men_men_n1345_));
  OAI210     u1296(.A0(men_men_n1345_), .A1(men_men_n1344_), .B0(men_men_n495_), .Y(men_men_n1346_));
  NO2        u1297(.A(men_men_n872_), .B(men_men_n50_), .Y(men_men_n1347_));
  NO2        u1298(.A(men_men_n247_), .B(men_men_n64_), .Y(men_men_n1348_));
  OA210      u1299(.A0(men_men_n1348_), .A1(men_men_n1347_), .B0(men_men_n411_), .Y(men_men_n1349_));
  NA2        u1300(.A(men_men_n57_), .B(x3), .Y(men_men_n1350_));
  AOI210     u1301(.A0(men_men_n981_), .A1(men_men_n1350_), .B0(men_men_n684_), .Y(men_men_n1351_));
  OAI210     u1302(.A0(men_men_n1351_), .A1(men_men_n1349_), .B0(men_men_n1020_), .Y(men_men_n1352_));
  NA2        u1303(.A(men_men_n1309_), .B(men_men_n68_), .Y(men_men_n1353_));
  NO2        u1304(.A(men_men_n1256_), .B(x0), .Y(men_men_n1354_));
  AOI210     u1305(.A0(men_men_n1354_), .A1(men_men_n607_), .B0(x8), .Y(men_men_n1355_));
  NO2        u1306(.A(men_men_n432_), .B(men_men_n81_), .Y(men_men_n1356_));
  NO2        u1307(.A(men_men_n932_), .B(men_men_n71_), .Y(men_men_n1357_));
  NA2        u1308(.A(men_men_n1357_), .B(men_men_n1356_), .Y(men_men_n1358_));
  NO2        u1309(.A(men_men_n979_), .B(x6), .Y(men_men_n1359_));
  NA4        u1310(.A(men_men_n1359_), .B(men_men_n597_), .C(men_men_n157_), .D(men_men_n415_), .Y(men_men_n1360_));
  AN4        u1311(.A(men_men_n1360_), .B(men_men_n1358_), .C(men_men_n1355_), .D(men_men_n1353_), .Y(men_men_n1361_));
  NA4        u1312(.A(men_men_n1361_), .B(men_men_n1352_), .C(men_men_n1346_), .D(men_men_n1340_), .Y(men_men_n1362_));
  NA2        u1313(.A(men_men_n163_), .B(men_men_n736_), .Y(men_men_n1363_));
  NO2        u1314(.A(men_men_n652_), .B(x2), .Y(men_men_n1364_));
  OAI210     u1315(.A0(men_men_n68_), .A1(men_men_n53_), .B0(men_men_n142_), .Y(men_men_n1365_));
  OAI210     u1316(.A0(men_men_n1364_), .A1(men_men_n85_), .B0(men_men_n1365_), .Y(men_men_n1366_));
  AOI210     u1317(.A0(men_men_n1366_), .A1(men_men_n1363_), .B0(men_men_n322_), .Y(men_men_n1367_));
  NO3        u1318(.A(men_men_n1319_), .B(men_men_n266_), .C(men_men_n247_), .Y(men_men_n1368_));
  NA3        u1319(.A(men_men_n57_), .B(x1), .C(x0), .Y(men_men_n1369_));
  NA3        u1320(.A(men_men_n71_), .B(x5), .C(x2), .Y(men_men_n1370_));
  NA4        u1321(.A(x7), .B(x3), .C(men_men_n53_), .D(x0), .Y(men_men_n1371_));
  OAI220     u1322(.A0(men_men_n1371_), .A1(x6), .B0(men_men_n1370_), .B1(men_men_n1369_), .Y(men_men_n1372_));
  NO2        u1323(.A(men_men_n1372_), .B(men_men_n1368_), .Y(men_men_n1373_));
  NAi21      u1324(.An(men_men_n116_), .B(men_men_n745_), .Y(men_men_n1374_));
  NA4        u1325(.A(men_men_n1374_), .B(men_men_n320_), .C(men_men_n290_), .D(men_men_n627_), .Y(men_men_n1375_));
  OAI220     u1326(.A0(men_men_n325_), .A1(x7), .B0(men_men_n128_), .B1(men_men_n71_), .Y(men_men_n1376_));
  NA3        u1327(.A(men_men_n1376_), .B(men_men_n789_), .C(men_men_n1097_), .Y(men_men_n1377_));
  NA2        u1328(.A(men_men_n82_), .B(men_men_n50_), .Y(men_men_n1378_));
  AO210      u1329(.A0(men_men_n1378_), .A1(men_men_n315_), .B0(men_men_n155_), .Y(men_men_n1379_));
  NA4        u1330(.A(men_men_n1379_), .B(men_men_n1377_), .C(men_men_n1375_), .D(men_men_n1373_), .Y(men_men_n1380_));
  OAI210     u1331(.A0(men_men_n1380_), .A1(men_men_n1367_), .B0(men_men_n56_), .Y(men_men_n1381_));
  AOI210     u1332(.A0(men_men_n692_), .A1(x4), .B0(men_men_n958_), .Y(men_men_n1382_));
  OAI220     u1333(.A0(men_men_n1382_), .A1(men_men_n301_), .B0(men_men_n1024_), .B1(men_men_n946_), .Y(men_men_n1383_));
  NA2        u1334(.A(men_men_n833_), .B(men_men_n408_), .Y(men_men_n1384_));
  OAI210     u1335(.A0(men_men_n1356_), .A1(men_men_n1348_), .B0(men_men_n291_), .Y(men_men_n1385_));
  OAI210     u1336(.A0(men_men_n1384_), .A1(men_men_n845_), .B0(men_men_n1385_), .Y(men_men_n1386_));
  OAI210     u1337(.A0(men_men_n1386_), .A1(men_men_n1383_), .B0(x6), .Y(men_men_n1387_));
  NO2        u1338(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n1388_));
  NO2        u1339(.A(x7), .B(x5), .Y(men_men_n1389_));
  AOI220     u1340(.A0(men_men_n854_), .A1(men_men_n1388_), .B0(men_men_n541_), .B1(men_men_n1389_), .Y(men_men_n1390_));
  NA2        u1341(.A(men_men_n761_), .B(men_men_n291_), .Y(men_men_n1391_));
  NA3        u1342(.A(men_men_n619_), .B(men_men_n293_), .C(men_men_n242_), .Y(men_men_n1392_));
  NA2        u1343(.A(men_men_n1392_), .B(men_men_n1390_), .Y(men_men_n1393_));
  NA2        u1344(.A(men_men_n1393_), .B(men_men_n426_), .Y(men_men_n1394_));
  AOI210     u1345(.A0(men_men_n380_), .A1(men_men_n341_), .B0(men_men_n55_), .Y(men_men_n1395_));
  NA4        u1346(.A(men_men_n1395_), .B(men_men_n1394_), .C(men_men_n1387_), .D(men_men_n1381_), .Y(men_men_n1396_));
  AO220      u1347(.A0(men_men_n1396_), .A1(men_men_n1362_), .B0(men_men_n1331_), .B1(men_men_n1325_), .Y(men16));
  NO2        u1348(.A(x4), .B(men_men_n59_), .Y(men_men_n1398_));
  NA2        u1349(.A(men_men_n665_), .B(men_men_n538_), .Y(men_men_n1399_));
  NA3        u1350(.A(men_men_n231_), .B(men_men_n433_), .C(men_men_n958_), .Y(men_men_n1400_));
  NA2        u1351(.A(men_men_n131_), .B(men_men_n207_), .Y(men_men_n1401_));
  AOI210     u1352(.A0(men_men_n1400_), .A1(men_men_n1399_), .B0(men_men_n1401_), .Y(men_men_n1402_));
  NO3        u1353(.A(x8), .B(x6), .C(men_men_n50_), .Y(men_men_n1403_));
  NO2        u1354(.A(men_men_n734_), .B(men_men_n185_), .Y(men_men_n1404_));
  OAI210     u1355(.A0(men_men_n1403_), .A1(men_men_n239_), .B0(men_men_n1404_), .Y(men_men_n1405_));
  NO2        u1356(.A(men_men_n159_), .B(x5), .Y(men_men_n1406_));
  NA2        u1357(.A(men_men_n1406_), .B(men_men_n1364_), .Y(men_men_n1407_));
  NA3        u1358(.A(men_men_n582_), .B(men_men_n540_), .C(men_men_n479_), .Y(men_men_n1408_));
  NA3        u1359(.A(men_men_n1408_), .B(men_men_n1407_), .C(men_men_n1405_), .Y(men_men_n1409_));
  OAI210     u1360(.A0(men_men_n1409_), .A1(men_men_n1402_), .B0(men_men_n1398_), .Y(men_men_n1410_));
  OAI210     u1361(.A0(men_men_n1277_), .A1(men_men_n925_), .B0(men_men_n423_), .Y(men_men_n1411_));
  NO2        u1362(.A(men_men_n322_), .B(x7), .Y(men_men_n1412_));
  NA2        u1363(.A(men_men_n1412_), .B(x0), .Y(men_men_n1413_));
  AOI210     u1364(.A0(men_men_n1413_), .A1(men_men_n1411_), .B0(men_men_n641_), .Y(men_men_n1414_));
  NA2        u1365(.A(men_men_n1077_), .B(men_men_n198_), .Y(men_men_n1415_));
  NA2        u1366(.A(men_men_n55_), .B(men_men_n108_), .Y(men_men_n1416_));
  NA2        u1367(.A(men_men_n1416_), .B(men_men_n686_), .Y(men_men_n1417_));
  NA2        u1368(.A(men_men_n379_), .B(men_men_n1081_), .Y(men_men_n1418_));
  OA220      u1369(.A0(men_men_n1418_), .A1(men_men_n1417_), .B0(men_men_n1415_), .B1(men_men_n635_), .Y(men_men_n1419_));
  OAI210     u1370(.A0(men_men_n1419_), .A1(men_men_n656_), .B0(men_men_n500_), .Y(men_men_n1420_));
  INV        u1371(.A(men_men_n1020_), .Y(men_men_n1421_));
  NO2        u1372(.A(men_men_n1421_), .B(men_men_n62_), .Y(men_men_n1422_));
  AOI220     u1373(.A0(men_men_n1422_), .A1(men_men_n270_), .B0(men_men_n1262_), .B1(men_men_n126_), .Y(men_men_n1423_));
  NA2        u1374(.A(men_men_n640_), .B(men_men_n364_), .Y(men_men_n1424_));
  NA3        u1375(.A(men_men_n466_), .B(men_men_n589_), .C(men_men_n192_), .Y(men_men_n1425_));
  OAI220     u1376(.A0(men_men_n1425_), .A1(men_men_n1424_), .B0(men_men_n1423_), .B1(men_men_n311_), .Y(men_men_n1426_));
  NO3        u1377(.A(men_men_n1426_), .B(men_men_n1420_), .C(men_men_n1414_), .Y(men_men_n1427_));
  NO3        u1378(.A(x6), .B(x4), .C(x3), .Y(men_men_n1428_));
  NA2        u1379(.A(men_men_n1428_), .B(men_men_n537_), .Y(men_men_n1429_));
  NA4        u1380(.A(men_men_n710_), .B(men_men_n185_), .C(men_men_n58_), .D(x6), .Y(men_men_n1430_));
  AOI210     u1381(.A0(men_men_n1430_), .A1(men_men_n1429_), .B0(men_men_n54_), .Y(men_men_n1431_));
  NO2        u1382(.A(men_men_n722_), .B(x3), .Y(men_men_n1432_));
  NO3        u1383(.A(men_men_n502_), .B(men_men_n220_), .C(men_men_n75_), .Y(men_men_n1433_));
  NO2        u1384(.A(men_men_n761_), .B(men_men_n514_), .Y(men_men_n1434_));
  NO3        u1385(.A(men_men_n1434_), .B(men_men_n260_), .C(men_men_n154_), .Y(men_men_n1435_));
  NO3        u1386(.A(men_men_n1435_), .B(men_men_n1433_), .C(men_men_n1431_), .Y(men_men_n1436_));
  NA2        u1387(.A(men_men_n409_), .B(men_men_n958_), .Y(men_men_n1437_));
  NA4        u1388(.A(men_men_n485_), .B(men_men_n372_), .C(men_men_n222_), .D(x6), .Y(men_men_n1438_));
  OAI210     u1389(.A0(men_men_n722_), .A1(men_men_n1437_), .B0(men_men_n1438_), .Y(men_men_n1439_));
  NA2        u1390(.A(men_men_n908_), .B(men_men_n1308_), .Y(men_men_n1440_));
  NA2        u1391(.A(men_men_n731_), .B(x7), .Y(men_men_n1441_));
  OAI210     u1392(.A0(men_men_n1441_), .A1(men_men_n391_), .B0(men_men_n1440_), .Y(men_men_n1442_));
  NA2        u1393(.A(men_men_n277_), .B(x2), .Y(men_men_n1443_));
  NO3        u1394(.A(men_men_n1443_), .B(men_men_n597_), .C(men_men_n72_), .Y(men_men_n1444_));
  OA210      u1395(.A0(men_men_n1261_), .A1(men_men_n58_), .B0(men_men_n778_), .Y(men_men_n1445_));
  AOI210     u1396(.A0(men_men_n582_), .A1(men_men_n50_), .B0(men_men_n592_), .Y(men_men_n1446_));
  OAI210     u1397(.A0(men_men_n926_), .A1(men_men_n945_), .B0(men_men_n386_), .Y(men_men_n1447_));
  OAI220     u1398(.A0(men_men_n1447_), .A1(men_men_n1446_), .B0(men_men_n1445_), .B1(men_men_n190_), .Y(men_men_n1448_));
  NO4        u1399(.A(men_men_n1448_), .B(men_men_n1444_), .C(men_men_n1442_), .D(men_men_n1439_), .Y(men_men_n1449_));
  OA220      u1400(.A0(men_men_n1449_), .A1(men_men_n446_), .B0(men_men_n1436_), .B1(men_men_n205_), .Y(men_men_n1450_));
  NO2        u1401(.A(men_men_n921_), .B(men_men_n55_), .Y(men_men_n1451_));
  NA2        u1402(.A(men_men_n420_), .B(men_men_n804_), .Y(men_men_n1452_));
  NO2        u1403(.A(men_men_n1452_), .B(men_men_n1451_), .Y(men_men_n1453_));
  NO3        u1404(.A(men_men_n959_), .B(men_men_n334_), .C(x8), .Y(men_men_n1454_));
  OAI210     u1405(.A0(men_men_n1454_), .A1(men_men_n1453_), .B0(x6), .Y(men_men_n1455_));
  NO2        u1406(.A(men_men_n1092_), .B(men_men_n1055_), .Y(men_men_n1456_));
  NA2        u1407(.A(men_men_n190_), .B(x7), .Y(men_men_n1457_));
  OAI220     u1408(.A0(men_men_n1457_), .A1(men_men_n1456_), .B0(men_men_n763_), .B1(men_men_n87_), .Y(men_men_n1458_));
  NA2        u1409(.A(men_men_n1458_), .B(men_men_n926_), .Y(men_men_n1459_));
  NA2        u1410(.A(men_men_n874_), .B(men_men_n71_), .Y(men_men_n1460_));
  OAI210     u1411(.A0(men_men_n1460_), .A1(men_men_n157_), .B0(men_men_n1009_), .Y(men_men_n1461_));
  AOI210     u1412(.A0(men_men_n502_), .A1(men_men_n57_), .B0(men_men_n635_), .Y(men_men_n1462_));
  NA2        u1413(.A(men_men_n1462_), .B(men_men_n1461_), .Y(men_men_n1463_));
  NA3        u1414(.A(men_men_n1463_), .B(men_men_n1459_), .C(men_men_n1455_), .Y(men_men_n1464_));
  NO2        u1415(.A(men_men_n642_), .B(x6), .Y(men_men_n1465_));
  OAI210     u1416(.A0(men_men_n386_), .A1(men_men_n84_), .B0(men_men_n384_), .Y(men_men_n1466_));
  OA210      u1417(.A0(men_men_n1466_), .A1(men_men_n1465_), .B0(men_men_n129_), .Y(men_men_n1467_));
  NO3        u1418(.A(men_men_n448_), .B(men_men_n389_), .C(x7), .Y(men_men_n1468_));
  NO3        u1419(.A(men_men_n159_), .B(men_men_n75_), .C(x2), .Y(men_men_n1469_));
  NO3        u1420(.A(men_men_n1469_), .B(men_men_n1468_), .C(men_men_n1467_), .Y(men_men_n1470_));
  NO2        u1421(.A(men_men_n57_), .B(men_men_n108_), .Y(men_men_n1471_));
  AOI220     u1422(.A0(men_men_n763_), .A1(men_men_n774_), .B0(men_men_n517_), .B1(men_men_n281_), .Y(men_men_n1472_));
  NO2        u1423(.A(men_men_n1472_), .B(men_men_n1308_), .Y(men_men_n1473_));
  NO3        u1424(.A(men_men_n537_), .B(men_men_n172_), .C(men_men_n1055_), .Y(men_men_n1474_));
  NA2        u1425(.A(men_men_n945_), .B(x4), .Y(men_men_n1475_));
  OAI220     u1426(.A0(men_men_n1475_), .A1(men_men_n691_), .B0(men_men_n650_), .B1(men_men_n613_), .Y(men_men_n1476_));
  NO3        u1427(.A(men_men_n1476_), .B(men_men_n1474_), .C(men_men_n1473_), .Y(men_men_n1477_));
  OAI210     u1428(.A0(men_men_n1470_), .A1(x5), .B0(men_men_n1477_), .Y(men_men_n1478_));
  AOI220     u1429(.A0(men_men_n1478_), .A1(men_men_n99_), .B0(men_men_n1464_), .B1(men_men_n341_), .Y(men_men_n1479_));
  NA4        u1430(.A(men_men_n1479_), .B(men_men_n1450_), .C(men_men_n1427_), .D(men_men_n1410_), .Y(men17));
  NO4        u1431(.A(men_men_n604_), .B(men_men_n704_), .C(men_men_n102_), .D(men_men_n101_), .Y(men_men_n1481_));
  NO2        u1432(.A(men_men_n125_), .B(men_men_n1167_), .Y(men_men_n1482_));
  AOI220     u1433(.A0(men_men_n1482_), .A1(men_men_n716_), .B0(men_men_n1481_), .B1(men_men_n508_), .Y(men_men_n1483_));
  NA2        u1434(.A(men_men_n163_), .B(men_men_n78_), .Y(men_men_n1484_));
  NOi21      u1435(.An(men_men_n384_), .B(men_men_n84_), .Y(men_men_n1485_));
  OAI210     u1436(.A0(men_men_n627_), .A1(men_men_n55_), .B0(men_men_n1485_), .Y(men_men_n1486_));
  NA2        u1437(.A(men_men_n1220_), .B(men_men_n1015_), .Y(men_men_n1487_));
  NA4        u1438(.A(men_men_n1487_), .B(men_men_n1486_), .C(men_men_n734_), .D(men_men_n57_), .Y(men_men_n1488_));
  OAI210     u1439(.A0(men_men_n710_), .A1(x8), .B0(men_men_n1308_), .Y(men_men_n1489_));
  NA3        u1440(.A(men_men_n1489_), .B(men_men_n1246_), .C(men_men_n402_), .Y(men_men_n1490_));
  NA3        u1441(.A(men_men_n396_), .B(men_men_n270_), .C(men_men_n588_), .Y(men_men_n1491_));
  OA210      u1442(.A0(men_men_n1319_), .A1(men_men_n1160_), .B0(men_men_n753_), .Y(men_men_n1492_));
  NA4        u1443(.A(men_men_n1492_), .B(men_men_n1491_), .C(men_men_n1490_), .D(men_men_n1488_), .Y(men_men_n1493_));
  NA3        u1444(.A(men_men_n162_), .B(men_men_n633_), .C(men_men_n1055_), .Y(men_men_n1494_));
  AOI210     u1445(.A0(men_men_n1083_), .A1(men_men_n307_), .B0(men_men_n59_), .Y(men_men_n1495_));
  NA2        u1446(.A(men_men_n1495_), .B(men_men_n1494_), .Y(men_men_n1496_));
  AOI210     u1447(.A0(men_men_n1493_), .A1(x1), .B0(men_men_n1496_), .Y(men_men_n1497_));
  NO2        u1448(.A(men_men_n984_), .B(men_men_n502_), .Y(men_men_n1498_));
  OAI210     u1449(.A0(men_men_n1498_), .A1(men_men_n1067_), .B0(men_men_n610_), .Y(men_men_n1499_));
  NO3        u1450(.A(men_men_n635_), .B(men_men_n557_), .C(men_men_n528_), .Y(men_men_n1500_));
  OAI210     u1451(.A0(men_men_n1500_), .A1(men_men_n907_), .B0(men_men_n1432_), .Y(men_men_n1501_));
  AOI210     u1452(.A0(men_men_n1501_), .A1(men_men_n1499_), .B0(x8), .Y(men_men_n1502_));
  NA3        u1453(.A(men_men_n635_), .B(men_men_n273_), .C(men_men_n122_), .Y(men_men_n1503_));
  NO2        u1454(.A(men_men_n142_), .B(men_men_n140_), .Y(men_men_n1504_));
  NO3        u1455(.A(men_men_n902_), .B(men_men_n774_), .C(men_men_n704_), .Y(men_men_n1505_));
  AOI210     u1456(.A0(men_men_n1505_), .A1(men_men_n1504_), .B0(x0), .Y(men_men_n1506_));
  OAI210     u1457(.A0(men_men_n1503_), .A1(men_men_n249_), .B0(men_men_n1506_), .Y(men_men_n1507_));
  NO2        u1458(.A(men_men_n1507_), .B(men_men_n1502_), .Y(men_men_n1508_));
  OAI220     u1459(.A0(men_men_n1508_), .A1(men_men_n1497_), .B0(men_men_n1484_), .B1(men_men_n1483_), .Y(men18));
  AOI210     u1460(.A0(x8), .A1(x0), .B0(x5), .Y(men_men_n1510_));
  NOi31      u1461(.An(men_men_n307_), .B(men_men_n1510_), .C(men_men_n1054_), .Y(men_men_n1511_));
  NA2        u1462(.A(men_men_n604_), .B(men_men_n59_), .Y(men_men_n1512_));
  AOI210     u1463(.A0(men_men_n1415_), .A1(men_men_n352_), .B0(men_men_n1512_), .Y(men_men_n1513_));
  NO2        u1464(.A(men_men_n620_), .B(men_men_n775_), .Y(men_men_n1514_));
  NO4        u1465(.A(men_men_n256_), .B(men_men_n814_), .C(men_men_n153_), .D(men_men_n70_), .Y(men_men_n1515_));
  NO4        u1466(.A(men_men_n1515_), .B(men_men_n1514_), .C(men_men_n1513_), .D(men_men_n1511_), .Y(men_men_n1516_));
  NA3        u1467(.A(men_men_n523_), .B(men_men_n216_), .C(x0), .Y(men_men_n1517_));
  NAi21      u1468(.An(men_men_n390_), .B(men_men_n1517_), .Y(men_men_n1518_));
  NO2        u1469(.A(men_men_n892_), .B(x5), .Y(men_men_n1519_));
  AOI210     u1470(.A0(men_men_n1145_), .A1(x5), .B0(men_men_n1519_), .Y(men_men_n1520_));
  OA220      u1471(.A0(men_men_n523_), .A1(men_men_n334_), .B0(men_men_n402_), .B1(x5), .Y(men_men_n1521_));
  OAI220     u1472(.A0(men_men_n1521_), .A1(men_men_n295_), .B0(men_men_n1520_), .B1(men_men_n214_), .Y(men_men_n1522_));
  AOI210     u1473(.A0(men_men_n1518_), .A1(men_men_n293_), .B0(men_men_n1522_), .Y(men_men_n1523_));
  AOI210     u1474(.A0(men_men_n1523_), .A1(men_men_n1516_), .B0(x6), .Y(men_men_n1524_));
  NA3        u1475(.A(men_men_n527_), .B(men_men_n423_), .C(x2), .Y(men_men_n1525_));
  NA3        u1476(.A(men_men_n1054_), .B(men_men_n51_), .C(men_men_n57_), .Y(men_men_n1526_));
  AOI210     u1477(.A0(men_men_n1526_), .A1(men_men_n1525_), .B0(men_men_n789_), .Y(men_men_n1527_));
  AOI210     u1478(.A0(men_men_n427_), .A1(men_men_n136_), .B0(men_men_n787_), .Y(men_men_n1528_));
  NA2        u1479(.A(men_men_n270_), .B(x6), .Y(men_men_n1529_));
  OAI210     u1480(.A0(men_men_n178_), .A1(men_men_n110_), .B0(men_men_n1151_), .Y(men_men_n1530_));
  OAI220     u1481(.A0(men_men_n1530_), .A1(men_men_n1529_), .B0(men_men_n1528_), .B1(men_men_n745_), .Y(men_men_n1531_));
  OAI210     u1482(.A0(men_men_n1531_), .A1(men_men_n1527_), .B0(men_men_n53_), .Y(men_men_n1532_));
  NO2        u1483(.A(men_men_n690_), .B(men_men_n263_), .Y(men_men_n1533_));
  NO2        u1484(.A(men_men_n266_), .B(x3), .Y(men_men_n1534_));
  NO3        u1485(.A(men_men_n437_), .B(men_men_n604_), .C(men_men_n838_), .Y(men_men_n1535_));
  OAI210     u1486(.A0(men_men_n1535_), .A1(men_men_n1533_), .B0(men_men_n1534_), .Y(men_men_n1536_));
  AOI210     u1487(.A0(men_men_n1154_), .A1(men_men_n619_), .B0(x4), .Y(men_men_n1537_));
  OAI210     u1488(.A0(men_men_n557_), .A1(men_men_n604_), .B0(men_men_n59_), .Y(men_men_n1538_));
  OAI210     u1489(.A0(men_men_n627_), .A1(men_men_n652_), .B0(men_men_n1538_), .Y(men_men_n1539_));
  AO220      u1490(.A0(men_men_n1265_), .A1(men_men_n734_), .B0(men_men_n558_), .B1(men_men_n357_), .Y(men_men_n1540_));
  AOI220     u1491(.A0(men_men_n1540_), .A1(x1), .B0(men_men_n1539_), .B1(men_men_n160_), .Y(men_men_n1541_));
  NA4        u1492(.A(men_men_n1541_), .B(men_men_n1537_), .C(men_men_n1536_), .D(men_men_n1532_), .Y(men_men_n1542_));
  NO3        u1493(.A(men_men_n1074_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n1543_));
  OAI210     u1494(.A0(men_men_n1543_), .A1(men_men_n657_), .B0(men_men_n108_), .Y(men_men_n1544_));
  AOI210     u1495(.A0(men_men_n1544_), .A1(men_men_n563_), .B0(men_men_n789_), .Y(men_men_n1545_));
  NA3        u1496(.A(men_men_n1213_), .B(men_men_n190_), .C(men_men_n139_), .Y(men_men_n1546_));
  NA3        u1497(.A(men_men_n1077_), .B(men_men_n777_), .C(men_men_n345_), .Y(men_men_n1547_));
  NA2        u1498(.A(men_men_n170_), .B(men_men_n774_), .Y(men_men_n1548_));
  OAI210     u1499(.A0(men_men_n1548_), .A1(men_men_n1322_), .B0(men_men_n1547_), .Y(men_men_n1549_));
  AOI210     u1500(.A0(men_men_n1546_), .A1(men_men_n177_), .B0(men_men_n1549_), .Y(men_men_n1550_));
  OAI210     u1501(.A0(men_men_n1550_), .A1(men_men_n546_), .B0(x4), .Y(men_men_n1551_));
  OAI220     u1502(.A0(men_men_n1551_), .A1(men_men_n1545_), .B0(men_men_n1542_), .B1(men_men_n1524_), .Y(men_men_n1552_));
  NO2        u1503(.A(men_men_n145_), .B(men_men_n123_), .Y(men_men_n1553_));
  NO2        u1504(.A(men_men_n190_), .B(men_men_n804_), .Y(men_men_n1554_));
  AOI210     u1505(.A0(men_men_n605_), .A1(men_men_n514_), .B0(men_men_n1554_), .Y(men_men_n1555_));
  NO2        u1506(.A(men_men_n1555_), .B(x6), .Y(men_men_n1556_));
  NO2        u1507(.A(men_men_n389_), .B(men_men_n255_), .Y(men_men_n1557_));
  NO2        u1508(.A(men_men_n129_), .B(men_men_n736_), .Y(men_men_n1558_));
  NO2        u1509(.A(men_men_n959_), .B(men_men_n588_), .Y(men_men_n1559_));
  AO220      u1510(.A0(men_men_n1559_), .A1(men_men_n1558_), .B0(men_men_n1557_), .B1(men_men_n125_), .Y(men_men_n1560_));
  NO3        u1511(.A(men_men_n1560_), .B(men_men_n1556_), .C(men_men_n1553_), .Y(men_men_n1561_));
  NA2        u1512(.A(men_men_n1074_), .B(x3), .Y(men_men_n1562_));
  NA2        u1513(.A(men_men_n1359_), .B(men_men_n131_), .Y(men_men_n1563_));
  OAI220     u1514(.A0(men_men_n1563_), .A1(men_men_n1562_), .B0(men_men_n1561_), .B1(x3), .Y(men_men_n1564_));
  NO3        u1515(.A(men_men_n1005_), .B(men_men_n690_), .C(men_men_n329_), .Y(men_men_n1565_));
  AO210      u1516(.A0(men_men_n1034_), .A1(men_men_n300_), .B0(men_men_n1565_), .Y(men_men_n1566_));
  AOI220     u1517(.A0(men_men_n1566_), .A1(x8), .B0(men_men_n1359_), .B1(men_men_n438_), .Y(men_men_n1567_));
  NA2        u1518(.A(men_men_n749_), .B(men_men_n321_), .Y(men_men_n1568_));
  NO4        u1519(.A(men_men_n370_), .B(men_men_n203_), .C(men_men_n340_), .D(x2), .Y(men_men_n1569_));
  NA2        u1520(.A(men_men_n1416_), .B(men_men_n110_), .Y(men_men_n1570_));
  NO3        u1521(.A(men_men_n1214_), .B(men_men_n998_), .C(men_men_n1151_), .Y(men_men_n1571_));
  AOI210     u1522(.A0(men_men_n1571_), .A1(men_men_n1570_), .B0(men_men_n1569_), .Y(men_men_n1572_));
  OA220      u1523(.A0(men_men_n1572_), .A1(men_men_n959_), .B0(men_men_n1568_), .B1(men_men_n572_), .Y(men_men_n1573_));
  OAI210     u1524(.A0(men_men_n1567_), .A1(men_men_n412_), .B0(men_men_n1573_), .Y(men_men_n1574_));
  AOI210     u1525(.A0(men_men_n1564_), .A1(men_men_n136_), .B0(men_men_n1574_), .Y(men_men_n1575_));
  NA2        u1526(.A(men_men_n1575_), .B(men_men_n1552_), .Y(men19));
  NO2        u1527(.A(men_men_n1460_), .B(men_men_n259_), .Y(men_men_n1577_));
  NA2        u1528(.A(men_men_n652_), .B(x3), .Y(men_men_n1578_));
  OAI210     u1529(.A0(men_men_n153_), .A1(men_men_n109_), .B0(men_men_n81_), .Y(men_men_n1579_));
  NA3        u1530(.A(men_men_n1579_), .B(men_men_n1578_), .C(men_men_n242_), .Y(men_men_n1580_));
  NO2        u1531(.A(men_men_n1317_), .B(men_men_n170_), .Y(men_men_n1581_));
  AOI210     u1532(.A0(men_men_n1481_), .A1(men_men_n355_), .B0(men_men_n1581_), .Y(men_men_n1582_));
  AOI210     u1533(.A0(men_men_n1582_), .A1(men_men_n1580_), .B0(men_men_n56_), .Y(men_men_n1583_));
  NO2        u1534(.A(men_men_n863_), .B(men_men_n1227_), .Y(men_men_n1584_));
  OAI210     u1535(.A0(men_men_n1583_), .A1(men_men_n1577_), .B0(men_men_n1584_), .Y(men_men_n1585_));
  NOi21      u1536(.An(men_men_n614_), .B(men_men_n656_), .Y(men_men_n1586_));
  AOI210     u1537(.A0(men_men_n355_), .A1(x6), .B0(men_men_n122_), .Y(men_men_n1587_));
  NO3        u1538(.A(men_men_n1587_), .B(men_men_n758_), .C(men_men_n126_), .Y(men_men_n1588_));
  NA2        u1539(.A(men_men_n1208_), .B(men_men_n123_), .Y(men_men_n1589_));
  NO4        u1540(.A(men_men_n1589_), .B(men_men_n1005_), .C(men_men_n892_), .D(men_men_n77_), .Y(men_men_n1590_));
  NO3        u1541(.A(men_men_n1590_), .B(men_men_n1588_), .C(men_men_n1031_), .Y(men_men_n1591_));
  NO2        u1542(.A(men_men_n546_), .B(men_men_n623_), .Y(men_men_n1592_));
  NA2        u1543(.A(men_men_n1261_), .B(men_men_n50_), .Y(men_men_n1593_));
  NO3        u1544(.A(men_men_n521_), .B(men_men_n309_), .C(men_men_n64_), .Y(men_men_n1594_));
  AOI220     u1545(.A0(men_men_n1594_), .A1(men_men_n1593_), .B0(men_men_n1592_), .B1(men_men_n777_), .Y(men_men_n1595_));
  OAI210     u1546(.A0(men_men_n1591_), .A1(men_men_n57_), .B0(men_men_n1595_), .Y(men_men_n1596_));
  AOI210     u1547(.A0(men_men_n1596_), .A1(men_men_n774_), .B0(men_men_n1586_), .Y(men_men_n1597_));
  AOI210     u1548(.A0(men_men_n824_), .A1(men_men_n736_), .B0(men_men_n764_), .Y(men_men_n1598_));
  NO2        u1549(.A(men_men_n1598_), .B(x4), .Y(men_men_n1599_));
  NA3        u1550(.A(men_men_n734_), .B(men_men_n258_), .C(x7), .Y(men_men_n1600_));
  AOI220     u1551(.A0(men_men_n1412_), .A1(men_men_n789_), .B0(men_men_n704_), .B1(men_men_n1167_), .Y(men_men_n1601_));
  AOI210     u1552(.A0(men_men_n1601_), .A1(men_men_n1600_), .B0(men_men_n506_), .Y(men_men_n1602_));
  OAI210     u1553(.A0(men_men_n1602_), .A1(men_men_n1599_), .B0(men_men_n814_), .Y(men_men_n1603_));
  NO2        u1554(.A(men_men_n745_), .B(men_men_n325_), .Y(men_men_n1604_));
  NO2        u1555(.A(men_men_n153_), .B(men_men_n1030_), .Y(men_men_n1605_));
  AOI220     u1556(.A0(men_men_n1605_), .A1(men_men_n1277_), .B0(men_men_n1604_), .B1(men_men_n480_), .Y(men_men_n1606_));
  AO210      u1557(.A0(men_men_n1606_), .A1(men_men_n1603_), .B0(x1), .Y(men_men_n1607_));
  NA3        u1558(.A(men_men_n635_), .B(men_men_n1055_), .C(men_men_n1200_), .Y(men_men_n1608_));
  NA2        u1559(.A(men_men_n146_), .B(men_men_n111_), .Y(men_men_n1609_));
  NOi21      u1560(.An(x1), .B(x6), .Y(men_men_n1610_));
  NA2        u1561(.A(men_men_n1610_), .B(men_men_n84_), .Y(men_men_n1611_));
  NA3        u1562(.A(men_men_n1611_), .B(men_men_n1609_), .C(men_men_n1608_), .Y(men_men_n1612_));
  AOI220     u1563(.A0(men_men_n1612_), .A1(x3), .B0(men_men_n1215_), .B1(men_men_n385_), .Y(men_men_n1613_));
  NA3        u1564(.A(men_men_n1220_), .B(men_men_n799_), .C(men_men_n606_), .Y(men_men_n1614_));
  AOI220     u1565(.A0(men_men_n1265_), .A1(men_men_n122_), .B0(men_men_n921_), .B1(men_men_n816_), .Y(men_men_n1615_));
  AOI210     u1566(.A0(men_men_n1615_), .A1(men_men_n1614_), .B0(men_men_n325_), .Y(men_men_n1616_));
  NA3        u1567(.A(men_men_n1208_), .B(men_men_n386_), .C(men_men_n110_), .Y(men_men_n1617_));
  NO2        u1568(.A(men_men_n1617_), .B(men_men_n969_), .Y(men_men_n1618_));
  NO3        u1569(.A(men_men_n621_), .B(men_men_n520_), .C(men_men_n1233_), .Y(men_men_n1619_));
  NO3        u1570(.A(men_men_n1619_), .B(men_men_n1618_), .C(men_men_n1616_), .Y(men_men_n1620_));
  OAI210     u1571(.A0(men_men_n1613_), .A1(men_men_n850_), .B0(men_men_n1620_), .Y(men_men_n1621_));
  NO2        u1572(.A(men_men_n557_), .B(men_men_n68_), .Y(men_men_n1622_));
  OAI220     u1573(.A0(men_men_n1622_), .A1(men_men_n1578_), .B0(men_men_n308_), .B1(men_men_n900_), .Y(men_men_n1623_));
  AOI220     u1574(.A0(men_men_n1623_), .A1(men_men_n56_), .B0(men_men_n1364_), .B1(men_men_n731_), .Y(men_men_n1624_));
  NO2        u1575(.A(men_men_n54_), .B(men_men_n71_), .Y(men_men_n1625_));
  AO220      u1576(.A0(men_men_n1625_), .A1(men_men_n1005_), .B0(men_men_n816_), .B1(men_men_n958_), .Y(men_men_n1626_));
  NA2        u1577(.A(men_men_n1191_), .B(men_men_n362_), .Y(men_men_n1627_));
  NO2        u1578(.A(men_men_n998_), .B(men_men_n1610_), .Y(men_men_n1628_));
  NA2        u1579(.A(men_men_n502_), .B(men_men_n731_), .Y(men_men_n1629_));
  OAI210     u1580(.A0(men_men_n1629_), .A1(men_men_n1628_), .B0(men_men_n1627_), .Y(men_men_n1630_));
  AOI210     u1581(.A0(men_men_n1626_), .A1(x2), .B0(men_men_n1630_), .Y(men_men_n1631_));
  OAI220     u1582(.A0(men_men_n1631_), .A1(men_men_n153_), .B0(men_men_n1624_), .B1(men_men_n54_), .Y(men_men_n1632_));
  OAI210     u1583(.A0(men_men_n1632_), .A1(men_men_n1621_), .B0(x8), .Y(men_men_n1633_));
  NA4        u1584(.A(men_men_n1633_), .B(men_men_n1607_), .C(men_men_n1597_), .D(men_men_n1585_), .Y(men20));
  NA2        u1585(.A(men_men_n480_), .B(men_men_n416_), .Y(men_men_n1635_));
  NO2        u1586(.A(men_men_n1635_), .B(men_men_n87_), .Y(men_men_n1636_));
  AOI210     u1587(.A0(men_men_n1059_), .A1(men_men_n62_), .B0(men_men_n1592_), .Y(men_men_n1637_));
  AOI210     u1588(.A0(men_men_n993_), .A1(men_men_n351_), .B0(men_men_n1198_), .Y(men_men_n1638_));
  OAI210     u1589(.A0(men_men_n1637_), .A1(men_men_n686_), .B0(men_men_n1638_), .Y(men_men_n1639_));
  OAI210     u1590(.A0(men_men_n1639_), .A1(men_men_n1636_), .B0(men_men_n1114_), .Y(men_men_n1640_));
  NAi21      u1591(.An(men_men_n553_), .B(men_men_n404_), .Y(men_men_n1641_));
  NA3        u1592(.A(men_men_n1641_), .B(men_men_n991_), .C(men_men_n958_), .Y(men_men_n1642_));
  NA3        u1593(.A(men_men_n1113_), .B(men_men_n281_), .C(men_men_n587_), .Y(men_men_n1643_));
  AOI210     u1594(.A0(men_men_n1643_), .A1(men_men_n1642_), .B0(men_men_n1308_), .Y(men_men_n1644_));
  NO2        u1595(.A(men_men_n749_), .B(men_men_n979_), .Y(men_men_n1645_));
  NA2        u1596(.A(men_men_n1644_), .B(men_men_n329_), .Y(men_men_n1646_));
  NO4        u1597(.A(men_men_n550_), .B(men_men_n237_), .C(x5), .D(x2), .Y(men_men_n1647_));
  NA2        u1598(.A(men_men_n321_), .B(men_men_n93_), .Y(men_men_n1648_));
  NA2        u1599(.A(men_men_n330_), .B(men_men_n108_), .Y(men_men_n1649_));
  INV        u1600(.A(men_men_n426_), .Y(men_men_n1650_));
  OAI220     u1601(.A0(men_men_n1650_), .A1(men_men_n1649_), .B0(men_men_n1648_), .B1(men_men_n276_), .Y(men_men_n1651_));
  OAI210     u1602(.A0(men_men_n1651_), .A1(men_men_n1647_), .B0(men_men_n222_), .Y(men_men_n1652_));
  NO2        u1603(.A(men_men_n670_), .B(men_men_n610_), .Y(men_men_n1653_));
  NA2        u1604(.A(men_men_n959_), .B(men_men_n50_), .Y(men_men_n1654_));
  NO3        u1605(.A(men_men_n1654_), .B(men_men_n368_), .C(men_men_n230_), .Y(men_men_n1655_));
  NA4        u1606(.A(men_men_n341_), .B(men_men_n239_), .C(men_men_n804_), .D(men_men_n64_), .Y(men_men_n1656_));
  OAI220     u1607(.A0(men_men_n1656_), .A1(men_men_n680_), .B0(men_men_n1475_), .B1(men_men_n1043_), .Y(men_men_n1657_));
  AOI210     u1608(.A0(men_men_n1655_), .A1(men_men_n1653_), .B0(men_men_n1657_), .Y(men_men_n1658_));
  NA4        u1609(.A(men_men_n1658_), .B(men_men_n1652_), .C(men_men_n1646_), .D(men_men_n1640_), .Y(men21));
  OAI210     u1610(.A0(men_men_n409_), .A1(men_men_n54_), .B0(x7), .Y(men_men_n1660_));
  OAI220     u1611(.A0(men_men_n1660_), .A1(men_men_n1297_), .B0(men_men_n1060_), .B1(men_men_n96_), .Y(men_men_n1661_));
  NA2        u1612(.A(men_men_n1661_), .B(men_men_n78_), .Y(men_men_n1662_));
  NA2        u1613(.A(men_men_n293_), .B(men_men_n861_), .Y(men_men_n1663_));
  AOI220     u1614(.A0(men_men_n1663_), .A1(men_men_n311_), .B0(men_men_n572_), .B1(men_men_n464_), .Y(men_men_n1664_));
  NA2        u1615(.A(men_men_n945_), .B(men_men_n275_), .Y(men_men_n1665_));
  NA2        u1616(.A(men_men_n541_), .B(men_men_n465_), .Y(men_men_n1666_));
  NA4        u1617(.A(men_men_n1666_), .B(men_men_n1665_), .C(men_men_n1391_), .D(men_men_n56_), .Y(men_men_n1667_));
  NO2        u1618(.A(men_men_n777_), .B(men_men_n437_), .Y(men_men_n1668_));
  NO3        u1619(.A(men_men_n1668_), .B(men_men_n723_), .C(men_men_n251_), .Y(men_men_n1669_));
  NOi31      u1620(.An(men_men_n193_), .B(men_men_n635_), .C(men_men_n1097_), .Y(men_men_n1670_));
  NO4        u1621(.A(men_men_n1670_), .B(men_men_n1669_), .C(men_men_n1667_), .D(men_men_n1664_), .Y(men_men_n1671_));
  NO3        u1622(.A(men_men_n437_), .B(men_men_n279_), .C(men_men_n52_), .Y(men_men_n1672_));
  OA210      u1623(.A0(men_men_n1672_), .A1(men_men_n889_), .B0(x3), .Y(men_men_n1673_));
  OAI210     u1624(.A0(men_men_n788_), .A1(men_men_n592_), .B0(men_men_n343_), .Y(men_men_n1674_));
  NO2        u1625(.A(men_men_n70_), .B(x2), .Y(men_men_n1675_));
  OAI210     u1626(.A0(men_men_n177_), .A1(x0), .B0(men_men_n1675_), .Y(men_men_n1676_));
  NA2        u1627(.A(men_men_n143_), .B(men_men_n108_), .Y(men_men_n1677_));
  NA3        u1628(.A(men_men_n1677_), .B(men_men_n1676_), .C(men_men_n1674_), .Y(men_men_n1678_));
  OAI210     u1629(.A0(men_men_n1678_), .A1(men_men_n1673_), .B0(x8), .Y(men_men_n1679_));
  NO3        u1630(.A(men_men_n775_), .B(men_men_n624_), .C(men_men_n588_), .Y(men_men_n1680_));
  NA2        u1631(.A(men_men_n55_), .B(men_men_n50_), .Y(men_men_n1681_));
  MUX2       u1632(.S(men_men_n604_), .A(men_men_n1681_), .B(men_men_n107_), .Y(men_men_n1682_));
  AOI210     u1633(.A0(men_men_n1369_), .A1(men_men_n240_), .B0(men_men_n1682_), .Y(men_men_n1683_));
  OAI210     u1634(.A0(men_men_n648_), .A1(men_men_n587_), .B0(x4), .Y(men_men_n1684_));
  NO3        u1635(.A(men_men_n1684_), .B(men_men_n1683_), .C(men_men_n1680_), .Y(men_men_n1685_));
  AO220      u1636(.A0(men_men_n1685_), .A1(men_men_n1679_), .B0(men_men_n1671_), .B1(men_men_n1662_), .Y(men_men_n1686_));
  AO220      u1637(.A0(men_men_n636_), .A1(men_men_n325_), .B0(men_men_n593_), .B1(x8), .Y(men_men_n1687_));
  NO2        u1638(.A(men_men_n863_), .B(x0), .Y(men_men_n1688_));
  NO3        u1639(.A(men_men_n1688_), .B(men_men_n551_), .C(men_men_n88_), .Y(men_men_n1689_));
  NO2        u1640(.A(men_men_n159_), .B(x2), .Y(men_men_n1690_));
  NO3        u1641(.A(men_men_n381_), .B(men_men_n256_), .C(men_men_n185_), .Y(men_men_n1691_));
  AOI210     u1642(.A0(men_men_n1690_), .A1(men_men_n68_), .B0(men_men_n1691_), .Y(men_men_n1692_));
  OAI210     u1643(.A0(men_men_n1689_), .A1(men_men_n402_), .B0(men_men_n1692_), .Y(men_men_n1693_));
  AOI220     u1644(.A0(men_men_n1693_), .A1(x5), .B0(men_men_n1687_), .B1(men_men_n749_), .Y(men_men_n1694_));
  AOI210     u1645(.A0(men_men_n1694_), .A1(men_men_n1686_), .B0(men_men_n71_), .Y(men_men_n1695_));
  NO2        u1646(.A(men_men_n912_), .B(men_men_n168_), .Y(men_men_n1696_));
  NOi41      u1647(.An(men_men_n1443_), .B(men_men_n1510_), .C(men_men_n1166_), .D(men_men_n854_), .Y(men_men_n1697_));
  NA2        u1648(.A(men_men_n1697_), .B(men_men_n1696_), .Y(men_men_n1698_));
  NO2        u1649(.A(men_men_n78_), .B(x4), .Y(men_men_n1699_));
  OAI210     u1650(.A0(men_men_n291_), .A1(men_men_n157_), .B0(men_men_n1699_), .Y(men_men_n1700_));
  OAI210     u1651(.A0(men_men_n411_), .A1(men_men_n427_), .B0(men_men_n230_), .Y(men_men_n1701_));
  NO2        u1652(.A(men_men_n258_), .B(men_men_n50_), .Y(men_men_n1702_));
  NO2        u1653(.A(men_men_n1702_), .B(men_men_n57_), .Y(men_men_n1703_));
  NA2        u1654(.A(men_men_n1703_), .B(men_men_n1701_), .Y(men_men_n1704_));
  AOI210     u1655(.A0(men_men_n1700_), .A1(men_men_n1698_), .B0(men_men_n1704_), .Y(men_men_n1705_));
  NA2        u1656(.A(men_men_n761_), .B(men_men_n553_), .Y(men_men_n1706_));
  AO210      u1657(.A0(men_men_n1706_), .A1(men_men_n969_), .B0(men_men_n50_), .Y(men_men_n1707_));
  NO2        u1658(.A(men_men_n1641_), .B(men_men_n1227_), .Y(men_men_n1708_));
  AOI220     u1659(.A0(men_men_n1708_), .A1(men_men_n1176_), .B0(men_men_n1336_), .B1(men_men_n1054_), .Y(men_men_n1709_));
  AOI210     u1660(.A0(men_men_n1709_), .A1(men_men_n1707_), .B0(men_men_n110_), .Y(men_men_n1710_));
  NA2        u1661(.A(men_men_n300_), .B(men_men_n108_), .Y(men_men_n1711_));
  NA2        u1662(.A(men_men_n899_), .B(men_men_n55_), .Y(men_men_n1712_));
  NO2        u1663(.A(men_men_n675_), .B(men_men_n1063_), .Y(men_men_n1713_));
  NO3        u1664(.A(men_men_n1713_), .B(men_men_n1710_), .C(men_men_n1705_), .Y(men_men_n1714_));
  NO2        u1665(.A(men_men_n1714_), .B(x6), .Y(men_men_n1715_));
  AOI210     u1666(.A0(men_men_n613_), .A1(men_men_n1063_), .B0(men_men_n1510_), .Y(men_men_n1716_));
  OAI210     u1667(.A0(men_men_n1716_), .A1(men_men_n693_), .B0(men_men_n56_), .Y(men_men_n1717_));
  NO2        u1668(.A(men_men_n751_), .B(men_men_n54_), .Y(men_men_n1718_));
  NO4        u1669(.A(men_men_n967_), .B(men_men_n279_), .C(men_men_n774_), .D(men_men_n758_), .Y(men_men_n1719_));
  NO2        u1670(.A(men_men_n868_), .B(x5), .Y(men_men_n1720_));
  NO4        u1671(.A(men_men_n1720_), .B(men_men_n1719_), .C(men_men_n1718_), .D(men_men_n952_), .Y(men_men_n1721_));
  AOI210     u1672(.A0(men_men_n1721_), .A1(men_men_n1717_), .B0(men_men_n50_), .Y(men_men_n1722_));
  NA2        u1673(.A(men_men_n159_), .B(men_men_n108_), .Y(men_men_n1723_));
  OA220      u1674(.A0(men_men_n1723_), .A1(men_men_n441_), .B0(men_men_n470_), .B1(men_men_n749_), .Y(men_men_n1724_));
  NA3        u1675(.A(men_men_n55_), .B(x2), .C(x0), .Y(men_men_n1725_));
  AOI220     u1676(.A0(men_men_n1725_), .A1(men_men_n170_), .B0(men_men_n868_), .B1(men_men_n155_), .Y(men_men_n1726_));
  NO2        u1677(.A(men_men_n686_), .B(men_men_n258_), .Y(men_men_n1727_));
  NO3        u1678(.A(men_men_n246_), .B(men_men_n228_), .C(men_men_n362_), .Y(men_men_n1728_));
  NO3        u1679(.A(men_men_n1728_), .B(men_men_n1727_), .C(men_men_n1726_), .Y(men_men_n1729_));
  OAI220     u1680(.A0(men_men_n1729_), .A1(men_men_n56_), .B0(men_men_n1724_), .B1(men_men_n702_), .Y(men_men_n1730_));
  OAI210     u1681(.A0(men_men_n1730_), .A1(men_men_n1722_), .B0(men_men_n116_), .Y(men_men_n1731_));
  NO2        u1682(.A(men_men_n618_), .B(men_men_n306_), .Y(men_men_n1732_));
  AOI210     u1683(.A0(men_men_n611_), .A1(x5), .B0(men_men_n1732_), .Y(men_men_n1733_));
  NO2        u1684(.A(men_men_n1733_), .B(men_men_n110_), .Y(men_men_n1734_));
  NA2        u1685(.A(men_men_n710_), .B(men_men_n81_), .Y(men_men_n1735_));
  NA3        u1686(.A(men_men_n1735_), .B(men_men_n434_), .C(men_men_n57_), .Y(men_men_n1736_));
  OAI210     u1687(.A0(men_men_n1712_), .A1(men_men_n1711_), .B0(men_men_n1736_), .Y(men_men_n1737_));
  OAI210     u1688(.A0(men_men_n1737_), .A1(men_men_n1734_), .B0(x1), .Y(men_men_n1738_));
  NO4        u1689(.A(men_men_n420_), .B(men_men_n78_), .C(men_men_n147_), .D(x3), .Y(men_men_n1739_));
  NO2        u1690(.A(men_men_n330_), .B(men_men_n112_), .Y(men_men_n1740_));
  OAI210     u1691(.A0(men_men_n1739_), .A1(men_men_n1309_), .B0(men_men_n1740_), .Y(men_men_n1741_));
  NO2        u1692(.A(men_men_n60_), .B(men_men_n108_), .Y(men_men_n1742_));
  NO4        u1693(.A(men_men_n1711_), .B(men_men_n967_), .C(men_men_n670_), .D(men_men_n50_), .Y(men_men_n1743_));
  AOI210     u1694(.A0(men_men_n1742_), .A1(men_men_n1554_), .B0(men_men_n1743_), .Y(men_men_n1744_));
  NA4        u1695(.A(men_men_n1744_), .B(men_men_n1741_), .C(men_men_n1738_), .D(men_men_n1731_), .Y(men_men_n1745_));
  NO3        u1696(.A(men_men_n1745_), .B(men_men_n1715_), .C(men_men_n1695_), .Y(men22));
  AOI210     u1697(.A0(men_men_n527_), .A1(men_men_n71_), .B0(men_men_n473_), .Y(men_men_n1747_));
  NO2        u1698(.A(men_men_n1203_), .B(men_men_n557_), .Y(men_men_n1748_));
  AOI210     u1699(.A0(x5), .A1(x2), .B0(x8), .Y(men_men_n1749_));
  NA2        u1700(.A(men_men_n1749_), .B(men_men_n59_), .Y(men_men_n1750_));
  OAI220     u1701(.A0(men_men_n1750_), .A1(men_men_n1748_), .B0(men_men_n1747_), .B1(men_men_n402_), .Y(men_men_n1751_));
  NA2        u1702(.A(men_men_n587_), .B(men_men_n87_), .Y(men_men_n1752_));
  NA2        u1703(.A(men_men_n276_), .B(men_men_n77_), .Y(men_men_n1753_));
  OA220      u1704(.A0(men_men_n1753_), .A1(men_men_n1752_), .B0(men_men_n847_), .B1(men_men_n1015_), .Y(men_men_n1754_));
  NO3        u1705(.A(men_men_n1256_), .B(men_men_n87_), .C(x0), .Y(men_men_n1755_));
  OAI210     u1706(.A0(men_men_n402_), .A1(men_men_n205_), .B0(x4), .Y(men_men_n1756_));
  NO2        u1707(.A(men_men_n1756_), .B(men_men_n1755_), .Y(men_men_n1757_));
  OAI210     u1708(.A0(men_men_n1754_), .A1(men_men_n198_), .B0(men_men_n1757_), .Y(men_men_n1758_));
  AOI210     u1709(.A0(men_men_n1751_), .A1(men_men_n53_), .B0(men_men_n1758_), .Y(men_men_n1759_));
  NA2        u1710(.A(men_men_n304_), .B(men_men_n309_), .Y(men_men_n1760_));
  NA3        u1711(.A(men_men_n1760_), .B(men_men_n222_), .C(men_men_n308_), .Y(men_men_n1761_));
  NA2        u1712(.A(men_men_n582_), .B(men_men_n245_), .Y(men_men_n1762_));
  NO3        u1713(.A(men_men_n502_), .B(men_men_n266_), .C(men_men_n214_), .Y(men_men_n1763_));
  NA2        u1714(.A(men_men_n1762_), .B(men_men_n1761_), .Y(men_men_n1764_));
  NO2        u1715(.A(men_men_n470_), .B(men_men_n260_), .Y(men_men_n1765_));
  NO2        u1716(.A(men_men_n1256_), .B(x3), .Y(men_men_n1766_));
  AOI210     u1717(.A0(men_men_n1766_), .A1(men_men_n351_), .B0(men_men_n1765_), .Y(men_men_n1767_));
  OAI210     u1718(.A0(men_men_n1092_), .A1(men_men_n187_), .B0(men_men_n56_), .Y(men_men_n1768_));
  NA3        u1719(.A(men_men_n55_), .B(men_men_n71_), .C(x0), .Y(men_men_n1769_));
  OAI220     u1720(.A0(men_men_n1769_), .A1(men_men_n1063_), .B0(men_men_n368_), .B1(men_men_n213_), .Y(men_men_n1770_));
  NO2        u1721(.A(men_men_n1770_), .B(men_men_n1768_), .Y(men_men_n1771_));
  OAI210     u1722(.A0(men_men_n1767_), .A1(men_men_n258_), .B0(men_men_n1771_), .Y(men_men_n1772_));
  AOI210     u1723(.A0(men_men_n1764_), .A1(men_men_n108_), .B0(men_men_n1772_), .Y(men_men_n1773_));
  AOI210     u1724(.A0(men_men_n956_), .A1(men_men_n776_), .B0(men_men_n872_), .Y(men_men_n1774_));
  NO2        u1725(.A(men_men_n806_), .B(men_men_n159_), .Y(men_men_n1775_));
  OAI210     u1726(.A0(men_men_n1775_), .A1(men_men_n1774_), .B0(men_men_n617_), .Y(men_men_n1776_));
  OA210      u1727(.A0(men_men_n1773_), .A1(men_men_n1759_), .B0(men_men_n1776_), .Y(men_men_n1777_));
  OAI210     u1728(.A0(men_men_n1185_), .A1(men_men_n709_), .B0(men_men_n697_), .Y(men_men_n1778_));
  NO2        u1729(.A(men_men_n356_), .B(x0), .Y(men_men_n1779_));
  NA3        u1730(.A(men_men_n1779_), .B(men_men_n351_), .C(men_men_n56_), .Y(men_men_n1780_));
  AOI210     u1731(.A0(men_men_n1780_), .A1(men_men_n1778_), .B0(men_men_n402_), .Y(men_men_n1781_));
  NO3        u1732(.A(men_men_n170_), .B(men_men_n159_), .C(men_men_n62_), .Y(men_men_n1782_));
  OAI210     u1733(.A0(men_men_n1782_), .A1(men_men_n422_), .B0(men_men_n110_), .Y(men_men_n1783_));
  NA2        u1734(.A(men_men_n139_), .B(men_men_n789_), .Y(men_men_n1784_));
  NA2        u1735(.A(men_men_n420_), .B(x3), .Y(men_men_n1785_));
  NAi31      u1736(.An(men_men_n1785_), .B(men_men_n1784_), .C(men_men_n1570_), .Y(men_men_n1786_));
  NO3        u1737(.A(men_men_n863_), .B(men_men_n469_), .C(men_men_n110_), .Y(men_men_n1787_));
  NO2        u1738(.A(men_men_n1094_), .B(men_men_n140_), .Y(men_men_n1788_));
  NO3        u1739(.A(men_men_n902_), .B(men_men_n416_), .C(men_men_n305_), .Y(men_men_n1789_));
  AOI220     u1740(.A0(men_men_n1789_), .A1(men_men_n1788_), .B0(men_men_n1787_), .B1(men_men_n1779_), .Y(men_men_n1790_));
  NA3        u1741(.A(men_men_n416_), .B(men_men_n93_), .C(men_men_n81_), .Y(men_men_n1791_));
  AOI210     u1742(.A0(men_men_n613_), .A1(men_men_n459_), .B0(men_men_n499_), .Y(men_men_n1792_));
  NA2        u1743(.A(men_men_n1187_), .B(x3), .Y(men_men_n1793_));
  OAI210     u1744(.A0(men_men_n1793_), .A1(men_men_n1792_), .B0(men_men_n1791_), .Y(men_men_n1794_));
  NA3        u1745(.A(men_men_n56_), .B(men_men_n50_), .C(x0), .Y(men_men_n1795_));
  NOi21      u1746(.An(men_men_n83_), .B(men_men_n734_), .Y(men_men_n1796_));
  NA3        u1747(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n1797_));
  NA3        u1748(.A(men_men_n1797_), .B(men_men_n998_), .C(men_men_n267_), .Y(men_men_n1798_));
  OAI220     u1749(.A0(men_men_n1798_), .A1(men_men_n1796_), .B0(men_men_n1066_), .B1(men_men_n1795_), .Y(men_men_n1799_));
  AOI220     u1750(.A0(men_men_n1799_), .A1(men_men_n1077_), .B0(men_men_n1794_), .B1(men_men_n351_), .Y(men_men_n1800_));
  NA4        u1751(.A(men_men_n1800_), .B(men_men_n1790_), .C(men_men_n1786_), .D(men_men_n1783_), .Y(men_men_n1801_));
  AOI210     u1752(.A0(men_men_n1801_), .A1(x7), .B0(men_men_n1781_), .Y(men_men_n1802_));
  OAI210     u1753(.A0(men_men_n1777_), .A1(x7), .B0(men_men_n1802_), .Y(men23));
  OR2        u1754(.A(men_men_n521_), .B(men_men_n222_), .Y(men_men_n1804_));
  NA2        u1755(.A(men_men_n1804_), .B(men_men_n1645_), .Y(men_men_n1805_));
  NO3        u1756(.A(men_men_n847_), .B(men_men_n596_), .C(men_men_n492_), .Y(men_men_n1806_));
  NO3        u1757(.A(men_men_n960_), .B(men_men_n148_), .C(men_men_n117_), .Y(men_men_n1807_));
  AOI210     u1758(.A0(men_men_n1807_), .A1(men_men_n1037_), .B0(men_men_n1806_), .Y(men_men_n1808_));
  OAI210     u1759(.A0(men_men_n1805_), .A1(men_men_n153_), .B0(men_men_n1808_), .Y(men_men_n1809_));
  NA2        u1760(.A(men_men_n1809_), .B(men_men_n55_), .Y(men_men_n1810_));
  NO2        u1761(.A(men_men_n967_), .B(men_men_n519_), .Y(men_men_n1811_));
  AO220      u1762(.A0(men_men_n1293_), .A1(men_men_n181_), .B0(men_men_n1005_), .B1(men_men_n749_), .Y(men_men_n1812_));
  OAI210     u1763(.A0(men_men_n1812_), .A1(men_men_n1811_), .B0(men_men_n593_), .Y(men_men_n1813_));
  NA2        u1764(.A(men_men_n178_), .B(men_men_n168_), .Y(men_men_n1814_));
  NA2        u1765(.A(men_men_n408_), .B(men_men_n160_), .Y(men_men_n1815_));
  AOI210     u1766(.A0(men_men_n1815_), .A1(men_men_n1814_), .B0(men_men_n237_), .Y(men_men_n1816_));
  NA3        u1767(.A(men_men_n872_), .B(men_men_n427_), .C(men_men_n258_), .Y(men_men_n1817_));
  AOI210     u1768(.A0(men_men_n1817_), .A1(men_men_n504_), .B0(men_men_n386_), .Y(men_men_n1818_));
  OAI210     u1769(.A0(men_men_n1818_), .A1(men_men_n1816_), .B0(men_men_n300_), .Y(men_men_n1819_));
  NA3        u1770(.A(men_men_n57_), .B(x4), .C(x3), .Y(men_men_n1820_));
  NO3        u1771(.A(men_men_n1820_), .B(men_men_n746_), .C(men_men_n139_), .Y(men_men_n1821_));
  AOI210     u1772(.A0(men_men_n925_), .A1(men_men_n141_), .B0(men_men_n1821_), .Y(men_men_n1822_));
  NA4        u1773(.A(men_men_n1822_), .B(men_men_n1819_), .C(men_men_n1813_), .D(men_men_n1810_), .Y(men24));
  NO2        u1774(.A(men_men_n242_), .B(x1), .Y(men_men_n1824_));
  NA2        u1775(.A(men_men_n341_), .B(men_men_n496_), .Y(men_men_n1825_));
  NAi21      u1776(.An(men_men_n1824_), .B(men_men_n1825_), .Y(men_men_n1826_));
  NO3        u1777(.A(men_men_n546_), .B(men_men_n689_), .C(men_men_n155_), .Y(men_men_n1827_));
  AOI210     u1778(.A0(men_men_n1826_), .A1(men_men_n93_), .B0(men_men_n1827_), .Y(men_men_n1828_));
  NA2        u1779(.A(men_men_n102_), .B(x8), .Y(men_men_n1829_));
  NO3        u1780(.A(men_men_n1074_), .B(men_men_n1350_), .C(men_men_n1055_), .Y(men_men_n1830_));
  AOI210     u1781(.A0(men_men_n991_), .A1(men_men_n56_), .B0(men_men_n1465_), .Y(men_men_n1831_));
  AO220      u1782(.A0(men_men_n1831_), .A1(men_men_n1830_), .B0(men_men_n1279_), .B1(men_men_n329_), .Y(men_men_n1832_));
  NA2        u1783(.A(men_men_n459_), .B(x8), .Y(men_men_n1833_));
  NA2        u1784(.A(men_men_n671_), .B(men_men_n125_), .Y(men_men_n1834_));
  OAI220     u1785(.A0(men_men_n1834_), .A1(men_men_n1452_), .B0(men_men_n1833_), .B1(men_men_n845_), .Y(men_men_n1835_));
  AOI220     u1786(.A0(men_men_n1835_), .A1(men_men_n1702_), .B0(men_men_n1832_), .B1(men_men_n1037_), .Y(men_men_n1836_));
  OAI210     u1787(.A0(men_men_n1829_), .A1(men_men_n1828_), .B0(men_men_n1836_), .Y(men25));
  NA2        u1788(.A(men_men_n330_), .B(men_men_n59_), .Y(men_men_n1838_));
  NO2        u1789(.A(men_men_n1838_), .B(men_men_n322_), .Y(men_men_n1839_));
  OAI210     u1790(.A0(men_men_n1839_), .A1(men_men_n1192_), .B0(men_men_n116_), .Y(men_men_n1840_));
  INV        u1791(.A(men_men_n1288_), .Y(men_men_n1841_));
  NO2        u1792(.A(men_men_n745_), .B(men_men_n55_), .Y(men_men_n1842_));
  AOI220     u1793(.A0(men_men_n1842_), .A1(men_men_n1841_), .B0(men_men_n1604_), .B1(men_men_n1193_), .Y(men_men_n1843_));
  AOI210     u1794(.A0(men_men_n1843_), .A1(men_men_n1840_), .B0(men_men_n684_), .Y(men_men_n1844_));
  NO3        u1795(.A(men_men_n1049_), .B(men_men_n142_), .C(men_men_n78_), .Y(men_men_n1845_));
  OAI210     u1796(.A0(men_men_n198_), .A1(men_men_n276_), .B0(men_men_n331_), .Y(men_men_n1846_));
  OAI210     u1797(.A0(men_men_n1846_), .A1(men_men_n1845_), .B0(men_men_n1191_), .Y(men_men_n1847_));
  NO2        u1798(.A(men_men_n1403_), .B(men_men_n452_), .Y(men_men_n1848_));
  NO3        u1799(.A(men_men_n1848_), .B(men_men_n537_), .C(men_men_n99_), .Y(men_men_n1849_));
  NA2        u1800(.A(men_men_n514_), .B(men_men_n55_), .Y(men_men_n1850_));
  OAI220     u1801(.A0(men_men_n1850_), .A1(men_men_n242_), .B0(men_men_n590_), .B1(men_men_n276_), .Y(men_men_n1851_));
  OAI210     u1802(.A0(men_men_n1851_), .A1(men_men_n1849_), .B0(men_men_n640_), .Y(men_men_n1852_));
  AOI220     u1803(.A0(men_men_n1765_), .A1(men_men_n1145_), .B0(men_men_n1504_), .B1(men_men_n382_), .Y(men_men_n1853_));
  NA3        u1804(.A(men_men_n1853_), .B(men_men_n1852_), .C(men_men_n1847_), .Y(men_men_n1854_));
  AO210      u1805(.A0(men_men_n1854_), .A1(men_men_n108_), .B0(men_men_n1844_), .Y(men26));
  NA2        u1806(.A(men_men_n774_), .B(men_men_n50_), .Y(men_men_n1856_));
  OAI220     u1807(.A0(men_men_n306_), .A1(men_men_n251_), .B0(men_men_n1856_), .B1(x7), .Y(men_men_n1857_));
  AOI220     u1808(.A0(men_men_n1857_), .A1(men_men_n93_), .B0(men_men_n1309_), .B1(men_men_n1151_), .Y(men_men_n1858_));
  NA2        u1809(.A(men_men_n628_), .B(men_men_n582_), .Y(men_men_n1859_));
  OAI210     u1810(.A0(men_men_n636_), .A1(men_men_n628_), .B0(men_men_n749_), .Y(men_men_n1860_));
  AOI210     u1811(.A0(men_men_n1859_), .A1(men_men_n1214_), .B0(men_men_n1860_), .Y(men_men_n1861_));
  NA2        u1812(.A(men_men_n1028_), .B(men_men_n588_), .Y(men_men_n1862_));
  NO2        u1813(.A(men_men_n1862_), .B(men_men_n1261_), .Y(men_men_n1863_));
  AOI210     u1814(.A0(men_men_n1788_), .A1(men_men_n1471_), .B0(men_men_n1863_), .Y(men_men_n1864_));
  NO2        u1815(.A(men_men_n1094_), .B(men_men_n75_), .Y(men_men_n1865_));
  NA2        u1816(.A(men_men_n814_), .B(men_men_n177_), .Y(men_men_n1866_));
  NO2        u1817(.A(men_men_n1866_), .B(men_men_n542_), .Y(men_men_n1867_));
  AOI210     u1818(.A0(men_men_n1865_), .A1(men_men_n589_), .B0(men_men_n1867_), .Y(men_men_n1868_));
  OAI220     u1819(.A0(men_men_n1868_), .A1(men_men_n108_), .B0(men_men_n1864_), .B1(men_men_n53_), .Y(men_men_n1869_));
  NA2        u1820(.A(men_men_n605_), .B(men_men_n514_), .Y(men_men_n1870_));
  NO2        u1821(.A(men_men_n132_), .B(men_men_n129_), .Y(men_men_n1871_));
  NA2        u1822(.A(men_men_n1871_), .B(men_men_n122_), .Y(men_men_n1872_));
  NA2        u1823(.A(men_men_n749_), .B(x3), .Y(men_men_n1873_));
  AOI210     u1824(.A0(men_men_n1872_), .A1(men_men_n1870_), .B0(men_men_n1873_), .Y(men_men_n1874_));
  NO2        u1825(.A(men_men_n1015_), .B(x3), .Y(men_men_n1875_));
  AOI210     u1826(.A0(men_men_n450_), .A1(men_men_n108_), .B0(men_men_n1875_), .Y(men_men_n1876_));
  NA3        u1827(.A(men_men_n573_), .B(men_men_n51_), .C(men_men_n56_), .Y(men_men_n1877_));
  AOI210     u1828(.A0(men_men_n1653_), .A1(men_men_n1067_), .B0(x0), .Y(men_men_n1878_));
  OAI210     u1829(.A0(men_men_n1877_), .A1(men_men_n1876_), .B0(men_men_n1878_), .Y(men_men_n1879_));
  NO4        u1830(.A(men_men_n1879_), .B(men_men_n1874_), .C(men_men_n1869_), .D(men_men_n1861_), .Y(men_men_n1880_));
  AOI210     u1831(.A0(x8), .A1(x6), .B0(x5), .Y(men_men_n1881_));
  AO220      u1832(.A0(men_men_n1881_), .A1(men_men_n144_), .B0(men_men_n596_), .B1(men_men_n139_), .Y(men_men_n1882_));
  NA2        u1833(.A(men_men_n1882_), .B(men_men_n451_), .Y(men_men_n1883_));
  NO2        u1834(.A(men_men_n759_), .B(men_men_n144_), .Y(men_men_n1884_));
  NA3        u1835(.A(men_men_n1884_), .B(men_men_n1675_), .C(men_men_n133_), .Y(men_men_n1885_));
  NO2        u1836(.A(men_men_n402_), .B(men_men_n1389_), .Y(men_men_n1886_));
  NA2        u1837(.A(men_men_n1886_), .B(men_men_n450_), .Y(men_men_n1887_));
  NA3        u1838(.A(men_men_n376_), .B(men_men_n861_), .C(men_men_n255_), .Y(men_men_n1888_));
  NA4        u1839(.A(men_men_n1888_), .B(men_men_n1887_), .C(men_men_n1885_), .D(men_men_n1883_), .Y(men_men_n1889_));
  INV        u1840(.A(men_men_n497_), .Y(men_men_n1890_));
  NO2        u1841(.A(men_men_n1890_), .B(men_men_n117_), .Y(men_men_n1891_));
  NA3        u1842(.A(men_men_n816_), .B(men_men_n1015_), .C(x7), .Y(men_men_n1892_));
  AOI210     u1843(.A0(men_men_n345_), .A1(men_men_n216_), .B0(men_men_n1892_), .Y(men_men_n1893_));
  OAI220     u1844(.A0(men_men_n905_), .A1(men_men_n306_), .B0(men_men_n648_), .B1(men_men_n689_), .Y(men_men_n1894_));
  NO3        u1845(.A(men_men_n1894_), .B(men_men_n1893_), .C(men_men_n1891_), .Y(men_men_n1895_));
  NA3        u1846(.A(men_men_n671_), .B(men_men_n192_), .C(men_men_n958_), .Y(men_men_n1896_));
  NA2        u1847(.A(men_men_n1896_), .B(men_men_n648_), .Y(men_men_n1897_));
  NA2        u1848(.A(men_men_n139_), .B(men_men_n131_), .Y(men_men_n1898_));
  OAI210     u1849(.A0(men_men_n1898_), .A1(men_men_n1438_), .B0(x0), .Y(men_men_n1899_));
  AOI210     u1850(.A0(men_men_n1897_), .A1(men_men_n1428_), .B0(men_men_n1899_), .Y(men_men_n1900_));
  OAI210     u1851(.A0(men_men_n1895_), .A1(men_men_n53_), .B0(men_men_n1900_), .Y(men_men_n1901_));
  AOI210     u1852(.A0(men_men_n1889_), .A1(x4), .B0(men_men_n1901_), .Y(men_men_n1902_));
  OA220      u1853(.A0(men_men_n1902_), .A1(men_men_n1880_), .B0(men_men_n1858_), .B1(men_men_n109_), .Y(men27));
  NA2        u1854(.A(men_men_n1155_), .B(men_men_n450_), .Y(men_men_n1904_));
  NO2        u1855(.A(men_men_n1904_), .B(men_men_n301_), .Y(men_men_n1905_));
  NA2        u1856(.A(men_men_n921_), .B(men_men_n816_), .Y(men_men_n1906_));
  NA3        u1857(.A(men_men_n822_), .B(men_men_n365_), .C(men_men_n1030_), .Y(men_men_n1907_));
  AOI210     u1858(.A0(men_men_n1907_), .A1(men_men_n1906_), .B0(men_men_n216_), .Y(men_men_n1908_));
  OAI210     u1859(.A0(men_men_n1908_), .A1(men_men_n1905_), .B0(men_men_n705_), .Y(men_men_n1909_));
  XO2        u1860(.A(x8), .B(x4), .Y(men_men_n1910_));
  NO3        u1861(.A(men_men_n1910_), .B(men_men_n450_), .C(men_men_n170_), .Y(men_men_n1911_));
  OA210      u1862(.A0(men_men_n1911_), .A1(men_men_n1262_), .B0(men_men_n279_), .Y(men_men_n1912_));
  NO2        u1863(.A(men_men_n397_), .B(men_men_n164_), .Y(men_men_n1913_));
  OAI210     u1864(.A0(men_men_n1913_), .A1(men_men_n1912_), .B0(men_men_n1129_), .Y(men_men_n1914_));
  AOI210     u1865(.A0(men_men_n636_), .A1(men_men_n56_), .B0(men_men_n1865_), .Y(men_men_n1915_));
  OAI220     u1866(.A0(men_men_n1915_), .A1(men_men_n1261_), .B0(men_men_n1213_), .B1(men_men_n207_), .Y(men_men_n1916_));
  NO2        u1867(.A(men_men_n702_), .B(men_men_n142_), .Y(men_men_n1917_));
  NO2        u1868(.A(men_men_n1197_), .B(men_men_n258_), .Y(men_men_n1918_));
  AOI220     u1869(.A0(men_men_n1918_), .A1(men_men_n1917_), .B0(men_men_n1916_), .B1(men_men_n541_), .Y(men_men_n1919_));
  NA3        u1870(.A(men_men_n1919_), .B(men_men_n1914_), .C(men_men_n1909_), .Y(men28));
  NO3        u1871(.A(men_men_n1910_), .B(men_men_n1398_), .C(men_men_n146_), .Y(men_men_n1921_));
  OAI210     u1872(.A0(men_men_n1921_), .A1(men_men_n1281_), .B0(men_men_n588_), .Y(men_men_n1922_));
  NA3        u1873(.A(men_men_n1193_), .B(men_men_n899_), .C(x7), .Y(men_men_n1923_));
  NA3        u1874(.A(men_men_n499_), .B(men_men_n78_), .C(men_men_n610_), .Y(men_men_n1924_));
  NA3        u1875(.A(men_men_n1924_), .B(men_men_n1923_), .C(men_men_n1922_), .Y(men_men_n1925_));
  NA2        u1876(.A(men_men_n1256_), .B(men_men_n448_), .Y(men_men_n1926_));
  NA3        u1877(.A(men_men_n1926_), .B(men_men_n1417_), .C(men_men_n415_), .Y(men_men_n1927_));
  NO2        u1878(.A(men_men_n309_), .B(x4), .Y(men_men_n1928_));
  AOI220     u1879(.A0(men_men_n1928_), .A1(men_men_n1875_), .B0(men_men_n1130_), .B1(men_men_n679_), .Y(men_men_n1929_));
  NA2        u1880(.A(men_men_n1929_), .B(men_men_n1927_), .Y(men_men_n1930_));
  NO2        u1881(.A(men_men_n1256_), .B(men_men_n1233_), .Y(men_men_n1931_));
  NO4        u1882(.A(x6), .B(men_men_n56_), .C(x2), .D(x0), .Y(men_men_n1932_));
  OAI210     u1883(.A0(men_men_n1932_), .A1(men_men_n1931_), .B0(men_men_n1054_), .Y(men_men_n1933_));
  NA2        u1884(.A(men_men_n1187_), .B(men_men_n108_), .Y(men_men_n1934_));
  NA2        u1885(.A(men_men_n1090_), .B(men_men_n107_), .Y(men_men_n1935_));
  OAI210     u1886(.A0(men_men_n1935_), .A1(men_men_n1934_), .B0(men_men_n1933_), .Y(men_men_n1936_));
  OAI210     u1887(.A0(men_men_n1936_), .A1(men_men_n1930_), .B0(x7), .Y(men_men_n1937_));
  NO2        u1888(.A(men_men_n389_), .B(x7), .Y(men_men_n1938_));
  NO3        u1889(.A(men_men_n402_), .B(men_men_n273_), .C(men_men_n123_), .Y(men_men_n1939_));
  INV        u1890(.A(men_men_n81_), .Y(men_men_n1940_));
  OAI220     u1891(.A0(men_men_n1940_), .A1(men_men_n1939_), .B0(men_men_n1938_), .B1(men_men_n111_), .Y(men_men_n1941_));
  NA2        u1892(.A(men_men_n1797_), .B(men_men_n659_), .Y(men_men_n1942_));
  NO2        u1893(.A(men_men_n1850_), .B(men_men_n77_), .Y(men_men_n1943_));
  AOI220     u1894(.A0(men_men_n1943_), .A1(men_men_n1942_), .B0(men_men_n481_), .B1(men_men_n50_), .Y(men_men_n1944_));
  AOI210     u1895(.A0(men_men_n1944_), .A1(men_men_n1941_), .B0(men_men_n59_), .Y(men_men_n1945_));
  AOI220     u1896(.A0(men_men_n1403_), .A1(men_men_n677_), .B0(men_men_n414_), .B1(men_men_n459_), .Y(men_men_n1946_));
  OAI210     u1897(.A0(men_men_n1946_), .A1(men_men_n142_), .B0(x1), .Y(men_men_n1947_));
  NO2        u1898(.A(men_men_n1947_), .B(men_men_n1945_), .Y(men_men_n1948_));
  AOI210     u1899(.A0(men_men_n1589_), .A1(men_men_n402_), .B0(men_men_n669_), .Y(men_men_n1949_));
  NO2        u1900(.A(men_men_n402_), .B(x5), .Y(men_men_n1950_));
  NO2        u1901(.A(men_men_n1950_), .B(men_men_n228_), .Y(men_men_n1951_));
  NO2        u1902(.A(men_men_n1951_), .B(men_men_n1949_), .Y(men_men_n1952_));
  NOi21      u1903(.An(men_men_n710_), .B(men_men_n1005_), .Y(men_men_n1953_));
  NA3        u1904(.A(men_men_n1953_), .B(men_men_n1090_), .C(men_men_n872_), .Y(men_men_n1954_));
  OAI210     u1905(.A0(men_men_n1370_), .A1(men_men_n1681_), .B0(men_men_n1954_), .Y(men_men_n1955_));
  OAI210     u1906(.A0(men_men_n1955_), .A1(men_men_n1952_), .B0(men_men_n1129_), .Y(men_men_n1956_));
  OAI210     u1907(.A0(men_men_n448_), .A1(men_men_n51_), .B0(men_men_n1024_), .Y(men_men_n1957_));
  AOI220     u1908(.A0(men_men_n1957_), .A1(men_men_n465_), .B0(men_men_n448_), .B1(men_men_n390_), .Y(men_men_n1958_));
  NO2        u1909(.A(men_men_n1958_), .B(men_men_n153_), .Y(men_men_n1959_));
  NA2        u1910(.A(men_men_n162_), .B(men_men_n71_), .Y(men_men_n1960_));
  OAI210     u1911(.A0(men_men_n1862_), .A1(men_men_n1960_), .B0(men_men_n53_), .Y(men_men_n1961_));
  OAI220     u1912(.A0(men_men_n690_), .A1(men_men_n263_), .B0(men_men_n686_), .B1(x6), .Y(men_men_n1962_));
  NO2        u1913(.A(men_men_n304_), .B(x4), .Y(men_men_n1963_));
  AOI220     u1914(.A0(men_men_n1963_), .A1(men_men_n365_), .B0(men_men_n1962_), .B1(x4), .Y(men_men_n1964_));
  NO3        u1915(.A(men_men_n1964_), .B(men_men_n325_), .C(x5), .Y(men_men_n1965_));
  NO2        u1916(.A(men_men_n710_), .B(men_men_n57_), .Y(men_men_n1966_));
  OAI210     u1917(.A0(men_men_n1966_), .A1(men_men_n1917_), .B0(men_men_n450_), .Y(men_men_n1967_));
  AOI220     u1918(.A0(men_men_n667_), .A1(men_men_n736_), .B0(men_men_n497_), .B1(men_men_n238_), .Y(men_men_n1968_));
  AOI210     u1919(.A0(men_men_n1968_), .A1(men_men_n1967_), .B0(men_men_n258_), .Y(men_men_n1969_));
  NO4        u1920(.A(men_men_n1969_), .B(men_men_n1965_), .C(men_men_n1961_), .D(men_men_n1959_), .Y(men_men_n1970_));
  AOI220     u1921(.A0(men_men_n1970_), .A1(men_men_n1956_), .B0(men_men_n1948_), .B1(men_men_n1937_), .Y(men_men_n1971_));
  AOI210     u1922(.A0(men_men_n1925_), .A1(x3), .B0(men_men_n1971_), .Y(men29));
  OAI210     u1923(.A0(men_men_n558_), .A1(men_men_n264_), .B0(men_men_n731_), .Y(men_men_n1973_));
  NA2        u1924(.A(men_men_n751_), .B(men_men_n1054_), .Y(men_men_n1974_));
  AO210      u1925(.A0(men_men_n1168_), .A1(men_men_n1177_), .B0(men_men_n1974_), .Y(men_men_n1975_));
  AOI210     u1926(.A0(men_men_n182_), .A1(men_men_n166_), .B0(men_men_n710_), .Y(men_men_n1976_));
  AOI210     u1927(.A0(men_men_n1432_), .A1(men_men_n78_), .B0(men_men_n1976_), .Y(men_men_n1977_));
  NA3        u1928(.A(men_men_n1977_), .B(men_men_n1975_), .C(men_men_n1973_), .Y(men_men_n1978_));
  NO3        u1929(.A(men_men_n669_), .B(men_men_n1151_), .C(men_men_n50_), .Y(men_men_n1979_));
  NO3        u1930(.A(men_men_n1979_), .B(men_men_n1255_), .C(men_men_n558_), .Y(men_men_n1980_));
  NO2        u1931(.A(men_men_n446_), .B(men_men_n58_), .Y(men_men_n1981_));
  AOI220     u1932(.A0(men_men_n1981_), .A1(men_men_n1214_), .B0(men_men_n674_), .B1(men_men_n1388_), .Y(men_men_n1982_));
  OAI210     u1933(.A0(men_men_n1980_), .A1(men_men_n546_), .B0(men_men_n1982_), .Y(men_men_n1983_));
  AOI210     u1934(.A0(men_men_n1978_), .A1(x6), .B0(men_men_n1983_), .Y(men_men_n1984_));
  OAI210     u1935(.A0(x8), .A1(x4), .B0(x5), .Y(men_men_n1985_));
  NA2        u1936(.A(men_men_n1985_), .B(men_men_n112_), .Y(men_men_n1986_));
  NA2        u1937(.A(men_men_n304_), .B(men_men_n146_), .Y(men_men_n1987_));
  NA4        u1938(.A(men_men_n1987_), .B(men_men_n1986_), .C(men_men_n668_), .D(men_men_n64_), .Y(men_men_n1988_));
  AOI210     u1939(.A0(men_men_n1328_), .A1(men_men_n273_), .B0(men_men_n1732_), .Y(men_men_n1989_));
  AOI210     u1940(.A0(men_men_n1989_), .A1(men_men_n1988_), .B0(men_men_n892_), .Y(men_men_n1990_));
  NA4        u1941(.A(men_men_n669_), .B(men_men_n309_), .C(men_men_n182_), .D(men_men_n166_), .Y(men_men_n1991_));
  NA3        u1942(.A(men_men_n634_), .B(men_men_n297_), .C(men_men_n804_), .Y(men_men_n1992_));
  AOI210     u1943(.A0(men_men_n1992_), .A1(men_men_n1991_), .B0(men_men_n1214_), .Y(men_men_n1993_));
  OAI210     u1944(.A0(men_men_n899_), .A1(x8), .B0(x7), .Y(men_men_n1994_));
  NO2        u1945(.A(men_men_n1994_), .B(men_men_n127_), .Y(men_men_n1995_));
  OA210      u1946(.A0(men_men_n872_), .A1(men_men_n276_), .B0(men_men_n1985_), .Y(men_men_n1996_));
  OAI220     u1947(.A0(men_men_n1996_), .A1(men_men_n590_), .B0(men_men_n1512_), .B1(men_men_n397_), .Y(men_men_n1997_));
  NO4        u1948(.A(men_men_n1997_), .B(men_men_n1995_), .C(men_men_n1993_), .D(men_men_n1990_), .Y(men_men_n1998_));
  OAI210     u1949(.A0(men_men_n1984_), .A1(x2), .B0(men_men_n1998_), .Y(men_men_n1999_));
  NA3        u1950(.A(x6), .B(men_men_n50_), .C(x2), .Y(men_men_n2000_));
  OAI210     u1951(.A0(men_men_n1233_), .A1(men_men_n355_), .B0(men_men_n2000_), .Y(men_men_n2001_));
  NO3        u1952(.A(men_men_n448_), .B(x3), .C(x0), .Y(men_men_n2002_));
  AO220      u1953(.A0(men_men_n2002_), .A1(x5), .B0(men_men_n1932_), .B1(men_men_n81_), .Y(men_men_n2003_));
  AOI210     u1954(.A0(men_men_n2001_), .A1(men_men_n345_), .B0(men_men_n2003_), .Y(men_men_n2004_));
  NO3        u1955(.A(men_men_n703_), .B(men_men_n366_), .C(men_men_n140_), .Y(men_men_n2005_));
  AOI210     u1956(.A0(men_men_n730_), .A1(men_men_n617_), .B0(men_men_n2005_), .Y(men_men_n2006_));
  OAI210     u1957(.A0(men_men_n2004_), .A1(x7), .B0(men_men_n2006_), .Y(men_men_n2007_));
  AOI210     u1958(.A0(men_men_n1100_), .A1(men_men_n402_), .B0(men_men_n1416_), .Y(men_men_n2008_));
  NO2        u1959(.A(men_men_n146_), .B(x2), .Y(men_men_n2009_));
  OA210      u1960(.A0(men_men_n2009_), .A1(men_men_n632_), .B0(men_men_n669_), .Y(men_men_n2010_));
  OAI210     u1961(.A0(men_men_n2010_), .A1(men_men_n2008_), .B0(men_men_n68_), .Y(men_men_n2011_));
  NO2        u1962(.A(men_men_n198_), .B(men_men_n85_), .Y(men_men_n2012_));
  OAI210     u1963(.A0(men_men_n2012_), .A1(men_men_n790_), .B0(men_men_n1109_), .Y(men_men_n2013_));
  NA3        u1964(.A(men_men_n1950_), .B(men_men_n231_), .C(men_men_n83_), .Y(men_men_n2014_));
  NA3        u1965(.A(men_men_n2014_), .B(men_men_n2013_), .C(men_men_n2011_), .Y(men_men_n2015_));
  AOI210     u1966(.A0(men_men_n2007_), .A1(x8), .B0(men_men_n2015_), .Y(men_men_n2016_));
  OAI210     u1967(.A0(men_men_n446_), .A1(men_men_n247_), .B0(men_men_n969_), .Y(men_men_n2017_));
  OAI210     u1968(.A0(men_men_n2017_), .A1(men_men_n1130_), .B0(men_men_n679_), .Y(men_men_n2018_));
  NO3        u1969(.A(men_men_n1028_), .B(men_men_n356_), .C(men_men_n147_), .Y(men_men_n2019_));
  NA3        u1970(.A(men_men_n2019_), .B(men_men_n1308_), .C(men_men_n50_), .Y(men_men_n2020_));
  NO2        u1971(.A(men_men_n133_), .B(men_men_n93_), .Y(men_men_n2021_));
  AOI220     u1972(.A0(men_men_n2021_), .A1(men_men_n591_), .B0(men_men_n1931_), .B1(men_men_n362_), .Y(men_men_n2022_));
  NOi31      u1973(.An(men_men_n1131_), .B(men_men_n1881_), .C(men_men_n627_), .Y(men_men_n2023_));
  NA2        u1974(.A(men_men_n172_), .B(x4), .Y(men_men_n2024_));
  NO3        u1975(.A(men_men_n1485_), .B(men_men_n242_), .C(men_men_n71_), .Y(men_men_n2025_));
  AOI210     u1976(.A0(men_men_n2025_), .A1(men_men_n2024_), .B0(men_men_n2023_), .Y(men_men_n2026_));
  NA4        u1977(.A(men_men_n2026_), .B(men_men_n2022_), .C(men_men_n2020_), .D(men_men_n2018_), .Y(men_men_n2027_));
  NO4        u1978(.A(men_men_n1233_), .B(men_men_n170_), .C(men_men_n55_), .D(men_men_n71_), .Y(men_men_n2028_));
  NO4        u1979(.A(men_men_n1208_), .B(men_men_n506_), .C(men_men_n1388_), .D(men_men_n108_), .Y(men_men_n2029_));
  OAI210     u1980(.A0(men_men_n2029_), .A1(men_men_n2028_), .B0(men_men_n110_), .Y(men_men_n2030_));
  AOI210     u1981(.A0(men_men_n308_), .A1(x4), .B0(men_men_n192_), .Y(men_men_n2031_));
  OAI210     u1982(.A0(men_men_n2031_), .A1(men_men_n1981_), .B0(men_men_n725_), .Y(men_men_n2032_));
  OR3        u1983(.A(men_men_n1753_), .B(men_men_n1441_), .C(men_men_n1092_), .Y(men_men_n2033_));
  NA2        u1984(.A(men_men_n1932_), .B(men_men_n811_), .Y(men_men_n2034_));
  OA220      u1985(.A0(men_men_n2034_), .A1(men_men_n247_), .B0(men_men_n583_), .B1(men_men_n1795_), .Y(men_men_n2035_));
  NA4        u1986(.A(men_men_n2035_), .B(men_men_n2033_), .C(men_men_n2032_), .D(men_men_n2030_), .Y(men_men_n2036_));
  AOI210     u1987(.A0(men_men_n2027_), .A1(men_men_n293_), .B0(men_men_n2036_), .Y(men_men_n2037_));
  OAI210     u1988(.A0(men_men_n2016_), .A1(x1), .B0(men_men_n2037_), .Y(men_men_n2038_));
  AO210      u1989(.A0(men_men_n1999_), .A1(x1), .B0(men_men_n2038_), .Y(men30));
  NO3        u1990(.A(men_men_n1779_), .B(men_men_n579_), .C(men_men_n99_), .Y(men_men_n2040_));
  NO3        u1991(.A(men_men_n1149_), .B(men_men_n136_), .C(men_men_n386_), .Y(men_men_n2041_));
  AOI210     u1992(.A0(men_men_n725_), .A1(men_men_n255_), .B0(men_men_n2041_), .Y(men_men_n2042_));
  AOI210     u1993(.A0(men_men_n2042_), .A1(men_men_n2040_), .B0(men_men_n56_), .Y(men_men_n2043_));
  NA2        u1994(.A(men_men_n816_), .B(men_men_n343_), .Y(men_men_n2044_));
  NA2        u1995(.A(men_men_n2044_), .B(men_men_n1371_), .Y(men_men_n2045_));
  OAI210     u1996(.A0(men_men_n2045_), .A1(men_men_n2043_), .B0(men_men_n110_), .Y(men_men_n2046_));
  OAI210     u1997(.A0(men_men_n1005_), .A1(men_men_n573_), .B0(men_men_n679_), .Y(men_men_n2047_));
  AOI220     u1998(.A0(men_men_n451_), .A1(men_men_n945_), .B0(men_men_n329_), .B1(men_men_n459_), .Y(men_men_n2048_));
  AOI210     u1999(.A0(men_men_n2048_), .A1(men_men_n2047_), .B0(men_men_n258_), .Y(men_men_n2049_));
  NO3        u2000(.A(men_men_n282_), .B(men_men_n124_), .C(x0), .Y(men_men_n2050_));
  AOI210     u2001(.A0(men_men_n508_), .A1(x6), .B0(men_men_n2050_), .Y(men_men_n2051_));
  AOI220     u2002(.A0(men_men_n1145_), .A1(men_men_n426_), .B0(men_men_n763_), .B1(men_men_n92_), .Y(men_men_n2052_));
  OAI220     u2003(.A0(men_men_n2052_), .A1(men_men_n247_), .B0(men_men_n2051_), .B1(men_men_n54_), .Y(men_men_n2053_));
  NA2        u2004(.A(men_men_n163_), .B(men_men_n71_), .Y(men_men_n2054_));
  AO210      u2005(.A0(men_men_n572_), .A1(men_men_n522_), .B0(x5), .Y(men_men_n2055_));
  AOI210     u2006(.A0(men_men_n2054_), .A1(men_men_n722_), .B0(men_men_n2055_), .Y(men_men_n2056_));
  AOI210     u2007(.A0(men_men_n1610_), .A1(men_men_n50_), .B0(men_men_n459_), .Y(men_men_n2057_));
  NA2        u2008(.A(men_men_n197_), .B(x2), .Y(men_men_n2058_));
  OA220      u2009(.A0(men_men_n2058_), .A1(men_men_n2057_), .B0(men_men_n277_), .B1(x6), .Y(men_men_n2059_));
  OAI210     u2010(.A0(x7), .A1(x6), .B0(x1), .Y(men_men_n2060_));
  NA3        u2011(.A(men_men_n57_), .B(x4), .C(men_men_n59_), .Y(men_men_n2061_));
  AOI220     u2012(.A0(men_men_n2061_), .A1(men_men_n1378_), .B0(men_men_n2060_), .B1(men_men_n1820_), .Y(men_men_n2062_));
  NO3        u2013(.A(men_men_n1374_), .B(men_men_n345_), .C(men_men_n1030_), .Y(men_men_n2063_));
  NO2        u2014(.A(men_men_n520_), .B(men_men_n865_), .Y(men_men_n2064_));
  NOi21      u2015(.An(men_men_n2064_), .B(men_men_n850_), .Y(men_men_n2065_));
  NO3        u2016(.A(men_men_n1308_), .B(men_men_n233_), .C(men_men_n652_), .Y(men_men_n2066_));
  NO4        u2017(.A(men_men_n2066_), .B(men_men_n2065_), .C(men_men_n2063_), .D(men_men_n2062_), .Y(men_men_n2067_));
  OAI210     u2018(.A0(men_men_n2059_), .A1(men_men_n758_), .B0(men_men_n2067_), .Y(men_men_n2068_));
  NO4        u2019(.A(men_men_n2068_), .B(men_men_n2056_), .C(men_men_n2053_), .D(men_men_n2049_), .Y(men_men_n2069_));
  AOI210     u2020(.A0(men_men_n2069_), .A1(men_men_n2046_), .B0(x8), .Y(men_men_n2070_));
  NO3        u2021(.A(men_men_n495_), .B(men_men_n787_), .C(men_men_n53_), .Y(men_men_n2071_));
  OAI220     u2022(.A0(men_men_n1795_), .A1(men_men_n345_), .B0(men_men_n487_), .B1(men_men_n587_), .Y(men_men_n2072_));
  OAI210     u2023(.A0(men_men_n2072_), .A1(men_men_n2071_), .B0(x6), .Y(men_men_n2073_));
  OAI210     u2024(.A0(men_men_n1045_), .A1(men_men_n541_), .B0(men_men_n816_), .Y(men_men_n2074_));
  OAI210     u2025(.A0(men_men_n1742_), .A1(men_men_n332_), .B0(men_men_n126_), .Y(men_men_n2075_));
  AOI210     u2026(.A0(men_men_n381_), .A1(men_men_n230_), .B0(men_men_n72_), .Y(men_men_n2076_));
  AOI210     u2027(.A0(men_men_n1005_), .A1(men_men_n749_), .B0(men_men_n2076_), .Y(men_men_n2077_));
  NA4        u2028(.A(men_men_n2077_), .B(men_men_n2075_), .C(men_men_n2074_), .D(men_men_n2073_), .Y(men_men_n2078_));
  NA2        u2029(.A(men_men_n1097_), .B(men_men_n59_), .Y(men_men_n2079_));
  AOI210     u2030(.A0(men_men_n926_), .A1(men_men_n496_), .B0(men_men_n685_), .Y(men_men_n2080_));
  OAI220     u2031(.A0(men_men_n2080_), .A1(men_men_n308_), .B0(men_men_n2079_), .B1(men_men_n486_), .Y(men_men_n2081_));
  AOI210     u2032(.A0(men_men_n2078_), .A1(x8), .B0(men_men_n2081_), .Y(men_men_n2082_));
  NO2        u2033(.A(men_men_n2082_), .B(men_men_n57_), .Y(men_men_n2083_));
  NA2        u2034(.A(men_men_n437_), .B(men_men_n850_), .Y(men_men_n2084_));
  NO2        u2035(.A(men_men_n925_), .B(men_men_n665_), .Y(men_men_n2085_));
  AOI210     u2036(.A0(men_men_n2085_), .A1(men_men_n2084_), .B0(men_men_n448_), .Y(men_men_n2086_));
  NO3        u2037(.A(men_men_n640_), .B(men_men_n411_), .C(men_men_n1149_), .Y(men_men_n2087_));
  NO3        u2038(.A(men_men_n2087_), .B(men_men_n1261_), .C(men_men_n1388_), .Y(men_men_n2088_));
  AOI210     u2039(.A0(men_men_n305_), .A1(x1), .B0(men_men_n147_), .Y(men_men_n2089_));
  NO2        u2040(.A(men_men_n311_), .B(x5), .Y(men_men_n2090_));
  NO2        u2041(.A(men_men_n2090_), .B(men_men_n858_), .Y(men_men_n2091_));
  OAI220     u2042(.A0(men_men_n2091_), .A1(men_men_n1064_), .B0(men_men_n2089_), .B1(men_men_n207_), .Y(men_men_n2092_));
  NO3        u2043(.A(men_men_n2092_), .B(men_men_n2088_), .C(men_men_n2086_), .Y(men_men_n2093_));
  NA2        u2044(.A(men_men_n967_), .B(men_men_n82_), .Y(men_men_n2094_));
  AO210      u2045(.A0(men_men_n2094_), .A1(men_men_n1611_), .B0(x3), .Y(men_men_n2095_));
  NO2        u2046(.A(men_men_n219_), .B(men_men_n56_), .Y(men_men_n2096_));
  OAI220     u2047(.A0(men_men_n381_), .A1(men_men_n1261_), .B0(men_men_n356_), .B1(men_men_n233_), .Y(men_men_n2097_));
  AOI220     u2048(.A0(men_men_n2097_), .A1(x2), .B0(men_men_n2096_), .B1(men_men_n1625_), .Y(men_men_n2098_));
  AOI210     u2049(.A0(men_men_n2098_), .A1(men_men_n2095_), .B0(men_men_n263_), .Y(men_men_n2099_));
  NO3        u2050(.A(men_men_n821_), .B(men_men_n704_), .C(men_men_n166_), .Y(men_men_n2100_));
  OAI210     u2051(.A0(men_men_n2100_), .A1(men_men_n2676_), .B0(men_men_n154_), .Y(men_men_n2101_));
  NA3        u2052(.A(x5), .B(x4), .C(men_men_n59_), .Y(men_men_n2102_));
  AOI210     u2053(.A0(men_men_n2102_), .A1(men_men_n1316_), .B0(men_men_n542_), .Y(men_men_n2103_));
  AOI210     u2054(.A0(men_men_n1336_), .A1(x2), .B0(men_men_n2103_), .Y(men_men_n2104_));
  AOI210     u2055(.A0(men_men_n2104_), .A1(men_men_n2101_), .B0(men_men_n50_), .Y(men_men_n2105_));
  NA3        u2056(.A(men_men_n1482_), .B(men_men_n1140_), .C(men_men_n479_), .Y(men_men_n2106_));
  AOI210     u2057(.A0(men_men_n2106_), .A1(men_men_n2094_), .B0(men_men_n613_), .Y(men_men_n2107_));
  AOI210     u2058(.A0(men_men_n1030_), .A1(x1), .B0(men_men_n1328_), .Y(men_men_n2108_));
  OAI220     u2059(.A0(men_men_n309_), .A1(x4), .B0(men_men_n51_), .B1(x6), .Y(men_men_n2109_));
  NO2        u2060(.A(men_men_n122_), .B(men_men_n112_), .Y(men_men_n2110_));
  AOI220     u2061(.A0(men_men_n2110_), .A1(men_men_n2109_), .B0(men_men_n1170_), .B1(men_men_n627_), .Y(men_men_n2111_));
  OAI210     u2062(.A0(men_men_n2108_), .A1(men_men_n490_), .B0(men_men_n2111_), .Y(men_men_n2112_));
  NO4        u2063(.A(men_men_n2112_), .B(men_men_n2107_), .C(men_men_n2105_), .D(men_men_n2099_), .Y(men_men_n2113_));
  OAI210     u2064(.A0(men_men_n2093_), .A1(men_men_n133_), .B0(men_men_n2113_), .Y(men_men_n2114_));
  NO3        u2065(.A(men_men_n2114_), .B(men_men_n2083_), .C(men_men_n2070_), .Y(men31));
  NA2        u2066(.A(men_men_n991_), .B(men_men_n357_), .Y(men_men_n2116_));
  NO2        u2067(.A(men_men_n452_), .B(men_men_n679_), .Y(men_men_n2117_));
  AOI210     u2068(.A0(men_men_n2117_), .A1(men_men_n2116_), .B0(men_men_n58_), .Y(men_men_n2118_));
  NO2        u2069(.A(men_men_n789_), .B(men_men_n56_), .Y(men_men_n2119_));
  AOI220     u2070(.A0(men_men_n2119_), .A1(x2), .B0(men_men_n91_), .B1(x0), .Y(men_men_n2120_));
  NA3        u2071(.A(men_men_n2120_), .B(men_men_n2034_), .C(men_men_n1859_), .Y(men_men_n2121_));
  OAI210     u2072(.A0(men_men_n2121_), .A1(men_men_n2118_), .B0(men_men_n53_), .Y(men_men_n2122_));
  INV        u2073(.A(men_men_n679_), .Y(men_men_n2123_));
  NO3        u2074(.A(men_men_n1963_), .B(men_men_n1932_), .C(men_men_n893_), .Y(men_men_n2124_));
  OA220      u2075(.A0(men_men_n2124_), .A1(men_men_n479_), .B0(men_men_n2123_), .B1(men_men_n1475_), .Y(men_men_n2125_));
  AOI210     u2076(.A0(men_men_n2125_), .A1(men_men_n2122_), .B0(men_men_n108_), .Y(men_men_n2126_));
  NO2        u2077(.A(men_men_n502_), .B(men_men_n75_), .Y(men_men_n2127_));
  NA2        u2078(.A(men_men_n448_), .B(men_men_n57_), .Y(men_men_n2128_));
  AOI210     u2079(.A0(men_men_n308_), .A1(men_men_n86_), .B0(men_men_n2128_), .Y(men_men_n2129_));
  OAI210     u2080(.A0(men_men_n2129_), .A1(men_men_n2127_), .B0(men_men_n774_), .Y(men_men_n2130_));
  NO4        u2081(.A(men_men_n1166_), .B(men_men_n366_), .C(men_men_n1610_), .D(men_men_n67_), .Y(men_men_n2131_));
  AOI210     u2082(.A0(men_men_n1648_), .A1(men_men_n1363_), .B0(men_men_n446_), .Y(men_men_n2132_));
  OAI220     u2083(.A0(men_men_n1317_), .A1(men_men_n959_), .B0(men_men_n776_), .B1(men_men_n117_), .Y(men_men_n2133_));
  NO3        u2084(.A(men_men_n2133_), .B(men_men_n2132_), .C(men_men_n2131_), .Y(men_men_n2134_));
  AOI210     u2085(.A0(men_men_n2134_), .A1(men_men_n2130_), .B0(x5), .Y(men_men_n2135_));
  AOI220     u2086(.A0(men_men_n450_), .A1(men_men_n627_), .B0(men_men_n573_), .B1(men_men_n63_), .Y(men_men_n2136_));
  AOI210     u2087(.A0(men_men_n2136_), .A1(men_men_n583_), .B0(men_men_n1233_), .Y(men_men_n2137_));
  AOI220     u2088(.A0(men_men_n968_), .A1(men_men_n736_), .B0(men_men_n1149_), .B1(men_men_n121_), .Y(men_men_n2138_));
  OAI220     u2089(.A0(men_men_n2138_), .A1(men_men_n389_), .B0(men_men_n486_), .B1(men_men_n775_), .Y(men_men_n2139_));
  NO4        u2090(.A(men_men_n2139_), .B(men_men_n2137_), .C(men_men_n2135_), .D(men_men_n2126_), .Y(men_men_n2140_));
  NA2        u2091(.A(men_men_n496_), .B(men_men_n59_), .Y(men_men_n2141_));
  AOI210     u2092(.A0(men_men_n546_), .A1(men_men_n2141_), .B0(men_men_n139_), .Y(men_men_n2142_));
  OAI210     u2093(.A0(men_men_n104_), .A1(men_men_n276_), .B0(men_men_n2079_), .Y(men_men_n2143_));
  OAI210     u2094(.A0(men_men_n2143_), .A1(men_men_n2142_), .B0(x7), .Y(men_men_n2144_));
  NO3        u2095(.A(men_men_n381_), .B(men_men_n55_), .C(x7), .Y(men_men_n2145_));
  OA210      u2096(.A0(men_men_n2145_), .A1(men_men_n1327_), .B0(men_men_n101_), .Y(men_men_n2146_));
  NA2        u2097(.A(men_men_n1094_), .B(men_men_n92_), .Y(men_men_n2147_));
  AOI210     u2098(.A0(men_men_n905_), .A1(men_men_n112_), .B0(men_men_n2147_), .Y(men_men_n2148_));
  NA2        u2099(.A(men_men_n1557_), .B(x6), .Y(men_men_n2149_));
  AOI210     u2100(.A0(men_men_n2149_), .A1(men_men_n292_), .B0(men_men_n108_), .Y(men_men_n2150_));
  NA2        u2101(.A(men_men_n1193_), .B(men_men_n321_), .Y(men_men_n2151_));
  AOI210     u2102(.A0(men_men_n2151_), .A1(men_men_n648_), .B0(men_men_n53_), .Y(men_men_n2152_));
  NO4        u2103(.A(men_men_n2152_), .B(men_men_n2150_), .C(men_men_n2148_), .D(men_men_n2146_), .Y(men_men_n2153_));
  AOI210     u2104(.A0(men_men_n2153_), .A1(men_men_n2144_), .B0(men_men_n689_), .Y(men_men_n2154_));
  NOi21      u2105(.An(men_men_n1769_), .B(men_men_n1068_), .Y(men_men_n2155_));
  OAI220     u2106(.A0(men_men_n2155_), .A1(men_men_n1934_), .B0(men_men_n927_), .B1(men_men_n2141_), .Y(men_men_n2156_));
  NA2        u2107(.A(men_men_n2156_), .B(x3), .Y(men_men_n2157_));
  AOI220     u2108(.A0(men_men_n1398_), .A1(x8), .B0(men_men_n60_), .B1(x1), .Y(men_men_n2158_));
  NO3        u2109(.A(men_men_n2158_), .B(men_men_n1121_), .C(x6), .Y(men_men_n2159_));
  AOI220     u2110(.A0(men_men_n617_), .A1(men_men_n411_), .B0(men_men_n496_), .B1(men_men_n78_), .Y(men_men_n2160_));
  NA2        u2111(.A(men_men_n118_), .B(men_men_n533_), .Y(men_men_n2161_));
  OAI220     u2112(.A0(men_men_n2161_), .A1(men_men_n1934_), .B0(men_men_n2160_), .B1(x4), .Y(men_men_n2162_));
  NO2        u2113(.A(men_men_n2162_), .B(men_men_n2159_), .Y(men_men_n2163_));
  AOI210     u2114(.A0(men_men_n2163_), .A1(men_men_n2157_), .B0(men_men_n185_), .Y(men_men_n2164_));
  NO4        u2115(.A(men_men_n618_), .B(men_men_n591_), .C(men_men_n705_), .D(men_men_n704_), .Y(men_men_n2165_));
  OAI210     u2116(.A0(men_men_n2165_), .A1(men_men_n1086_), .B0(x3), .Y(men_men_n2166_));
  NO4        u2117(.A(men_men_n807_), .B(men_men_n1233_), .C(men_men_n774_), .D(x5), .Y(men_men_n2167_));
  NO3        u2118(.A(x6), .B(men_men_n56_), .C(x1), .Y(men_men_n2168_));
  NA2        u2119(.A(men_men_n2168_), .B(men_men_n288_), .Y(men_men_n2169_));
  OAI210     u2120(.A0(men_men_n1904_), .A1(men_men_n381_), .B0(men_men_n2169_), .Y(men_men_n2170_));
  NA4        u2121(.A(men_men_n640_), .B(men_men_n178_), .C(x6), .D(men_men_n108_), .Y(men_men_n2171_));
  NO2        u2122(.A(men_men_n859_), .B(men_men_n251_), .Y(men_men_n2172_));
  NOi41      u2123(.An(men_men_n2171_), .B(men_men_n2172_), .C(men_men_n2170_), .D(men_men_n2167_), .Y(men_men_n2173_));
  AOI210     u2124(.A0(men_men_n2173_), .A1(men_men_n2166_), .B0(men_men_n537_), .Y(men_men_n2174_));
  OAI210     u2125(.A0(men_men_n617_), .A1(men_men_n473_), .B0(men_men_n945_), .Y(men_men_n2175_));
  NO3        u2126(.A(men_men_n376_), .B(men_men_n77_), .C(men_men_n53_), .Y(men_men_n2176_));
  NO3        u2127(.A(men_men_n465_), .B(men_men_n351_), .C(men_men_n50_), .Y(men_men_n2177_));
  OAI210     u2128(.A0(men_men_n2177_), .A1(men_men_n2176_), .B0(men_men_n1167_), .Y(men_men_n2178_));
  AOI210     u2129(.A0(men_men_n2178_), .A1(men_men_n2175_), .B0(men_men_n395_), .Y(men_men_n2179_));
  NO2        u2130(.A(men_men_n216_), .B(men_men_n542_), .Y(men_men_n2180_));
  OAI210     u2131(.A0(men_men_n136_), .A1(x2), .B0(men_men_n2180_), .Y(men_men_n2181_));
  NA3        u2132(.A(men_men_n411_), .B(men_men_n330_), .C(men_men_n77_), .Y(men_men_n2182_));
  OA210      u2133(.A0(men_men_n246_), .A1(men_men_n229_), .B0(men_men_n2182_), .Y(men_men_n2183_));
  AOI210     u2134(.A0(men_men_n2183_), .A1(men_men_n2181_), .B0(men_men_n64_), .Y(men_men_n2184_));
  NA2        u2135(.A(men_men_n122_), .B(men_men_n57_), .Y(men_men_n2185_));
  AOI220     u2136(.A0(men_men_n1589_), .A1(men_men_n912_), .B0(men_men_n275_), .B1(x4), .Y(men_men_n2186_));
  AOI220     u2137(.A0(men_men_n1641_), .A1(men_men_n619_), .B0(men_men_n723_), .B1(men_men_n774_), .Y(men_men_n2187_));
  OAI220     u2138(.A0(men_men_n2187_), .A1(men_men_n2185_), .B0(men_men_n2186_), .B1(men_men_n190_), .Y(men_men_n2188_));
  OR3        u2139(.A(men_men_n2188_), .B(men_men_n2184_), .C(men_men_n2179_), .Y(men_men_n2189_));
  NO4        u2140(.A(men_men_n2189_), .B(men_men_n2174_), .C(men_men_n2164_), .D(men_men_n2154_), .Y(men_men_n2190_));
  OAI210     u2141(.A0(men_men_n2140_), .A1(x3), .B0(men_men_n2190_), .Y(men32));
  OAI210     u2142(.A0(men_men_n566_), .A1(men_men_n53_), .B0(men_men_n416_), .Y(men_men_n2192_));
  NA2        u2143(.A(men_men_n517_), .B(x2), .Y(men_men_n2193_));
  AOI210     u2144(.A0(men_men_n2193_), .A1(men_men_n2192_), .B0(men_men_n57_), .Y(men_men_n2194_));
  OAI210     u2145(.A0(men_men_n2194_), .A1(men_men_n790_), .B0(men_men_n56_), .Y(men_men_n2195_));
  OAI210     u2146(.A0(men_men_n1712_), .A1(men_men_n1460_), .B0(men_men_n1484_), .Y(men_men_n2196_));
  AOI210     u2147(.A0(men_men_n2119_), .A1(men_men_n279_), .B0(men_men_n2196_), .Y(men_men_n2197_));
  AOI210     u2148(.A0(men_men_n2197_), .A1(men_men_n2195_), .B0(men_men_n50_), .Y(men_men_n2198_));
  NA3        u2149(.A(men_men_n1558_), .B(men_men_n805_), .C(men_men_n291_), .Y(men_men_n2199_));
  NA2        u2150(.A(men_men_n746_), .B(men_men_n550_), .Y(men_men_n2200_));
  OAI220     u2151(.A0(men_men_n1063_), .A1(men_men_n231_), .B0(men_men_n686_), .B1(men_men_n207_), .Y(men_men_n2201_));
  NO3        u2152(.A(men_men_n377_), .B(men_men_n576_), .C(men_men_n811_), .Y(men_men_n2202_));
  NO3        u2153(.A(men_men_n1374_), .B(men_men_n587_), .C(men_men_n273_), .Y(men_men_n2203_));
  NO4        u2154(.A(men_men_n2203_), .B(men_men_n2202_), .C(men_men_n2201_), .D(men_men_n2200_), .Y(men_men_n2204_));
  AOI210     u2155(.A0(men_men_n2204_), .A1(men_men_n2199_), .B0(men_men_n140_), .Y(men_men_n2205_));
  OAI220     u2156(.A0(men_men_n404_), .A1(x7), .B0(men_men_n304_), .B1(men_men_n297_), .Y(men_men_n2206_));
  NA2        u2157(.A(men_men_n2206_), .B(men_men_n967_), .Y(men_men_n2207_));
  NO2        u2158(.A(men_men_n553_), .B(men_men_n865_), .Y(men_men_n2208_));
  AOI220     u2159(.A0(men_men_n2208_), .A1(men_men_n1884_), .B0(men_men_n534_), .B1(men_men_n129_), .Y(men_men_n2209_));
  AOI210     u2160(.A0(men_men_n2209_), .A1(men_men_n2207_), .B0(men_men_n110_), .Y(men_men_n2210_));
  NA3        u2161(.A(men_men_n1327_), .B(men_men_n1151_), .C(men_men_n117_), .Y(men_men_n2211_));
  AOI220     u2162(.A0(men_men_n1364_), .A1(men_men_n705_), .B0(men_men_n1247_), .B1(men_men_n1052_), .Y(men_men_n2212_));
  AOI210     u2163(.A0(men_men_n2212_), .A1(men_men_n2211_), .B0(men_men_n56_), .Y(men_men_n2213_));
  NA2        u2164(.A(men_men_n967_), .B(men_men_n57_), .Y(men_men_n2214_));
  NOi21      u2165(.An(men_men_n2214_), .B(men_men_n129_), .Y(men_men_n2215_));
  NA2        u2166(.A(men_men_n1020_), .B(men_men_n251_), .Y(men_men_n2216_));
  NO3        u2167(.A(men_men_n2216_), .B(men_men_n2215_), .C(men_men_n59_), .Y(men_men_n2217_));
  OR4        u2168(.A(men_men_n2217_), .B(men_men_n2213_), .C(men_men_n2210_), .D(men_men_n2205_), .Y(men_men_n2218_));
  OAI210     u2169(.A0(men_men_n2218_), .A1(men_men_n2198_), .B0(men_men_n108_), .Y(men_men_n2219_));
  NO3        u2170(.A(men_men_n1233_), .B(men_men_n144_), .C(men_men_n125_), .Y(men_men_n2220_));
  NO2        u2171(.A(men_men_n384_), .B(men_men_n55_), .Y(men_men_n2221_));
  NA2        u2172(.A(men_men_n2221_), .B(men_men_n116_), .Y(men_men_n2222_));
  OAI210     u2173(.A0(men_men_n636_), .A1(men_men_n593_), .B0(men_men_n816_), .Y(men_men_n2223_));
  NA2        u2174(.A(men_men_n2223_), .B(men_men_n2222_), .Y(men_men_n2224_));
  OAI210     u2175(.A0(men_men_n2224_), .A1(men_men_n2220_), .B0(x3), .Y(men_men_n2225_));
  OAI210     u2176(.A0(men_men_n899_), .A1(men_men_n273_), .B0(men_men_n50_), .Y(men_men_n2226_));
  AOI210     u2177(.A0(men_men_n62_), .A1(men_men_n110_), .B0(men_men_n2226_), .Y(men_men_n2227_));
  OAI210     u2178(.A0(men_men_n2227_), .A1(men_men_n1865_), .B0(men_men_n704_), .Y(men_men_n2228_));
  NO3        u2179(.A(men_men_n306_), .B(men_men_n172_), .C(men_men_n123_), .Y(men_men_n2229_));
  NO3        u2180(.A(men_men_n805_), .B(men_men_n364_), .C(men_men_n140_), .Y(men_men_n2230_));
  OAI210     u2181(.A0(men_men_n2230_), .A1(men_men_n2229_), .B0(men_men_n59_), .Y(men_men_n2231_));
  NA2        u2182(.A(men_men_n1155_), .B(men_men_n71_), .Y(men_men_n2232_));
  NO2        u2183(.A(men_men_n1938_), .B(men_men_n593_), .Y(men_men_n2233_));
  AOI210     u2184(.A0(men_men_n2233_), .A1(men_men_n1866_), .B0(men_men_n2232_), .Y(men_men_n2234_));
  NO2        u2185(.A(men_men_n276_), .B(men_men_n57_), .Y(men_men_n2235_));
  NO2        u2186(.A(men_men_n2235_), .B(men_men_n1012_), .Y(men_men_n2236_));
  NOi31      u2187(.An(men_men_n725_), .B(men_men_n2236_), .C(men_men_n282_), .Y(men_men_n2237_));
  NO3        u2188(.A(men_men_n1319_), .B(men_men_n216_), .C(men_men_n258_), .Y(men_men_n2238_));
  NO4        u2189(.A(men_men_n2238_), .B(men_men_n2237_), .C(men_men_n2234_), .D(x1), .Y(men_men_n2239_));
  NA4        u2190(.A(men_men_n2239_), .B(men_men_n2231_), .C(men_men_n2228_), .D(men_men_n2225_), .Y(men_men_n2240_));
  AO210      u2191(.A0(men_men_n1100_), .A1(men_men_n399_), .B0(men_men_n1015_), .Y(men_men_n2241_));
  NA3        u2192(.A(men_men_n1910_), .B(men_men_n557_), .C(men_men_n276_), .Y(men_men_n2242_));
  AOI210     u2193(.A0(men_men_n2242_), .A1(men_men_n2241_), .B0(men_men_n306_), .Y(men_men_n2243_));
  NA4        u2194(.A(men_men_n1270_), .B(men_men_n531_), .C(men_men_n389_), .D(men_men_n231_), .Y(men_men_n2244_));
  NO3        u2195(.A(men_men_n1441_), .B(men_men_n1015_), .C(x2), .Y(men_men_n2245_));
  NO2        u2196(.A(men_men_n1256_), .B(men_men_n387_), .Y(men_men_n2246_));
  NO2        u2197(.A(men_men_n1838_), .B(men_men_n64_), .Y(men_men_n2247_));
  NO4        u2198(.A(men_men_n2247_), .B(men_men_n2246_), .C(men_men_n2245_), .D(men_men_n53_), .Y(men_men_n2248_));
  NO3        u2199(.A(men_men_n469_), .B(men_men_n1094_), .C(men_men_n122_), .Y(men_men_n2249_));
  OAI220     u2200(.A0(men_men_n689_), .A1(men_men_n172_), .B0(men_men_n356_), .B1(men_men_n140_), .Y(men_men_n2250_));
  OAI210     u2201(.A0(men_men_n2250_), .A1(men_men_n2249_), .B0(men_men_n68_), .Y(men_men_n2251_));
  NO2        u2202(.A(men_men_n1985_), .B(men_men_n368_), .Y(men_men_n2252_));
  OAI210     u2203(.A0(men_men_n1871_), .A1(men_men_n611_), .B0(men_men_n2252_), .Y(men_men_n2253_));
  NA4        u2204(.A(men_men_n2253_), .B(men_men_n2251_), .C(men_men_n2248_), .D(men_men_n2244_), .Y(men_men_n2254_));
  OAI210     u2205(.A0(men_men_n2254_), .A1(men_men_n2243_), .B0(men_men_n2240_), .Y(men_men_n2255_));
  NO3        u2206(.A(men_men_n1220_), .B(men_men_n107_), .C(men_men_n71_), .Y(men_men_n2256_));
  NO2        u2207(.A(men_men_n566_), .B(men_men_n372_), .Y(men_men_n2257_));
  OAI210     u2208(.A0(men_men_n2256_), .A1(men_men_n1422_), .B0(men_men_n2257_), .Y(men_men_n2258_));
  NO3        u2209(.A(x8), .B(men_men_n71_), .C(x2), .Y(men_men_n2259_));
  OAI220     u2210(.A0(men_men_n2259_), .A1(men_men_n627_), .B0(men_men_n1432_), .B1(men_men_n91_), .Y(men_men_n2260_));
  AOI220     u2211(.A0(men_men_n558_), .A1(men_men_n816_), .B0(men_men_n679_), .B1(men_men_n256_), .Y(men_men_n2261_));
  AOI210     u2212(.A0(men_men_n2261_), .A1(men_men_n2260_), .B0(men_men_n266_), .Y(men_men_n2262_));
  NA2        u2213(.A(men_men_n1020_), .B(men_men_n1149_), .Y(men_men_n2263_));
  AOI210     u2214(.A0(men_men_n675_), .A1(men_men_n689_), .B0(men_men_n2263_), .Y(men_men_n2264_));
  AOI210     u2215(.A0(men_men_n591_), .A1(men_men_n627_), .B0(men_men_n695_), .Y(men_men_n2265_));
  NO2        u2216(.A(men_men_n2265_), .B(men_men_n1820_), .Y(men_men_n2266_));
  NO2        u2217(.A(men_men_n453_), .B(men_men_n434_), .Y(men_men_n2267_));
  NOi31      u2218(.An(men_men_n1504_), .B(men_men_n2267_), .C(men_men_n591_), .Y(men_men_n2268_));
  NO4        u2219(.A(men_men_n2268_), .B(men_men_n2266_), .C(men_men_n2264_), .D(men_men_n2262_), .Y(men_men_n2269_));
  NA4        u2220(.A(men_men_n2269_), .B(men_men_n2258_), .C(men_men_n2255_), .D(men_men_n2219_), .Y(men33));
  OAI210     u2221(.A0(men_men_n812_), .A1(x1), .B0(men_men_n201_), .Y(men_men_n2271_));
  OAI210     u2222(.A0(men_men_n2090_), .A1(men_men_n177_), .B0(men_men_n330_), .Y(men_men_n2272_));
  OAI220     u2223(.A0(men_men_n1081_), .A1(men_men_n811_), .B0(men_men_n1675_), .B1(men_men_n355_), .Y(men_men_n2273_));
  NA3        u2224(.A(men_men_n2273_), .B(men_men_n2272_), .C(men_men_n639_), .Y(men_men_n2274_));
  AOI210     u2225(.A0(men_men_n2271_), .A1(x5), .B0(men_men_n2274_), .Y(men_men_n2275_));
  NA2        u2226(.A(men_men_n230_), .B(men_men_n76_), .Y(men_men_n2276_));
  NA4        u2227(.A(men_men_n1749_), .B(men_men_n567_), .C(men_men_n247_), .D(x4), .Y(men_men_n2277_));
  AOI210     u2228(.A0(men_men_n2277_), .A1(men_men_n2276_), .B0(men_men_n355_), .Y(men_men_n2278_));
  OAI210     u2229(.A0(men_men_n437_), .A1(men_men_n270_), .B0(men_men_n53_), .Y(men_men_n2279_));
  AOI210     u2230(.A0(men_men_n2279_), .A1(men_men_n439_), .B0(men_men_n64_), .Y(men_men_n2280_));
  NA2        u2231(.A(men_men_n1663_), .B(men_men_n71_), .Y(men_men_n2281_));
  NO3        u2232(.A(men_men_n2281_), .B(men_men_n2280_), .C(men_men_n2278_), .Y(men_men_n2282_));
  OAI210     u2233(.A0(men_men_n2275_), .A1(x4), .B0(men_men_n2282_), .Y(men_men_n2283_));
  OAI210     u2234(.A0(men_men_n142_), .A1(x5), .B0(men_men_n240_), .Y(men_men_n2284_));
  NO2        u2235(.A(men_men_n967_), .B(men_men_n228_), .Y(men_men_n2285_));
  NA2        u2236(.A(men_men_n642_), .B(x7), .Y(men_men_n2286_));
  NO2        u2237(.A(men_men_n2286_), .B(men_men_n2285_), .Y(men_men_n2287_));
  AOI210     u2238(.A0(men_men_n2284_), .A1(men_men_n1028_), .B0(men_men_n2287_), .Y(men_men_n2288_));
  NA2        u2239(.A(men_men_n212_), .B(men_men_n958_), .Y(men_men_n2289_));
  AOI210     u2240(.A0(men_men_n2289_), .A1(men_men_n2214_), .B0(men_men_n214_), .Y(men_men_n2290_));
  NO2        u2241(.A(men_men_n1649_), .B(men_men_n959_), .Y(men_men_n2291_));
  OAI210     u2242(.A0(men_men_n865_), .A1(men_men_n51_), .B0(x6), .Y(men_men_n2292_));
  NO2        u2243(.A(men_men_n621_), .B(men_men_n508_), .Y(men_men_n2293_));
  NO4        u2244(.A(men_men_n2293_), .B(men_men_n2292_), .C(men_men_n2291_), .D(men_men_n2290_), .Y(men_men_n2294_));
  OAI210     u2245(.A0(men_men_n2288_), .A1(men_men_n50_), .B0(men_men_n2294_), .Y(men_men_n2295_));
  NA3        u2246(.A(men_men_n2295_), .B(men_men_n2283_), .C(men_men_n59_), .Y(men_men_n2296_));
  NA2        u2247(.A(men_men_n538_), .B(men_men_n109_), .Y(men_men_n2297_));
  NO3        u2248(.A(men_men_n1570_), .B(men_men_n376_), .C(x4), .Y(men_men_n2298_));
  AOI210     u2249(.A0(men_men_n2298_), .A1(men_men_n2297_), .B0(men_men_n440_), .Y(men_men_n2299_));
  NA2        u2250(.A(men_men_n814_), .B(men_men_n108_), .Y(men_men_n2300_));
  NA2        u2251(.A(men_men_n2300_), .B(men_men_n464_), .Y(men_men_n2301_));
  NO2        u2252(.A(men_men_n710_), .B(men_men_n377_), .Y(men_men_n2302_));
  NA2        u2253(.A(men_men_n504_), .B(men_men_n53_), .Y(men_men_n2303_));
  AOI210     u2254(.A0(men_men_n2302_), .A1(men_men_n2301_), .B0(men_men_n2303_), .Y(men_men_n2304_));
  OAI210     u2255(.A0(men_men_n2299_), .A1(men_men_n59_), .B0(men_men_n2304_), .Y(men_men_n2305_));
  AOI220     u2256(.A0(men_men_n689_), .A1(men_men_n237_), .B0(men_men_n389_), .B1(men_men_n231_), .Y(men_men_n2306_));
  NA2        u2257(.A(men_men_n732_), .B(men_men_n979_), .Y(men_men_n2307_));
  OAI210     u2258(.A0(men_men_n2307_), .A1(men_men_n2306_), .B0(men_men_n305_), .Y(men_men_n2308_));
  AOI210     u2259(.A0(men_men_n2119_), .A1(men_men_n215_), .B0(men_men_n53_), .Y(men_men_n2309_));
  NO2        u2260(.A(men_men_n140_), .B(men_men_n340_), .Y(men_men_n2310_));
  AOI220     u2261(.A0(men_men_n2310_), .A1(men_men_n998_), .B0(men_men_n674_), .B1(men_men_n355_), .Y(men_men_n2311_));
  NA2        u2262(.A(men_men_n448_), .B(men_men_n502_), .Y(men_men_n2312_));
  NO3        u2263(.A(men_men_n2312_), .B(men_men_n1034_), .C(men_men_n182_), .Y(men_men_n2313_));
  AOI210     u2264(.A0(men_men_n1796_), .A1(men_men_n1193_), .B0(men_men_n2313_), .Y(men_men_n2314_));
  NA4        u2265(.A(men_men_n2314_), .B(men_men_n2311_), .C(men_men_n2309_), .D(men_men_n2308_), .Y(men_men_n2315_));
  NA3        u2266(.A(men_men_n2315_), .B(men_men_n2305_), .C(men_men_n57_), .Y(men_men_n2316_));
  NAi21      u2267(.An(men_men_n1195_), .B(men_men_n492_), .Y(men_men_n2317_));
  NA4        u2268(.A(men_men_n642_), .B(men_men_n1308_), .C(men_men_n473_), .D(men_men_n50_), .Y(men_men_n2318_));
  OAI210     u2269(.A0(men_men_n2310_), .A1(men_men_n2064_), .B0(x2), .Y(men_men_n2319_));
  NA4        u2270(.A(men_men_n288_), .B(men_men_n155_), .C(men_men_n277_), .D(men_men_n122_), .Y(men_men_n2320_));
  NA3        u2271(.A(men_men_n2320_), .B(men_men_n2319_), .C(men_men_n2318_), .Y(men_men_n2321_));
  AO220      u2272(.A0(men_men_n2321_), .A1(x0), .B0(men_men_n2317_), .B1(men_men_n137_), .Y(men_men_n2322_));
  NA3        u2273(.A(men_men_n774_), .B(men_men_n355_), .C(men_men_n60_), .Y(men_men_n2323_));
  NO2        u2274(.A(men_men_n2259_), .B(men_men_n415_), .Y(men_men_n2324_));
  NA2        u2275(.A(men_men_n640_), .B(men_men_n520_), .Y(men_men_n2325_));
  OAI220     u2276(.A0(men_men_n2325_), .A1(men_men_n2324_), .B0(men_men_n2323_), .B1(men_men_n71_), .Y(men_men_n2326_));
  OAI210     u2277(.A0(men_men_n1534_), .A1(men_men_n351_), .B0(men_men_n111_), .Y(men_men_n2327_));
  AOI210     u2278(.A0(men_men_n591_), .A1(men_men_n469_), .B0(men_men_n137_), .Y(men_men_n2328_));
  OAI210     u2279(.A0(men_men_n2328_), .A1(men_men_n389_), .B0(men_men_n2327_), .Y(men_men_n2329_));
  OAI210     u2280(.A0(men_men_n2329_), .A1(men_men_n2326_), .B0(men_men_n102_), .Y(men_men_n2330_));
  NA2        u2281(.A(men_men_n130_), .B(men_men_n384_), .Y(men_men_n2331_));
  NA2        u2282(.A(men_men_n2331_), .B(men_men_n1824_), .Y(men_men_n2332_));
  NA2        u2283(.A(men_men_n1192_), .B(men_men_n711_), .Y(men_men_n2333_));
  AOI220     u2284(.A0(men_men_n2221_), .A1(men_men_n296_), .B0(men_men_n1364_), .B1(men_men_n1173_), .Y(men_men_n2334_));
  NA4        u2285(.A(men_men_n2334_), .B(men_men_n2333_), .C(men_men_n2332_), .D(men_men_n2330_), .Y(men_men_n2335_));
  AOI210     u2286(.A0(men_men_n2322_), .A1(x7), .B0(men_men_n2335_), .Y(men_men_n2336_));
  NA3        u2287(.A(men_men_n2336_), .B(men_men_n2316_), .C(men_men_n2296_), .Y(men34));
  NA2        u2288(.A(men_men_n434_), .B(x4), .Y(men_men_n2338_));
  NO2        u2289(.A(men_men_n1963_), .B(men_men_n858_), .Y(men_men_n2339_));
  AOI210     u2290(.A0(men_men_n2339_), .A1(men_men_n2338_), .B0(men_men_n322_), .Y(men_men_n2340_));
  NA2        u2291(.A(men_men_n288_), .B(men_men_n123_), .Y(men_men_n2341_));
  NO2        u2292(.A(men_men_n977_), .B(men_men_n2341_), .Y(men_men_n2342_));
  AOI210     u2293(.A0(men_men_n2044_), .A1(men_men_n546_), .B0(men_men_n139_), .Y(men_men_n2343_));
  NA2        u2294(.A(men_men_n1963_), .B(x0), .Y(men_men_n2344_));
  OAI210     u2295(.A0(men_men_n1833_), .A1(men_men_n981_), .B0(men_men_n2344_), .Y(men_men_n2345_));
  NO4        u2296(.A(men_men_n2345_), .B(men_men_n2343_), .C(men_men_n2342_), .D(men_men_n2340_), .Y(men_men_n2346_));
  NO2        u2297(.A(men_men_n2346_), .B(men_men_n479_), .Y(men_men_n2347_));
  NA2        u2298(.A(men_men_n734_), .B(x8), .Y(men_men_n2348_));
  AO210      u2299(.A0(men_men_n2348_), .A1(men_men_n489_), .B0(men_men_n664_), .Y(men_men_n2349_));
  NA2        u2300(.A(men_men_n674_), .B(men_men_n632_), .Y(men_men_n2350_));
  AOI210     u2301(.A0(men_men_n2350_), .A1(men_men_n2349_), .B0(men_men_n266_), .Y(men_men_n2351_));
  OAI210     u2302(.A0(men_men_n122_), .A1(men_men_n1055_), .B0(men_men_n1471_), .Y(men_men_n2352_));
  OAI210     u2303(.A0(men_men_n1610_), .A1(men_men_n58_), .B0(men_men_n2352_), .Y(men_men_n2353_));
  NA3        u2304(.A(men_men_n2353_), .B(men_men_n341_), .C(x8), .Y(men_men_n2354_));
  NA2        u2305(.A(men_men_n1592_), .B(men_men_n329_), .Y(men_men_n2355_));
  NA2        u2306(.A(men_men_n668_), .B(men_men_n322_), .Y(men_men_n2356_));
  NA2        u2307(.A(men_men_n133_), .B(x0), .Y(men_men_n2357_));
  NAi31      u2308(.An(men_men_n2357_), .B(men_men_n2356_), .C(men_men_n799_), .Y(men_men_n2358_));
  NA3        u2309(.A(men_men_n1605_), .B(men_men_n1406_), .C(men_men_n50_), .Y(men_men_n2359_));
  NA4        u2310(.A(men_men_n2359_), .B(men_men_n2358_), .C(men_men_n2355_), .D(men_men_n2354_), .Y(men_men_n2360_));
  NA2        u2311(.A(men_men_n1113_), .B(men_men_n749_), .Y(men_men_n2361_));
  NA3        u2312(.A(men_men_n1151_), .B(men_men_n166_), .C(men_men_n1097_), .Y(men_men_n2362_));
  AOI210     u2313(.A0(men_men_n2362_), .A1(men_men_n2361_), .B0(men_men_n759_), .Y(men_men_n2363_));
  AOI210     u2314(.A0(men_men_n1779_), .A1(men_men_n129_), .B0(men_men_n2363_), .Y(men_men_n2364_));
  AOI210     u2315(.A0(men_men_n558_), .A1(men_men_n816_), .B0(men_men_n255_), .Y(men_men_n2365_));
  OAI220     u2316(.A0(men_men_n2365_), .A1(men_men_n59_), .B0(men_men_n1124_), .B1(men_men_n55_), .Y(men_men_n2366_));
  NA3        u2317(.A(men_men_n2366_), .B(men_men_n734_), .C(men_men_n56_), .Y(men_men_n2367_));
  OAI210     u2318(.A0(men_men_n2364_), .A1(men_men_n140_), .B0(men_men_n2367_), .Y(men_men_n2368_));
  NO4        u2319(.A(men_men_n2368_), .B(men_men_n2360_), .C(men_men_n2351_), .D(men_men_n2347_), .Y(men_men_n2369_));
  NO2        u2320(.A(men_men_n312_), .B(men_men_n958_), .Y(men_men_n2370_));
  NO3        u2321(.A(men_men_n2370_), .B(men_men_n446_), .C(men_men_n329_), .Y(men_men_n2371_));
  NA2        u2322(.A(men_men_n784_), .B(men_men_n159_), .Y(men_men_n2372_));
  NO2        u2323(.A(men_men_n2235_), .B(men_men_n305_), .Y(men_men_n2373_));
  OAI220     u2324(.A0(men_men_n2373_), .A1(men_men_n1562_), .B0(men_men_n2372_), .B1(men_men_n1177_), .Y(men_men_n2374_));
  OAI210     u2325(.A0(men_men_n2374_), .A1(men_men_n2371_), .B0(x2), .Y(men_men_n2375_));
  OAI210     u2326(.A0(men_men_n868_), .A1(men_men_n372_), .B0(men_men_n2375_), .Y(men_men_n2376_));
  NA2        u2327(.A(men_men_n315_), .B(x4), .Y(men_men_n2377_));
  OAI220     u2328(.A0(men_men_n745_), .A1(men_men_n55_), .B0(men_men_n281_), .B1(men_men_n107_), .Y(men_men_n2378_));
  NO4        u2329(.A(men_men_n450_), .B(men_men_n77_), .C(x7), .D(x3), .Y(men_men_n2379_));
  NO2        u2330(.A(men_men_n1113_), .B(men_men_n289_), .Y(men_men_n2380_));
  NO4        u2331(.A(men_men_n2380_), .B(men_men_n2379_), .C(men_men_n2378_), .D(men_men_n2377_), .Y(men_men_n2381_));
  NA2        u2332(.A(men_men_n1247_), .B(men_men_n1054_), .Y(men_men_n2382_));
  NA3        u2333(.A(men_men_n1403_), .B(men_men_n258_), .C(x7), .Y(men_men_n2383_));
  NA2        u2334(.A(men_men_n2383_), .B(men_men_n2382_), .Y(men_men_n2384_));
  OAI210     u2335(.A0(men_men_n2384_), .A1(men_men_n2381_), .B0(men_men_n163_), .Y(men_men_n2385_));
  NA3        u2336(.A(men_men_n863_), .B(men_men_n87_), .C(x0), .Y(men_men_n2386_));
  NA4        u2337(.A(men_men_n2386_), .B(men_men_n1155_), .C(men_men_n298_), .D(men_men_n589_), .Y(men_men_n2387_));
  NA2        u2338(.A(men_men_n1159_), .B(men_men_n679_), .Y(men_men_n2388_));
  OAI210     u2339(.A0(men_men_n2388_), .A1(men_men_n267_), .B0(men_men_n2171_), .Y(men_men_n2389_));
  AOI220     u2340(.A0(men_men_n2389_), .A1(x7), .B0(men_men_n1019_), .B1(men_men_n665_), .Y(men_men_n2390_));
  OAI210     u2341(.A0(men_men_n2057_), .A1(men_men_n263_), .B0(men_men_n737_), .Y(men_men_n2391_));
  AOI220     u2342(.A0(men_men_n411_), .A1(x8), .B0(men_men_n92_), .B1(x2), .Y(men_men_n2392_));
  AOI210     u2343(.A0(men_men_n271_), .A1(men_men_n53_), .B0(men_men_n657_), .Y(men_men_n2393_));
  OAI220     u2344(.A0(men_men_n2393_), .A1(men_men_n97_), .B0(men_men_n2392_), .B1(men_men_n1350_), .Y(men_men_n2394_));
  AOI220     u2345(.A0(men_men_n2394_), .A1(men_men_n1328_), .B0(men_men_n2391_), .B1(men_men_n1519_), .Y(men_men_n2395_));
  NA4        u2346(.A(men_men_n2395_), .B(men_men_n2390_), .C(men_men_n2387_), .D(men_men_n2385_), .Y(men_men_n2396_));
  AOI210     u2347(.A0(men_men_n2376_), .A1(men_men_n816_), .B0(men_men_n2396_), .Y(men_men_n2397_));
  OAI210     u2348(.A0(men_men_n2369_), .A1(x2), .B0(men_men_n2397_), .Y(men35));
  NA2        u2349(.A(men_men_n508_), .B(men_men_n178_), .Y(men_men_n2399_));
  AOI220     u2350(.A0(men_men_n640_), .A1(men_men_n55_), .B0(men_men_n774_), .B1(men_men_n1227_), .Y(men_men_n2400_));
  AOI210     u2351(.A0(men_men_n2400_), .A1(men_men_n2399_), .B0(men_men_n71_), .Y(men_men_n2401_));
  NO3        u2352(.A(men_men_n516_), .B(men_men_n469_), .C(men_men_n340_), .Y(men_men_n2402_));
  OAI210     u2353(.A0(men_men_n2402_), .A1(men_men_n2401_), .B0(x2), .Y(men_men_n2403_));
  AOI210     u2354(.A0(men_men_n216_), .A1(x0), .B0(men_men_n275_), .Y(men_men_n2404_));
  OAI220     u2355(.A0(men_men_n2404_), .A1(men_men_n670_), .B0(men_men_n198_), .B1(x4), .Y(men_men_n2405_));
  NA2        u2356(.A(men_men_n2405_), .B(men_men_n137_), .Y(men_men_n2406_));
  NA3        u2357(.A(men_men_n411_), .B(x8), .C(men_men_n71_), .Y(men_men_n2407_));
  AOI210     u2358(.A0(men_men_n2407_), .A1(men_men_n1725_), .B0(men_men_n689_), .Y(men_men_n2408_));
  OAI210     u2359(.A0(men_men_n2323_), .A1(x6), .B0(men_men_n748_), .Y(men_men_n2409_));
  NO2        u2360(.A(men_men_n2409_), .B(men_men_n2408_), .Y(men_men_n2410_));
  NA3        u2361(.A(men_men_n2410_), .B(men_men_n2406_), .C(men_men_n2403_), .Y(men_men_n2411_));
  NAi21      u2362(.An(men_men_n1690_), .B(men_men_n1304_), .Y(men_men_n2412_));
  NA2        u2363(.A(men_men_n214_), .B(men_men_n576_), .Y(men_men_n2413_));
  NO2        u2364(.A(men_men_n434_), .B(men_men_n427_), .Y(men_men_n2414_));
  AOI220     u2365(.A0(men_men_n2414_), .A1(men_men_n2413_), .B0(men_men_n2412_), .B1(men_men_n56_), .Y(men_men_n2415_));
  NA2        u2366(.A(men_men_n763_), .B(men_men_n702_), .Y(men_men_n2416_));
  NO3        u2367(.A(men_men_n684_), .B(men_men_n55_), .C(x6), .Y(men_men_n2417_));
  OAI210     u2368(.A0(men_men_n2417_), .A1(men_men_n711_), .B0(men_men_n219_), .Y(men_men_n2418_));
  NA2        u2369(.A(men_men_n1336_), .B(men_men_n63_), .Y(men_men_n2419_));
  OAI210     u2370(.A0(men_men_n1077_), .A1(x6), .B0(men_men_n474_), .Y(men_men_n2420_));
  NA3        u2371(.A(men_men_n2420_), .B(men_men_n2419_), .C(men_men_n2418_), .Y(men_men_n2421_));
  NA3        u2372(.A(men_men_n1278_), .B(men_men_n751_), .C(x3), .Y(men_men_n2422_));
  NO3        u2373(.A(men_men_n2422_), .B(men_men_n686_), .C(men_men_n207_), .Y(men_men_n2423_));
  AOI210     u2374(.A0(men_men_n2421_), .A1(men_men_n50_), .B0(men_men_n2423_), .Y(men_men_n2424_));
  OAI210     u2375(.A0(men_men_n2416_), .A1(men_men_n2415_), .B0(men_men_n2424_), .Y(men_men_n2425_));
  AOI210     u2376(.A0(men_men_n2411_), .A1(men_men_n57_), .B0(men_men_n2425_), .Y(men_men_n2426_));
  NA2        u2377(.A(men_men_n967_), .B(men_men_n63_), .Y(men_men_n2427_));
  NO3        u2378(.A(men_men_n1077_), .B(men_men_n566_), .C(men_men_n123_), .Y(men_men_n2428_));
  NA2        u2379(.A(men_men_n156_), .B(men_men_n2428_), .Y(men_men_n2429_));
  AOI210     u2380(.A0(men_men_n2429_), .A1(men_men_n2427_), .B0(men_men_n50_), .Y(men_men_n2430_));
  NA4        u2381(.A(men_men_n469_), .B(men_men_n231_), .C(men_men_n874_), .D(men_men_n104_), .Y(men_men_n2431_));
  OAI210     u2382(.A0(men_men_n967_), .A1(men_men_n256_), .B0(men_men_n752_), .Y(men_men_n2432_));
  OAI210     u2383(.A0(men_men_n256_), .A1(men_men_n588_), .B0(men_men_n2168_), .Y(men_men_n2433_));
  NA3        u2384(.A(men_men_n2433_), .B(men_men_n2432_), .C(men_men_n2431_), .Y(men_men_n2434_));
  OAI210     u2385(.A0(men_men_n2434_), .A1(men_men_n2430_), .B0(men_men_n59_), .Y(men_men_n2435_));
  AOI210     u2386(.A0(men_men_n863_), .A1(men_men_n537_), .B0(men_men_n1910_), .Y(men_men_n2436_));
  AOI210     u2387(.A0(men_men_n566_), .A1(men_men_n610_), .B0(men_men_n2436_), .Y(men_men_n2437_));
  NO4        u2388(.A(men_men_n959_), .B(men_men_n566_), .C(men_men_n364_), .D(men_men_n409_), .Y(men_men_n2438_));
  XN2        u2389(.A(x4), .B(x3), .Y(men_men_n2439_));
  NO3        u2390(.A(men_men_n2439_), .B(men_men_n669_), .C(men_men_n311_), .Y(men_men_n2440_));
  NO3        u2391(.A(men_men_n2440_), .B(men_men_n2438_), .C(men_men_n1469_), .Y(men_men_n2441_));
  OAI210     u2392(.A0(men_men_n2437_), .A1(x3), .B0(men_men_n2441_), .Y(men_men_n2442_));
  NO3        u2393(.A(men_men_n745_), .B(men_men_n865_), .C(men_men_n276_), .Y(men_men_n2443_));
  OAI210     u2394(.A0(men_men_n2443_), .A1(men_men_n1469_), .B0(men_men_n50_), .Y(men_men_n2444_));
  INV        u2395(.A(men_men_n2444_), .Y(men_men_n2445_));
  AOI210     u2396(.A0(men_men_n2442_), .A1(men_men_n591_), .B0(men_men_n2445_), .Y(men_men_n2446_));
  AOI210     u2397(.A0(men_men_n1441_), .A1(men_men_n647_), .B0(men_men_n686_), .Y(men_men_n2447_));
  NO2        u2398(.A(men_men_n874_), .B(men_men_n56_), .Y(men_men_n2448_));
  OAI210     u2399(.A0(men_men_n1966_), .A1(men_men_n610_), .B0(men_men_n2259_), .Y(men_men_n2449_));
  OAI210     u2400(.A0(men_men_n2348_), .A1(men_men_n2448_), .B0(men_men_n2449_), .Y(men_men_n2450_));
  OAI210     u2401(.A0(men_men_n2450_), .A1(men_men_n2447_), .B0(men_men_n92_), .Y(men_men_n2451_));
  NO2        u2402(.A(men_men_n856_), .B(men_men_n666_), .Y(men_men_n2452_));
  NO2        u2403(.A(men_men_n289_), .B(x6), .Y(men_men_n2453_));
  OAI210     u2404(.A0(men_men_n2452_), .A1(men_men_n1787_), .B0(men_men_n2453_), .Y(men_men_n2454_));
  NA4        u2405(.A(men_men_n2454_), .B(men_men_n2451_), .C(men_men_n2446_), .D(men_men_n2435_), .Y(men_men_n2455_));
  NA4        u2406(.A(men_men_n618_), .B(men_men_n689_), .C(men_men_n433_), .D(x6), .Y(men_men_n2456_));
  AOI210     u2407(.A0(men_men_n2456_), .A1(men_men_n428_), .B0(x1), .Y(men_men_n2457_));
  NO2        u2408(.A(men_men_n732_), .B(men_men_n686_), .Y(men_men_n2458_));
  OAI210     u2409(.A0(men_men_n469_), .A1(men_men_n167_), .B0(men_men_n796_), .Y(men_men_n2459_));
  AOI210     u2410(.A0(men_men_n2459_), .A1(men_men_n1024_), .B0(men_men_n53_), .Y(men_men_n2460_));
  NO3        u2411(.A(men_men_n2460_), .B(men_men_n2458_), .C(men_men_n2457_), .Y(men_men_n2461_));
  NA3        u2412(.A(men_men_n1443_), .B(men_men_n1279_), .C(men_men_n820_), .Y(men_men_n2462_));
  AOI220     u2413(.A0(men_men_n1953_), .A1(men_men_n137_), .B0(men_men_n420_), .B1(men_men_n126_), .Y(men_men_n2463_));
  AOI210     u2414(.A0(men_men_n2463_), .A1(men_men_n2462_), .B0(men_men_n1512_), .Y(men_men_n2464_));
  NO2        u2415(.A(men_men_n640_), .B(x3), .Y(men_men_n2465_));
  NO3        u2416(.A(men_men_n697_), .B(men_men_n1610_), .C(x2), .Y(men_men_n2466_));
  AOI220     u2417(.A0(men_men_n2466_), .A1(men_men_n2465_), .B0(men_men_n1926_), .B1(men_men_n770_), .Y(men_men_n2467_));
  NA3        u2418(.A(x6), .B(x4), .C(x0), .Y(men_men_n2468_));
  OAI220     u2419(.A0(men_men_n2468_), .A1(men_men_n197_), .B0(men_men_n684_), .B1(men_men_n533_), .Y(men_men_n2469_));
  OAI220     u2420(.A0(men_men_n1317_), .A1(x8), .B0(men_men_n376_), .B1(men_men_n354_), .Y(men_men_n2470_));
  AOI220     u2421(.A0(men_men_n2470_), .A1(men_men_n420_), .B0(men_men_n2469_), .B1(men_men_n920_), .Y(men_men_n2471_));
  OAI210     u2422(.A0(men_men_n2467_), .A1(men_men_n1168_), .B0(men_men_n2471_), .Y(men_men_n2472_));
  NO2        u2423(.A(men_men_n2472_), .B(men_men_n2464_), .Y(men_men_n2473_));
  OAI210     u2424(.A0(men_men_n2461_), .A1(men_men_n315_), .B0(men_men_n2473_), .Y(men_men_n2474_));
  AOI210     u2425(.A0(men_men_n2455_), .A1(x5), .B0(men_men_n2474_), .Y(men_men_n2475_));
  OAI210     u2426(.A0(men_men_n2426_), .A1(x5), .B0(men_men_n2475_), .Y(men36));
  NO2        u2427(.A(men_men_n865_), .B(men_men_n304_), .Y(men_men_n2477_));
  NO3        u2428(.A(men_men_n122_), .B(men_men_n1055_), .C(men_men_n55_), .Y(men_men_n2478_));
  NO3        u2429(.A(men_men_n2478_), .B(men_men_n1985_), .C(men_men_n1077_), .Y(men_men_n2479_));
  OAI210     u2430(.A0(men_men_n2479_), .A1(men_men_n2477_), .B0(men_men_n110_), .Y(men_men_n2480_));
  OR4        u2431(.A(men_men_n960_), .B(men_men_n807_), .C(men_men_n379_), .D(men_men_n496_), .Y(men_men_n2481_));
  INV        u2432(.A(men_men_n1009_), .Y(men_men_n2482_));
  OAI210     u2433(.A0(men_men_n2221_), .A1(men_men_n2482_), .B0(men_men_n281_), .Y(men_men_n2483_));
  NA3        u2434(.A(men_men_n448_), .B(men_men_n228_), .C(men_men_n121_), .Y(men_men_n2484_));
  NA4        u2435(.A(men_men_n2484_), .B(men_men_n2483_), .C(men_men_n2481_), .D(men_men_n2480_), .Y(men_men_n2485_));
  NO2        u2436(.A(men_men_n998_), .B(x8), .Y(men_men_n2486_));
  NO3        u2437(.A(men_men_n2486_), .B(men_men_n995_), .C(men_men_n542_), .Y(men_men_n2487_));
  AOI220     u2438(.A0(men_men_n305_), .A1(x1), .B0(men_men_n136_), .B1(x6), .Y(men_men_n2488_));
  AOI210     u2439(.A0(men_men_n1097_), .A1(x6), .B0(men_men_n424_), .Y(men_men_n2489_));
  OAI220     u2440(.A0(men_men_n2489_), .A1(men_men_n363_), .B0(men_men_n2488_), .B1(men_men_n470_), .Y(men_men_n2490_));
  OAI210     u2441(.A0(men_men_n2490_), .A1(men_men_n2487_), .B0(men_men_n469_), .Y(men_men_n2491_));
  NA2        u2442(.A(men_men_n674_), .B(men_men_n496_), .Y(men_men_n2492_));
  AOI210     u2443(.A0(men_men_n2492_), .A1(men_men_n654_), .B0(men_men_n267_), .Y(men_men_n2493_));
  NO3        u2444(.A(men_men_n1881_), .B(men_men_n1609_), .C(men_men_n277_), .Y(men_men_n2494_));
  NO2        u2445(.A(men_men_n2427_), .B(men_men_n230_), .Y(men_men_n2495_));
  NO4        u2446(.A(men_men_n2495_), .B(men_men_n2494_), .C(men_men_n2493_), .D(men_men_n422_), .Y(men_men_n2496_));
  OAI210     u2447(.A0(men_men_n642_), .A1(men_men_n806_), .B0(men_men_n985_), .Y(men_men_n2497_));
  OAI220     u2448(.A0(men_men_n1654_), .A1(men_men_n1649_), .B0(men_men_n985_), .B1(men_men_n1097_), .Y(men_men_n2498_));
  AOI220     u2449(.A0(men_men_n2498_), .A1(men_men_n120_), .B0(men_men_n2497_), .B1(men_men_n632_), .Y(men_men_n2499_));
  NA3        u2450(.A(men_men_n2499_), .B(men_men_n2496_), .C(men_men_n2491_), .Y(men_men_n2500_));
  AOI210     u2451(.A0(men_men_n2485_), .A1(men_men_n341_), .B0(men_men_n2500_), .Y(men_men_n2501_));
  OAI210     u2452(.A0(men_men_n596_), .A1(men_men_n521_), .B0(men_men_n167_), .Y(men_men_n2502_));
  OAI210     u2453(.A0(men_men_n2000_), .A1(men_men_n70_), .B0(men_men_n2502_), .Y(men_men_n2503_));
  OAI210     u2454(.A0(men_men_n499_), .A1(men_men_n239_), .B0(men_men_n256_), .Y(men_men_n2504_));
  NO2        u2455(.A(men_men_n2009_), .B(men_men_n174_), .Y(men_men_n2505_));
  NA2        u2456(.A(men_men_n1214_), .B(men_men_n55_), .Y(men_men_n2506_));
  OAI210     u2457(.A0(men_men_n2506_), .A1(men_men_n2505_), .B0(men_men_n2504_), .Y(men_men_n2507_));
  OAI210     u2458(.A0(men_men_n2507_), .A1(men_men_n2503_), .B0(men_men_n899_), .Y(men_men_n2508_));
  AOI210     u2459(.A0(men_men_n107_), .A1(men_men_n110_), .B0(men_men_n343_), .Y(men_men_n2509_));
  NA2        u2460(.A(men_men_n674_), .B(men_men_n1610_), .Y(men_men_n2510_));
  OAI220     u2461(.A0(men_men_n2510_), .A1(men_men_n2509_), .B0(men_men_n748_), .B1(men_men_n1261_), .Y(men_men_n2511_));
  NO2        u2462(.A(men_men_n1406_), .B(men_men_n582_), .Y(men_men_n2512_));
  NO3        u2463(.A(men_men_n2512_), .B(men_men_n1795_), .C(men_men_n697_), .Y(men_men_n2513_));
  NOi31      u2464(.An(men_men_n2021_), .B(men_men_n2312_), .C(men_men_n758_), .Y(men_men_n2514_));
  NO3        u2465(.A(men_men_n2514_), .B(men_men_n2513_), .C(men_men_n2511_), .Y(men_men_n2515_));
  AOI210     u2466(.A0(men_men_n2515_), .A1(men_men_n2508_), .B0(x7), .Y(men_men_n2516_));
  NA2        u2467(.A(men_men_n136_), .B(men_men_n63_), .Y(men_men_n2517_));
  AOI210     u2468(.A0(men_men_n591_), .A1(men_men_n627_), .B0(men_men_n1193_), .Y(men_men_n2518_));
  NA3        u2469(.A(men_men_n2518_), .B(men_men_n2517_), .C(men_men_n892_), .Y(men_men_n2519_));
  NA2        u2470(.A(men_men_n2519_), .B(men_men_n508_), .Y(men_men_n2520_));
  AOI220     u2471(.A0(men_men_n1749_), .A1(men_men_n259_), .B0(men_men_n1054_), .B1(men_men_n126_), .Y(men_men_n2521_));
  NO2        u2472(.A(men_men_n2521_), .B(men_men_n448_), .Y(men_men_n2522_));
  NO2        u2473(.A(men_men_n409_), .B(men_men_n228_), .Y(men_men_n2523_));
  NO3        u2474(.A(men_men_n2523_), .B(men_men_n1283_), .C(men_men_n59_), .Y(men_men_n2524_));
  NO2        u2475(.A(men_men_n1231_), .B(x6), .Y(men_men_n2525_));
  NA3        u2476(.A(men_men_n1681_), .B(men_men_n281_), .C(men_men_n271_), .Y(men_men_n2526_));
  NA2        u2477(.A(men_men_n2526_), .B(men_men_n1635_), .Y(men_men_n2527_));
  NO4        u2478(.A(men_men_n2527_), .B(men_men_n2525_), .C(men_men_n2524_), .D(men_men_n2522_), .Y(men_men_n2528_));
  AOI210     u2479(.A0(men_men_n2528_), .A1(men_men_n2520_), .B0(men_men_n458_), .Y(men_men_n2529_));
  NO3        u2480(.A(men_men_n2439_), .B(men_men_n905_), .C(men_men_n507_), .Y(men_men_n2530_));
  AOI210     u2481(.A0(men_men_n1281_), .A1(men_men_n270_), .B0(men_men_n2530_), .Y(men_men_n2531_));
  OAI210     u2482(.A0(men_men_n872_), .A1(men_men_n276_), .B0(men_men_n399_), .Y(men_men_n2532_));
  NA2        u2483(.A(men_men_n1214_), .B(men_men_n172_), .Y(men_men_n2533_));
  NO2        u2484(.A(men_men_n617_), .B(men_men_n110_), .Y(men_men_n2534_));
  AO210      u2485(.A0(men_men_n2534_), .A1(men_men_n2533_), .B0(men_men_n1765_), .Y(men_men_n2535_));
  NO2        u2486(.A(men_men_n465_), .B(men_men_n421_), .Y(men_men_n2536_));
  AOI220     u2487(.A0(men_men_n2536_), .A1(men_men_n2535_), .B0(men_men_n2532_), .B1(men_men_n296_), .Y(men_men_n2537_));
  OAI210     u2488(.A0(men_men_n2531_), .A1(x1), .B0(men_men_n2537_), .Y(men_men_n2538_));
  NO3        u2489(.A(men_men_n2538_), .B(men_men_n2529_), .C(men_men_n2516_), .Y(men_men_n2539_));
  OAI210     u2490(.A0(men_men_n2501_), .A1(men_men_n57_), .B0(men_men_n2539_), .Y(men37));
  NA3        u2491(.A(men_men_n1074_), .B(men_men_n139_), .C(x3), .Y(men_men_n2541_));
  NA3        u2492(.A(men_men_n784_), .B(men_men_n159_), .C(men_men_n50_), .Y(men_men_n2542_));
  AOI210     u2493(.A0(men_men_n2542_), .A1(men_men_n2541_), .B0(men_men_n690_), .Y(men_men_n2543_));
  NO3        u2494(.A(men_men_n1074_), .B(men_men_n379_), .C(men_men_n515_), .Y(men_men_n2544_));
  OAI210     u2495(.A0(men_men_n2544_), .A1(men_men_n2543_), .B0(men_men_n56_), .Y(men_men_n2545_));
  AOI220     u2496(.A0(men_men_n605_), .A1(men_men_n749_), .B0(men_men_n469_), .B1(men_men_n1054_), .Y(men_men_n2546_));
  NO2        u2497(.A(men_men_n669_), .B(men_men_n181_), .Y(men_men_n2547_));
  OAI220     u2498(.A0(men_men_n2547_), .A1(men_men_n841_), .B0(men_men_n2546_), .B1(men_men_n110_), .Y(men_men_n2548_));
  NA2        u2499(.A(men_men_n2548_), .B(men_men_n71_), .Y(men_men_n2549_));
  NA2        u2500(.A(men_men_n1195_), .B(men_men_n1077_), .Y(men_men_n2550_));
  OAI210     u2501(.A0(men_men_n1216_), .A1(men_men_n191_), .B0(men_men_n459_), .Y(men_men_n2551_));
  NA4        u2502(.A(men_men_n2551_), .B(men_men_n2550_), .C(men_men_n2549_), .D(men_men_n2545_), .Y(men_men_n2552_));
  NA2        u2503(.A(men_men_n427_), .B(men_men_n136_), .Y(men_men_n2553_));
  NO2        u2504(.A(men_men_n1712_), .B(men_men_n109_), .Y(men_men_n2554_));
  AOI210     u2505(.A0(men_men_n1987_), .A1(men_men_n866_), .B0(men_men_n2554_), .Y(men_men_n2555_));
  OAI220     u2506(.A0(men_men_n2555_), .A1(men_men_n51_), .B0(men_men_n1611_), .B1(men_men_n2553_), .Y(men_men_n2556_));
  AOI210     u2507(.A0(men_men_n2552_), .A1(men_men_n68_), .B0(men_men_n2556_), .Y(men_men_n2557_));
  OAI210     u2508(.A0(men_men_n271_), .A1(men_men_n1101_), .B0(men_men_n490_), .Y(men_men_n2558_));
  NA3        u2509(.A(men_men_n2558_), .B(men_men_n267_), .C(men_men_n1055_), .Y(men_men_n2559_));
  OAI210     u2510(.A0(men_men_n231_), .A1(men_men_n219_), .B0(men_men_n1725_), .Y(men_men_n2560_));
  NA2        u2511(.A(men_men_n349_), .B(men_men_n275_), .Y(men_men_n2561_));
  NA3        u2512(.A(men_men_n405_), .B(men_men_n820_), .C(men_men_n110_), .Y(men_men_n2562_));
  NO2        u2513(.A(men_men_n534_), .B(men_men_n56_), .Y(men_men_n2563_));
  NA3        u2514(.A(men_men_n2563_), .B(men_men_n2562_), .C(men_men_n2561_), .Y(men_men_n2564_));
  AOI210     u2515(.A0(men_men_n2560_), .A1(men_men_n515_), .B0(men_men_n2564_), .Y(men_men_n2565_));
  NO2        u2516(.A(men_men_n1186_), .B(men_men_n276_), .Y(men_men_n2566_));
  OAI210     u2517(.A0(men_men_n296_), .A1(men_men_n265_), .B0(men_men_n2566_), .Y(men_men_n2567_));
  OAI210     u2518(.A0(men_men_n671_), .A1(men_men_n137_), .B0(x3), .Y(men_men_n2568_));
  AOI210     u2519(.A0(men_men_n671_), .A1(men_men_n368_), .B0(men_men_n2568_), .Y(men_men_n2569_));
  AOI210     u2520(.A0(men_men_n1610_), .A1(men_men_n50_), .B0(men_men_n349_), .Y(men_men_n2570_));
  OAI210     u2521(.A0(men_men_n2570_), .A1(men_men_n404_), .B0(men_men_n56_), .Y(men_men_n2571_));
  NO2        u2522(.A(men_men_n2571_), .B(men_men_n2569_), .Y(men_men_n2572_));
  AOI220     u2523(.A0(men_men_n2572_), .A1(men_men_n2567_), .B0(men_men_n2565_), .B1(men_men_n2559_), .Y(men_men_n2573_));
  OAI210     u2524(.A0(men_men_n2573_), .A1(men_men_n1763_), .B0(men_men_n102_), .Y(men_men_n2574_));
  NO2        u2525(.A(men_men_n2232_), .B(men_men_n55_), .Y(men_men_n2575_));
  OAI210     u2526(.A0(men_men_n2575_), .A1(men_men_n111_), .B0(men_men_n1824_), .Y(men_men_n2576_));
  NA2        u2527(.A(men_men_n178_), .B(men_men_n108_), .Y(men_men_n2577_));
  NA2        u2528(.A(men_men_n689_), .B(x6), .Y(men_men_n2578_));
  AOI210     u2529(.A0(men_men_n2578_), .A1(men_men_n489_), .B0(men_men_n2577_), .Y(men_men_n2579_));
  AOI210     u2530(.A0(men_men_n356_), .A1(men_men_n139_), .B0(men_men_n140_), .Y(men_men_n2580_));
  OAI210     u2531(.A0(men_men_n2580_), .A1(men_men_n2579_), .B0(men_men_n349_), .Y(men_men_n2581_));
  AOI210     u2532(.A0(men_men_n618_), .A1(men_men_n437_), .B0(men_men_n1293_), .Y(men_men_n2582_));
  NO3        u2533(.A(men_men_n2582_), .B(men_men_n267_), .C(men_men_n63_), .Y(men_men_n2583_));
  OAI220     u2534(.A0(men_men_n2348_), .A1(men_men_n487_), .B0(men_men_n2102_), .B1(men_men_n389_), .Y(men_men_n2584_));
  OAI210     u2535(.A0(men_men_n2584_), .A1(men_men_n2583_), .B0(men_men_n53_), .Y(men_men_n2585_));
  NO4        u2536(.A(men_men_n2357_), .B(men_men_n938_), .C(men_men_n438_), .D(men_men_n222_), .Y(men_men_n2586_));
  NO4        u2537(.A(men_men_n734_), .B(men_men_n606_), .C(men_men_n446_), .D(men_men_n1063_), .Y(men_men_n2587_));
  NO3        u2538(.A(men_men_n2587_), .B(men_men_n2586_), .C(men_men_n1069_), .Y(men_men_n2588_));
  NA4        u2539(.A(men_men_n2588_), .B(men_men_n2585_), .C(men_men_n2581_), .D(men_men_n2576_), .Y(men_men_n2589_));
  NO2        u2540(.A(men_men_n251_), .B(men_men_n84_), .Y(men_men_n2590_));
  NO2        u2541(.A(men_men_n279_), .B(men_men_n774_), .Y(men_men_n2591_));
  NO3        u2542(.A(men_men_n2591_), .B(men_men_n1214_), .C(men_men_n1233_), .Y(men_men_n2592_));
  OAI220     u2543(.A0(men_men_n2592_), .A1(men_men_n2590_), .B0(men_men_n469_), .B1(men_men_n85_), .Y(men_men_n2593_));
  OR2        u2544(.A(men_men_n944_), .B(men_men_n751_), .Y(men_men_n2594_));
  NA2        u2545(.A(men_men_n1227_), .B(men_men_n55_), .Y(men_men_n2595_));
  NOi21      u2546(.An(men_men_n2595_), .B(men_men_n390_), .Y(men_men_n2596_));
  AOI210     u2547(.A0(men_men_n2596_), .A1(men_men_n2594_), .B0(x1), .Y(men_men_n2597_));
  NA2        u2548(.A(men_men_n266_), .B(men_men_n84_), .Y(men_men_n2598_));
  AOI210     u2549(.A0(men_men_n1562_), .A1(men_men_n404_), .B0(men_men_n2598_), .Y(men_men_n2599_));
  NA2        u2550(.A(men_men_n1113_), .B(men_men_n62_), .Y(men_men_n2600_));
  NA2        u2551(.A(men_men_n1159_), .B(men_men_n174_), .Y(men_men_n2601_));
  OAI210     u2552(.A0(men_men_n2600_), .A1(men_men_n314_), .B0(men_men_n2601_), .Y(men_men_n2602_));
  NO3        u2553(.A(men_men_n2602_), .B(men_men_n2599_), .C(men_men_n2597_), .Y(men_men_n2603_));
  OAI210     u2554(.A0(men_men_n2603_), .A1(x6), .B0(men_men_n2593_), .Y(men_men_n2604_));
  AOI220     u2555(.A0(men_men_n2604_), .A1(men_men_n1471_), .B0(men_men_n2589_), .B1(men_men_n57_), .Y(men_men_n2605_));
  NA3        u2556(.A(men_men_n2605_), .B(men_men_n2574_), .C(men_men_n2557_), .Y(men38));
  AOI210     u2557(.A0(men_men_n1666_), .A1(men_men_n187_), .B0(men_men_n979_), .Y(men_men_n2607_));
  AOI210     u2558(.A0(men_men_n1231_), .A1(men_men_n581_), .B0(men_men_n1094_), .Y(men_men_n2608_));
  AOI210     u2559(.A0(men_men_n2595_), .A1(men_men_n1856_), .B0(men_men_n230_), .Y(men_men_n2609_));
  NO3        u2560(.A(men_men_n1303_), .B(men_men_n322_), .C(x8), .Y(men_men_n2610_));
  NO4        u2561(.A(men_men_n2610_), .B(men_men_n2609_), .C(men_men_n2608_), .D(men_men_n2607_), .Y(men_men_n2611_));
  NO2        u2562(.A(men_men_n2611_), .B(x6), .Y(men_men_n2612_));
  NA4        u2563(.A(men_men_n381_), .B(men_men_n258_), .C(men_men_n190_), .D(x8), .Y(men_men_n2613_));
  NA2        u2564(.A(men_men_n403_), .B(men_men_n108_), .Y(men_men_n2614_));
  AOI210     u2565(.A0(men_men_n2614_), .A1(men_men_n2613_), .B0(men_men_n140_), .Y(men_men_n2615_));
  AOI210     u2566(.A0(men_men_n438_), .A1(men_men_n408_), .B0(men_men_n1735_), .Y(men_men_n2616_));
  NO2        u2567(.A(men_men_n2616_), .B(men_men_n190_), .Y(men_men_n2617_));
  OAI210     u2568(.A0(men_men_n2617_), .A1(men_men_n2615_), .B0(x6), .Y(men_men_n2618_));
  NO2        u2569(.A(men_men_n248_), .B(men_men_n774_), .Y(men_men_n2619_));
  NO3        u2570(.A(men_men_n2619_), .B(men_men_n1690_), .C(men_men_n258_), .Y(men_men_n2620_));
  NO3        u2571(.A(x3), .B(men_men_n53_), .C(x0), .Y(men_men_n2621_));
  OAI210     u2572(.A0(men_men_n527_), .A1(x2), .B0(men_men_n2621_), .Y(men_men_n2622_));
  NA3        u2573(.A(men_men_n437_), .B(men_men_n427_), .C(men_men_n295_), .Y(men_men_n2623_));
  NA3        u2574(.A(men_men_n2623_), .B(men_men_n2622_), .C(men_men_n1814_), .Y(men_men_n2624_));
  OAI210     u2575(.A0(men_men_n2624_), .A1(men_men_n2620_), .B0(men_men_n816_), .Y(men_men_n2625_));
  NO2        u2576(.A(men_men_n606_), .B(men_men_n277_), .Y(men_men_n2626_));
  AN3        u2577(.A(men_men_n821_), .B(men_men_n784_), .C(x0), .Y(men_men_n2627_));
  OAI210     u2578(.A0(men_men_n2627_), .A1(men_men_n2626_), .B0(men_men_n330_), .Y(men_men_n2628_));
  OAI220     u2579(.A0(men_men_n606_), .A1(men_men_n277_), .B0(men_men_n820_), .B1(men_men_n93_), .Y(men_men_n2629_));
  OAI210     u2580(.A0(men_men_n689_), .A1(x0), .B0(men_men_n51_), .Y(men_men_n2630_));
  AOI210     u2581(.A0(men_men_n587_), .A1(x4), .B0(men_men_n229_), .Y(men_men_n2631_));
  AOI220     u2582(.A0(men_men_n2631_), .A1(men_men_n2630_), .B0(men_men_n2629_), .B1(men_men_n405_), .Y(men_men_n2632_));
  NA4        u2583(.A(men_men_n2632_), .B(men_men_n2628_), .C(men_men_n2625_), .D(men_men_n2618_), .Y(men_men_n2633_));
  OAI210     u2584(.A0(men_men_n2633_), .A1(men_men_n2612_), .B0(x7), .Y(men_men_n2634_));
  AOI210     u2585(.A0(men_men_n377_), .A1(x1), .B0(men_men_n1239_), .Y(men_men_n2635_));
  NO2        u2586(.A(men_men_n2635_), .B(men_men_n51_), .Y(men_men_n2636_));
  AOI210     u2587(.A0(men_men_n92_), .A1(men_men_n71_), .B0(men_men_n2259_), .Y(men_men_n2637_));
  NA2        u2588(.A(men_men_n389_), .B(x3), .Y(men_men_n2638_));
  NO2        u2589(.A(men_men_n1755_), .B(men_men_n534_), .Y(men_men_n2639_));
  OAI210     u2590(.A0(men_men_n2638_), .A1(men_men_n2637_), .B0(men_men_n2639_), .Y(men_men_n2640_));
  OAI210     u2591(.A0(men_men_n2640_), .A1(men_men_n2636_), .B0(x4), .Y(men_men_n2641_));
  NO2        u2592(.A(men_men_n1766_), .B(men_men_n463_), .Y(men_men_n2642_));
  NO3        u2593(.A(men_men_n2642_), .B(men_men_n404_), .C(men_men_n120_), .Y(men_men_n2643_));
  AOI210     u2594(.A0(men_men_n1063_), .A1(men_men_n242_), .B0(men_men_n397_), .Y(men_men_n2644_));
  AO210      u2595(.A0(men_men_n1309_), .A1(x6), .B0(men_men_n2644_), .Y(men_men_n2645_));
  NO2        u2596(.A(men_men_n1428_), .B(men_men_n137_), .Y(men_men_n2646_));
  NA2        u2597(.A(men_men_n1963_), .B(men_men_n325_), .Y(men_men_n2647_));
  OAI220     u2598(.A0(men_men_n2647_), .A1(men_men_n1082_), .B0(men_men_n2646_), .B1(men_men_n1838_), .Y(men_men_n2648_));
  NO3        u2599(.A(men_men_n2648_), .B(men_men_n2645_), .C(men_men_n2643_), .Y(men_men_n2649_));
  AOI210     u2600(.A0(men_men_n2649_), .A1(men_men_n2641_), .B0(men_men_n108_), .Y(men_men_n2650_));
  NA3        u2601(.A(men_men_n1953_), .B(men_men_n606_), .C(men_men_n163_), .Y(men_men_n2651_));
  NO2        u2602(.A(men_men_n2651_), .B(men_men_n231_), .Y(men_men_n2652_));
  AOI210     u2603(.A0(men_men_n508_), .A1(men_men_n496_), .B0(men_men_n685_), .Y(men_men_n2653_));
  OAI220     u2604(.A0(men_men_n2653_), .A1(men_men_n470_), .B0(men_men_n198_), .B1(men_men_n119_), .Y(men_men_n2654_));
  OAI210     u2605(.A0(men_men_n2654_), .A1(men_men_n2652_), .B0(x0), .Y(men_men_n2655_));
  NA3        u2606(.A(men_men_n408_), .B(men_men_n820_), .C(men_men_n277_), .Y(men_men_n2656_));
  AOI210     u2607(.A0(men_men_n2656_), .A1(men_men_n717_), .B0(men_men_n2216_), .Y(men_men_n2657_));
  NA2        u2608(.A(men_men_n1131_), .B(men_men_n958_), .Y(men_men_n2658_));
  NA4        u2609(.A(men_men_n684_), .B(men_men_n606_), .C(men_men_n178_), .D(x3), .Y(men_men_n2659_));
  AOI210     u2610(.A0(men_men_n2659_), .A1(men_men_n2658_), .B0(men_men_n502_), .Y(men_men_n2660_));
  NO4        u2611(.A(men_men_n1421_), .B(men_men_n523_), .C(men_men_n1233_), .D(men_men_n774_), .Y(men_men_n2661_));
  OAI220     u2612(.A0(men_men_n1785_), .A1(men_men_n2300_), .B0(men_men_n229_), .B1(men_men_n149_), .Y(men_men_n2662_));
  NO4        u2613(.A(men_men_n2662_), .B(men_men_n2661_), .C(men_men_n2660_), .D(men_men_n2657_), .Y(men_men_n2663_));
  NA2        u2614(.A(men_men_n2663_), .B(men_men_n2655_), .Y(men_men_n2664_));
  OAI210     u2615(.A0(men_men_n2664_), .A1(men_men_n2650_), .B0(men_men_n57_), .Y(men_men_n2665_));
  AOI210     u2616(.A0(men_men_n1825_), .A1(men_men_n277_), .B0(men_men_n686_), .Y(men_men_n2666_));
  OAI210     u2617(.A0(men_men_n1762_), .A1(men_men_n214_), .B0(men_men_n498_), .Y(men_men_n2667_));
  OAI210     u2618(.A0(men_men_n2667_), .A1(men_men_n2666_), .B0(men_men_n634_), .Y(men_men_n2668_));
  OAI220     u2619(.A0(men_men_n1769_), .A1(men_men_n277_), .B0(men_men_n257_), .B1(men_men_n104_), .Y(men_men_n2669_));
  NA2        u2620(.A(men_men_n1875_), .B(men_men_n357_), .Y(men_men_n2670_));
  OAI220     u2621(.A0(men_men_n2670_), .A1(men_men_n642_), .B0(men_men_n696_), .B1(men_men_n149_), .Y(men_men_n2671_));
  AOI210     u2622(.A0(men_men_n2669_), .A1(men_men_n998_), .B0(men_men_n2671_), .Y(men_men_n2672_));
  NA4        u2623(.A(men_men_n2672_), .B(men_men_n2668_), .C(men_men_n2665_), .D(men_men_n2634_), .Y(men39));
  INV        u2624(.A(men_men_n123_), .Y(men_men_n2676_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
  VOTADOR g14(.A(ori14), .B(mai14), .C(men14), .Y(z14));
  VOTADOR g15(.A(ori15), .B(mai15), .C(men15), .Y(z15));
  VOTADOR g16(.A(ori16), .B(mai16), .C(men16), .Y(z16));
  VOTADOR g17(.A(ori17), .B(mai17), .C(men17), .Y(z17));
  VOTADOR g18(.A(ori18), .B(mai18), .C(men18), .Y(z18));
  VOTADOR g19(.A(ori19), .B(mai19), .C(men19), .Y(z19));
  VOTADOR g20(.A(ori20), .B(mai20), .C(men20), .Y(z20));
  VOTADOR g21(.A(ori21), .B(mai21), .C(men21), .Y(z21));
  VOTADOR g22(.A(ori22), .B(mai22), .C(men22), .Y(z22));
  VOTADOR g23(.A(ori23), .B(mai23), .C(men23), .Y(z23));
  VOTADOR g24(.A(ori24), .B(mai24), .C(men24), .Y(z24));
  VOTADOR g25(.A(ori25), .B(mai25), .C(men25), .Y(z25));
  VOTADOR g26(.A(ori26), .B(mai26), .C(men26), .Y(z26));
  VOTADOR g27(.A(ori27), .B(mai27), .C(men27), .Y(z27));
  VOTADOR g28(.A(ori28), .B(mai28), .C(men28), .Y(z28));
  VOTADOR g29(.A(ori29), .B(mai29), .C(men29), .Y(z29));
  VOTADOR g30(.A(ori30), .B(mai30), .C(men30), .Y(z30));
  VOTADOR g31(.A(ori31), .B(mai31), .C(men31), .Y(z31));
  VOTADOR g32(.A(ori32), .B(mai32), .C(men32), .Y(z32));
  VOTADOR g33(.A(ori33), .B(mai33), .C(men33), .Y(z33));
  VOTADOR g34(.A(ori34), .B(mai34), .C(men34), .Y(z34));
  VOTADOR g35(.A(ori35), .B(mai35), .C(men35), .Y(z35));
  VOTADOR g36(.A(ori36), .B(mai36), .C(men36), .Y(z36));
  VOTADOR g37(.A(ori37), .B(mai37), .C(men37), .Y(z37));
  VOTADOR g38(.A(ori38), .B(mai38), .C(men38), .Y(z38));
  VOTADOR g39(.A(ori39), .B(mai39), .C(men39), .Y(z39));
endmodule