//Benchmark atmr_alu4_1266_0.0156

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n893_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1110_, men_men_n1111_, men_men_n1112_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NA3        o034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n57_));
  NO2        o035(.A(i_1_), .B(i_6_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  OAI210     o037(.A0(ori_ori_n59_), .A1(ori_ori_n58_), .B0(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n61_));
  NAi21      o039(.An(i_2_), .B(i_7_), .Y(ori_ori_n62_));
  INV        o040(.A(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NA3        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .C(ori_ori_n31_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_1_), .B(i_10_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(i_6_), .Y(ori_ori_n67_));
  NAi31      o045(.An(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n61_), .Y(ori_ori_n68_));
  NA2        o046(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_1_), .B(i_6_), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n71_), .B(ori_ori_n25_), .Y(ori_ori_n72_));
  INV        o050(.A(i_0_), .Y(ori_ori_n73_));
  NAi21      o051(.An(i_5_), .B(i_10_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_5_), .B(i_9_), .Y(ori_ori_n75_));
  AOI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n73_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  OAI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n68_), .B0(i_0_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_12_), .B(i_5_), .Y(ori_ori_n80_));
  NA2        o058(.A(i_2_), .B(i_8_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n81_), .B(ori_ori_n58_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_9_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_3_), .B(i_7_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(ori_ori_n63_), .Y(ori_ori_n85_));
  INV        o063(.A(i_6_), .Y(ori_ori_n86_));
  OR4        o064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NO2        o066(.A(i_2_), .B(i_7_), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n88_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  OAI210     o068(.A0(ori_ori_n85_), .A1(ori_ori_n82_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NAi21      o069(.An(i_6_), .B(i_10_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_6_), .B(i_9_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n93_), .A1(ori_ori_n92_), .B0(ori_ori_n63_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_2_), .B(i_6_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n96_), .B(ori_ori_n94_), .Y(ori_ori_n97_));
  AOI210     o075(.A0(ori_ori_n97_), .A1(ori_ori_n91_), .B0(ori_ori_n80_), .Y(ori_ori_n98_));
  AN3        o076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n99_));
  NAi21      o077(.An(i_6_), .B(i_11_), .Y(ori_ori_n100_));
  NO2        o078(.A(i_5_), .B(i_8_), .Y(ori_ori_n101_));
  NOi21      o079(.An(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  AOI220     o080(.A0(ori_ori_n102_), .A1(ori_ori_n62_), .B0(ori_ori_n99_), .B1(ori_ori_n32_), .Y(ori_ori_n103_));
  INV        o081(.A(i_7_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n46_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o083(.A(i_0_), .B(i_5_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n86_), .Y(ori_ori_n107_));
  NA2        o085(.A(i_12_), .B(i_3_), .Y(ori_ori_n108_));
  INV        o086(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NA3        o087(.A(ori_ori_n109_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n110_));
  NAi21      o088(.An(i_7_), .B(i_11_), .Y(ori_ori_n111_));
  NO3        o089(.A(ori_ori_n111_), .B(ori_ori_n92_), .C(ori_ori_n53_), .Y(ori_ori_n112_));
  AN2        o090(.A(i_2_), .B(i_10_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(i_7_), .Y(ori_ori_n114_));
  OR2        o092(.A(ori_ori_n80_), .B(ori_ori_n58_), .Y(ori_ori_n115_));
  NO2        o093(.A(i_8_), .B(ori_ori_n104_), .Y(ori_ori_n116_));
  NO3        o094(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(ori_ori_n114_), .Y(ori_ori_n117_));
  NA2        o095(.A(i_12_), .B(i_7_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n63_), .B(ori_ori_n26_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(i_0_), .Y(ori_ori_n120_));
  NA2        o098(.A(i_11_), .B(i_12_), .Y(ori_ori_n121_));
  OAI210     o099(.A0(ori_ori_n120_), .A1(ori_ori_n118_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n122_), .B(ori_ori_n117_), .Y(ori_ori_n123_));
  NAi41      o101(.An(ori_ori_n112_), .B(ori_ori_n123_), .C(ori_ori_n110_), .D(ori_ori_n103_), .Y(ori_ori_n124_));
  NOi21      o102(.An(i_1_), .B(i_5_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(i_11_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n127_));
  NA2        o105(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n129_), .B(ori_ori_n46_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n93_), .B(ori_ori_n92_), .Y(ori_ori_n131_));
  NAi21      o109(.An(i_3_), .B(i_8_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n62_), .Y(ori_ori_n133_));
  NOi31      o111(.An(ori_ori_n133_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_1_), .B(ori_ori_n86_), .Y(ori_ori_n135_));
  NO2        o113(.A(i_6_), .B(i_5_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(i_3_), .Y(ori_ori_n137_));
  AO210      o115(.A0(ori_ori_n137_), .A1(ori_ori_n47_), .B0(ori_ori_n135_), .Y(ori_ori_n138_));
  OAI220     o116(.A0(ori_ori_n138_), .A1(ori_ori_n111_), .B0(ori_ori_n134_), .B1(ori_ori_n126_), .Y(ori_ori_n139_));
  NO3        o117(.A(ori_ori_n139_), .B(ori_ori_n124_), .C(ori_ori_n98_), .Y(ori_ori_n140_));
  NA3        o118(.A(ori_ori_n140_), .B(ori_ori_n79_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o119(.A(ori_ori_n63_), .B(ori_ori_n37_), .Y(ori_ori_n142_));
  INV        o120(.A(i_6_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(ori_ori_n142_), .Y(ori_ori_n144_));
  NA4        o122(.A(ori_ori_n144_), .B(ori_ori_n77_), .C(ori_ori_n69_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o123(.A(i_8_), .B(i_7_), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n146_), .B(i_6_), .Y(ori_ori_n147_));
  NO2        o125(.A(i_12_), .B(i_13_), .Y(ori_ori_n148_));
  NAi21      o126(.An(i_5_), .B(i_11_), .Y(ori_ori_n149_));
  NOi21      o127(.An(ori_ori_n148_), .B(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o128(.A(i_0_), .B(i_1_), .Y(ori_ori_n151_));
  NA2        o129(.A(i_2_), .B(i_3_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n152_), .B(i_4_), .Y(ori_ori_n153_));
  NA3        o131(.A(ori_ori_n153_), .B(ori_ori_n151_), .C(ori_ori_n150_), .Y(ori_ori_n154_));
  AN2        o132(.A(ori_ori_n148_), .B(ori_ori_n83_), .Y(ori_ori_n155_));
  NA2        o133(.A(i_1_), .B(i_5_), .Y(ori_ori_n156_));
  OR2        o134(.A(i_0_), .B(i_1_), .Y(ori_ori_n157_));
  NO3        o135(.A(ori_ori_n157_), .B(ori_ori_n80_), .C(i_13_), .Y(ori_ori_n158_));
  NAi32      o136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n159_));
  NAi21      o137(.An(ori_ori_n159_), .B(ori_ori_n158_), .Y(ori_ori_n160_));
  NOi21      o138(.An(i_4_), .B(i_10_), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n161_), .B(ori_ori_n40_), .Y(ori_ori_n162_));
  NO3        o140(.A(ori_ori_n73_), .B(i_2_), .C(i_1_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n160_), .B(ori_ori_n147_), .Y(ori_ori_n164_));
  NOi21      o142(.An(i_4_), .B(i_9_), .Y(ori_ori_n165_));
  NOi21      o143(.An(i_11_), .B(i_13_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n166_), .B(ori_ori_n165_), .Y(ori_ori_n167_));
  NO2        o145(.A(i_4_), .B(i_5_), .Y(ori_ori_n168_));
  NAi21      o146(.An(i_12_), .B(i_11_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n169_), .B(i_13_), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n73_), .B(ori_ori_n63_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(ori_ori_n46_), .Y(ori_ori_n172_));
  NA2        o150(.A(i_3_), .B(i_5_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n174_));
  NO2        o152(.A(i_13_), .B(i_10_), .Y(ori_ori_n175_));
  NA3        o153(.A(ori_ori_n175_), .B(ori_ori_n174_), .C(ori_ori_n44_), .Y(ori_ori_n176_));
  NO2        o154(.A(i_2_), .B(i_1_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n177_), .B(i_3_), .Y(ori_ori_n178_));
  NAi21      o156(.An(i_4_), .B(i_12_), .Y(ori_ori_n179_));
  INV        o157(.A(i_8_), .Y(ori_ori_n180_));
  NO3        o158(.A(i_3_), .B(ori_ori_n86_), .C(ori_ori_n48_), .Y(ori_ori_n181_));
  NA2        o159(.A(ori_ori_n181_), .B(ori_ori_n116_), .Y(ori_ori_n182_));
  NO3        o160(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n183_));
  NO3        o161(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n184_));
  NA2        o162(.A(i_12_), .B(ori_ori_n184_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n185_), .B(ori_ori_n182_), .Y(ori_ori_n186_));
  NO2        o164(.A(i_3_), .B(i_8_), .Y(ori_ori_n187_));
  NO3        o165(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n188_));
  NA3        o166(.A(ori_ori_n188_), .B(ori_ori_n187_), .C(ori_ori_n40_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n106_), .B(ori_ori_n58_), .Y(ori_ori_n190_));
  INV        o168(.A(ori_ori_n190_), .Y(ori_ori_n191_));
  NO2        o169(.A(i_13_), .B(i_9_), .Y(ori_ori_n192_));
  NAi21      o170(.An(i_12_), .B(i_3_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n191_), .B(ori_ori_n189_), .Y(ori_ori_n195_));
  AOI210     o173(.A0(ori_ori_n195_), .A1(i_7_), .B0(ori_ori_n186_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n196_), .B(i_4_), .Y(ori_ori_n197_));
  NAi21      o175(.An(i_12_), .B(i_7_), .Y(ori_ori_n198_));
  NA3        o176(.A(i_13_), .B(ori_ori_n180_), .C(i_10_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .Y(ori_ori_n200_));
  NA2        o178(.A(i_0_), .B(i_5_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n201_), .B(ori_ori_n107_), .Y(ori_ori_n202_));
  OAI220     o180(.A0(ori_ori_n202_), .A1(ori_ori_n178_), .B0(ori_ori_n172_), .B1(ori_ori_n137_), .Y(ori_ori_n203_));
  NAi31      o181(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n73_), .B(ori_ori_n26_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n46_), .B(ori_ori_n63_), .Y(ori_ori_n207_));
  INV        o185(.A(i_13_), .Y(ori_ori_n208_));
  NO2        o186(.A(i_12_), .B(ori_ori_n208_), .Y(ori_ori_n209_));
  NA3        o187(.A(ori_ori_n209_), .B(ori_ori_n183_), .C(ori_ori_n181_), .Y(ori_ori_n210_));
  INV        o188(.A(ori_ori_n210_), .Y(ori_ori_n211_));
  AOI220     o189(.A0(ori_ori_n211_), .A1(ori_ori_n146_), .B0(ori_ori_n203_), .B1(ori_ori_n200_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n213_));
  OR2        o191(.A(i_8_), .B(i_7_), .Y(ori_ori_n214_));
  INV        o192(.A(i_12_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n44_), .B(ori_ori_n215_), .Y(ori_ori_n216_));
  NO3        o194(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n217_));
  NA2        o195(.A(i_2_), .B(i_1_), .Y(ori_ori_n218_));
  NO3        o196(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n219_));
  NAi21      o197(.An(i_4_), .B(i_3_), .Y(ori_ori_n220_));
  NO2        o198(.A(i_0_), .B(i_6_), .Y(ori_ori_n221_));
  NOi41      o199(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n222_));
  NA2        o200(.A(ori_ori_n222_), .B(ori_ori_n221_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n218_), .B(ori_ori_n173_), .Y(ori_ori_n224_));
  NO2        o202(.A(i_11_), .B(ori_ori_n208_), .Y(ori_ori_n225_));
  NOi21      o203(.An(i_1_), .B(i_6_), .Y(ori_ori_n226_));
  NAi21      o204(.An(i_3_), .B(i_7_), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n215_), .B(i_9_), .Y(ori_ori_n228_));
  OR4        o206(.A(ori_ori_n228_), .B(ori_ori_n227_), .C(ori_ori_n226_), .D(ori_ori_n174_), .Y(ori_ori_n229_));
  NA2        o207(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n230_));
  NA2        o208(.A(i_3_), .B(i_9_), .Y(ori_ori_n231_));
  NAi21      o209(.An(i_7_), .B(i_10_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n232_), .B(ori_ori_n231_), .Y(ori_ori_n233_));
  NA3        o211(.A(ori_ori_n233_), .B(ori_ori_n230_), .C(ori_ori_n64_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n234_), .B(ori_ori_n229_), .Y(ori_ori_n235_));
  INV        o213(.A(ori_ori_n147_), .Y(ori_ori_n236_));
  NA2        o214(.A(ori_ori_n215_), .B(i_13_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n237_), .B(ori_ori_n75_), .Y(ori_ori_n238_));
  AOI220     o216(.A0(ori_ori_n238_), .A1(ori_ori_n236_), .B0(ori_ori_n235_), .B1(ori_ori_n225_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n214_), .B(ori_ori_n37_), .Y(ori_ori_n240_));
  NA2        o218(.A(i_12_), .B(i_6_), .Y(ori_ori_n241_));
  OR2        o219(.A(i_13_), .B(i_9_), .Y(ori_ori_n242_));
  NO3        o220(.A(ori_ori_n242_), .B(ori_ori_n241_), .C(ori_ori_n48_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n220_), .B(i_2_), .Y(ori_ori_n244_));
  NA3        o222(.A(ori_ori_n244_), .B(ori_ori_n243_), .C(ori_ori_n44_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n225_), .B(i_9_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n230_), .B(ori_ori_n64_), .Y(ori_ori_n247_));
  OAI210     o225(.A0(ori_ori_n247_), .A1(ori_ori_n246_), .B0(ori_ori_n245_), .Y(ori_ori_n248_));
  NO3        o226(.A(i_11_), .B(ori_ori_n208_), .C(ori_ori_n25_), .Y(ori_ori_n249_));
  NO2        o227(.A(ori_ori_n227_), .B(i_8_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n248_), .B(ori_ori_n240_), .Y(ori_ori_n251_));
  NA3        o229(.A(ori_ori_n251_), .B(ori_ori_n239_), .C(ori_ori_n212_), .Y(ori_ori_n252_));
  NO3        o230(.A(i_12_), .B(ori_ori_n208_), .C(ori_ori_n37_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n218_), .B(i_0_), .Y(ori_ori_n254_));
  NO2        o232(.A(i_2_), .B(ori_ori_n104_), .Y(ori_ori_n255_));
  AN2        o233(.A(i_3_), .B(i_10_), .Y(ori_ori_n256_));
  NO2        o234(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n252_), .B(ori_ori_n197_), .C(ori_ori_n164_), .Y(ori_ori_n259_));
  NO3        o237(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n260_));
  NO2        o238(.A(i_2_), .B(i_3_), .Y(ori_ori_n261_));
  OR2        o239(.A(i_0_), .B(i_5_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n157_), .B(ori_ori_n46_), .Y(ori_ori_n263_));
  NO2        o241(.A(i_12_), .B(i_10_), .Y(ori_ori_n264_));
  NOi21      o242(.An(i_5_), .B(i_0_), .Y(ori_ori_n265_));
  NA4        o243(.A(ori_ori_n84_), .B(ori_ori_n36_), .C(ori_ori_n86_), .D(i_8_), .Y(ori_ori_n266_));
  NO2        o244(.A(i_6_), .B(i_8_), .Y(ori_ori_n267_));
  NO2        o245(.A(i_1_), .B(i_7_), .Y(ori_ori_n268_));
  NOi21      o246(.An(ori_ori_n156_), .B(ori_ori_n107_), .Y(ori_ori_n269_));
  NO2        o247(.A(ori_ori_n269_), .B(ori_ori_n128_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(i_3_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n180_), .B(i_9_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n272_), .B(ori_ori_n190_), .Y(ori_ori_n273_));
  NO2        o251(.A(ori_ori_n273_), .B(ori_ori_n46_), .Y(ori_ori_n274_));
  INV        o252(.A(ori_ori_n274_), .Y(ori_ori_n275_));
  AOI210     o253(.A0(ori_ori_n275_), .A1(ori_ori_n271_), .B0(ori_ori_n162_), .Y(ori_ori_n276_));
  INV        o254(.A(ori_ori_n276_), .Y(ori_ori_n277_));
  NOi32      o255(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n278_));
  INV        o256(.A(ori_ori_n278_), .Y(ori_ori_n279_));
  NAi21      o257(.An(i_0_), .B(i_6_), .Y(ori_ori_n280_));
  NAi21      o258(.An(i_1_), .B(i_5_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n281_), .B(ori_ori_n280_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n25_), .Y(ori_ori_n283_));
  OAI210     o261(.A0(ori_ori_n283_), .A1(ori_ori_n159_), .B0(ori_ori_n223_), .Y(ori_ori_n284_));
  NAi41      o262(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n285_));
  OAI220     o263(.A0(ori_ori_n285_), .A1(ori_ori_n281_), .B0(ori_ori_n204_), .B1(ori_ori_n159_), .Y(ori_ori_n286_));
  AOI210     o264(.A0(ori_ori_n285_), .A1(ori_ori_n159_), .B0(ori_ori_n157_), .Y(ori_ori_n287_));
  NOi32      o265(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n288_));
  NAi21      o266(.An(i_6_), .B(i_1_), .Y(ori_ori_n289_));
  NA3        o267(.A(ori_ori_n289_), .B(ori_ori_n288_), .C(ori_ori_n46_), .Y(ori_ori_n290_));
  NO2        o268(.A(ori_ori_n290_), .B(i_0_), .Y(ori_ori_n291_));
  OR3        o269(.A(ori_ori_n291_), .B(ori_ori_n287_), .C(ori_ori_n286_), .Y(ori_ori_n292_));
  NO2        o270(.A(i_1_), .B(ori_ori_n104_), .Y(ori_ori_n293_));
  NAi21      o271(.An(i_3_), .B(i_4_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n294_), .B(i_9_), .Y(ori_ori_n295_));
  AN2        o273(.A(i_6_), .B(i_7_), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n296_), .A1(ori_ori_n293_), .B0(ori_ori_n295_), .Y(ori_ori_n297_));
  NA2        o275(.A(i_2_), .B(i_7_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n294_), .B(i_10_), .Y(ori_ori_n299_));
  NA3        o277(.A(ori_ori_n299_), .B(ori_ori_n298_), .C(ori_ori_n221_), .Y(ori_ori_n300_));
  AOI210     o278(.A0(ori_ori_n300_), .A1(ori_ori_n297_), .B0(ori_ori_n174_), .Y(ori_ori_n301_));
  AOI210     o279(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n302_));
  OAI210     o280(.A0(ori_ori_n302_), .A1(ori_ori_n177_), .B0(ori_ori_n299_), .Y(ori_ori_n303_));
  AOI220     o281(.A0(ori_ori_n299_), .A1(ori_ori_n268_), .B0(ori_ori_n217_), .B1(ori_ori_n177_), .Y(ori_ori_n304_));
  AOI210     o282(.A0(ori_ori_n304_), .A1(ori_ori_n303_), .B0(i_5_), .Y(ori_ori_n305_));
  NO4        o283(.A(ori_ori_n305_), .B(ori_ori_n301_), .C(ori_ori_n292_), .D(ori_ori_n284_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n306_), .B(ori_ori_n279_), .Y(ori_ori_n307_));
  NO2        o285(.A(ori_ori_n59_), .B(ori_ori_n25_), .Y(ori_ori_n308_));
  AN2        o286(.A(i_12_), .B(i_5_), .Y(ori_ori_n309_));
  NO2        o287(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n310_), .B(ori_ori_n309_), .Y(ori_ori_n311_));
  NO2        o289(.A(i_11_), .B(i_6_), .Y(ori_ori_n312_));
  NA3        o290(.A(ori_ori_n312_), .B(ori_ori_n263_), .C(ori_ori_n208_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n313_), .B(ori_ori_n311_), .Y(ori_ori_n314_));
  NO2        o292(.A(i_5_), .B(i_10_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n316_));
  NO2        o294(.A(ori_ori_n154_), .B(ori_ori_n86_), .Y(ori_ori_n317_));
  OAI210     o295(.A0(ori_ori_n317_), .A1(ori_ori_n314_), .B0(ori_ori_n316_), .Y(ori_ori_n318_));
  NO3        o296(.A(ori_ori_n86_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n319_));
  NO2        o297(.A(i_11_), .B(i_12_), .Y(ori_ori_n320_));
  NAi21      o298(.An(i_13_), .B(i_0_), .Y(ori_ori_n321_));
  INV        o299(.A(ori_ori_n318_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n44_), .B(ori_ori_n208_), .Y(ori_ori_n323_));
  NO3        o301(.A(i_1_), .B(i_12_), .C(ori_ori_n86_), .Y(ori_ori_n324_));
  NO2        o302(.A(i_0_), .B(i_11_), .Y(ori_ori_n325_));
  AN2        o303(.A(i_1_), .B(i_6_), .Y(ori_ori_n326_));
  NOi21      o304(.An(i_2_), .B(i_12_), .Y(ori_ori_n327_));
  NAi21      o305(.An(i_9_), .B(i_4_), .Y(ori_ori_n328_));
  OR2        o306(.A(i_13_), .B(i_10_), .Y(ori_ori_n329_));
  NO3        o307(.A(ori_ori_n329_), .B(ori_ori_n121_), .C(ori_ori_n328_), .Y(ori_ori_n330_));
  NO2        o308(.A(ori_ori_n167_), .B(ori_ori_n127_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n104_), .B(ori_ori_n25_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n253_), .B(ori_ori_n332_), .Y(ori_ori_n333_));
  NO2        o311(.A(ori_ori_n333_), .B(ori_ori_n269_), .Y(ori_ori_n334_));
  INV        o312(.A(ori_ori_n334_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n335_), .B(ori_ori_n26_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n173_), .B(ori_ori_n86_), .Y(ori_ori_n337_));
  NA2        o315(.A(ori_ori_n180_), .B(i_10_), .Y(ori_ori_n338_));
  NA3        o316(.A(ori_ori_n230_), .B(ori_ori_n64_), .C(i_2_), .Y(ori_ori_n339_));
  NO2        o317(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  NO2        o318(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n341_));
  INV        o319(.A(ori_ori_n340_), .Y(ori_ori_n342_));
  NO2        o320(.A(ori_ori_n342_), .B(ori_ori_n246_), .Y(ori_ori_n343_));
  NO4        o321(.A(ori_ori_n343_), .B(ori_ori_n336_), .C(ori_ori_n322_), .D(ori_ori_n307_), .Y(ori_ori_n344_));
  NO2        o322(.A(ori_ori_n63_), .B(i_4_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n73_), .B(i_13_), .Y(ori_ori_n346_));
  NA3        o324(.A(ori_ori_n346_), .B(ori_ori_n345_), .C(i_2_), .Y(ori_ori_n347_));
  NO2        o325(.A(i_10_), .B(i_9_), .Y(ori_ori_n348_));
  NAi21      o326(.An(i_12_), .B(i_8_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n349_), .B(i_3_), .Y(ori_ori_n350_));
  NA2        o328(.A(ori_ori_n350_), .B(ori_ori_n348_), .Y(ori_ori_n351_));
  NO2        o329(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n352_), .B(ori_ori_n107_), .Y(ori_ori_n353_));
  OAI220     o331(.A0(ori_ori_n353_), .A1(ori_ori_n189_), .B0(ori_ori_n351_), .B1(ori_ori_n347_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n258_), .B(i_0_), .Y(ori_ori_n355_));
  NO3        o333(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n241_), .B(ori_ori_n100_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n357_), .B(ori_ori_n356_), .Y(ori_ori_n358_));
  NA2        o336(.A(i_8_), .B(i_9_), .Y(ori_ori_n359_));
  AOI210     o337(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n360_));
  OR2        o338(.A(ori_ori_n360_), .B(ori_ori_n359_), .Y(ori_ori_n361_));
  NA2        o339(.A(ori_ori_n253_), .B(ori_ori_n190_), .Y(ori_ori_n362_));
  OAI220     o340(.A0(ori_ori_n362_), .A1(ori_ori_n361_), .B0(ori_ori_n358_), .B1(ori_ori_n355_), .Y(ori_ori_n363_));
  NA2        o341(.A(ori_ori_n225_), .B(ori_ori_n257_), .Y(ori_ori_n364_));
  NO3        o342(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n365_));
  INV        o343(.A(ori_ori_n365_), .Y(ori_ori_n366_));
  NA3        o344(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n367_));
  NA4        o345(.A(ori_ori_n149_), .B(ori_ori_n119_), .C(ori_ori_n80_), .D(ori_ori_n23_), .Y(ori_ori_n368_));
  OAI220     o346(.A0(ori_ori_n368_), .A1(ori_ori_n367_), .B0(ori_ori_n366_), .B1(ori_ori_n364_), .Y(ori_ori_n369_));
  NO3        o347(.A(ori_ori_n369_), .B(ori_ori_n363_), .C(ori_ori_n354_), .Y(ori_ori_n370_));
  OR2        o348(.A(ori_ori_n273_), .B(ori_ori_n104_), .Y(ori_ori_n371_));
  OR2        o349(.A(ori_ori_n371_), .B(ori_ori_n162_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n99_), .B(i_13_), .Y(ori_ori_n373_));
  NA2        o351(.A(ori_ori_n337_), .B(ori_ori_n308_), .Y(ori_ori_n374_));
  NO2        o352(.A(i_2_), .B(i_13_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n374_), .B(ori_ori_n373_), .Y(ori_ori_n376_));
  NO3        o354(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n377_));
  NO2        o355(.A(i_6_), .B(i_7_), .Y(ori_ori_n378_));
  NO2        o356(.A(i_11_), .B(i_1_), .Y(ori_ori_n379_));
  OR2        o357(.A(i_11_), .B(i_8_), .Y(ori_ori_n380_));
  NOi21      o358(.An(i_2_), .B(i_7_), .Y(ori_ori_n381_));
  NO2        o359(.A(i_3_), .B(ori_ori_n180_), .Y(ori_ori_n382_));
  NO2        o360(.A(i_6_), .B(i_10_), .Y(ori_ori_n383_));
  NA3        o361(.A(ori_ori_n222_), .B(ori_ori_n166_), .C(ori_ori_n136_), .Y(ori_ori_n384_));
  NA2        o362(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n157_), .B(i_3_), .Y(ori_ori_n386_));
  NAi31      o364(.An(ori_ori_n385_), .B(ori_ori_n386_), .C(ori_ori_n209_), .Y(ori_ori_n387_));
  NA3        o365(.A(ori_ori_n316_), .B(ori_ori_n171_), .C(ori_ori_n153_), .Y(ori_ori_n388_));
  NA3        o366(.A(ori_ori_n388_), .B(ori_ori_n387_), .C(ori_ori_n384_), .Y(ori_ori_n389_));
  NO2        o367(.A(ori_ori_n389_), .B(ori_ori_n376_), .Y(ori_ori_n390_));
  NA2        o368(.A(ori_ori_n356_), .B(ori_ori_n309_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n365_), .B(ori_ori_n315_), .Y(ori_ori_n392_));
  NAi21      o370(.An(ori_ori_n199_), .B(ori_ori_n320_), .Y(ori_ori_n393_));
  NA2        o371(.A(ori_ori_n268_), .B(ori_ori_n201_), .Y(ori_ori_n394_));
  NO2        o372(.A(ori_ori_n394_), .B(ori_ori_n393_), .Y(ori_ori_n395_));
  NA2        o373(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n396_));
  NA2        o374(.A(ori_ori_n260_), .B(ori_ori_n217_), .Y(ori_ori_n397_));
  OAI220     o375(.A0(ori_ori_n397_), .A1(ori_ori_n339_), .B0(ori_ori_n396_), .B1(ori_ori_n373_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n395_), .Y(ori_ori_n399_));
  NA4        o377(.A(ori_ori_n399_), .B(ori_ori_n390_), .C(ori_ori_n372_), .D(ori_ori_n370_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n126_), .B(ori_ori_n115_), .Y(ori_ori_n401_));
  AN2        o379(.A(ori_ori_n401_), .B(ori_ori_n356_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n402_), .B(ori_ori_n258_), .Y(ori_ori_n403_));
  NA4        o381(.A(ori_ori_n346_), .B(ori_ori_n345_), .C(ori_ori_n187_), .D(i_2_), .Y(ori_ori_n404_));
  INV        o382(.A(ori_ori_n404_), .Y(ori_ori_n405_));
  NA2        o383(.A(ori_ori_n309_), .B(ori_ori_n208_), .Y(ori_ori_n406_));
  NA2        o384(.A(ori_ori_n278_), .B(ori_ori_n73_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n296_), .B(ori_ori_n288_), .Y(ori_ori_n408_));
  OR2        o386(.A(ori_ori_n406_), .B(ori_ori_n408_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n410_));
  AOI210     o388(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n330_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n411_), .B(ori_ori_n409_), .Y(ori_ori_n412_));
  AOI210     o390(.A0(ori_ori_n405_), .A1(ori_ori_n188_), .B0(ori_ori_n412_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n230_), .B(ori_ori_n64_), .Y(ori_ori_n414_));
  OAI210     o392(.A0(i_8_), .A1(ori_ori_n414_), .B0(ori_ori_n138_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(ori_ori_n331_), .Y(ori_ori_n416_));
  NA3        o394(.A(ori_ori_n416_), .B(ori_ori_n413_), .C(ori_ori_n403_), .Y(ori_ori_n417_));
  NO2        o395(.A(i_12_), .B(ori_ori_n180_), .Y(ori_ori_n418_));
  NO2        o396(.A(i_8_), .B(i_7_), .Y(ori_ori_n419_));
  NA2        o397(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n420_));
  NO2        o398(.A(ori_ori_n420_), .B(i_6_), .Y(ori_ori_n421_));
  AOI220     o399(.A0(ori_ori_n337_), .A1(ori_ori_n263_), .B0(ori_ori_n224_), .B1(ori_ori_n221_), .Y(ori_ori_n422_));
  OAI220     o400(.A0(ori_ori_n422_), .A1(ori_ori_n237_), .B0(ori_ori_n373_), .B1(ori_ori_n137_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n423_), .B(ori_ori_n240_), .Y(ori_ori_n424_));
  NA3        o402(.A(ori_ori_n256_), .B(ori_ori_n168_), .C(ori_ori_n99_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n205_), .B(ori_ori_n44_), .Y(ori_ori_n426_));
  NO2        o404(.A(ori_ori_n157_), .B(i_5_), .Y(ori_ori_n427_));
  NA3        o405(.A(ori_ori_n427_), .B(ori_ori_n323_), .C(ori_ori_n261_), .Y(ori_ori_n428_));
  OAI210     o406(.A0(ori_ori_n428_), .A1(ori_ori_n426_), .B0(ori_ori_n425_), .Y(ori_ori_n429_));
  NA2        o407(.A(ori_ori_n429_), .B(ori_ori_n365_), .Y(ori_ori_n430_));
  NA2        o408(.A(ori_ori_n430_), .B(ori_ori_n424_), .Y(ori_ori_n431_));
  NA3        o409(.A(ori_ori_n201_), .B(ori_ori_n71_), .C(ori_ori_n44_), .Y(ori_ori_n432_));
  NA2        o410(.A(ori_ori_n253_), .B(ori_ori_n84_), .Y(ori_ori_n433_));
  NO2        o411(.A(ori_ori_n432_), .B(ori_ori_n433_), .Y(ori_ori_n434_));
  NA2        o412(.A(ori_ori_n207_), .B(ori_ori_n206_), .Y(ori_ori_n435_));
  NA2        o413(.A(ori_ori_n348_), .B(ori_ori_n205_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n435_), .B(ori_ori_n436_), .Y(ori_ori_n437_));
  AOI210     o415(.A0(ori_ori_n289_), .A1(ori_ori_n46_), .B0(ori_ori_n293_), .Y(ori_ori_n438_));
  NA2        o416(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n439_));
  NA3        o417(.A(ori_ori_n418_), .B(ori_ori_n249_), .C(ori_ori_n439_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n438_), .B(ori_ori_n440_), .Y(ori_ori_n441_));
  NO3        o419(.A(ori_ori_n441_), .B(ori_ori_n437_), .C(ori_ori_n434_), .Y(ori_ori_n442_));
  NO4        o420(.A(ori_ori_n226_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n443_));
  NO3        o421(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n444_));
  NO2        o422(.A(ori_ori_n329_), .B(i_1_), .Y(ori_ori_n445_));
  NOi31      o423(.An(ori_ori_n445_), .B(ori_ori_n357_), .C(ori_ori_n73_), .Y(ori_ori_n446_));
  NOi21      o424(.An(i_10_), .B(i_6_), .Y(ori_ori_n447_));
  NO2        o425(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n448_));
  AOI220     o426(.A0(ori_ori_n253_), .A1(ori_ori_n448_), .B0(ori_ori_n249_), .B1(ori_ori_n447_), .Y(ori_ori_n449_));
  NO2        o427(.A(ori_ori_n449_), .B(ori_ori_n355_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n118_), .B(ori_ori_n23_), .Y(ori_ori_n451_));
  NO2        o429(.A(ori_ori_n183_), .B(ori_ori_n37_), .Y(ori_ori_n452_));
  NOi31      o430(.An(ori_ori_n150_), .B(ori_ori_n452_), .C(ori_ori_n266_), .Y(ori_ori_n453_));
  NO2        o431(.A(ori_ori_n453_), .B(ori_ori_n450_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n407_), .B(ori_ori_n304_), .Y(ori_ori_n455_));
  INV        o433(.A(ori_ori_n261_), .Y(ori_ori_n456_));
  NO2        o434(.A(i_12_), .B(ori_ori_n86_), .Y(ori_ori_n457_));
  NA3        o435(.A(ori_ori_n457_), .B(ori_ori_n249_), .C(ori_ori_n439_), .Y(ori_ori_n458_));
  NA3        o436(.A(ori_ori_n312_), .B(ori_ori_n253_), .C(ori_ori_n201_), .Y(ori_ori_n459_));
  AOI210     o437(.A0(ori_ori_n459_), .A1(ori_ori_n458_), .B0(ori_ori_n456_), .Y(ori_ori_n460_));
  OR2        o438(.A(i_2_), .B(i_5_), .Y(ori_ori_n461_));
  OR2        o439(.A(ori_ori_n461_), .B(ori_ori_n326_), .Y(ori_ori_n462_));
  AOI210     o440(.A0(ori_ori_n298_), .A1(ori_ori_n221_), .B0(ori_ori_n183_), .Y(ori_ori_n463_));
  AOI210     o441(.A0(ori_ori_n463_), .A1(ori_ori_n462_), .B0(ori_ori_n393_), .Y(ori_ori_n464_));
  NO3        o442(.A(ori_ori_n464_), .B(ori_ori_n460_), .C(ori_ori_n455_), .Y(ori_ori_n465_));
  NA3        o443(.A(ori_ori_n465_), .B(ori_ori_n454_), .C(ori_ori_n442_), .Y(ori_ori_n466_));
  NO4        o444(.A(ori_ori_n466_), .B(ori_ori_n431_), .C(ori_ori_n417_), .D(ori_ori_n400_), .Y(ori_ori_n467_));
  NA4        o445(.A(ori_ori_n467_), .B(ori_ori_n344_), .C(ori_ori_n277_), .D(ori_ori_n259_), .Y(ori7));
  NO2        o446(.A(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n469_));
  NO2        o447(.A(ori_ori_n111_), .B(ori_ori_n92_), .Y(ori_ori_n470_));
  NA2        o448(.A(ori_ori_n310_), .B(ori_ori_n470_), .Y(ori_ori_n471_));
  NA2        o449(.A(ori_ori_n383_), .B(ori_ori_n84_), .Y(ori_ori_n472_));
  NA2        o450(.A(i_11_), .B(ori_ori_n180_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n148_), .B(ori_ori_n473_), .Y(ori_ori_n474_));
  OAI210     o452(.A0(ori_ori_n474_), .A1(ori_ori_n472_), .B0(ori_ori_n471_), .Y(ori_ori_n475_));
  NA3        o453(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n476_));
  NO2        o454(.A(ori_ori_n215_), .B(i_4_), .Y(ori_ori_n477_));
  NA2        o455(.A(ori_ori_n477_), .B(i_8_), .Y(ori_ori_n478_));
  NO2        o456(.A(ori_ori_n108_), .B(ori_ori_n476_), .Y(ori_ori_n479_));
  NA2        o457(.A(i_2_), .B(ori_ori_n86_), .Y(ori_ori_n480_));
  OAI210     o458(.A0(ori_ori_n89_), .A1(ori_ori_n187_), .B0(ori_ori_n188_), .Y(ori_ori_n481_));
  NO2        o459(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n482_));
  NA2        o460(.A(i_4_), .B(i_8_), .Y(ori_ori_n483_));
  AOI210     o461(.A0(ori_ori_n483_), .A1(ori_ori_n256_), .B0(ori_ori_n482_), .Y(ori_ori_n484_));
  OAI220     o462(.A0(ori_ori_n484_), .A1(ori_ori_n480_), .B0(ori_ori_n481_), .B1(i_13_), .Y(ori_ori_n485_));
  NO4        o463(.A(ori_ori_n485_), .B(ori_ori_n479_), .C(ori_ori_n475_), .D(ori_ori_n469_), .Y(ori_ori_n486_));
  AOI210     o464(.A0(ori_ori_n132_), .A1(ori_ori_n62_), .B0(i_10_), .Y(ori_ori_n487_));
  AOI210     o465(.A0(ori_ori_n487_), .A1(ori_ori_n215_), .B0(ori_ori_n161_), .Y(ori_ori_n488_));
  OR2        o466(.A(i_6_), .B(i_10_), .Y(ori_ori_n489_));
  NO2        o467(.A(ori_ori_n489_), .B(ori_ori_n23_), .Y(ori_ori_n490_));
  OR3        o468(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n491_));
  NO3        o469(.A(ori_ori_n491_), .B(i_8_), .C(ori_ori_n31_), .Y(ori_ori_n492_));
  INV        o470(.A(ori_ori_n184_), .Y(ori_ori_n493_));
  NO2        o471(.A(ori_ori_n492_), .B(ori_ori_n490_), .Y(ori_ori_n494_));
  OA220      o472(.A0(ori_ori_n494_), .A1(ori_ori_n456_), .B0(ori_ori_n488_), .B1(ori_ori_n242_), .Y(ori_ori_n495_));
  AOI210     o473(.A0(ori_ori_n495_), .A1(ori_ori_n486_), .B0(ori_ori_n63_), .Y(ori_ori_n496_));
  NOi21      o474(.An(i_11_), .B(i_7_), .Y(ori_ori_n497_));
  AO210      o475(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n498_));
  NO2        o476(.A(ori_ori_n498_), .B(ori_ori_n497_), .Y(ori_ori_n499_));
  NA2        o477(.A(ori_ori_n499_), .B(ori_ori_n192_), .Y(ori_ori_n500_));
  NA3        o478(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n501_));
  NAi31      o479(.An(ori_ori_n501_), .B(ori_ori_n198_), .C(i_11_), .Y(ori_ori_n502_));
  AOI210     o480(.A0(ori_ori_n502_), .A1(ori_ori_n500_), .B0(ori_ori_n63_), .Y(ori_ori_n503_));
  NA2        o481(.A(ori_ori_n88_), .B(ori_ori_n63_), .Y(ori_ori_n504_));
  AO210      o482(.A0(ori_ori_n504_), .A1(ori_ori_n304_), .B0(ori_ori_n41_), .Y(ori_ori_n505_));
  NO3        o483(.A(ori_ori_n232_), .B(ori_ori_n193_), .C(ori_ori_n473_), .Y(ori_ori_n506_));
  OAI210     o484(.A0(ori_ori_n506_), .A1(ori_ori_n209_), .B0(ori_ori_n63_), .Y(ori_ori_n507_));
  NA2        o485(.A(ori_ori_n327_), .B(ori_ori_n31_), .Y(ori_ori_n508_));
  OR2        o486(.A(ori_ori_n193_), .B(ori_ori_n111_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n509_), .B(ori_ori_n508_), .Y(ori_ori_n510_));
  NO2        o488(.A(i_1_), .B(i_4_), .Y(ori_ori_n511_));
  NA2        o489(.A(ori_ori_n511_), .B(ori_ori_n510_), .Y(ori_ori_n512_));
  NO2        o490(.A(i_1_), .B(i_12_), .Y(ori_ori_n513_));
  NA3        o491(.A(ori_ori_n513_), .B(ori_ori_n113_), .C(ori_ori_n24_), .Y(ori_ori_n514_));
  BUFFER     o492(.A(ori_ori_n514_), .Y(ori_ori_n515_));
  NA4        o493(.A(ori_ori_n515_), .B(ori_ori_n512_), .C(ori_ori_n507_), .D(ori_ori_n505_), .Y(ori_ori_n516_));
  OAI210     o494(.A0(ori_ori_n516_), .A1(ori_ori_n503_), .B0(i_6_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n501_), .B(ori_ori_n111_), .Y(ori_ori_n518_));
  NA2        o496(.A(ori_ori_n518_), .B(ori_ori_n457_), .Y(ori_ori_n519_));
  NO2        o497(.A(ori_ori_n215_), .B(ori_ori_n86_), .Y(ori_ori_n520_));
  NO2        o498(.A(ori_ori_n520_), .B(i_11_), .Y(ori_ori_n521_));
  NA2        o499(.A(ori_ori_n519_), .B(ori_ori_n358_), .Y(ori_ori_n522_));
  NO3        o500(.A(ori_ori_n489_), .B(ori_ori_n214_), .C(ori_ori_n23_), .Y(ori_ori_n523_));
  AOI210     o501(.A0(i_1_), .A1(ori_ori_n233_), .B0(ori_ori_n523_), .Y(ori_ori_n524_));
  NO2        o502(.A(ori_ori_n524_), .B(ori_ori_n44_), .Y(ori_ori_n525_));
  NA3        o503(.A(ori_ori_n419_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n526_));
  INV        o504(.A(i_2_), .Y(ori_ori_n527_));
  NA2        o505(.A(ori_ori_n142_), .B(i_9_), .Y(ori_ori_n528_));
  NA3        o506(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n529_));
  NO2        o507(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n530_));
  NA3        o508(.A(ori_ori_n530_), .B(ori_ori_n241_), .C(ori_ori_n44_), .Y(ori_ori_n531_));
  OAI220     o509(.A0(ori_ori_n531_), .A1(ori_ori_n529_), .B0(ori_ori_n528_), .B1(ori_ori_n527_), .Y(ori_ori_n532_));
  AOI210     o510(.A0(ori_ori_n379_), .A1(ori_ori_n332_), .B0(ori_ori_n219_), .Y(ori_ori_n533_));
  NO2        o511(.A(ori_ori_n533_), .B(ori_ori_n480_), .Y(ori_ori_n534_));
  NAi21      o512(.An(ori_ori_n526_), .B(ori_ori_n94_), .Y(ori_ori_n535_));
  NA2        o513(.A(ori_ori_n530_), .B(ori_ori_n241_), .Y(ori_ori_n536_));
  NO2        o514(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n537_));
  NA2        o515(.A(ori_ori_n537_), .B(ori_ori_n24_), .Y(ori_ori_n538_));
  OAI210     o516(.A0(ori_ori_n538_), .A1(ori_ori_n536_), .B0(ori_ori_n535_), .Y(ori_ori_n539_));
  OR3        o517(.A(ori_ori_n539_), .B(ori_ori_n534_), .C(ori_ori_n532_), .Y(ori_ori_n540_));
  NO3        o518(.A(ori_ori_n540_), .B(ori_ori_n525_), .C(ori_ori_n522_), .Y(ori_ori_n541_));
  NO2        o519(.A(ori_ori_n215_), .B(ori_ori_n104_), .Y(ori_ori_n542_));
  NO2        o520(.A(ori_ori_n542_), .B(ori_ori_n497_), .Y(ori_ori_n543_));
  NA2        o521(.A(ori_ori_n543_), .B(i_1_), .Y(ori_ori_n544_));
  NO2        o522(.A(ori_ori_n544_), .B(ori_ori_n491_), .Y(ori_ori_n545_));
  NO2        o523(.A(ori_ori_n328_), .B(ori_ori_n86_), .Y(ori_ori_n546_));
  NA2        o524(.A(ori_ori_n545_), .B(ori_ori_n46_), .Y(ori_ori_n547_));
  NA2        o525(.A(i_3_), .B(ori_ori_n180_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n548_), .B(ori_ori_n118_), .Y(ori_ori_n549_));
  AN2        o527(.A(ori_ori_n549_), .B(ori_ori_n421_), .Y(ori_ori_n550_));
  NO2        o528(.A(ori_ori_n214_), .B(ori_ori_n44_), .Y(ori_ori_n551_));
  NO3        o529(.A(ori_ori_n551_), .B(ori_ori_n258_), .C(ori_ori_n216_), .Y(ori_ori_n552_));
  NO2        o530(.A(ori_ori_n121_), .B(ori_ori_n37_), .Y(ori_ori_n553_));
  NO2        o531(.A(ori_ori_n553_), .B(i_6_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n86_), .B(i_9_), .Y(ori_ori_n555_));
  NO2        o533(.A(ori_ori_n555_), .B(ori_ori_n63_), .Y(ori_ori_n556_));
  NO2        o534(.A(ori_ori_n556_), .B(ori_ori_n513_), .Y(ori_ori_n557_));
  NO4        o535(.A(ori_ori_n557_), .B(ori_ori_n554_), .C(ori_ori_n552_), .D(i_4_), .Y(ori_ori_n558_));
  NA2        o536(.A(i_1_), .B(i_3_), .Y(ori_ori_n559_));
  NO2        o537(.A(ori_ori_n359_), .B(ori_ori_n95_), .Y(ori_ori_n560_));
  AOI210     o538(.A0(ori_ori_n551_), .A1(ori_ori_n447_), .B0(ori_ori_n560_), .Y(ori_ori_n561_));
  NO2        o539(.A(ori_ori_n561_), .B(ori_ori_n559_), .Y(ori_ori_n562_));
  NO3        o540(.A(ori_ori_n562_), .B(ori_ori_n558_), .C(ori_ori_n550_), .Y(ori_ori_n563_));
  NA4        o541(.A(ori_ori_n563_), .B(ori_ori_n547_), .C(ori_ori_n541_), .D(ori_ori_n517_), .Y(ori_ori_n564_));
  AN2        o542(.A(ori_ori_n222_), .B(ori_ori_n86_), .Y(ori_ori_n565_));
  NA2        o543(.A(ori_ori_n296_), .B(ori_ori_n295_), .Y(ori_ori_n566_));
  NA3        o544(.A(ori_ori_n383_), .B(ori_ori_n410_), .C(ori_ori_n46_), .Y(ori_ori_n567_));
  NO3        o545(.A(ori_ori_n381_), .B(ori_ori_n483_), .C(ori_ori_n86_), .Y(ori_ori_n568_));
  NA2        o546(.A(ori_ori_n568_), .B(ori_ori_n25_), .Y(ori_ori_n569_));
  NA3        o547(.A(ori_ori_n161_), .B(ori_ori_n84_), .C(ori_ori_n86_), .Y(ori_ori_n570_));
  NA4        o548(.A(ori_ori_n570_), .B(ori_ori_n569_), .C(ori_ori_n567_), .D(ori_ori_n566_), .Y(ori_ori_n571_));
  OAI210     o549(.A0(ori_ori_n571_), .A1(ori_ori_n565_), .B0(i_1_), .Y(ori_ori_n572_));
  AOI210     o550(.A0(ori_ori_n241_), .A1(ori_ori_n100_), .B0(i_1_), .Y(ori_ori_n573_));
  NO2        o551(.A(ori_ori_n294_), .B(i_2_), .Y(ori_ori_n574_));
  NA2        o552(.A(ori_ori_n574_), .B(ori_ori_n573_), .Y(ori_ori_n575_));
  AOI210     o553(.A0(ori_ori_n575_), .A1(ori_ori_n572_), .B0(i_13_), .Y(ori_ori_n576_));
  OR2        o554(.A(i_11_), .B(i_7_), .Y(ori_ori_n577_));
  NA3        o555(.A(ori_ori_n577_), .B(ori_ori_n109_), .C(ori_ori_n142_), .Y(ori_ori_n578_));
  AOI220     o556(.A0(ori_ori_n375_), .A1(ori_ori_n161_), .B0(ori_ori_n352_), .B1(ori_ori_n142_), .Y(ori_ori_n579_));
  OAI210     o557(.A0(ori_ori_n579_), .A1(ori_ori_n44_), .B0(ori_ori_n578_), .Y(ori_ori_n580_));
  AOI210     o558(.A0(ori_ori_n529_), .A1(ori_ori_n54_), .B0(i_12_), .Y(ori_ori_n581_));
  NO2        o559(.A(ori_ori_n381_), .B(ori_ori_n24_), .Y(ori_ori_n582_));
  AOI220     o560(.A0(ori_ori_n582_), .A1(ori_ori_n546_), .B0(ori_ori_n222_), .B1(ori_ori_n135_), .Y(ori_ori_n583_));
  OAI220     o561(.A0(ori_ori_n583_), .A1(ori_ori_n41_), .B0(ori_ori_n893_), .B1(ori_ori_n95_), .Y(ori_ori_n584_));
  AOI210     o562(.A0(ori_ori_n580_), .A1(ori_ori_n267_), .B0(ori_ori_n584_), .Y(ori_ori_n585_));
  INV        o563(.A(ori_ori_n118_), .Y(ori_ori_n586_));
  AOI220     o564(.A0(ori_ori_n586_), .A1(ori_ori_n72_), .B0(ori_ori_n312_), .B1(ori_ori_n530_), .Y(ori_ori_n587_));
  NO2        o565(.A(ori_ori_n587_), .B(ori_ori_n220_), .Y(ori_ori_n588_));
  AOI210     o566(.A0(ori_ori_n349_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n589_));
  NOi31      o567(.An(ori_ori_n589_), .B(ori_ori_n472_), .C(ori_ori_n44_), .Y(ori_ori_n590_));
  NA2        o568(.A(ori_ori_n131_), .B(i_13_), .Y(ori_ori_n591_));
  NO2        o569(.A(ori_ori_n529_), .B(ori_ori_n118_), .Y(ori_ori_n592_));
  INV        o570(.A(ori_ori_n592_), .Y(ori_ori_n593_));
  OAI220     o571(.A0(ori_ori_n593_), .A1(ori_ori_n71_), .B0(ori_ori_n591_), .B1(ori_ori_n573_), .Y(ori_ori_n594_));
  NO3        o572(.A(ori_ori_n71_), .B(ori_ori_n32_), .C(ori_ori_n104_), .Y(ori_ori_n595_));
  NA2        o573(.A(ori_ori_n26_), .B(ori_ori_n180_), .Y(ori_ori_n596_));
  NA2        o574(.A(ori_ori_n596_), .B(i_7_), .Y(ori_ori_n597_));
  NO3        o575(.A(ori_ori_n381_), .B(ori_ori_n215_), .C(ori_ori_n86_), .Y(ori_ori_n598_));
  AOI210     o576(.A0(ori_ori_n598_), .A1(ori_ori_n597_), .B0(ori_ori_n595_), .Y(ori_ori_n599_));
  AOI220     o577(.A0(ori_ori_n312_), .A1(ori_ori_n530_), .B0(ori_ori_n94_), .B1(ori_ori_n105_), .Y(ori_ori_n600_));
  OAI220     o578(.A0(ori_ori_n600_), .A1(ori_ori_n478_), .B0(ori_ori_n599_), .B1(ori_ori_n493_), .Y(ori_ori_n601_));
  NO4        o579(.A(ori_ori_n601_), .B(ori_ori_n594_), .C(ori_ori_n590_), .D(ori_ori_n588_), .Y(ori_ori_n602_));
  OR2        o580(.A(i_11_), .B(i_6_), .Y(ori_ori_n603_));
  NA3        o581(.A(ori_ori_n477_), .B(ori_ori_n596_), .C(i_7_), .Y(ori_ori_n604_));
  AOI210     o582(.A0(ori_ori_n604_), .A1(ori_ori_n593_), .B0(ori_ori_n603_), .Y(ori_ori_n605_));
  NA3        o583(.A(ori_ori_n327_), .B(ori_ori_n482_), .C(ori_ori_n100_), .Y(ori_ori_n606_));
  NA2        o584(.A(ori_ori_n521_), .B(i_13_), .Y(ori_ori_n607_));
  NA2        o585(.A(ori_ori_n105_), .B(ori_ori_n596_), .Y(ori_ori_n608_));
  NAi21      o586(.An(i_11_), .B(i_12_), .Y(ori_ori_n609_));
  NOi41      o587(.An(ori_ori_n114_), .B(ori_ori_n609_), .C(i_13_), .D(ori_ori_n86_), .Y(ori_ori_n610_));
  NO3        o588(.A(ori_ori_n381_), .B(ori_ori_n457_), .C(ori_ori_n483_), .Y(ori_ori_n611_));
  AOI220     o589(.A0(ori_ori_n611_), .A1(ori_ori_n260_), .B0(ori_ori_n610_), .B1(ori_ori_n608_), .Y(ori_ori_n612_));
  NA3        o590(.A(ori_ori_n612_), .B(ori_ori_n607_), .C(ori_ori_n606_), .Y(ori_ori_n613_));
  OAI210     o591(.A0(ori_ori_n613_), .A1(ori_ori_n605_), .B0(ori_ori_n63_), .Y(ori_ori_n614_));
  NO2        o592(.A(i_2_), .B(i_12_), .Y(ori_ori_n615_));
  NA2        o593(.A(ori_ori_n293_), .B(ori_ori_n615_), .Y(ori_ori_n616_));
  NA2        o594(.A(i_8_), .B(ori_ori_n25_), .Y(ori_ori_n617_));
  NO3        o595(.A(ori_ori_n617_), .B(ori_ori_n310_), .C(ori_ori_n477_), .Y(ori_ori_n618_));
  OAI210     o596(.A0(ori_ori_n618_), .A1(ori_ori_n295_), .B0(ori_ori_n293_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n132_), .B(i_2_), .Y(ori_ori_n620_));
  NA2        o598(.A(ori_ori_n620_), .B(ori_ori_n513_), .Y(ori_ori_n621_));
  NA3        o599(.A(ori_ori_n621_), .B(ori_ori_n619_), .C(ori_ori_n616_), .Y(ori_ori_n622_));
  NA3        o600(.A(ori_ori_n622_), .B(ori_ori_n45_), .C(ori_ori_n208_), .Y(ori_ori_n623_));
  NA4        o601(.A(ori_ori_n623_), .B(ori_ori_n614_), .C(ori_ori_n602_), .D(ori_ori_n585_), .Y(ori_ori_n624_));
  OR4        o602(.A(ori_ori_n624_), .B(ori_ori_n576_), .C(ori_ori_n564_), .D(ori_ori_n496_), .Y(ori5));
  NA2        o603(.A(ori_ori_n543_), .B(ori_ori_n244_), .Y(ori_ori_n626_));
  AN2        o604(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n627_));
  NA3        o605(.A(ori_ori_n627_), .B(ori_ori_n615_), .C(ori_ori_n111_), .Y(ori_ori_n628_));
  NO2        o606(.A(ori_ori_n478_), .B(i_11_), .Y(ori_ori_n629_));
  NA2        o607(.A(ori_ori_n89_), .B(ori_ori_n629_), .Y(ori_ori_n630_));
  NA3        o608(.A(ori_ori_n630_), .B(ori_ori_n628_), .C(ori_ori_n626_), .Y(ori_ori_n631_));
  NO3        o609(.A(i_11_), .B(ori_ori_n215_), .C(i_13_), .Y(ori_ori_n632_));
  NO2        o610(.A(ori_ori_n128_), .B(ori_ori_n23_), .Y(ori_ori_n633_));
  NA2        o611(.A(i_12_), .B(i_8_), .Y(ori_ori_n634_));
  OAI210     o612(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n634_), .Y(ori_ori_n635_));
  INV        o613(.A(ori_ori_n348_), .Y(ori_ori_n636_));
  AOI220     o614(.A0(ori_ori_n261_), .A1(ori_ori_n451_), .B0(ori_ori_n635_), .B1(ori_ori_n633_), .Y(ori_ori_n637_));
  INV        o615(.A(ori_ori_n637_), .Y(ori_ori_n638_));
  NO2        o616(.A(ori_ori_n638_), .B(ori_ori_n631_), .Y(ori_ori_n639_));
  INV        o617(.A(ori_ori_n166_), .Y(ori_ori_n640_));
  INV        o618(.A(ori_ori_n222_), .Y(ori_ori_n641_));
  OAI210     o619(.A0(ori_ori_n574_), .A1(ori_ori_n350_), .B0(ori_ori_n114_), .Y(ori_ori_n642_));
  AOI210     o620(.A0(ori_ori_n642_), .A1(ori_ori_n641_), .B0(ori_ori_n640_), .Y(ori_ori_n643_));
  NO2        o621(.A(ori_ori_n359_), .B(ori_ori_n26_), .Y(ori_ori_n644_));
  NO2        o622(.A(ori_ori_n644_), .B(ori_ori_n332_), .Y(ori_ori_n645_));
  NA2        o623(.A(ori_ori_n645_), .B(i_2_), .Y(ori_ori_n646_));
  INV        o624(.A(ori_ori_n646_), .Y(ori_ori_n647_));
  AOI210     o625(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n329_), .Y(ori_ori_n648_));
  AOI210     o626(.A0(ori_ori_n648_), .A1(ori_ori_n647_), .B0(ori_ori_n643_), .Y(ori_ori_n649_));
  NO2        o627(.A(ori_ori_n179_), .B(ori_ori_n129_), .Y(ori_ori_n650_));
  OAI210     o628(.A0(ori_ori_n650_), .A1(ori_ori_n633_), .B0(i_2_), .Y(ori_ori_n651_));
  INV        o629(.A(ori_ori_n167_), .Y(ori_ori_n652_));
  NO3        o630(.A(ori_ori_n498_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n653_));
  AOI210     o631(.A0(ori_ori_n652_), .A1(ori_ori_n89_), .B0(ori_ori_n653_), .Y(ori_ori_n654_));
  AOI210     o632(.A0(ori_ori_n654_), .A1(ori_ori_n651_), .B0(ori_ori_n180_), .Y(ori_ori_n655_));
  OA210      o633(.A0(ori_ori_n499_), .A1(ori_ori_n130_), .B0(i_13_), .Y(ori_ori_n656_));
  NA2        o634(.A(ori_ori_n184_), .B(ori_ori_n187_), .Y(ori_ori_n657_));
  NA2        o635(.A(ori_ori_n155_), .B(ori_ori_n473_), .Y(ori_ori_n658_));
  AOI210     o636(.A0(ori_ori_n658_), .A1(ori_ori_n657_), .B0(ori_ori_n298_), .Y(ori_ori_n659_));
  AOI210     o637(.A0(ori_ori_n193_), .A1(ori_ori_n152_), .B0(ori_ori_n410_), .Y(ori_ori_n660_));
  NA2        o638(.A(ori_ori_n660_), .B(ori_ori_n332_), .Y(ori_ori_n661_));
  NO2        o639(.A(ori_ori_n105_), .B(ori_ori_n44_), .Y(ori_ori_n662_));
  INV        o640(.A(ori_ori_n255_), .Y(ori_ori_n663_));
  NA4        o641(.A(ori_ori_n663_), .B(ori_ori_n256_), .C(ori_ori_n128_), .D(ori_ori_n42_), .Y(ori_ori_n664_));
  OAI210     o642(.A0(ori_ori_n664_), .A1(ori_ori_n662_), .B0(ori_ori_n661_), .Y(ori_ori_n665_));
  NO4        o643(.A(ori_ori_n665_), .B(ori_ori_n659_), .C(ori_ori_n656_), .D(ori_ori_n655_), .Y(ori_ori_n666_));
  NA2        o644(.A(ori_ori_n451_), .B(ori_ori_n28_), .Y(ori_ori_n667_));
  NA2        o645(.A(ori_ori_n632_), .B(ori_ori_n250_), .Y(ori_ori_n668_));
  NA2        o646(.A(ori_ori_n668_), .B(ori_ori_n667_), .Y(ori_ori_n669_));
  NO2        o647(.A(ori_ori_n62_), .B(i_12_), .Y(ori_ori_n670_));
  NO2        o648(.A(ori_ori_n670_), .B(ori_ori_n130_), .Y(ori_ori_n671_));
  NO2        o649(.A(ori_ori_n671_), .B(ori_ori_n473_), .Y(ori_ori_n672_));
  AOI220     o650(.A0(ori_ori_n672_), .A1(ori_ori_n36_), .B0(ori_ori_n669_), .B1(ori_ori_n46_), .Y(ori_ori_n673_));
  NA4        o651(.A(ori_ori_n673_), .B(ori_ori_n666_), .C(ori_ori_n649_), .D(ori_ori_n639_), .Y(ori6));
  NA4        o652(.A(ori_ori_n315_), .B(ori_ori_n382_), .C(ori_ori_n71_), .D(ori_ori_n104_), .Y(ori_ori_n675_));
  INV        o653(.A(ori_ori_n675_), .Y(ori_ori_n676_));
  NO2        o654(.A(ori_ori_n204_), .B(ori_ori_n385_), .Y(ori_ori_n677_));
  NO2        o655(.A(i_11_), .B(i_9_), .Y(ori_ori_n678_));
  NO2        o656(.A(ori_ori_n676_), .B(ori_ori_n265_), .Y(ori_ori_n679_));
  OR2        o657(.A(ori_ori_n679_), .B(i_12_), .Y(ori_ori_n680_));
  NA2        o658(.A(ori_ori_n299_), .B(ori_ori_n268_), .Y(ori_ori_n681_));
  NA2        o659(.A(ori_ori_n457_), .B(ori_ori_n63_), .Y(ori_ori_n682_));
  BUFFER     o660(.A(ori_ori_n504_), .Y(ori_ori_n683_));
  NA3        o661(.A(ori_ori_n683_), .B(ori_ori_n682_), .C(ori_ori_n681_), .Y(ori_ori_n684_));
  INV        o662(.A(ori_ori_n182_), .Y(ori_ori_n685_));
  AOI220     o663(.A0(ori_ori_n685_), .A1(ori_ori_n678_), .B0(ori_ori_n684_), .B1(ori_ori_n73_), .Y(ori_ori_n686_));
  INV        o664(.A(ori_ori_n264_), .Y(ori_ori_n687_));
  NA2        o665(.A(ori_ori_n75_), .B(ori_ori_n135_), .Y(ori_ori_n688_));
  INV        o666(.A(ori_ori_n128_), .Y(ori_ori_n689_));
  NA2        o667(.A(ori_ori_n689_), .B(ori_ori_n46_), .Y(ori_ori_n690_));
  AOI210     o668(.A0(ori_ori_n690_), .A1(ori_ori_n688_), .B0(ori_ori_n687_), .Y(ori_ori_n691_));
  NO3        o669(.A(ori_ori_n226_), .B(ori_ori_n136_), .C(i_9_), .Y(ori_ori_n692_));
  NA2        o670(.A(ori_ori_n692_), .B(ori_ori_n670_), .Y(ori_ori_n693_));
  AOI210     o671(.A0(ori_ori_n693_), .A1(ori_ori_n408_), .B0(ori_ori_n174_), .Y(ori_ori_n694_));
  NO2        o672(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n695_));
  NAi32      o673(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n696_));
  NO2        o674(.A(ori_ori_n603_), .B(ori_ori_n696_), .Y(ori_ori_n697_));
  OR3        o675(.A(ori_ori_n697_), .B(ori_ori_n694_), .C(ori_ori_n691_), .Y(ori_ori_n698_));
  NO2        o676(.A(ori_ori_n577_), .B(i_2_), .Y(ori_ori_n699_));
  NA2        o677(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n700_));
  NO2        o678(.A(ori_ori_n700_), .B(ori_ori_n326_), .Y(ori_ori_n701_));
  NA2        o679(.A(ori_ori_n701_), .B(ori_ori_n699_), .Y(ori_ori_n702_));
  OR2        o680(.A(ori_ori_n499_), .B(ori_ori_n350_), .Y(ori_ori_n703_));
  NA3        o681(.A(ori_ori_n703_), .B(ori_ori_n151_), .C(ori_ori_n69_), .Y(ori_ori_n704_));
  AO210      o682(.A0(ori_ori_n392_), .A1(ori_ori_n636_), .B0(ori_ori_n36_), .Y(ori_ori_n705_));
  NA3        o683(.A(ori_ori_n705_), .B(ori_ori_n704_), .C(ori_ori_n702_), .Y(ori_ori_n706_));
  OAI210     o684(.A0(ori_ori_n520_), .A1(i_11_), .B0(ori_ori_n87_), .Y(ori_ori_n707_));
  AOI220     o685(.A0(ori_ori_n707_), .A1(ori_ori_n444_), .B0(ori_ori_n677_), .B1(ori_ori_n597_), .Y(ori_ori_n708_));
  NA3        o686(.A(ori_ori_n298_), .B(ori_ori_n217_), .C(ori_ori_n151_), .Y(ori_ori_n709_));
  NA2        o687(.A(ori_ori_n319_), .B(ori_ori_n70_), .Y(ori_ori_n710_));
  NA4        o688(.A(ori_ori_n710_), .B(ori_ori_n709_), .C(ori_ori_n708_), .D(ori_ori_n481_), .Y(ori_ori_n711_));
  AO210      o689(.A0(ori_ori_n410_), .A1(ori_ori_n46_), .B0(ori_ori_n88_), .Y(ori_ori_n712_));
  NA3        o690(.A(ori_ori_n712_), .B(ori_ori_n383_), .C(ori_ori_n201_), .Y(ori_ori_n713_));
  AOI210     o691(.A0(ori_ori_n350_), .A1(ori_ori_n348_), .B0(ori_ori_n443_), .Y(ori_ori_n714_));
  NO2        o692(.A(ori_ori_n489_), .B(ori_ori_n105_), .Y(ori_ori_n715_));
  OAI210     o693(.A0(ori_ori_n715_), .A1(ori_ori_n115_), .B0(ori_ori_n325_), .Y(ori_ori_n716_));
  NA2        o694(.A(ori_ori_n221_), .B(ori_ori_n46_), .Y(ori_ori_n717_));
  INV        o695(.A(ori_ori_n462_), .Y(ori_ori_n718_));
  NA3        o696(.A(ori_ori_n718_), .B(ori_ori_n264_), .C(i_7_), .Y(ori_ori_n719_));
  NA4        o697(.A(ori_ori_n719_), .B(ori_ori_n716_), .C(ori_ori_n714_), .D(ori_ori_n713_), .Y(ori_ori_n720_));
  NO4        o698(.A(ori_ori_n720_), .B(ori_ori_n711_), .C(ori_ori_n706_), .D(ori_ori_n698_), .Y(ori_ori_n721_));
  NA4        o699(.A(ori_ori_n721_), .B(ori_ori_n686_), .C(ori_ori_n680_), .D(ori_ori_n306_), .Y(ori3));
  NA2        o700(.A(i_12_), .B(i_10_), .Y(ori_ori_n723_));
  NO2        o701(.A(i_11_), .B(ori_ori_n215_), .Y(ori_ori_n724_));
  NA3        o702(.A(ori_ori_n709_), .B(ori_ori_n481_), .C(ori_ori_n297_), .Y(ori_ori_n725_));
  NA2        o703(.A(ori_ori_n725_), .B(ori_ori_n40_), .Y(ori_ori_n726_));
  NOi21      o704(.An(ori_ori_n99_), .B(ori_ori_n645_), .Y(ori_ori_n727_));
  NO3        o705(.A(ori_ori_n509_), .B(ori_ori_n359_), .C(ori_ori_n135_), .Y(ori_ori_n728_));
  NA2        o706(.A(ori_ori_n327_), .B(ori_ori_n45_), .Y(ori_ori_n729_));
  AN2        o707(.A(ori_ori_n357_), .B(ori_ori_n55_), .Y(ori_ori_n730_));
  NO3        o708(.A(ori_ori_n730_), .B(ori_ori_n728_), .C(ori_ori_n727_), .Y(ori_ori_n731_));
  AOI210     o709(.A0(ori_ori_n731_), .A1(ori_ori_n726_), .B0(ori_ori_n48_), .Y(ori_ori_n732_));
  NO4        o710(.A(ori_ori_n302_), .B(ori_ori_n309_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n174_), .B(ori_ori_n447_), .Y(ori_ori_n734_));
  NOi21      o712(.An(ori_ori_n734_), .B(ori_ori_n733_), .Y(ori_ori_n735_));
  NO2        o713(.A(ori_ori_n735_), .B(ori_ori_n63_), .Y(ori_ori_n736_));
  NOi21      o714(.An(i_5_), .B(i_9_), .Y(ori_ori_n737_));
  NA2        o715(.A(ori_ori_n737_), .B(ori_ori_n346_), .Y(ori_ori_n738_));
  BUFFER     o716(.A(ori_ori_n241_), .Y(ori_ori_n739_));
  AOI210     o717(.A0(ori_ori_n739_), .A1(ori_ori_n379_), .B0(ori_ori_n568_), .Y(ori_ori_n740_));
  NO2        o718(.A(ori_ori_n740_), .B(ori_ori_n738_), .Y(ori_ori_n741_));
  NO3        o719(.A(ori_ori_n741_), .B(ori_ori_n736_), .C(ori_ori_n732_), .Y(ori_ori_n742_));
  NA2        o720(.A(ori_ori_n174_), .B(ori_ori_n24_), .Y(ori_ori_n743_));
  NO2        o721(.A(ori_ori_n553_), .B(ori_ori_n470_), .Y(ori_ori_n744_));
  NO2        o722(.A(ori_ori_n744_), .B(ori_ori_n743_), .Y(ori_ori_n745_));
  NAi21      o723(.An(ori_ori_n162_), .B(ori_ori_n341_), .Y(ori_ori_n746_));
  NO2        o724(.A(ori_ori_n746_), .B(ori_ori_n717_), .Y(ori_ori_n747_));
  NO2        o725(.A(ori_ori_n747_), .B(ori_ori_n745_), .Y(ori_ori_n748_));
  NA2        o726(.A(ori_ori_n448_), .B(i_0_), .Y(ori_ori_n749_));
  NO3        o727(.A(ori_ori_n749_), .B(ori_ori_n311_), .C(ori_ori_n89_), .Y(ori_ori_n750_));
  NO4        o728(.A(ori_ori_n461_), .B(ori_ori_n198_), .C(ori_ori_n329_), .D(ori_ori_n326_), .Y(ori_ori_n751_));
  AOI210     o729(.A0(ori_ori_n751_), .A1(i_11_), .B0(ori_ori_n750_), .Y(ori_ori_n752_));
  INV        o730(.A(ori_ori_n378_), .Y(ori_ori_n753_));
  NA2        o731(.A(ori_ori_n632_), .B(ori_ori_n265_), .Y(ori_ori_n754_));
  AOI210     o732(.A0(ori_ori_n383_), .A1(ori_ori_n89_), .B0(ori_ori_n58_), .Y(ori_ori_n755_));
  NO2        o733(.A(ori_ori_n755_), .B(ori_ori_n754_), .Y(ori_ori_n756_));
  NO2        o734(.A(ori_ori_n228_), .B(ori_ori_n156_), .Y(ori_ori_n757_));
  NA2        o735(.A(i_0_), .B(i_10_), .Y(ori_ori_n758_));
  INV        o736(.A(ori_ori_n420_), .Y(ori_ori_n759_));
  NO4        o737(.A(ori_ori_n118_), .B(ori_ori_n58_), .C(ori_ori_n548_), .D(i_5_), .Y(ori_ori_n760_));
  AO220      o738(.A0(ori_ori_n760_), .A1(ori_ori_n759_), .B0(ori_ori_n757_), .B1(i_6_), .Y(ori_ori_n761_));
  NO2        o739(.A(ori_ori_n761_), .B(ori_ori_n756_), .Y(ori_ori_n762_));
  NA3        o740(.A(ori_ori_n762_), .B(ori_ori_n752_), .C(ori_ori_n748_), .Y(ori_ori_n763_));
  NO2        o741(.A(ori_ori_n106_), .B(ori_ori_n37_), .Y(ori_ori_n764_));
  NA2        o742(.A(i_11_), .B(i_9_), .Y(ori_ori_n765_));
  NO3        o743(.A(i_12_), .B(ori_ori_n765_), .C(ori_ori_n480_), .Y(ori_ori_n766_));
  AN2        o744(.A(ori_ori_n766_), .B(ori_ori_n764_), .Y(ori_ori_n767_));
  NO2        o745(.A(ori_ori_n48_), .B(i_7_), .Y(ori_ori_n768_));
  NA2        o746(.A(ori_ori_n316_), .B(ori_ori_n171_), .Y(ori_ori_n769_));
  NA2        o747(.A(ori_ori_n769_), .B(ori_ori_n160_), .Y(ori_ori_n770_));
  NO2        o748(.A(ori_ori_n765_), .B(ori_ori_n73_), .Y(ori_ori_n771_));
  NO2        o749(.A(ori_ori_n169_), .B(i_0_), .Y(ori_ori_n772_));
  INV        o750(.A(ori_ori_n324_), .Y(ori_ori_n773_));
  NO2        o751(.A(ori_ori_n773_), .B(ori_ori_n738_), .Y(ori_ori_n774_));
  NO3        o752(.A(ori_ori_n774_), .B(ori_ori_n770_), .C(ori_ori_n767_), .Y(ori_ori_n775_));
  NA2        o753(.A(ori_ori_n537_), .B(ori_ori_n125_), .Y(ori_ori_n776_));
  NO2        o754(.A(i_6_), .B(ori_ori_n776_), .Y(ori_ori_n777_));
  AOI210     o755(.A0(ori_ori_n349_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n778_));
  NA2        o756(.A(ori_ori_n166_), .B(ori_ori_n106_), .Y(ori_ori_n779_));
  NOi32      o757(.An(ori_ori_n778_), .Bn(ori_ori_n177_), .C(ori_ori_n779_), .Y(ori_ori_n780_));
  NA2        o758(.A(ori_ori_n482_), .B(ori_ori_n265_), .Y(ori_ori_n781_));
  NO2        o759(.A(ori_ori_n781_), .B(ori_ori_n729_), .Y(ori_ori_n782_));
  NO3        o760(.A(ori_ori_n782_), .B(ori_ori_n780_), .C(ori_ori_n777_), .Y(ori_ori_n783_));
  NOi21      o761(.An(i_7_), .B(i_5_), .Y(ori_ori_n784_));
  NOi31      o762(.An(ori_ori_n784_), .B(i_0_), .C(ori_ori_n609_), .Y(ori_ori_n785_));
  NA3        o763(.A(ori_ori_n785_), .B(ori_ori_n310_), .C(i_6_), .Y(ori_ori_n786_));
  BUFFER     o764(.A(ori_ori_n786_), .Y(ori_ori_n787_));
  INV        o765(.A(ori_ori_n262_), .Y(ori_ori_n788_));
  NA3        o766(.A(ori_ori_n787_), .B(ori_ori_n783_), .C(ori_ori_n775_), .Y(ori_ori_n789_));
  NO2        o767(.A(ori_ori_n723_), .B(ori_ori_n261_), .Y(ori_ori_n790_));
  OA210      o768(.A0(ori_ori_n378_), .A1(ori_ori_n207_), .B0(ori_ori_n377_), .Y(ori_ori_n791_));
  NA2        o769(.A(ori_ori_n790_), .B(ori_ori_n771_), .Y(ori_ori_n792_));
  NA3        o770(.A(ori_ori_n377_), .B(ori_ori_n327_), .C(ori_ori_n45_), .Y(ori_ori_n793_));
  OAI210     o771(.A0(ori_ori_n746_), .A1(ori_ori_n753_), .B0(ori_ori_n793_), .Y(ori_ori_n794_));
  NA2        o772(.A(ori_ori_n771_), .B(ori_ori_n256_), .Y(ori_ori_n795_));
  OAI210     o773(.A0(i_2_), .A1(ori_ori_n176_), .B0(ori_ori_n795_), .Y(ori_ori_n796_));
  AOI220     o774(.A0(ori_ori_n796_), .A1(ori_ori_n378_), .B0(ori_ori_n794_), .B1(ori_ori_n73_), .Y(ori_ori_n797_));
  NA3        o775(.A(ori_ori_n700_), .B(ori_ori_n308_), .C(ori_ori_n520_), .Y(ori_ori_n798_));
  NO2        o776(.A(ori_ori_n75_), .B(ori_ori_n634_), .Y(ori_ori_n799_));
  AOI220     o777(.A0(ori_ori_n799_), .A1(i_11_), .B0(ori_ori_n168_), .B1(ori_ori_n470_), .Y(ori_ori_n800_));
  AOI210     o778(.A0(ori_ori_n800_), .A1(ori_ori_n798_), .B0(ori_ori_n47_), .Y(ori_ori_n801_));
  NO3        o779(.A(ori_ori_n461_), .B(ori_ori_n280_), .C(ori_ori_n24_), .Y(ori_ori_n802_));
  AOI210     o780(.A0(ori_ori_n582_), .A1(ori_ori_n427_), .B0(ori_ori_n802_), .Y(ori_ori_n803_));
  NAi21      o781(.An(i_9_), .B(i_5_), .Y(ori_ori_n804_));
  NO2        o782(.A(ori_ori_n804_), .B(ori_ori_n321_), .Y(ori_ori_n805_));
  NA2        o783(.A(ori_ori_n805_), .B(ori_ori_n499_), .Y(ori_ori_n806_));
  OAI220     o784(.A0(ori_ori_n806_), .A1(ori_ori_n86_), .B0(ori_ori_n803_), .B1(ori_ori_n167_), .Y(ori_ori_n807_));
  NO3        o785(.A(ori_ori_n807_), .B(ori_ori_n801_), .C(ori_ori_n412_), .Y(ori_ori_n808_));
  NA3        o786(.A(ori_ori_n808_), .B(ori_ori_n797_), .C(ori_ori_n792_), .Y(ori_ori_n809_));
  NO3        o787(.A(ori_ori_n809_), .B(ori_ori_n789_), .C(ori_ori_n763_), .Y(ori_ori_n810_));
  NO2        o788(.A(i_0_), .B(ori_ori_n609_), .Y(ori_ori_n811_));
  AOI210     o789(.A0(ori_ori_n682_), .A1(ori_ori_n566_), .B0(ori_ori_n779_), .Y(ori_ori_n812_));
  INV        o790(.A(ori_ori_n812_), .Y(ori_ori_n813_));
  OAI210     o791(.A0(ori_ori_n221_), .A1(i_9_), .B0(ori_ori_n213_), .Y(ori_ori_n814_));
  AOI210     o792(.A0(ori_ori_n814_), .A1(ori_ori_n749_), .B0(ori_ori_n156_), .Y(ori_ori_n815_));
  INV        o793(.A(ori_ori_n815_), .Y(ori_ori_n816_));
  NA2        o794(.A(ori_ori_n816_), .B(ori_ori_n813_), .Y(ori_ori_n817_));
  NO3        o795(.A(ori_ori_n758_), .B(ori_ori_n737_), .C(ori_ori_n179_), .Y(ori_ori_n818_));
  AOI220     o796(.A0(ori_ori_n818_), .A1(i_11_), .B0(ori_ori_n446_), .B1(ori_ori_n75_), .Y(ori_ori_n819_));
  NO3        o797(.A(ori_ori_n194_), .B(ori_ori_n309_), .C(i_0_), .Y(ori_ori_n820_));
  OAI210     o798(.A0(ori_ori_n820_), .A1(ori_ori_n76_), .B0(i_13_), .Y(ori_ori_n821_));
  NA2        o799(.A(ori_ori_n821_), .B(ori_ori_n819_), .Y(ori_ori_n822_));
  NO2        o800(.A(ori_ori_n220_), .B(ori_ori_n95_), .Y(ori_ori_n823_));
  AOI210     o801(.A0(ori_ori_n823_), .A1(ori_ori_n811_), .B0(ori_ori_n112_), .Y(ori_ori_n824_));
  OR2        o802(.A(ori_ori_n824_), .B(i_5_), .Y(ori_ori_n825_));
  AOI210     o803(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n169_), .Y(ori_ori_n826_));
  NA2        o804(.A(ori_ori_n826_), .B(ori_ori_n791_), .Y(ori_ori_n827_));
  INV        o805(.A(ori_ori_n425_), .Y(ori_ori_n828_));
  NO3        o806(.A(ori_ori_n729_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n829_));
  NA2        o807(.A(ori_ori_n391_), .B(ori_ori_n384_), .Y(ori_ori_n830_));
  NO3        o808(.A(ori_ori_n830_), .B(ori_ori_n829_), .C(ori_ori_n828_), .Y(ori_ori_n831_));
  NA3        o809(.A(ori_ori_n315_), .B(ori_ori_n166_), .C(ori_ori_n165_), .Y(ori_ori_n832_));
  NA3        o810(.A(ori_ori_n768_), .B(ori_ori_n254_), .C(ori_ori_n213_), .Y(ori_ori_n833_));
  NA2        o811(.A(ori_ori_n833_), .B(ori_ori_n832_), .Y(ori_ori_n834_));
  NO3        o812(.A(ori_ori_n765_), .B(ori_ori_n201_), .C(ori_ori_n179_), .Y(ori_ori_n835_));
  NO2        o813(.A(ori_ori_n835_), .B(ori_ori_n834_), .Y(ori_ori_n836_));
  NA4        o814(.A(ori_ori_n836_), .B(ori_ori_n831_), .C(ori_ori_n827_), .D(ori_ori_n825_), .Y(ori_ori_n837_));
  NO2        o815(.A(ori_ori_n86_), .B(i_5_), .Y(ori_ori_n838_));
  NA3        o816(.A(ori_ori_n724_), .B(ori_ori_n113_), .C(ori_ori_n128_), .Y(ori_ori_n839_));
  INV        o817(.A(ori_ori_n839_), .Y(ori_ori_n840_));
  NA2        o818(.A(ori_ori_n840_), .B(ori_ori_n838_), .Y(ori_ori_n841_));
  NA3        o819(.A(ori_ori_n256_), .B(i_5_), .C(ori_ori_n180_), .Y(ori_ori_n842_));
  NAi31      o820(.An(ori_ori_n219_), .B(ori_ori_n842_), .C(ori_ori_n220_), .Y(ori_ori_n843_));
  NO4        o821(.A(ori_ori_n218_), .B(ori_ori_n194_), .C(i_0_), .D(i_12_), .Y(ori_ori_n844_));
  AOI220     o822(.A0(ori_ori_n844_), .A1(ori_ori_n843_), .B0(ori_ori_n676_), .B1(ori_ori_n170_), .Y(ori_ori_n845_));
  NA2        o823(.A(ori_ori_n784_), .B(ori_ori_n375_), .Y(ori_ori_n846_));
  NA2        o824(.A(ori_ori_n64_), .B(ori_ori_n104_), .Y(ori_ori_n847_));
  OAI220     o825(.A0(ori_ori_n847_), .A1(ori_ori_n842_), .B0(ori_ori_n846_), .B1(ori_ori_n556_), .Y(ori_ori_n848_));
  NA2        o826(.A(ori_ori_n848_), .B(ori_ori_n772_), .Y(ori_ori_n849_));
  NA3        o827(.A(ori_ori_n849_), .B(ori_ori_n845_), .C(ori_ori_n841_), .Y(ori_ori_n850_));
  NO4        o828(.A(ori_ori_n850_), .B(ori_ori_n837_), .C(ori_ori_n822_), .D(ori_ori_n817_), .Y(ori_ori_n851_));
  OAI210     o829(.A0(ori_ori_n699_), .A1(ori_ori_n695_), .B0(ori_ori_n37_), .Y(ori_ori_n852_));
  NA2        o830(.A(ori_ori_n852_), .B(ori_ori_n488_), .Y(ori_ori_n853_));
  NA2        o831(.A(ori_ori_n853_), .B(ori_ori_n192_), .Y(ori_ori_n854_));
  NA2        o832(.A(ori_ori_n175_), .B(ori_ori_n177_), .Y(ori_ori_n855_));
  AO210      o833(.A0(ori_ori_n577_), .A1(ori_ori_n33_), .B0(ori_ori_n855_), .Y(ori_ori_n856_));
  NAi31      o834(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n857_));
  AOI210     o835(.A0(ori_ori_n121_), .A1(ori_ori_n70_), .B0(ori_ori_n857_), .Y(ori_ori_n858_));
  NO2        o836(.A(ori_ori_n858_), .B(ori_ori_n523_), .Y(ori_ori_n859_));
  NA2        o837(.A(ori_ori_n859_), .B(ori_ori_n856_), .Y(ori_ori_n860_));
  NO2        o838(.A(ori_ori_n367_), .B(ori_ori_n241_), .Y(ori_ori_n861_));
  NO2        o839(.A(ori_ori_n861_), .B(ori_ori_n751_), .Y(ori_ori_n862_));
  INV        o840(.A(ori_ori_n862_), .Y(ori_ori_n863_));
  AOI210     o841(.A0(ori_ori_n860_), .A1(ori_ori_n48_), .B0(ori_ori_n863_), .Y(ori_ori_n864_));
  AOI210     o842(.A0(ori_ori_n864_), .A1(ori_ori_n854_), .B0(ori_ori_n73_), .Y(ori_ori_n865_));
  INV        o843(.A(ori_ori_n305_), .Y(ori_ori_n866_));
  NO2        o844(.A(ori_ori_n866_), .B(ori_ori_n640_), .Y(ori_ori_n867_));
  OAI210     o845(.A0(ori_ori_n80_), .A1(ori_ori_n54_), .B0(ori_ori_n111_), .Y(ori_ori_n868_));
  NA2        o846(.A(ori_ori_n868_), .B(ori_ori_n76_), .Y(ori_ori_n869_));
  AOI210     o847(.A0(ori_ori_n826_), .A1(ori_ori_n768_), .B0(ori_ori_n785_), .Y(ori_ori_n870_));
  AOI210     o848(.A0(ori_ori_n870_), .A1(ori_ori_n869_), .B0(ori_ori_n559_), .Y(ori_ori_n871_));
  INV        o849(.A(ori_ori_n871_), .Y(ori_ori_n872_));
  OAI210     o850(.A0(ori_ori_n243_), .A1(ori_ori_n158_), .B0(ori_ori_n89_), .Y(ori_ori_n873_));
  NA3        o851(.A(ori_ori_n644_), .B(ori_ori_n254_), .C(ori_ori_n80_), .Y(ori_ori_n874_));
  AOI210     o852(.A0(ori_ori_n874_), .A1(ori_ori_n873_), .B0(i_11_), .Y(ori_ori_n875_));
  NA2        o853(.A(ori_ori_n483_), .B(ori_ori_n198_), .Y(ori_ori_n876_));
  OAI210     o854(.A0(ori_ori_n876_), .A1(ori_ori_n778_), .B0(ori_ori_n192_), .Y(ori_ori_n877_));
  NA2        o855(.A(ori_ori_n163_), .B(i_5_), .Y(ori_ori_n878_));
  NO2        o856(.A(ori_ori_n877_), .B(ori_ori_n878_), .Y(ori_ori_n879_));
  NO3        o857(.A(ori_ori_n59_), .B(ori_ori_n58_), .C(i_4_), .Y(ori_ori_n880_));
  OAI210     o858(.A0(ori_ori_n788_), .A1(ori_ori_n257_), .B0(ori_ori_n880_), .Y(ori_ori_n881_));
  NO2        o859(.A(ori_ori_n881_), .B(ori_ori_n609_), .Y(ori_ori_n882_));
  NO4        o860(.A(ori_ori_n804_), .B(ori_ori_n380_), .C(ori_ori_n227_), .D(ori_ori_n226_), .Y(ori_ori_n883_));
  NO2        o861(.A(ori_ori_n883_), .B(ori_ori_n443_), .Y(ori_ori_n884_));
  INV        o862(.A(ori_ori_n286_), .Y(ori_ori_n885_));
  AOI210     o863(.A0(ori_ori_n885_), .A1(ori_ori_n884_), .B0(ori_ori_n41_), .Y(ori_ori_n886_));
  NO4        o864(.A(ori_ori_n886_), .B(ori_ori_n882_), .C(ori_ori_n879_), .D(ori_ori_n875_), .Y(ori_ori_n887_));
  OAI210     o865(.A0(ori_ori_n872_), .A1(i_4_), .B0(ori_ori_n887_), .Y(ori_ori_n888_));
  NO3        o866(.A(ori_ori_n888_), .B(ori_ori_n867_), .C(ori_ori_n865_), .Y(ori_ori_n889_));
  NA4        o867(.A(ori_ori_n889_), .B(ori_ori_n851_), .C(ori_ori_n810_), .D(ori_ori_n742_), .Y(ori4));
  INV        o868(.A(ori_ori_n581_), .Y(ori_ori_n893_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m0033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m0034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m0036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m0037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m0038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m0039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m0040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m0041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m0042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m0043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m0044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m0045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m0046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m0047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m0049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m0050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m0051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m0052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m0053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m0054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m0055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m0057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m0059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m0060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m0062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m0063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m0064(.A(i_6_), .Y(mai_mai_n87_));
  NO2        m0065(.A(i_2_), .B(i_7_), .Y(mai_mai_n88_));
  INV        m0066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OAI210     m0067(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NAi21      m0068(.An(i_6_), .B(i_10_), .Y(mai_mai_n91_));
  NA2        m0069(.A(i_6_), .B(i_9_), .Y(mai_mai_n92_));
  AOI210     m0070(.A0(mai_mai_n92_), .A1(mai_mai_n91_), .B0(mai_mai_n64_), .Y(mai_mai_n93_));
  NA2        m0071(.A(i_2_), .B(i_6_), .Y(mai_mai_n94_));
  NO3        m0072(.A(mai_mai_n94_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n95_));
  NO2        m0073(.A(mai_mai_n95_), .B(mai_mai_n93_), .Y(mai_mai_n96_));
  AOI210     m0074(.A0(mai_mai_n96_), .A1(mai_mai_n90_), .B0(mai_mai_n81_), .Y(mai_mai_n97_));
  AN3        m0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n98_));
  NAi21      m0076(.An(i_6_), .B(i_11_), .Y(mai_mai_n99_));
  NO2        m0077(.A(i_5_), .B(i_8_), .Y(mai_mai_n100_));
  NOi21      m0078(.An(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  AOI220     m0079(.A0(mai_mai_n101_), .A1(mai_mai_n63_), .B0(mai_mai_n98_), .B1(mai_mai_n32_), .Y(mai_mai_n102_));
  INV        m0080(.A(i_7_), .Y(mai_mai_n103_));
  NA2        m0081(.A(mai_mai_n47_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m0082(.A(i_0_), .B(i_5_), .Y(mai_mai_n105_));
  NO2        m0083(.A(mai_mai_n105_), .B(mai_mai_n87_), .Y(mai_mai_n106_));
  NA2        m0084(.A(i_12_), .B(i_3_), .Y(mai_mai_n107_));
  INV        m0085(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NA3        m0086(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n104_), .Y(mai_mai_n109_));
  NAi21      m0087(.An(i_7_), .B(i_11_), .Y(mai_mai_n110_));
  NO3        m0088(.A(mai_mai_n110_), .B(mai_mai_n91_), .C(mai_mai_n54_), .Y(mai_mai_n111_));
  AN2        m0089(.A(i_2_), .B(i_10_), .Y(mai_mai_n112_));
  NO2        m0090(.A(mai_mai_n112_), .B(i_7_), .Y(mai_mai_n113_));
  OR2        m0091(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n114_));
  NO2        m0092(.A(i_8_), .B(mai_mai_n103_), .Y(mai_mai_n115_));
  NO3        m0093(.A(mai_mai_n115_), .B(mai_mai_n114_), .C(mai_mai_n113_), .Y(mai_mai_n116_));
  NA2        m0094(.A(i_12_), .B(i_7_), .Y(mai_mai_n117_));
  NO2        m0095(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n118_));
  NA2        m0096(.A(mai_mai_n118_), .B(i_0_), .Y(mai_mai_n119_));
  NA2        m0097(.A(i_11_), .B(i_12_), .Y(mai_mai_n120_));
  OAI210     m0098(.A0(mai_mai_n119_), .A1(mai_mai_n117_), .B0(mai_mai_n120_), .Y(mai_mai_n121_));
  NO2        m0099(.A(mai_mai_n121_), .B(mai_mai_n116_), .Y(mai_mai_n122_));
  NAi41      m0100(.An(mai_mai_n111_), .B(mai_mai_n122_), .C(mai_mai_n109_), .D(mai_mai_n102_), .Y(mai_mai_n123_));
  NOi21      m0101(.An(i_1_), .B(i_5_), .Y(mai_mai_n124_));
  NA2        m0102(.A(mai_mai_n124_), .B(i_11_), .Y(mai_mai_n125_));
  NA2        m0103(.A(mai_mai_n103_), .B(mai_mai_n37_), .Y(mai_mai_n126_));
  NA2        m0104(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n127_));
  NA2        m0105(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NO2        m0106(.A(mai_mai_n128_), .B(mai_mai_n47_), .Y(mai_mai_n129_));
  NA2        m0107(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n130_));
  NAi21      m0108(.An(i_3_), .B(i_8_), .Y(mai_mai_n131_));
  NA2        m0109(.A(mai_mai_n131_), .B(mai_mai_n63_), .Y(mai_mai_n132_));
  NOi31      m0110(.An(mai_mai_n132_), .B(mai_mai_n130_), .C(mai_mai_n129_), .Y(mai_mai_n133_));
  NO2        m0111(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n134_));
  NO2        m0112(.A(i_6_), .B(i_5_), .Y(mai_mai_n135_));
  NA2        m0113(.A(mai_mai_n135_), .B(i_3_), .Y(mai_mai_n136_));
  AO210      m0114(.A0(mai_mai_n136_), .A1(mai_mai_n48_), .B0(mai_mai_n134_), .Y(mai_mai_n137_));
  OAI220     m0115(.A0(mai_mai_n137_), .A1(mai_mai_n110_), .B0(mai_mai_n133_), .B1(mai_mai_n125_), .Y(mai_mai_n138_));
  NO3        m0116(.A(mai_mai_n138_), .B(mai_mai_n123_), .C(mai_mai_n97_), .Y(mai_mai_n139_));
  NA3        m0117(.A(mai_mai_n139_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m0118(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n141_));
  NA2        m0119(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n142_));
  NA2        m0120(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  NA4        m0121(.A(mai_mai_n143_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0122(.A(i_8_), .B(i_7_), .Y(mai_mai_n145_));
  NA2        m0123(.A(mai_mai_n145_), .B(i_6_), .Y(mai_mai_n146_));
  NO2        m0124(.A(i_12_), .B(i_13_), .Y(mai_mai_n147_));
  NAi21      m0125(.An(i_5_), .B(i_11_), .Y(mai_mai_n148_));
  NOi21      m0126(.An(mai_mai_n147_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  NO2        m0127(.A(i_0_), .B(i_1_), .Y(mai_mai_n150_));
  NA2        m0128(.A(i_2_), .B(i_3_), .Y(mai_mai_n151_));
  NO2        m0129(.A(mai_mai_n151_), .B(i_4_), .Y(mai_mai_n152_));
  NA3        m0130(.A(mai_mai_n152_), .B(mai_mai_n150_), .C(mai_mai_n149_), .Y(mai_mai_n153_));
  AN2        m0131(.A(mai_mai_n147_), .B(mai_mai_n84_), .Y(mai_mai_n154_));
  NO2        m0132(.A(mai_mai_n154_), .B(mai_mai_n27_), .Y(mai_mai_n155_));
  NA2        m0133(.A(i_1_), .B(i_5_), .Y(mai_mai_n156_));
  NO2        m0134(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n157_));
  NA2        m0135(.A(mai_mai_n157_), .B(mai_mai_n36_), .Y(mai_mai_n158_));
  NO3        m0136(.A(mai_mai_n158_), .B(mai_mai_n156_), .C(mai_mai_n155_), .Y(mai_mai_n159_));
  OR2        m0137(.A(i_0_), .B(i_1_), .Y(mai_mai_n160_));
  NO3        m0138(.A(mai_mai_n160_), .B(mai_mai_n81_), .C(i_13_), .Y(mai_mai_n161_));
  NAi32      m0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n162_));
  NAi21      m0140(.An(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  NOi21      m0141(.An(i_4_), .B(i_10_), .Y(mai_mai_n164_));
  NA2        m0142(.A(mai_mai_n164_), .B(mai_mai_n40_), .Y(mai_mai_n165_));
  NO2        m0143(.A(i_3_), .B(i_5_), .Y(mai_mai_n166_));
  NO3        m0144(.A(mai_mai_n74_), .B(i_2_), .C(i_1_), .Y(mai_mai_n167_));
  NA2        m0145(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  OAI210     m0146(.A0(mai_mai_n168_), .A1(mai_mai_n165_), .B0(mai_mai_n163_), .Y(mai_mai_n169_));
  NO2        m0147(.A(mai_mai_n169_), .B(mai_mai_n159_), .Y(mai_mai_n170_));
  AOI210     m0148(.A0(mai_mai_n170_), .A1(mai_mai_n153_), .B0(mai_mai_n146_), .Y(mai_mai_n171_));
  NA3        m0149(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n172_));
  NA2        m0150(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n173_));
  NOi21      m0151(.An(i_4_), .B(i_9_), .Y(mai_mai_n174_));
  NOi21      m0152(.An(i_11_), .B(i_13_), .Y(mai_mai_n175_));
  NA2        m0153(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  OR2        m0154(.A(mai_mai_n176_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  NO2        m0155(.A(i_4_), .B(i_5_), .Y(mai_mai_n178_));
  NAi21      m0156(.An(i_12_), .B(i_11_), .Y(mai_mai_n179_));
  NO2        m0157(.A(mai_mai_n179_), .B(i_13_), .Y(mai_mai_n180_));
  NA3        m0158(.A(mai_mai_n180_), .B(mai_mai_n178_), .C(mai_mai_n84_), .Y(mai_mai_n181_));
  AOI210     m0159(.A0(mai_mai_n181_), .A1(mai_mai_n177_), .B0(mai_mai_n172_), .Y(mai_mai_n182_));
  NO2        m0160(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n183_));
  NA2        m0161(.A(mai_mai_n183_), .B(mai_mai_n47_), .Y(mai_mai_n184_));
  NA2        m0162(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n185_));
  NAi31      m0163(.An(mai_mai_n185_), .B(mai_mai_n154_), .C(i_11_), .Y(mai_mai_n186_));
  NA2        m0164(.A(i_3_), .B(i_5_), .Y(mai_mai_n187_));
  OR2        m0165(.A(mai_mai_n187_), .B(mai_mai_n176_), .Y(mai_mai_n188_));
  AOI210     m0166(.A0(mai_mai_n188_), .A1(mai_mai_n186_), .B0(mai_mai_n184_), .Y(mai_mai_n189_));
  NO2        m0167(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n190_));
  NO2        m0168(.A(i_13_), .B(i_10_), .Y(mai_mai_n191_));
  NA3        m0169(.A(mai_mai_n191_), .B(mai_mai_n190_), .C(mai_mai_n45_), .Y(mai_mai_n192_));
  NO2        m0170(.A(i_2_), .B(i_1_), .Y(mai_mai_n193_));
  NA2        m0171(.A(mai_mai_n193_), .B(i_3_), .Y(mai_mai_n194_));
  NAi21      m0172(.An(i_4_), .B(i_12_), .Y(mai_mai_n195_));
  NO4        m0173(.A(mai_mai_n195_), .B(mai_mai_n194_), .C(mai_mai_n192_), .D(mai_mai_n25_), .Y(mai_mai_n196_));
  NO3        m0174(.A(mai_mai_n196_), .B(mai_mai_n189_), .C(mai_mai_n182_), .Y(mai_mai_n197_));
  INV        m0175(.A(i_8_), .Y(mai_mai_n198_));
  NO2        m0176(.A(mai_mai_n198_), .B(i_7_), .Y(mai_mai_n199_));
  NA2        m0177(.A(mai_mai_n199_), .B(i_6_), .Y(mai_mai_n200_));
  NO3        m0178(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n201_));
  NA2        m0179(.A(mai_mai_n201_), .B(mai_mai_n115_), .Y(mai_mai_n202_));
  NO3        m0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n203_));
  NA3        m0181(.A(mai_mai_n203_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n204_));
  NO3        m0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n205_));
  OAI210     m0183(.A0(mai_mai_n98_), .A1(i_12_), .B0(mai_mai_n205_), .Y(mai_mai_n206_));
  AOI210     m0184(.A0(mai_mai_n206_), .A1(mai_mai_n204_), .B0(mai_mai_n202_), .Y(mai_mai_n207_));
  NO2        m0185(.A(i_3_), .B(i_8_), .Y(mai_mai_n208_));
  NO3        m0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n209_));
  NO2        m0187(.A(mai_mai_n105_), .B(mai_mai_n59_), .Y(mai_mai_n210_));
  NO2        m0188(.A(i_13_), .B(i_9_), .Y(mai_mai_n211_));
  NA3        m0189(.A(mai_mai_n211_), .B(i_6_), .C(mai_mai_n198_), .Y(mai_mai_n212_));
  NAi21      m0190(.An(i_12_), .B(i_3_), .Y(mai_mai_n213_));
  NO2        m0191(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n214_));
  NO3        m0192(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n215_));
  NA3        m0193(.A(mai_mai_n215_), .B(mai_mai_n214_), .C(i_10_), .Y(mai_mai_n216_));
  NO2        m0194(.A(mai_mai_n216_), .B(mai_mai_n212_), .Y(mai_mai_n217_));
  AOI210     m0195(.A0(mai_mai_n217_), .A1(i_7_), .B0(mai_mai_n207_), .Y(mai_mai_n218_));
  OAI220     m0196(.A0(mai_mai_n218_), .A1(i_4_), .B0(mai_mai_n200_), .B1(mai_mai_n197_), .Y(mai_mai_n219_));
  NAi21      m0197(.An(i_12_), .B(i_7_), .Y(mai_mai_n220_));
  NA3        m0198(.A(i_13_), .B(mai_mai_n198_), .C(i_10_), .Y(mai_mai_n221_));
  NA2        m0199(.A(i_0_), .B(i_5_), .Y(mai_mai_n222_));
  NAi31      m0200(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n223_));
  NO2        m0201(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n224_));
  NO2        m0202(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n225_));
  NO2        m0203(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n226_));
  NA3        m0204(.A(mai_mai_n226_), .B(mai_mai_n225_), .C(mai_mai_n224_), .Y(mai_mai_n227_));
  INV        m0205(.A(i_13_), .Y(mai_mai_n228_));
  NO2        m0206(.A(i_12_), .B(mai_mai_n228_), .Y(mai_mai_n229_));
  NO2        m0207(.A(mai_mai_n227_), .B(mai_mai_n223_), .Y(mai_mai_n230_));
  NA2        m0208(.A(mai_mai_n230_), .B(mai_mai_n145_), .Y(mai_mai_n231_));
  NO2        m0209(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n232_));
  NO2        m0210(.A(mai_mai_n187_), .B(i_4_), .Y(mai_mai_n233_));
  NA2        m0211(.A(mai_mai_n233_), .B(mai_mai_n232_), .Y(mai_mai_n234_));
  OR2        m0212(.A(i_8_), .B(i_7_), .Y(mai_mai_n235_));
  NO2        m0213(.A(mai_mai_n235_), .B(mai_mai_n87_), .Y(mai_mai_n236_));
  NO2        m0214(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n237_));
  NA2        m0215(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  INV        m0216(.A(i_12_), .Y(mai_mai_n239_));
  NO2        m0217(.A(mai_mai_n45_), .B(mai_mai_n239_), .Y(mai_mai_n240_));
  NO3        m0218(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n241_));
  NA2        m0219(.A(i_2_), .B(i_1_), .Y(mai_mai_n242_));
  NO2        m0220(.A(mai_mai_n238_), .B(mai_mai_n234_), .Y(mai_mai_n243_));
  NO3        m0221(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n244_));
  NAi21      m0222(.An(i_4_), .B(i_3_), .Y(mai_mai_n245_));
  NO2        m0223(.A(mai_mai_n245_), .B(mai_mai_n76_), .Y(mai_mai_n246_));
  NO2        m0224(.A(i_0_), .B(i_6_), .Y(mai_mai_n247_));
  NOi41      m0225(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n248_));
  NA2        m0226(.A(mai_mai_n248_), .B(mai_mai_n247_), .Y(mai_mai_n249_));
  NO2        m0227(.A(mai_mai_n242_), .B(mai_mai_n187_), .Y(mai_mai_n250_));
  NAi21      m0228(.An(mai_mai_n249_), .B(mai_mai_n250_), .Y(mai_mai_n251_));
  INV        m0229(.A(mai_mai_n251_), .Y(mai_mai_n252_));
  AOI220     m0230(.A0(mai_mai_n252_), .A1(mai_mai_n40_), .B0(mai_mai_n243_), .B1(mai_mai_n211_), .Y(mai_mai_n253_));
  NO2        m0231(.A(i_11_), .B(mai_mai_n228_), .Y(mai_mai_n254_));
  NOi21      m0232(.An(i_1_), .B(i_6_), .Y(mai_mai_n255_));
  NAi21      m0233(.An(i_3_), .B(i_7_), .Y(mai_mai_n256_));
  NA2        m0234(.A(mai_mai_n239_), .B(i_9_), .Y(mai_mai_n257_));
  OR4        m0235(.A(mai_mai_n257_), .B(mai_mai_n256_), .C(mai_mai_n255_), .D(mai_mai_n190_), .Y(mai_mai_n258_));
  NO2        m0236(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n259_));
  NO2        m0237(.A(i_12_), .B(i_3_), .Y(mai_mai_n260_));
  NA2        m0238(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n261_));
  NA2        m0239(.A(i_3_), .B(i_9_), .Y(mai_mai_n262_));
  NAi21      m0240(.An(i_7_), .B(i_10_), .Y(mai_mai_n263_));
  NO2        m0241(.A(mai_mai_n263_), .B(mai_mai_n262_), .Y(mai_mai_n264_));
  NA3        m0242(.A(mai_mai_n264_), .B(mai_mai_n261_), .C(mai_mai_n65_), .Y(mai_mai_n265_));
  NA2        m0243(.A(mai_mai_n265_), .B(mai_mai_n258_), .Y(mai_mai_n266_));
  NA3        m0244(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n267_));
  INV        m0245(.A(mai_mai_n146_), .Y(mai_mai_n268_));
  NA2        m0246(.A(mai_mai_n239_), .B(i_13_), .Y(mai_mai_n269_));
  NO2        m0247(.A(mai_mai_n269_), .B(mai_mai_n76_), .Y(mai_mai_n270_));
  AOI220     m0248(.A0(mai_mai_n270_), .A1(mai_mai_n268_), .B0(mai_mai_n266_), .B1(mai_mai_n254_), .Y(mai_mai_n271_));
  NO2        m0249(.A(mai_mai_n235_), .B(mai_mai_n37_), .Y(mai_mai_n272_));
  NA2        m0250(.A(i_12_), .B(i_6_), .Y(mai_mai_n273_));
  OR2        m0251(.A(i_13_), .B(i_9_), .Y(mai_mai_n274_));
  NO2        m0252(.A(mai_mai_n245_), .B(i_2_), .Y(mai_mai_n275_));
  NA2        m0253(.A(mai_mai_n254_), .B(i_9_), .Y(mai_mai_n276_));
  NA2        m0254(.A(mai_mai_n157_), .B(mai_mai_n64_), .Y(mai_mai_n277_));
  NO3        m0255(.A(i_11_), .B(mai_mai_n228_), .C(mai_mai_n25_), .Y(mai_mai_n278_));
  NO2        m0256(.A(mai_mai_n256_), .B(i_8_), .Y(mai_mai_n279_));
  NO2        m0257(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n280_));
  NA3        m0258(.A(mai_mai_n280_), .B(mai_mai_n279_), .C(mai_mai_n278_), .Y(mai_mai_n281_));
  NO3        m0259(.A(mai_mai_n26_), .B(mai_mai_n87_), .C(i_5_), .Y(mai_mai_n282_));
  NA3        m0260(.A(mai_mai_n282_), .B(mai_mai_n272_), .C(mai_mai_n229_), .Y(mai_mai_n283_));
  AOI210     m0261(.A0(mai_mai_n283_), .A1(mai_mai_n281_), .B0(mai_mai_n277_), .Y(mai_mai_n284_));
  INV        m0262(.A(mai_mai_n284_), .Y(mai_mai_n285_));
  NA4        m0263(.A(mai_mai_n285_), .B(mai_mai_n271_), .C(mai_mai_n253_), .D(mai_mai_n231_), .Y(mai_mai_n286_));
  NO3        m0264(.A(i_12_), .B(mai_mai_n228_), .C(mai_mai_n37_), .Y(mai_mai_n287_));
  INV        m0265(.A(mai_mai_n287_), .Y(mai_mai_n288_));
  NA2        m0266(.A(i_8_), .B(mai_mai_n103_), .Y(mai_mai_n289_));
  NOi21      m0267(.An(mai_mai_n166_), .B(mai_mai_n87_), .Y(mai_mai_n290_));
  NO3        m0268(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n291_));
  AOI220     m0269(.A0(mai_mai_n291_), .A1(mai_mai_n201_), .B0(mai_mai_n290_), .B1(mai_mai_n237_), .Y(mai_mai_n292_));
  NO2        m0270(.A(mai_mai_n292_), .B(mai_mai_n289_), .Y(mai_mai_n293_));
  NO3        m0271(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n294_));
  NO2        m0272(.A(mai_mai_n242_), .B(i_0_), .Y(mai_mai_n295_));
  AOI220     m0273(.A0(mai_mai_n295_), .A1(mai_mai_n199_), .B0(mai_mai_n294_), .B1(mai_mai_n145_), .Y(mai_mai_n296_));
  NA2        m0274(.A(mai_mai_n280_), .B(mai_mai_n26_), .Y(mai_mai_n297_));
  NO2        m0275(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  NA2        m0276(.A(i_0_), .B(i_1_), .Y(mai_mai_n299_));
  NO2        m0277(.A(mai_mai_n299_), .B(i_2_), .Y(mai_mai_n300_));
  NO2        m0278(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n301_));
  NA3        m0279(.A(mai_mai_n301_), .B(mai_mai_n300_), .C(mai_mai_n166_), .Y(mai_mai_n302_));
  OAI210     m0280(.A0(mai_mai_n168_), .A1(mai_mai_n146_), .B0(mai_mai_n302_), .Y(mai_mai_n303_));
  NO3        m0281(.A(mai_mai_n303_), .B(mai_mai_n298_), .C(mai_mai_n293_), .Y(mai_mai_n304_));
  NO2        m0282(.A(i_3_), .B(i_10_), .Y(mai_mai_n305_));
  NA3        m0283(.A(mai_mai_n305_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n306_));
  NO2        m0284(.A(i_2_), .B(mai_mai_n103_), .Y(mai_mai_n307_));
  NA2        m0285(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n308_));
  NO2        m0286(.A(mai_mai_n308_), .B(i_8_), .Y(mai_mai_n309_));
  NA2        m0287(.A(mai_mai_n309_), .B(mai_mai_n307_), .Y(mai_mai_n310_));
  AN2        m0288(.A(i_3_), .B(i_10_), .Y(mai_mai_n311_));
  NA4        m0289(.A(mai_mai_n311_), .B(mai_mai_n203_), .C(mai_mai_n180_), .D(mai_mai_n178_), .Y(mai_mai_n312_));
  NO2        m0290(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n313_));
  NO2        m0291(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n314_));
  OR2        m0292(.A(mai_mai_n310_), .B(mai_mai_n306_), .Y(mai_mai_n315_));
  OAI220     m0293(.A0(mai_mai_n315_), .A1(i_6_), .B0(mai_mai_n304_), .B1(mai_mai_n288_), .Y(mai_mai_n316_));
  NO4        m0294(.A(mai_mai_n316_), .B(mai_mai_n286_), .C(mai_mai_n219_), .D(mai_mai_n171_), .Y(mai_mai_n317_));
  NO3        m0295(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n318_));
  NO2        m0296(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n319_));
  NA2        m0297(.A(mai_mai_n295_), .B(mai_mai_n319_), .Y(mai_mai_n320_));
  NO3        m0298(.A(i_6_), .B(mai_mai_n198_), .C(i_7_), .Y(mai_mai_n321_));
  NA2        m0299(.A(mai_mai_n321_), .B(mai_mai_n203_), .Y(mai_mai_n322_));
  AOI210     m0300(.A0(mai_mai_n322_), .A1(mai_mai_n320_), .B0(mai_mai_n173_), .Y(mai_mai_n323_));
  NO2        m0301(.A(i_2_), .B(i_3_), .Y(mai_mai_n324_));
  OR2        m0302(.A(i_0_), .B(i_5_), .Y(mai_mai_n325_));
  NA2        m0303(.A(mai_mai_n222_), .B(mai_mai_n325_), .Y(mai_mai_n326_));
  NA4        m0304(.A(mai_mai_n326_), .B(mai_mai_n236_), .C(mai_mai_n324_), .D(i_1_), .Y(mai_mai_n327_));
  NA3        m0305(.A(mai_mai_n295_), .B(mai_mai_n290_), .C(mai_mai_n115_), .Y(mai_mai_n328_));
  NAi21      m0306(.An(i_8_), .B(i_7_), .Y(mai_mai_n329_));
  NO2        m0307(.A(mai_mai_n329_), .B(i_6_), .Y(mai_mai_n330_));
  NO2        m0308(.A(mai_mai_n160_), .B(mai_mai_n47_), .Y(mai_mai_n331_));
  NA3        m0309(.A(mai_mai_n331_), .B(mai_mai_n330_), .C(mai_mai_n166_), .Y(mai_mai_n332_));
  NA3        m0310(.A(mai_mai_n332_), .B(mai_mai_n328_), .C(mai_mai_n327_), .Y(mai_mai_n333_));
  OAI210     m0311(.A0(mai_mai_n333_), .A1(mai_mai_n323_), .B0(i_4_), .Y(mai_mai_n334_));
  NO2        m0312(.A(i_12_), .B(i_10_), .Y(mai_mai_n335_));
  NOi21      m0313(.An(i_5_), .B(i_0_), .Y(mai_mai_n336_));
  AOI210     m0314(.A0(i_2_), .A1(mai_mai_n49_), .B0(mai_mai_n103_), .Y(mai_mai_n337_));
  NO4        m0315(.A(mai_mai_n337_), .B(mai_mai_n308_), .C(mai_mai_n336_), .D(mai_mai_n131_), .Y(mai_mai_n338_));
  NA2        m0316(.A(mai_mai_n338_), .B(mai_mai_n335_), .Y(mai_mai_n339_));
  NO2        m0317(.A(i_6_), .B(i_8_), .Y(mai_mai_n340_));
  NOi21      m0318(.An(i_0_), .B(i_2_), .Y(mai_mai_n341_));
  AN2        m0319(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n342_));
  NO2        m0320(.A(i_1_), .B(i_7_), .Y(mai_mai_n343_));
  AO220      m0321(.A0(mai_mai_n343_), .A1(mai_mai_n342_), .B0(mai_mai_n330_), .B1(mai_mai_n237_), .Y(mai_mai_n344_));
  NA3        m0322(.A(mai_mai_n344_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n345_));
  NA3        m0323(.A(mai_mai_n345_), .B(mai_mai_n339_), .C(mai_mai_n334_), .Y(mai_mai_n346_));
  NO3        m0324(.A(mai_mai_n235_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n347_));
  NO3        m0325(.A(mai_mai_n329_), .B(i_2_), .C(i_1_), .Y(mai_mai_n348_));
  OAI210     m0326(.A0(mai_mai_n348_), .A1(mai_mai_n347_), .B0(i_6_), .Y(mai_mai_n349_));
  NA3        m0327(.A(mai_mai_n255_), .B(mai_mai_n307_), .C(mai_mai_n198_), .Y(mai_mai_n350_));
  AOI210     m0328(.A0(mai_mai_n350_), .A1(mai_mai_n349_), .B0(mai_mai_n326_), .Y(mai_mai_n351_));
  NOi21      m0329(.An(mai_mai_n156_), .B(mai_mai_n106_), .Y(mai_mai_n352_));
  NO2        m0330(.A(mai_mai_n352_), .B(mai_mai_n127_), .Y(mai_mai_n353_));
  OAI210     m0331(.A0(mai_mai_n353_), .A1(mai_mai_n351_), .B0(i_3_), .Y(mai_mai_n354_));
  INV        m0332(.A(mai_mai_n85_), .Y(mai_mai_n355_));
  NO2        m0333(.A(mai_mai_n299_), .B(mai_mai_n82_), .Y(mai_mai_n356_));
  NA2        m0334(.A(mai_mai_n356_), .B(mai_mai_n135_), .Y(mai_mai_n357_));
  NO2        m0335(.A(mai_mai_n94_), .B(mai_mai_n198_), .Y(mai_mai_n358_));
  NA2        m0336(.A(mai_mai_n358_), .B(mai_mai_n64_), .Y(mai_mai_n359_));
  AOI210     m0337(.A0(mai_mai_n359_), .A1(mai_mai_n357_), .B0(mai_mai_n355_), .Y(mai_mai_n360_));
  NO2        m0338(.A(mai_mai_n198_), .B(i_9_), .Y(mai_mai_n361_));
  NA2        m0339(.A(mai_mai_n361_), .B(mai_mai_n210_), .Y(mai_mai_n362_));
  NO2        m0340(.A(mai_mai_n362_), .B(mai_mai_n47_), .Y(mai_mai_n363_));
  NO3        m0341(.A(mai_mai_n363_), .B(mai_mai_n360_), .C(mai_mai_n298_), .Y(mai_mai_n364_));
  AOI210     m0342(.A0(mai_mai_n364_), .A1(mai_mai_n354_), .B0(mai_mai_n165_), .Y(mai_mai_n365_));
  AOI210     m0343(.A0(mai_mai_n346_), .A1(mai_mai_n318_), .B0(mai_mai_n365_), .Y(mai_mai_n366_));
  NOi32      m0344(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n367_));
  INV        m0345(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  NAi21      m0346(.An(i_0_), .B(i_6_), .Y(mai_mai_n369_));
  NAi21      m0347(.An(i_1_), .B(i_5_), .Y(mai_mai_n370_));
  NA2        m0348(.A(mai_mai_n370_), .B(mai_mai_n369_), .Y(mai_mai_n371_));
  NAi41      m0349(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n372_));
  OAI220     m0350(.A0(mai_mai_n372_), .A1(mai_mai_n370_), .B0(mai_mai_n223_), .B1(mai_mai_n162_), .Y(mai_mai_n373_));
  AOI210     m0351(.A0(mai_mai_n372_), .A1(mai_mai_n162_), .B0(mai_mai_n160_), .Y(mai_mai_n374_));
  NOi32      m0352(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n375_));
  NAi21      m0353(.An(i_6_), .B(i_1_), .Y(mai_mai_n376_));
  NA3        m0354(.A(mai_mai_n376_), .B(mai_mai_n375_), .C(mai_mai_n47_), .Y(mai_mai_n377_));
  NO2        m0355(.A(mai_mai_n377_), .B(i_0_), .Y(mai_mai_n378_));
  OR3        m0356(.A(mai_mai_n378_), .B(mai_mai_n374_), .C(mai_mai_n373_), .Y(mai_mai_n379_));
  NO2        m0357(.A(i_1_), .B(mai_mai_n103_), .Y(mai_mai_n380_));
  NAi21      m0358(.An(i_3_), .B(i_4_), .Y(mai_mai_n381_));
  NO2        m0359(.A(mai_mai_n381_), .B(i_9_), .Y(mai_mai_n382_));
  AN2        m0360(.A(i_6_), .B(i_7_), .Y(mai_mai_n383_));
  OAI210     m0361(.A0(mai_mai_n383_), .A1(mai_mai_n380_), .B0(mai_mai_n382_), .Y(mai_mai_n384_));
  NA2        m0362(.A(i_2_), .B(i_7_), .Y(mai_mai_n385_));
  NO2        m0363(.A(mai_mai_n381_), .B(i_10_), .Y(mai_mai_n386_));
  NA3        m0364(.A(mai_mai_n386_), .B(mai_mai_n385_), .C(mai_mai_n247_), .Y(mai_mai_n387_));
  AOI210     m0365(.A0(mai_mai_n387_), .A1(mai_mai_n384_), .B0(mai_mai_n190_), .Y(mai_mai_n388_));
  AOI210     m0366(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n389_));
  OAI210     m0367(.A0(mai_mai_n389_), .A1(mai_mai_n193_), .B0(mai_mai_n386_), .Y(mai_mai_n390_));
  AOI220     m0368(.A0(mai_mai_n386_), .A1(mai_mai_n343_), .B0(mai_mai_n241_), .B1(mai_mai_n193_), .Y(mai_mai_n391_));
  AOI210     m0369(.A0(mai_mai_n391_), .A1(mai_mai_n390_), .B0(i_5_), .Y(mai_mai_n392_));
  NO4        m0370(.A(mai_mai_n392_), .B(mai_mai_n388_), .C(mai_mai_n379_), .D(mai_mai_n1079_), .Y(mai_mai_n393_));
  NO2        m0371(.A(mai_mai_n393_), .B(mai_mai_n368_), .Y(mai_mai_n394_));
  NO2        m0372(.A(mai_mai_n60_), .B(mai_mai_n25_), .Y(mai_mai_n395_));
  AN2        m0373(.A(i_12_), .B(i_5_), .Y(mai_mai_n396_));
  NO2        m0374(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n397_));
  NA2        m0375(.A(mai_mai_n397_), .B(mai_mai_n396_), .Y(mai_mai_n398_));
  NO2        m0376(.A(i_11_), .B(i_6_), .Y(mai_mai_n399_));
  NA3        m0377(.A(mai_mai_n399_), .B(mai_mai_n331_), .C(mai_mai_n228_), .Y(mai_mai_n400_));
  NO2        m0378(.A(mai_mai_n400_), .B(mai_mai_n398_), .Y(mai_mai_n401_));
  NO2        m0379(.A(mai_mai_n245_), .B(i_5_), .Y(mai_mai_n402_));
  NO2        m0380(.A(i_5_), .B(i_10_), .Y(mai_mai_n403_));
  AOI220     m0381(.A0(mai_mai_n403_), .A1(mai_mai_n275_), .B0(mai_mai_n402_), .B1(mai_mai_n203_), .Y(mai_mai_n404_));
  NA2        m0382(.A(mai_mai_n147_), .B(mai_mai_n46_), .Y(mai_mai_n405_));
  NO2        m0383(.A(mai_mai_n405_), .B(mai_mai_n404_), .Y(mai_mai_n406_));
  OAI210     m0384(.A0(mai_mai_n406_), .A1(mai_mai_n401_), .B0(mai_mai_n395_), .Y(mai_mai_n407_));
  NO2        m0385(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n408_));
  NO3        m0386(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n409_));
  NO2        m0387(.A(i_3_), .B(mai_mai_n103_), .Y(mai_mai_n410_));
  NA4        m0388(.A(mai_mai_n305_), .B(mai_mai_n92_), .C(mai_mai_n76_), .D(mai_mai_n55_), .Y(mai_mai_n411_));
  NO2        m0389(.A(i_11_), .B(i_12_), .Y(mai_mai_n412_));
  NA2        m0390(.A(mai_mai_n412_), .B(mai_mai_n36_), .Y(mai_mai_n413_));
  NO2        m0391(.A(mai_mai_n411_), .B(mai_mai_n413_), .Y(mai_mai_n414_));
  NA2        m0392(.A(mai_mai_n403_), .B(mai_mai_n239_), .Y(mai_mai_n415_));
  NA3        m0393(.A(mai_mai_n115_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n416_));
  NO2        m0394(.A(mai_mai_n416_), .B(mai_mai_n223_), .Y(mai_mai_n417_));
  NAi21      m0395(.An(i_13_), .B(i_0_), .Y(mai_mai_n418_));
  NO2        m0396(.A(mai_mai_n418_), .B(mai_mai_n242_), .Y(mai_mai_n419_));
  OAI210     m0397(.A0(mai_mai_n417_), .A1(mai_mai_n414_), .B0(mai_mai_n419_), .Y(mai_mai_n420_));
  NA2        m0398(.A(mai_mai_n420_), .B(mai_mai_n407_), .Y(mai_mai_n421_));
  NO3        m0399(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n422_));
  NO2        m0400(.A(i_0_), .B(i_11_), .Y(mai_mai_n423_));
  INV        m0401(.A(i_5_), .Y(mai_mai_n424_));
  AN2        m0402(.A(i_1_), .B(i_6_), .Y(mai_mai_n425_));
  NOi21      m0403(.An(i_2_), .B(i_12_), .Y(mai_mai_n426_));
  NA2        m0404(.A(mai_mai_n426_), .B(mai_mai_n425_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n427_), .B(mai_mai_n424_), .Y(mai_mai_n428_));
  NA2        m0406(.A(mai_mai_n145_), .B(i_9_), .Y(mai_mai_n429_));
  NO2        m0407(.A(mai_mai_n429_), .B(i_4_), .Y(mai_mai_n430_));
  NA2        m0408(.A(mai_mai_n428_), .B(mai_mai_n430_), .Y(mai_mai_n431_));
  NAi21      m0409(.An(i_9_), .B(i_4_), .Y(mai_mai_n432_));
  OR2        m0410(.A(i_13_), .B(i_10_), .Y(mai_mai_n433_));
  NO3        m0411(.A(mai_mai_n433_), .B(mai_mai_n120_), .C(mai_mai_n432_), .Y(mai_mai_n434_));
  NO2        m0412(.A(mai_mai_n176_), .B(mai_mai_n126_), .Y(mai_mai_n435_));
  OR2        m0413(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n436_));
  NO2        m0414(.A(mai_mai_n103_), .B(mai_mai_n25_), .Y(mai_mai_n437_));
  NA2        m0415(.A(mai_mai_n287_), .B(mai_mai_n437_), .Y(mai_mai_n438_));
  NA2        m0416(.A(mai_mai_n280_), .B(mai_mai_n215_), .Y(mai_mai_n439_));
  OAI220     m0417(.A0(mai_mai_n439_), .A1(mai_mai_n436_), .B0(mai_mai_n438_), .B1(mai_mai_n352_), .Y(mai_mai_n440_));
  INV        m0418(.A(mai_mai_n440_), .Y(mai_mai_n441_));
  AOI210     m0419(.A0(mai_mai_n441_), .A1(mai_mai_n431_), .B0(mai_mai_n26_), .Y(mai_mai_n442_));
  NA2        m0420(.A(mai_mai_n328_), .B(mai_mai_n327_), .Y(mai_mai_n443_));
  AOI220     m0421(.A0(mai_mai_n301_), .A1(mai_mai_n291_), .B0(mai_mai_n295_), .B1(mai_mai_n319_), .Y(mai_mai_n444_));
  NO2        m0422(.A(mai_mai_n444_), .B(mai_mai_n173_), .Y(mai_mai_n445_));
  NO2        m0423(.A(mai_mai_n187_), .B(mai_mai_n87_), .Y(mai_mai_n446_));
  AOI220     m0424(.A0(mai_mai_n446_), .A1(mai_mai_n300_), .B0(mai_mai_n282_), .B1(mai_mai_n215_), .Y(mai_mai_n447_));
  NO2        m0425(.A(mai_mai_n447_), .B(mai_mai_n289_), .Y(mai_mai_n448_));
  NO3        m0426(.A(mai_mai_n448_), .B(mai_mai_n445_), .C(mai_mai_n443_), .Y(mai_mai_n449_));
  NA2        m0427(.A(mai_mai_n201_), .B(mai_mai_n98_), .Y(mai_mai_n450_));
  NA3        m0428(.A(mai_mai_n331_), .B(mai_mai_n166_), .C(mai_mai_n87_), .Y(mai_mai_n451_));
  AOI210     m0429(.A0(mai_mai_n451_), .A1(mai_mai_n450_), .B0(mai_mai_n329_), .Y(mai_mai_n452_));
  NA2        m0430(.A(mai_mai_n198_), .B(i_10_), .Y(mai_mai_n453_));
  NA3        m0431(.A(mai_mai_n261_), .B(mai_mai_n65_), .C(i_2_), .Y(mai_mai_n454_));
  NA2        m0432(.A(mai_mai_n301_), .B(mai_mai_n237_), .Y(mai_mai_n455_));
  OAI220     m0433(.A0(mai_mai_n455_), .A1(mai_mai_n187_), .B0(mai_mai_n454_), .B1(mai_mai_n453_), .Y(mai_mai_n456_));
  NO2        m0434(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n457_));
  NA3        m0435(.A(mai_mai_n343_), .B(mai_mai_n342_), .C(mai_mai_n457_), .Y(mai_mai_n458_));
  NA2        m0436(.A(mai_mai_n321_), .B(mai_mai_n326_), .Y(mai_mai_n459_));
  OAI210     m0437(.A0(mai_mai_n459_), .A1(mai_mai_n194_), .B0(mai_mai_n458_), .Y(mai_mai_n460_));
  NO3        m0438(.A(mai_mai_n460_), .B(mai_mai_n456_), .C(mai_mai_n452_), .Y(mai_mai_n461_));
  AOI210     m0439(.A0(mai_mai_n461_), .A1(mai_mai_n449_), .B0(mai_mai_n276_), .Y(mai_mai_n462_));
  NO4        m0440(.A(mai_mai_n462_), .B(mai_mai_n442_), .C(mai_mai_n421_), .D(mai_mai_n394_), .Y(mai_mai_n463_));
  NO2        m0441(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n464_));
  NO2        m0442(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n465_));
  NO2        m0443(.A(i_10_), .B(i_9_), .Y(mai_mai_n466_));
  NAi21      m0444(.An(i_12_), .B(i_8_), .Y(mai_mai_n467_));
  NO2        m0445(.A(mai_mai_n467_), .B(i_3_), .Y(mai_mai_n468_));
  NA2        m0446(.A(mai_mai_n314_), .B(i_0_), .Y(mai_mai_n469_));
  NO3        m0447(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n470_));
  NA2        m0448(.A(mai_mai_n273_), .B(mai_mai_n99_), .Y(mai_mai_n471_));
  NA2        m0449(.A(mai_mai_n471_), .B(mai_mai_n470_), .Y(mai_mai_n472_));
  NA2        m0450(.A(i_8_), .B(i_9_), .Y(mai_mai_n473_));
  AOI210     m0451(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n474_));
  OR2        m0452(.A(mai_mai_n474_), .B(mai_mai_n473_), .Y(mai_mai_n475_));
  NA2        m0453(.A(mai_mai_n287_), .B(mai_mai_n210_), .Y(mai_mai_n476_));
  NO2        m0454(.A(mai_mai_n476_), .B(mai_mai_n475_), .Y(mai_mai_n477_));
  NA2        m0455(.A(mai_mai_n254_), .B(mai_mai_n313_), .Y(mai_mai_n478_));
  NO3        m0456(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n479_));
  INV        m0457(.A(mai_mai_n479_), .Y(mai_mai_n480_));
  NA3        m0458(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n481_));
  NA4        m0459(.A(mai_mai_n148_), .B(mai_mai_n118_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n482_));
  OAI220     m0460(.A0(mai_mai_n482_), .A1(mai_mai_n481_), .B0(mai_mai_n480_), .B1(mai_mai_n478_), .Y(mai_mai_n483_));
  NO2        m0461(.A(mai_mai_n483_), .B(mai_mai_n477_), .Y(mai_mai_n484_));
  NA2        m0462(.A(mai_mai_n300_), .B(mai_mai_n110_), .Y(mai_mai_n485_));
  OR2        m0463(.A(mai_mai_n485_), .B(mai_mai_n212_), .Y(mai_mai_n486_));
  BUFFER     m0464(.A(mai_mai_n302_), .Y(mai_mai_n487_));
  OA220      m0465(.A0(mai_mai_n487_), .A1(mai_mai_n165_), .B0(mai_mai_n486_), .B1(mai_mai_n234_), .Y(mai_mai_n488_));
  NA2        m0466(.A(mai_mai_n98_), .B(i_13_), .Y(mai_mai_n489_));
  NO2        m0467(.A(i_2_), .B(i_13_), .Y(mai_mai_n490_));
  NO3        m0468(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n491_));
  NO2        m0469(.A(i_6_), .B(i_7_), .Y(mai_mai_n492_));
  NA2        m0470(.A(mai_mai_n492_), .B(mai_mai_n491_), .Y(mai_mai_n493_));
  NO2        m0471(.A(i_11_), .B(i_1_), .Y(mai_mai_n494_));
  NO2        m0472(.A(mai_mai_n74_), .B(i_3_), .Y(mai_mai_n495_));
  OR2        m0473(.A(i_11_), .B(i_8_), .Y(mai_mai_n496_));
  NOi21      m0474(.An(i_2_), .B(i_7_), .Y(mai_mai_n497_));
  NAi31      m0475(.An(mai_mai_n496_), .B(mai_mai_n497_), .C(mai_mai_n495_), .Y(mai_mai_n498_));
  NO2        m0476(.A(mai_mai_n433_), .B(i_6_), .Y(mai_mai_n499_));
  NA3        m0477(.A(mai_mai_n499_), .B(mai_mai_n464_), .C(mai_mai_n76_), .Y(mai_mai_n500_));
  NO2        m0478(.A(mai_mai_n500_), .B(mai_mai_n498_), .Y(mai_mai_n501_));
  NO2        m0479(.A(i_3_), .B(mai_mai_n198_), .Y(mai_mai_n502_));
  NO2        m0480(.A(i_6_), .B(i_10_), .Y(mai_mai_n503_));
  NA4        m0481(.A(mai_mai_n503_), .B(mai_mai_n318_), .C(mai_mai_n502_), .D(mai_mai_n239_), .Y(mai_mai_n504_));
  NO2        m0482(.A(mai_mai_n504_), .B(mai_mai_n158_), .Y(mai_mai_n505_));
  NA3        m0483(.A(mai_mai_n248_), .B(mai_mai_n175_), .C(mai_mai_n135_), .Y(mai_mai_n506_));
  NA2        m0484(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n507_));
  NO2        m0485(.A(mai_mai_n160_), .B(i_3_), .Y(mai_mai_n508_));
  NAi31      m0486(.An(mai_mai_n507_), .B(mai_mai_n508_), .C(mai_mai_n229_), .Y(mai_mai_n509_));
  NA3        m0487(.A(mai_mai_n408_), .B(mai_mai_n183_), .C(mai_mai_n152_), .Y(mai_mai_n510_));
  NA3        m0488(.A(mai_mai_n510_), .B(mai_mai_n509_), .C(mai_mai_n506_), .Y(mai_mai_n511_));
  NO3        m0489(.A(mai_mai_n511_), .B(mai_mai_n505_), .C(mai_mai_n501_), .Y(mai_mai_n512_));
  NA2        m0490(.A(mai_mai_n470_), .B(mai_mai_n396_), .Y(mai_mai_n513_));
  NA2        m0491(.A(mai_mai_n479_), .B(mai_mai_n403_), .Y(mai_mai_n514_));
  NO2        m0492(.A(mai_mai_n514_), .B(mai_mai_n227_), .Y(mai_mai_n515_));
  NAi21      m0493(.An(mai_mai_n221_), .B(mai_mai_n412_), .Y(mai_mai_n516_));
  NO2        m0494(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n517_));
  NO2        m0495(.A(i_0_), .B(mai_mai_n87_), .Y(mai_mai_n518_));
  NA3        m0496(.A(mai_mai_n518_), .B(mai_mai_n517_), .C(mai_mai_n145_), .Y(mai_mai_n519_));
  OR3        m0497(.A(mai_mai_n308_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n520_));
  NO2        m0498(.A(mai_mai_n520_), .B(mai_mai_n519_), .Y(mai_mai_n521_));
  NA2        m0499(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n522_));
  NA2        m0500(.A(mai_mai_n318_), .B(mai_mai_n241_), .Y(mai_mai_n523_));
  OAI220     m0501(.A0(mai_mai_n523_), .A1(mai_mai_n454_), .B0(mai_mai_n522_), .B1(mai_mai_n489_), .Y(mai_mai_n524_));
  NA4        m0502(.A(mai_mai_n311_), .B(mai_mai_n226_), .C(mai_mai_n74_), .D(mai_mai_n239_), .Y(mai_mai_n525_));
  NO2        m0503(.A(mai_mai_n525_), .B(mai_mai_n493_), .Y(mai_mai_n526_));
  NO4        m0504(.A(mai_mai_n526_), .B(mai_mai_n524_), .C(mai_mai_n521_), .D(mai_mai_n515_), .Y(mai_mai_n527_));
  NA4        m0505(.A(mai_mai_n527_), .B(mai_mai_n512_), .C(mai_mai_n488_), .D(mai_mai_n484_), .Y(mai_mai_n528_));
  NA3        m0506(.A(mai_mai_n311_), .B(mai_mai_n180_), .C(mai_mai_n178_), .Y(mai_mai_n529_));
  OAI210     m0507(.A0(mai_mai_n306_), .A1(mai_mai_n185_), .B0(mai_mai_n529_), .Y(mai_mai_n530_));
  AN2        m0508(.A(mai_mai_n291_), .B(mai_mai_n236_), .Y(mai_mai_n531_));
  NA2        m0509(.A(mai_mai_n531_), .B(mai_mai_n530_), .Y(mai_mai_n532_));
  NA2        m0510(.A(mai_mai_n318_), .B(mai_mai_n167_), .Y(mai_mai_n533_));
  OAI210     m0511(.A0(mai_mai_n533_), .A1(mai_mai_n234_), .B0(mai_mai_n312_), .Y(mai_mai_n534_));
  NA2        m0512(.A(mai_mai_n534_), .B(mai_mai_n330_), .Y(mai_mai_n535_));
  NA2        m0513(.A(mai_mai_n396_), .B(mai_mai_n228_), .Y(mai_mai_n536_));
  NA2        m0514(.A(mai_mai_n367_), .B(mai_mai_n74_), .Y(mai_mai_n537_));
  NA2        m0515(.A(mai_mai_n383_), .B(mai_mai_n375_), .Y(mai_mai_n538_));
  OR2        m0516(.A(mai_mai_n536_), .B(mai_mai_n538_), .Y(mai_mai_n539_));
  NO2        m0517(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n540_));
  NAi41      m0518(.An(mai_mai_n537_), .B(mai_mai_n503_), .C(mai_mai_n540_), .D(mai_mai_n47_), .Y(mai_mai_n541_));
  AOI210     m0519(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n434_), .Y(mai_mai_n542_));
  NA3        m0520(.A(mai_mai_n542_), .B(mai_mai_n541_), .C(mai_mai_n539_), .Y(mai_mai_n543_));
  INV        m0521(.A(mai_mai_n543_), .Y(mai_mai_n544_));
  INV        m0522(.A(mai_mai_n137_), .Y(mai_mai_n545_));
  AOI210     m0523(.A0(mai_mai_n199_), .A1(i_9_), .B0(mai_mai_n272_), .Y(mai_mai_n546_));
  NO2        m0524(.A(mai_mai_n546_), .B(mai_mai_n204_), .Y(mai_mai_n547_));
  OR2        m0525(.A(mai_mai_n187_), .B(i_4_), .Y(mai_mai_n548_));
  NO2        m0526(.A(mai_mai_n548_), .B(mai_mai_n87_), .Y(mai_mai_n549_));
  AOI220     m0527(.A0(mai_mai_n549_), .A1(mai_mai_n547_), .B0(mai_mai_n545_), .B1(mai_mai_n435_), .Y(mai_mai_n550_));
  NA4        m0528(.A(mai_mai_n550_), .B(mai_mai_n544_), .C(mai_mai_n535_), .D(mai_mai_n532_), .Y(mai_mai_n551_));
  NA2        m0529(.A(mai_mai_n402_), .B(mai_mai_n300_), .Y(mai_mai_n552_));
  OAI210     m0530(.A0(mai_mai_n398_), .A1(mai_mai_n172_), .B0(mai_mai_n552_), .Y(mai_mai_n553_));
  NO2        m0531(.A(i_12_), .B(mai_mai_n198_), .Y(mai_mai_n554_));
  NA2        m0532(.A(mai_mai_n554_), .B(mai_mai_n228_), .Y(mai_mai_n555_));
  NA3        m0533(.A(mai_mai_n503_), .B(mai_mai_n178_), .C(mai_mai_n27_), .Y(mai_mai_n556_));
  NO2        m0534(.A(mai_mai_n556_), .B(mai_mai_n555_), .Y(mai_mai_n557_));
  NOi31      m0535(.An(mai_mai_n321_), .B(mai_mai_n433_), .C(mai_mai_n38_), .Y(mai_mai_n558_));
  OAI210     m0536(.A0(mai_mai_n558_), .A1(mai_mai_n557_), .B0(mai_mai_n553_), .Y(mai_mai_n559_));
  NO2        m0537(.A(i_8_), .B(i_7_), .Y(mai_mai_n560_));
  OAI210     m0538(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n561_));
  NA2        m0539(.A(mai_mai_n561_), .B(mai_mai_n226_), .Y(mai_mai_n562_));
  AOI220     m0540(.A0(mai_mai_n331_), .A1(mai_mai_n40_), .B0(mai_mai_n237_), .B1(mai_mai_n211_), .Y(mai_mai_n563_));
  OAI220     m0541(.A0(mai_mai_n563_), .A1(mai_mai_n548_), .B0(mai_mai_n562_), .B1(mai_mai_n245_), .Y(mai_mai_n564_));
  NA2        m0542(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n565_));
  NO2        m0543(.A(mai_mai_n565_), .B(i_6_), .Y(mai_mai_n566_));
  NA3        m0544(.A(mai_mai_n566_), .B(mai_mai_n564_), .C(mai_mai_n560_), .Y(mai_mai_n567_));
  NOi31      m0545(.An(mai_mai_n295_), .B(mai_mai_n306_), .C(mai_mai_n185_), .Y(mai_mai_n568_));
  NO2        m0546(.A(mai_mai_n160_), .B(i_5_), .Y(mai_mai_n569_));
  NA2        m0547(.A(mai_mai_n568_), .B(mai_mai_n479_), .Y(mai_mai_n570_));
  NA3        m0548(.A(mai_mai_n570_), .B(mai_mai_n567_), .C(mai_mai_n559_), .Y(mai_mai_n571_));
  NA3        m0549(.A(mai_mai_n222_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n572_));
  NA2        m0550(.A(mai_mai_n287_), .B(mai_mai_n85_), .Y(mai_mai_n573_));
  AOI210     m0551(.A0(mai_mai_n572_), .A1(mai_mai_n357_), .B0(mai_mai_n573_), .Y(mai_mai_n574_));
  NA2        m0552(.A(mai_mai_n301_), .B(mai_mai_n291_), .Y(mai_mai_n575_));
  NO2        m0553(.A(mai_mai_n575_), .B(mai_mai_n177_), .Y(mai_mai_n576_));
  NA2        m0554(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n577_));
  NA2        m0555(.A(mai_mai_n466_), .B(mai_mai_n224_), .Y(mai_mai_n578_));
  NO2        m0556(.A(mai_mai_n577_), .B(mai_mai_n578_), .Y(mai_mai_n579_));
  AOI210     m0557(.A0(mai_mai_n376_), .A1(mai_mai_n47_), .B0(mai_mai_n380_), .Y(mai_mai_n580_));
  NA2        m0558(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n581_));
  NA3        m0559(.A(mai_mai_n554_), .B(mai_mai_n278_), .C(mai_mai_n581_), .Y(mai_mai_n582_));
  NO2        m0560(.A(mai_mai_n580_), .B(mai_mai_n582_), .Y(mai_mai_n583_));
  NO4        m0561(.A(mai_mai_n583_), .B(mai_mai_n579_), .C(mai_mai_n576_), .D(mai_mai_n574_), .Y(mai_mai_n584_));
  NO4        m0562(.A(mai_mai_n255_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n585_));
  NO3        m0563(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n586_));
  NO2        m0564(.A(mai_mai_n235_), .B(mai_mai_n36_), .Y(mai_mai_n587_));
  AN2        m0565(.A(mai_mai_n587_), .B(mai_mai_n586_), .Y(mai_mai_n588_));
  OA210      m0566(.A0(mai_mai_n588_), .A1(mai_mai_n585_), .B0(mai_mai_n367_), .Y(mai_mai_n589_));
  NO2        m0567(.A(mai_mai_n433_), .B(i_1_), .Y(mai_mai_n590_));
  NOi31      m0568(.An(mai_mai_n590_), .B(mai_mai_n471_), .C(mai_mai_n74_), .Y(mai_mai_n591_));
  AN4        m0569(.A(mai_mai_n591_), .B(mai_mai_n430_), .C(mai_mai_n517_), .D(i_2_), .Y(mai_mai_n592_));
  NO2        m0570(.A(mai_mai_n444_), .B(mai_mai_n181_), .Y(mai_mai_n593_));
  NO3        m0571(.A(mai_mai_n593_), .B(mai_mai_n592_), .C(mai_mai_n589_), .Y(mai_mai_n594_));
  NOi21      m0572(.An(i_10_), .B(i_6_), .Y(mai_mai_n595_));
  NO2        m0573(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n596_));
  NO2        m0574(.A(mai_mai_n117_), .B(mai_mai_n23_), .Y(mai_mai_n597_));
  NA2        m0575(.A(mai_mai_n321_), .B(mai_mai_n167_), .Y(mai_mai_n598_));
  AOI220     m0576(.A0(mai_mai_n598_), .A1(mai_mai_n455_), .B0(mai_mai_n188_), .B1(mai_mai_n186_), .Y(mai_mai_n599_));
  INV        m0577(.A(mai_mai_n599_), .Y(mai_mai_n600_));
  NO2        m0578(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n601_));
  NA2        m0579(.A(mai_mai_n178_), .B(i_0_), .Y(mai_mai_n602_));
  NO3        m0580(.A(mai_mai_n602_), .B(mai_mai_n349_), .C(mai_mai_n306_), .Y(mai_mai_n603_));
  OR2        m0581(.A(i_2_), .B(i_5_), .Y(mai_mai_n604_));
  OR2        m0582(.A(mai_mai_n604_), .B(mai_mai_n425_), .Y(mai_mai_n605_));
  AOI210     m0583(.A0(mai_mai_n385_), .A1(mai_mai_n247_), .B0(mai_mai_n203_), .Y(mai_mai_n606_));
  AOI210     m0584(.A0(mai_mai_n606_), .A1(mai_mai_n605_), .B0(mai_mai_n516_), .Y(mai_mai_n607_));
  NO2        m0585(.A(mai_mai_n607_), .B(mai_mai_n603_), .Y(mai_mai_n608_));
  NA4        m0586(.A(mai_mai_n608_), .B(mai_mai_n600_), .C(mai_mai_n594_), .D(mai_mai_n584_), .Y(mai_mai_n609_));
  NO4        m0587(.A(mai_mai_n609_), .B(mai_mai_n571_), .C(mai_mai_n551_), .D(mai_mai_n528_), .Y(mai_mai_n610_));
  NA4        m0588(.A(mai_mai_n610_), .B(mai_mai_n463_), .C(mai_mai_n366_), .D(mai_mai_n317_), .Y(mai7));
  NO2        m0589(.A(mai_mai_n94_), .B(mai_mai_n55_), .Y(mai_mai_n612_));
  NA2        m0590(.A(mai_mai_n503_), .B(mai_mai_n85_), .Y(mai_mai_n613_));
  NA2        m0591(.A(i_11_), .B(mai_mai_n198_), .Y(mai_mai_n614_));
  NA2        m0592(.A(mai_mai_n147_), .B(mai_mai_n614_), .Y(mai_mai_n615_));
  NO2        m0593(.A(mai_mai_n615_), .B(mai_mai_n613_), .Y(mai_mai_n616_));
  NA3        m0594(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n617_));
  NO2        m0595(.A(mai_mai_n239_), .B(i_4_), .Y(mai_mai_n618_));
  NA2        m0596(.A(mai_mai_n618_), .B(i_8_), .Y(mai_mai_n619_));
  NO2        m0597(.A(mai_mai_n107_), .B(mai_mai_n617_), .Y(mai_mai_n620_));
  NA2        m0598(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n621_));
  OAI210     m0599(.A0(mai_mai_n88_), .A1(mai_mai_n208_), .B0(mai_mai_n209_), .Y(mai_mai_n622_));
  NO2        m0600(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n623_));
  NA2        m0601(.A(i_4_), .B(i_8_), .Y(mai_mai_n624_));
  AOI210     m0602(.A0(mai_mai_n624_), .A1(mai_mai_n311_), .B0(mai_mai_n623_), .Y(mai_mai_n625_));
  OAI220     m0603(.A0(mai_mai_n625_), .A1(mai_mai_n621_), .B0(mai_mai_n622_), .B1(i_13_), .Y(mai_mai_n626_));
  NO4        m0604(.A(mai_mai_n626_), .B(mai_mai_n620_), .C(mai_mai_n616_), .D(mai_mai_n612_), .Y(mai_mai_n627_));
  AOI210     m0605(.A0(mai_mai_n131_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n628_));
  AOI210     m0606(.A0(mai_mai_n628_), .A1(mai_mai_n239_), .B0(mai_mai_n164_), .Y(mai_mai_n629_));
  OR2        m0607(.A(i_6_), .B(i_10_), .Y(mai_mai_n630_));
  NO2        m0608(.A(mai_mai_n630_), .B(mai_mai_n23_), .Y(mai_mai_n631_));
  OR3        m0609(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n632_));
  NO3        m0610(.A(mai_mai_n632_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n633_));
  INV        m0611(.A(mai_mai_n205_), .Y(mai_mai_n634_));
  OR2        m0612(.A(mai_mai_n629_), .B(mai_mai_n274_), .Y(mai_mai_n635_));
  AOI210     m0613(.A0(mai_mai_n635_), .A1(mai_mai_n627_), .B0(mai_mai_n64_), .Y(mai_mai_n636_));
  NOi21      m0614(.An(i_11_), .B(i_7_), .Y(mai_mai_n637_));
  AO210      m0615(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n638_));
  NO2        m0616(.A(mai_mai_n638_), .B(mai_mai_n637_), .Y(mai_mai_n639_));
  NA2        m0617(.A(mai_mai_n639_), .B(mai_mai_n211_), .Y(mai_mai_n640_));
  NA3        m0618(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n641_));
  NO2        m0619(.A(mai_mai_n640_), .B(mai_mai_n64_), .Y(mai_mai_n642_));
  OR2        m0620(.A(mai_mai_n391_), .B(mai_mai_n41_), .Y(mai_mai_n643_));
  NO3        m0621(.A(mai_mai_n263_), .B(mai_mai_n213_), .C(mai_mai_n614_), .Y(mai_mai_n644_));
  OAI210     m0622(.A0(mai_mai_n644_), .A1(mai_mai_n229_), .B0(mai_mai_n64_), .Y(mai_mai_n645_));
  NA2        m0623(.A(mai_mai_n426_), .B(mai_mai_n31_), .Y(mai_mai_n646_));
  OR2        m0624(.A(mai_mai_n213_), .B(mai_mai_n110_), .Y(mai_mai_n647_));
  NA2        m0625(.A(mai_mai_n647_), .B(mai_mai_n646_), .Y(mai_mai_n648_));
  NO2        m0626(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n649_));
  NO2        m0627(.A(mai_mai_n649_), .B(i_4_), .Y(mai_mai_n650_));
  NA2        m0628(.A(mai_mai_n650_), .B(mai_mai_n648_), .Y(mai_mai_n651_));
  NO2        m0629(.A(i_1_), .B(i_12_), .Y(mai_mai_n652_));
  NA3        m0630(.A(mai_mai_n651_), .B(mai_mai_n645_), .C(mai_mai_n643_), .Y(mai_mai_n653_));
  OAI210     m0631(.A0(mai_mai_n653_), .A1(mai_mai_n642_), .B0(i_6_), .Y(mai_mai_n654_));
  NO2        m0632(.A(mai_mai_n641_), .B(mai_mai_n110_), .Y(mai_mai_n655_));
  NA2        m0633(.A(mai_mai_n655_), .B(mai_mai_n601_), .Y(mai_mai_n656_));
  NO2        m0634(.A(i_6_), .B(i_11_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n656_), .B(mai_mai_n472_), .Y(mai_mai_n658_));
  NO4        m0636(.A(mai_mai_n220_), .B(mai_mai_n131_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n659_));
  NA2        m0637(.A(mai_mai_n659_), .B(mai_mai_n649_), .Y(mai_mai_n660_));
  NA2        m0638(.A(mai_mai_n239_), .B(i_6_), .Y(mai_mai_n661_));
  NO3        m0639(.A(mai_mai_n630_), .B(mai_mai_n235_), .C(mai_mai_n23_), .Y(mai_mai_n662_));
  AOI210     m0640(.A0(i_1_), .A1(mai_mai_n264_), .B0(mai_mai_n662_), .Y(mai_mai_n663_));
  OAI210     m0641(.A0(mai_mai_n663_), .A1(mai_mai_n45_), .B0(mai_mai_n660_), .Y(mai_mai_n664_));
  NA3        m0642(.A(mai_mai_n560_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n665_));
  NA2        m0643(.A(mai_mai_n141_), .B(i_9_), .Y(mai_mai_n666_));
  NA3        m0644(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n668_));
  NA3        m0646(.A(mai_mai_n668_), .B(mai_mai_n273_), .C(mai_mai_n45_), .Y(mai_mai_n669_));
  OAI220     m0647(.A0(mai_mai_n669_), .A1(mai_mai_n667_), .B0(mai_mai_n666_), .B1(mai_mai_n1078_), .Y(mai_mai_n670_));
  NA3        m0648(.A(mai_mai_n649_), .B(mai_mai_n324_), .C(i_6_), .Y(mai_mai_n671_));
  NO2        m0649(.A(mai_mai_n671_), .B(mai_mai_n23_), .Y(mai_mai_n672_));
  AOI210     m0650(.A0(mai_mai_n494_), .A1(mai_mai_n437_), .B0(mai_mai_n244_), .Y(mai_mai_n673_));
  NO2        m0651(.A(mai_mai_n673_), .B(mai_mai_n621_), .Y(mai_mai_n674_));
  NAi21      m0652(.An(mai_mai_n665_), .B(mai_mai_n93_), .Y(mai_mai_n675_));
  NA2        m0653(.A(mai_mai_n668_), .B(mai_mai_n273_), .Y(mai_mai_n676_));
  NO2        m0654(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n677_));
  NA2        m0655(.A(mai_mai_n677_), .B(mai_mai_n24_), .Y(mai_mai_n678_));
  OAI210     m0656(.A0(mai_mai_n678_), .A1(mai_mai_n676_), .B0(mai_mai_n675_), .Y(mai_mai_n679_));
  OR4        m0657(.A(mai_mai_n679_), .B(mai_mai_n674_), .C(mai_mai_n672_), .D(mai_mai_n670_), .Y(mai_mai_n680_));
  NO3        m0658(.A(mai_mai_n680_), .B(mai_mai_n664_), .C(mai_mai_n658_), .Y(mai_mai_n681_));
  NO2        m0659(.A(mai_mai_n239_), .B(mai_mai_n103_), .Y(mai_mai_n682_));
  NO2        m0660(.A(mai_mai_n682_), .B(mai_mai_n637_), .Y(mai_mai_n683_));
  NA2        m0661(.A(mai_mai_n683_), .B(i_1_), .Y(mai_mai_n684_));
  NO2        m0662(.A(mai_mai_n684_), .B(mai_mai_n632_), .Y(mai_mai_n685_));
  NO2        m0663(.A(mai_mai_n432_), .B(mai_mai_n87_), .Y(mai_mai_n686_));
  NA2        m0664(.A(mai_mai_n685_), .B(mai_mai_n47_), .Y(mai_mai_n687_));
  NA2        m0665(.A(i_3_), .B(mai_mai_n198_), .Y(mai_mai_n688_));
  NO2        m0666(.A(mai_mai_n688_), .B(mai_mai_n117_), .Y(mai_mai_n689_));
  AN2        m0667(.A(mai_mai_n689_), .B(mai_mai_n566_), .Y(mai_mai_n690_));
  NO2        m0668(.A(mai_mai_n235_), .B(mai_mai_n45_), .Y(mai_mai_n691_));
  NO3        m0669(.A(mai_mai_n691_), .B(mai_mai_n314_), .C(mai_mai_n240_), .Y(mai_mai_n692_));
  NO2        m0670(.A(mai_mai_n120_), .B(mai_mai_n37_), .Y(mai_mai_n693_));
  NO2        m0671(.A(mai_mai_n693_), .B(i_6_), .Y(mai_mai_n694_));
  NO2        m0672(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n695_));
  NO2        m0673(.A(mai_mai_n695_), .B(mai_mai_n64_), .Y(mai_mai_n696_));
  NO2        m0674(.A(mai_mai_n696_), .B(mai_mai_n652_), .Y(mai_mai_n697_));
  NO4        m0675(.A(mai_mai_n697_), .B(mai_mai_n694_), .C(mai_mai_n692_), .D(i_4_), .Y(mai_mai_n698_));
  NA2        m0676(.A(i_1_), .B(i_3_), .Y(mai_mai_n699_));
  NO2        m0677(.A(mai_mai_n473_), .B(mai_mai_n94_), .Y(mai_mai_n700_));
  AOI210     m0678(.A0(mai_mai_n691_), .A1(mai_mai_n595_), .B0(mai_mai_n700_), .Y(mai_mai_n701_));
  NO2        m0679(.A(mai_mai_n701_), .B(mai_mai_n699_), .Y(mai_mai_n702_));
  NO3        m0680(.A(mai_mai_n702_), .B(mai_mai_n698_), .C(mai_mai_n690_), .Y(mai_mai_n703_));
  NA4        m0681(.A(mai_mai_n703_), .B(mai_mai_n687_), .C(mai_mai_n681_), .D(mai_mai_n654_), .Y(mai_mai_n704_));
  NO3        m0682(.A(mai_mai_n496_), .B(i_3_), .C(i_7_), .Y(mai_mai_n705_));
  NOi21      m0683(.An(mai_mai_n705_), .B(i_10_), .Y(mai_mai_n706_));
  OA210      m0684(.A0(mai_mai_n706_), .A1(mai_mai_n248_), .B0(mai_mai_n87_), .Y(mai_mai_n707_));
  NA2        m0685(.A(mai_mai_n383_), .B(mai_mai_n382_), .Y(mai_mai_n708_));
  NA3        m0686(.A(mai_mai_n503_), .B(mai_mai_n540_), .C(mai_mai_n47_), .Y(mai_mai_n709_));
  NO3        m0687(.A(mai_mai_n497_), .B(mai_mai_n624_), .C(mai_mai_n87_), .Y(mai_mai_n710_));
  NA2        m0688(.A(mai_mai_n710_), .B(mai_mai_n25_), .Y(mai_mai_n711_));
  NA3        m0689(.A(mai_mai_n711_), .B(mai_mai_n709_), .C(mai_mai_n708_), .Y(mai_mai_n712_));
  OAI210     m0690(.A0(mai_mai_n712_), .A1(mai_mai_n707_), .B0(i_1_), .Y(mai_mai_n713_));
  AOI210     m0691(.A0(mai_mai_n273_), .A1(mai_mai_n99_), .B0(i_1_), .Y(mai_mai_n714_));
  NO2        m0692(.A(mai_mai_n381_), .B(i_2_), .Y(mai_mai_n715_));
  NA2        m0693(.A(mai_mai_n715_), .B(mai_mai_n714_), .Y(mai_mai_n716_));
  OAI210     m0694(.A0(mai_mai_n671_), .A1(mai_mai_n467_), .B0(mai_mai_n716_), .Y(mai_mai_n717_));
  INV        m0695(.A(mai_mai_n717_), .Y(mai_mai_n718_));
  AOI210     m0696(.A0(mai_mai_n718_), .A1(mai_mai_n713_), .B0(i_13_), .Y(mai_mai_n719_));
  OR2        m0697(.A(i_11_), .B(i_7_), .Y(mai_mai_n720_));
  AOI210     m0698(.A0(mai_mai_n667_), .A1(mai_mai_n55_), .B0(i_12_), .Y(mai_mai_n721_));
  NO2        m0699(.A(mai_mai_n497_), .B(mai_mai_n24_), .Y(mai_mai_n722_));
  AOI220     m0700(.A0(mai_mai_n722_), .A1(mai_mai_n686_), .B0(mai_mai_n248_), .B1(mai_mai_n134_), .Y(mai_mai_n723_));
  OAI220     m0701(.A0(mai_mai_n723_), .A1(mai_mai_n41_), .B0(mai_mai_n1077_), .B1(mai_mai_n94_), .Y(mai_mai_n724_));
  INV        m0702(.A(mai_mai_n724_), .Y(mai_mai_n725_));
  INV        m0703(.A(mai_mai_n117_), .Y(mai_mai_n726_));
  AOI220     m0704(.A0(mai_mai_n726_), .A1(mai_mai_n73_), .B0(mai_mai_n399_), .B1(mai_mai_n668_), .Y(mai_mai_n727_));
  NO2        m0705(.A(mai_mai_n727_), .B(mai_mai_n245_), .Y(mai_mai_n728_));
  AOI210     m0706(.A0(mai_mai_n467_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n729_));
  NOi31      m0707(.An(mai_mai_n729_), .B(mai_mai_n613_), .C(mai_mai_n45_), .Y(mai_mai_n730_));
  NA2        m0708(.A(mai_mai_n130_), .B(i_13_), .Y(mai_mai_n731_));
  NO2        m0709(.A(mai_mai_n667_), .B(mai_mai_n117_), .Y(mai_mai_n732_));
  INV        m0710(.A(mai_mai_n732_), .Y(mai_mai_n733_));
  OAI220     m0711(.A0(mai_mai_n733_), .A1(mai_mai_n72_), .B0(mai_mai_n731_), .B1(mai_mai_n714_), .Y(mai_mai_n734_));
  NA2        m0712(.A(mai_mai_n26_), .B(mai_mai_n198_), .Y(mai_mai_n735_));
  NA2        m0713(.A(mai_mai_n735_), .B(i_7_), .Y(mai_mai_n736_));
  NO3        m0714(.A(mai_mai_n497_), .B(mai_mai_n239_), .C(mai_mai_n87_), .Y(mai_mai_n737_));
  NA2        m0715(.A(mai_mai_n737_), .B(mai_mai_n736_), .Y(mai_mai_n738_));
  AOI220     m0716(.A0(mai_mai_n399_), .A1(mai_mai_n668_), .B0(mai_mai_n93_), .B1(mai_mai_n104_), .Y(mai_mai_n739_));
  OAI220     m0717(.A0(mai_mai_n739_), .A1(mai_mai_n619_), .B0(mai_mai_n738_), .B1(mai_mai_n634_), .Y(mai_mai_n740_));
  NO4        m0718(.A(mai_mai_n740_), .B(mai_mai_n734_), .C(mai_mai_n730_), .D(mai_mai_n728_), .Y(mai_mai_n741_));
  OR2        m0719(.A(i_11_), .B(i_6_), .Y(mai_mai_n742_));
  NA3        m0720(.A(mai_mai_n618_), .B(mai_mai_n735_), .C(i_7_), .Y(mai_mai_n743_));
  AOI210     m0721(.A0(mai_mai_n743_), .A1(mai_mai_n733_), .B0(mai_mai_n742_), .Y(mai_mai_n744_));
  NA3        m0722(.A(mai_mai_n426_), .B(mai_mai_n623_), .C(mai_mai_n99_), .Y(mai_mai_n745_));
  NA2        m0723(.A(mai_mai_n657_), .B(i_13_), .Y(mai_mai_n746_));
  NA2        m0724(.A(mai_mai_n104_), .B(mai_mai_n735_), .Y(mai_mai_n747_));
  NAi21      m0725(.An(i_11_), .B(i_12_), .Y(mai_mai_n748_));
  NOi41      m0726(.An(mai_mai_n113_), .B(mai_mai_n748_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n749_));
  NO3        m0727(.A(mai_mai_n497_), .B(mai_mai_n601_), .C(mai_mai_n624_), .Y(mai_mai_n750_));
  AOI220     m0728(.A0(mai_mai_n750_), .A1(mai_mai_n318_), .B0(mai_mai_n749_), .B1(mai_mai_n747_), .Y(mai_mai_n751_));
  NA3        m0729(.A(mai_mai_n751_), .B(mai_mai_n746_), .C(mai_mai_n745_), .Y(mai_mai_n752_));
  OAI210     m0730(.A0(mai_mai_n752_), .A1(mai_mai_n744_), .B0(mai_mai_n64_), .Y(mai_mai_n753_));
  NO2        m0731(.A(i_2_), .B(i_12_), .Y(mai_mai_n754_));
  NA2        m0732(.A(mai_mai_n380_), .B(mai_mai_n754_), .Y(mai_mai_n755_));
  NA2        m0733(.A(mai_mai_n382_), .B(mai_mai_n380_), .Y(mai_mai_n756_));
  NO2        m0734(.A(mai_mai_n131_), .B(i_2_), .Y(mai_mai_n757_));
  NA2        m0735(.A(mai_mai_n757_), .B(mai_mai_n652_), .Y(mai_mai_n758_));
  NA3        m0736(.A(mai_mai_n758_), .B(mai_mai_n756_), .C(mai_mai_n755_), .Y(mai_mai_n759_));
  NA3        m0737(.A(mai_mai_n759_), .B(mai_mai_n46_), .C(mai_mai_n228_), .Y(mai_mai_n760_));
  NA4        m0738(.A(mai_mai_n760_), .B(mai_mai_n753_), .C(mai_mai_n741_), .D(mai_mai_n725_), .Y(mai_mai_n761_));
  OR4        m0739(.A(mai_mai_n761_), .B(mai_mai_n719_), .C(mai_mai_n704_), .D(mai_mai_n636_), .Y(mai5));
  NA2        m0740(.A(mai_mai_n683_), .B(mai_mai_n275_), .Y(mai_mai_n763_));
  AN2        m0741(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n764_));
  NA3        m0742(.A(mai_mai_n764_), .B(mai_mai_n754_), .C(mai_mai_n110_), .Y(mai_mai_n765_));
  NO2        m0743(.A(mai_mai_n619_), .B(i_11_), .Y(mai_mai_n766_));
  NA2        m0744(.A(mai_mai_n88_), .B(mai_mai_n766_), .Y(mai_mai_n767_));
  NA3        m0745(.A(mai_mai_n767_), .B(mai_mai_n765_), .C(mai_mai_n763_), .Y(mai_mai_n768_));
  NO3        m0746(.A(i_11_), .B(mai_mai_n239_), .C(i_13_), .Y(mai_mai_n769_));
  NO2        m0747(.A(mai_mai_n127_), .B(mai_mai_n23_), .Y(mai_mai_n770_));
  NA2        m0748(.A(i_12_), .B(i_8_), .Y(mai_mai_n771_));
  OAI210     m0749(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n771_), .Y(mai_mai_n772_));
  INV        m0750(.A(mai_mai_n466_), .Y(mai_mai_n773_));
  AOI220     m0751(.A0(mai_mai_n324_), .A1(mai_mai_n597_), .B0(mai_mai_n772_), .B1(mai_mai_n770_), .Y(mai_mai_n774_));
  INV        m0752(.A(mai_mai_n774_), .Y(mai_mai_n775_));
  NO2        m0753(.A(mai_mai_n775_), .B(mai_mai_n768_), .Y(mai_mai_n776_));
  INV        m0754(.A(mai_mai_n175_), .Y(mai_mai_n777_));
  INV        m0755(.A(mai_mai_n248_), .Y(mai_mai_n778_));
  OAI210     m0756(.A0(mai_mai_n715_), .A1(mai_mai_n468_), .B0(mai_mai_n113_), .Y(mai_mai_n779_));
  AOI210     m0757(.A0(mai_mai_n779_), .A1(mai_mai_n778_), .B0(mai_mai_n777_), .Y(mai_mai_n780_));
  NO2        m0758(.A(mai_mai_n473_), .B(mai_mai_n26_), .Y(mai_mai_n781_));
  NO2        m0759(.A(mai_mai_n781_), .B(mai_mai_n437_), .Y(mai_mai_n782_));
  NA2        m0760(.A(mai_mai_n782_), .B(i_2_), .Y(mai_mai_n783_));
  INV        m0761(.A(mai_mai_n783_), .Y(mai_mai_n784_));
  AOI210     m0762(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n433_), .Y(mai_mai_n785_));
  AOI210     m0763(.A0(mai_mai_n785_), .A1(mai_mai_n784_), .B0(mai_mai_n780_), .Y(mai_mai_n786_));
  NO2        m0764(.A(mai_mai_n195_), .B(mai_mai_n128_), .Y(mai_mai_n787_));
  OAI210     m0765(.A0(mai_mai_n787_), .A1(mai_mai_n770_), .B0(i_2_), .Y(mai_mai_n788_));
  INV        m0766(.A(mai_mai_n176_), .Y(mai_mai_n789_));
  NO3        m0767(.A(mai_mai_n638_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n790_));
  AOI210     m0768(.A0(mai_mai_n789_), .A1(mai_mai_n88_), .B0(mai_mai_n790_), .Y(mai_mai_n791_));
  AOI210     m0769(.A0(mai_mai_n791_), .A1(mai_mai_n788_), .B0(mai_mai_n198_), .Y(mai_mai_n792_));
  OA210      m0770(.A0(mai_mai_n639_), .A1(mai_mai_n129_), .B0(i_13_), .Y(mai_mai_n793_));
  NA2        m0771(.A(mai_mai_n205_), .B(mai_mai_n208_), .Y(mai_mai_n794_));
  NA2        m0772(.A(mai_mai_n154_), .B(mai_mai_n614_), .Y(mai_mai_n795_));
  AOI210     m0773(.A0(mai_mai_n795_), .A1(mai_mai_n794_), .B0(mai_mai_n385_), .Y(mai_mai_n796_));
  AOI210     m0774(.A0(mai_mai_n213_), .A1(mai_mai_n151_), .B0(mai_mai_n540_), .Y(mai_mai_n797_));
  NA2        m0775(.A(mai_mai_n797_), .B(mai_mai_n437_), .Y(mai_mai_n798_));
  NO2        m0776(.A(mai_mai_n104_), .B(mai_mai_n45_), .Y(mai_mai_n799_));
  INV        m0777(.A(mai_mai_n307_), .Y(mai_mai_n800_));
  NA4        m0778(.A(mai_mai_n800_), .B(mai_mai_n311_), .C(mai_mai_n127_), .D(mai_mai_n43_), .Y(mai_mai_n801_));
  OAI210     m0779(.A0(mai_mai_n801_), .A1(mai_mai_n799_), .B0(mai_mai_n798_), .Y(mai_mai_n802_));
  NO4        m0780(.A(mai_mai_n802_), .B(mai_mai_n796_), .C(mai_mai_n793_), .D(mai_mai_n792_), .Y(mai_mai_n803_));
  NA2        m0781(.A(mai_mai_n597_), .B(mai_mai_n28_), .Y(mai_mai_n804_));
  NA2        m0782(.A(mai_mai_n769_), .B(mai_mai_n279_), .Y(mai_mai_n805_));
  NA2        m0783(.A(mai_mai_n805_), .B(mai_mai_n804_), .Y(mai_mai_n806_));
  NO2        m0784(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n807_));
  NO2        m0785(.A(mai_mai_n807_), .B(mai_mai_n129_), .Y(mai_mai_n808_));
  NO2        m0786(.A(mai_mai_n808_), .B(mai_mai_n614_), .Y(mai_mai_n809_));
  AOI220     m0787(.A0(mai_mai_n809_), .A1(mai_mai_n36_), .B0(mai_mai_n806_), .B1(mai_mai_n47_), .Y(mai_mai_n810_));
  NA4        m0788(.A(mai_mai_n810_), .B(mai_mai_n803_), .C(mai_mai_n786_), .D(mai_mai_n776_), .Y(mai6));
  NO3        m0789(.A(mai_mai_n259_), .B(mai_mai_n313_), .C(i_1_), .Y(mai_mai_n812_));
  NO2        m0790(.A(mai_mai_n190_), .B(mai_mai_n142_), .Y(mai_mai_n813_));
  OAI210     m0791(.A0(mai_mai_n813_), .A1(mai_mai_n812_), .B0(mai_mai_n757_), .Y(mai_mai_n814_));
  NO2        m0792(.A(mai_mai_n223_), .B(mai_mai_n507_), .Y(mai_mai_n815_));
  NO2        m0793(.A(i_11_), .B(i_9_), .Y(mai_mai_n816_));
  INV        m0794(.A(mai_mai_n336_), .Y(mai_mai_n817_));
  AO210      m0795(.A0(mai_mai_n817_), .A1(mai_mai_n814_), .B0(i_12_), .Y(mai_mai_n818_));
  NA2        m0796(.A(mai_mai_n386_), .B(mai_mai_n343_), .Y(mai_mai_n819_));
  NA2        m0797(.A(mai_mai_n601_), .B(mai_mai_n64_), .Y(mai_mai_n820_));
  NA2        m0798(.A(mai_mai_n706_), .B(mai_mai_n72_), .Y(mai_mai_n821_));
  NA3        m0799(.A(mai_mai_n821_), .B(mai_mai_n820_), .C(mai_mai_n819_), .Y(mai_mai_n822_));
  INV        m0800(.A(mai_mai_n202_), .Y(mai_mai_n823_));
  AOI220     m0801(.A0(mai_mai_n823_), .A1(mai_mai_n816_), .B0(mai_mai_n822_), .B1(mai_mai_n74_), .Y(mai_mai_n824_));
  INV        m0802(.A(mai_mai_n335_), .Y(mai_mai_n825_));
  NA2        m0803(.A(mai_mai_n76_), .B(mai_mai_n134_), .Y(mai_mai_n826_));
  INV        m0804(.A(mai_mai_n127_), .Y(mai_mai_n827_));
  NA2        m0805(.A(mai_mai_n827_), .B(mai_mai_n47_), .Y(mai_mai_n828_));
  AOI210     m0806(.A0(mai_mai_n828_), .A1(mai_mai_n826_), .B0(mai_mai_n825_), .Y(mai_mai_n829_));
  NO2        m0807(.A(mai_mai_n255_), .B(i_9_), .Y(mai_mai_n830_));
  NA2        m0808(.A(mai_mai_n830_), .B(mai_mai_n807_), .Y(mai_mai_n831_));
  AOI210     m0809(.A0(mai_mai_n831_), .A1(mai_mai_n538_), .B0(mai_mai_n190_), .Y(mai_mai_n832_));
  NO2        m0810(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n833_));
  NA3        m0811(.A(mai_mai_n833_), .B(mai_mai_n492_), .C(mai_mai_n403_), .Y(mai_mai_n834_));
  NAi32      m0812(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n835_));
  NO2        m0813(.A(mai_mai_n742_), .B(mai_mai_n835_), .Y(mai_mai_n836_));
  OAI210     m0814(.A0(mai_mai_n705_), .A1(mai_mai_n587_), .B0(mai_mai_n586_), .Y(mai_mai_n837_));
  NAi31      m0815(.An(mai_mai_n836_), .B(mai_mai_n837_), .C(mai_mai_n834_), .Y(mai_mai_n838_));
  OR3        m0816(.A(mai_mai_n838_), .B(mai_mai_n832_), .C(mai_mai_n829_), .Y(mai_mai_n839_));
  NO2        m0817(.A(mai_mai_n720_), .B(i_2_), .Y(mai_mai_n840_));
  NA2        m0818(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n841_));
  NO2        m0819(.A(mai_mai_n841_), .B(mai_mai_n425_), .Y(mai_mai_n842_));
  NA2        m0820(.A(mai_mai_n842_), .B(mai_mai_n840_), .Y(mai_mai_n843_));
  AO220      m0821(.A0(mai_mai_n371_), .A1(mai_mai_n361_), .B0(mai_mai_n409_), .B1(mai_mai_n614_), .Y(mai_mai_n844_));
  NA3        m0822(.A(mai_mai_n844_), .B(mai_mai_n260_), .C(i_7_), .Y(mai_mai_n845_));
  OR2        m0823(.A(mai_mai_n639_), .B(mai_mai_n468_), .Y(mai_mai_n846_));
  NA3        m0824(.A(mai_mai_n846_), .B(mai_mai_n150_), .C(mai_mai_n70_), .Y(mai_mai_n847_));
  AO210      m0825(.A0(mai_mai_n514_), .A1(mai_mai_n773_), .B0(mai_mai_n36_), .Y(mai_mai_n848_));
  NA4        m0826(.A(mai_mai_n848_), .B(mai_mai_n847_), .C(mai_mai_n845_), .D(mai_mai_n843_), .Y(mai_mai_n849_));
  NO2        m0827(.A(i_6_), .B(i_11_), .Y(mai_mai_n850_));
  AOI220     m0828(.A0(mai_mai_n850_), .A1(mai_mai_n586_), .B0(mai_mai_n815_), .B1(mai_mai_n736_), .Y(mai_mai_n851_));
  NA3        m0829(.A(mai_mai_n385_), .B(mai_mai_n241_), .C(mai_mai_n150_), .Y(mai_mai_n852_));
  NA2        m0830(.A(mai_mai_n409_), .B(mai_mai_n71_), .Y(mai_mai_n853_));
  NA4        m0831(.A(mai_mai_n853_), .B(mai_mai_n852_), .C(mai_mai_n851_), .D(mai_mai_n622_), .Y(mai_mai_n854_));
  AN2        m0832(.A(mai_mai_n540_), .B(mai_mai_n47_), .Y(mai_mai_n855_));
  NA3        m0833(.A(mai_mai_n855_), .B(mai_mai_n503_), .C(mai_mai_n222_), .Y(mai_mai_n856_));
  AOI210     m0834(.A0(mai_mai_n468_), .A1(mai_mai_n466_), .B0(mai_mai_n585_), .Y(mai_mai_n857_));
  NO2        m0835(.A(mai_mai_n630_), .B(mai_mai_n104_), .Y(mai_mai_n858_));
  OAI210     m0836(.A0(mai_mai_n858_), .A1(mai_mai_n114_), .B0(mai_mai_n423_), .Y(mai_mai_n859_));
  INV        m0837(.A(mai_mai_n605_), .Y(mai_mai_n860_));
  NA3        m0838(.A(mai_mai_n860_), .B(mai_mai_n335_), .C(i_7_), .Y(mai_mai_n861_));
  NA4        m0839(.A(mai_mai_n861_), .B(mai_mai_n859_), .C(mai_mai_n857_), .D(mai_mai_n856_), .Y(mai_mai_n862_));
  NO4        m0840(.A(mai_mai_n862_), .B(mai_mai_n854_), .C(mai_mai_n849_), .D(mai_mai_n839_), .Y(mai_mai_n863_));
  NA4        m0841(.A(mai_mai_n863_), .B(mai_mai_n824_), .C(mai_mai_n818_), .D(mai_mai_n393_), .Y(mai3));
  NA2        m0842(.A(i_12_), .B(i_10_), .Y(mai_mai_n865_));
  NA2        m0843(.A(i_6_), .B(i_7_), .Y(mai_mai_n866_));
  NO2        m0844(.A(mai_mai_n866_), .B(i_0_), .Y(mai_mai_n867_));
  NO2        m0845(.A(i_11_), .B(mai_mai_n239_), .Y(mai_mai_n868_));
  OAI210     m0846(.A0(mai_mai_n867_), .A1(mai_mai_n295_), .B0(mai_mai_n868_), .Y(mai_mai_n869_));
  NO2        m0847(.A(mai_mai_n869_), .B(mai_mai_n198_), .Y(mai_mai_n870_));
  NO3        m0848(.A(mai_mai_n469_), .B(mai_mai_n91_), .C(mai_mai_n45_), .Y(mai_mai_n871_));
  OA210      m0849(.A0(mai_mai_n871_), .A1(mai_mai_n870_), .B0(mai_mai_n178_), .Y(mai_mai_n872_));
  NA3        m0850(.A(mai_mai_n852_), .B(mai_mai_n622_), .C(mai_mai_n384_), .Y(mai_mai_n873_));
  NA2        m0851(.A(mai_mai_n873_), .B(mai_mai_n40_), .Y(mai_mai_n874_));
  NOi21      m0852(.An(mai_mai_n98_), .B(mai_mai_n782_), .Y(mai_mai_n875_));
  NO3        m0853(.A(mai_mai_n647_), .B(mai_mai_n473_), .C(mai_mai_n134_), .Y(mai_mai_n876_));
  NA2        m0854(.A(mai_mai_n426_), .B(mai_mai_n46_), .Y(mai_mai_n877_));
  AN2        m0855(.A(mai_mai_n471_), .B(mai_mai_n56_), .Y(mai_mai_n878_));
  NO3        m0856(.A(mai_mai_n878_), .B(mai_mai_n876_), .C(mai_mai_n875_), .Y(mai_mai_n879_));
  AOI210     m0857(.A0(mai_mai_n879_), .A1(mai_mai_n874_), .B0(mai_mai_n49_), .Y(mai_mai_n880_));
  NO4        m0858(.A(mai_mai_n389_), .B(mai_mai_n396_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n881_));
  NA2        m0859(.A(mai_mai_n190_), .B(mai_mai_n595_), .Y(mai_mai_n882_));
  NOi21      m0860(.An(mai_mai_n882_), .B(mai_mai_n881_), .Y(mai_mai_n883_));
  NA2        m0861(.A(mai_mai_n729_), .B(mai_mai_n695_), .Y(mai_mai_n884_));
  NA2        m0862(.A(mai_mai_n341_), .B(mai_mai_n457_), .Y(mai_mai_n885_));
  OAI220     m0863(.A0(mai_mai_n885_), .A1(mai_mai_n884_), .B0(mai_mai_n883_), .B1(mai_mai_n64_), .Y(mai_mai_n886_));
  NOi21      m0864(.An(i_5_), .B(i_9_), .Y(mai_mai_n887_));
  NA2        m0865(.A(mai_mai_n887_), .B(mai_mai_n465_), .Y(mai_mai_n888_));
  BUFFER     m0866(.A(mai_mai_n273_), .Y(mai_mai_n889_));
  AOI210     m0867(.A0(mai_mai_n889_), .A1(mai_mai_n494_), .B0(mai_mai_n710_), .Y(mai_mai_n890_));
  NO3        m0868(.A(mai_mai_n429_), .B(mai_mai_n273_), .C(mai_mai_n74_), .Y(mai_mai_n891_));
  NO2        m0869(.A(mai_mai_n179_), .B(mai_mai_n151_), .Y(mai_mai_n892_));
  AOI210     m0870(.A0(mai_mai_n892_), .A1(mai_mai_n247_), .B0(mai_mai_n891_), .Y(mai_mai_n893_));
  OAI220     m0871(.A0(mai_mai_n893_), .A1(mai_mai_n185_), .B0(mai_mai_n890_), .B1(mai_mai_n888_), .Y(mai_mai_n894_));
  NO4        m0872(.A(mai_mai_n894_), .B(mai_mai_n886_), .C(mai_mai_n880_), .D(mai_mai_n872_), .Y(mai_mai_n895_));
  NA2        m0873(.A(mai_mai_n190_), .B(mai_mai_n24_), .Y(mai_mai_n896_));
  NA2        m0874(.A(mai_mai_n318_), .B(mai_mai_n132_), .Y(mai_mai_n897_));
  NO2        m0875(.A(mai_mai_n897_), .B(mai_mai_n415_), .Y(mai_mai_n898_));
  INV        m0876(.A(mai_mai_n898_), .Y(mai_mai_n899_));
  NO2        m0877(.A(mai_mai_n403_), .B(mai_mai_n299_), .Y(mai_mai_n900_));
  NA2        m0878(.A(mai_mai_n900_), .B(mai_mai_n732_), .Y(mai_mai_n901_));
  NA2        m0879(.A(mai_mai_n596_), .B(i_0_), .Y(mai_mai_n902_));
  NO4        m0880(.A(mai_mai_n604_), .B(mai_mai_n220_), .C(mai_mai_n433_), .D(mai_mai_n425_), .Y(mai_mai_n903_));
  NA2        m0881(.A(mai_mai_n903_), .B(i_11_), .Y(mai_mai_n904_));
  AN2        m0882(.A(mai_mai_n98_), .B(mai_mai_n246_), .Y(mai_mai_n905_));
  NA2        m0883(.A(mai_mai_n769_), .B(mai_mai_n336_), .Y(mai_mai_n906_));
  AOI210     m0884(.A0(mai_mai_n503_), .A1(mai_mai_n88_), .B0(mai_mai_n59_), .Y(mai_mai_n907_));
  OAI220     m0885(.A0(mai_mai_n907_), .A1(mai_mai_n906_), .B0(mai_mai_n678_), .B1(mai_mai_n562_), .Y(mai_mai_n908_));
  NO2        m0886(.A(mai_mai_n257_), .B(mai_mai_n156_), .Y(mai_mai_n909_));
  NA2        m0887(.A(i_0_), .B(i_10_), .Y(mai_mai_n910_));
  OAI210     m0888(.A0(mai_mai_n910_), .A1(mai_mai_n87_), .B0(mai_mai_n565_), .Y(mai_mai_n911_));
  NO4        m0889(.A(mai_mai_n117_), .B(mai_mai_n59_), .C(mai_mai_n688_), .D(i_5_), .Y(mai_mai_n912_));
  AO220      m0890(.A0(mai_mai_n912_), .A1(mai_mai_n911_), .B0(mai_mai_n909_), .B1(i_6_), .Y(mai_mai_n913_));
  AOI220     m0891(.A0(mai_mai_n341_), .A1(mai_mai_n100_), .B0(mai_mai_n190_), .B1(mai_mai_n85_), .Y(mai_mai_n914_));
  NA2        m0892(.A(mai_mai_n590_), .B(i_4_), .Y(mai_mai_n915_));
  NA2        m0893(.A(mai_mai_n193_), .B(mai_mai_n208_), .Y(mai_mai_n916_));
  OAI220     m0894(.A0(mai_mai_n916_), .A1(mai_mai_n906_), .B0(mai_mai_n915_), .B1(mai_mai_n914_), .Y(mai_mai_n917_));
  NO4        m0895(.A(mai_mai_n917_), .B(mai_mai_n913_), .C(mai_mai_n908_), .D(mai_mai_n905_), .Y(mai_mai_n918_));
  NA4        m0896(.A(mai_mai_n918_), .B(mai_mai_n904_), .C(mai_mai_n901_), .D(mai_mai_n899_), .Y(mai_mai_n919_));
  NA2        m0897(.A(i_11_), .B(i_9_), .Y(mai_mai_n920_));
  NO2        m0898(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n921_));
  NA2        m0899(.A(mai_mai_n408_), .B(mai_mai_n183_), .Y(mai_mai_n922_));
  NA2        m0900(.A(mai_mai_n922_), .B(mai_mai_n163_), .Y(mai_mai_n923_));
  NO2        m0901(.A(mai_mai_n920_), .B(mai_mai_n74_), .Y(mai_mai_n924_));
  NO2        m0902(.A(mai_mai_n179_), .B(i_0_), .Y(mai_mai_n925_));
  INV        m0903(.A(mai_mai_n925_), .Y(mai_mai_n926_));
  NA2        m0904(.A(mai_mai_n492_), .B(mai_mai_n233_), .Y(mai_mai_n927_));
  AOI210     m0905(.A0(mai_mai_n383_), .A1(mai_mai_n42_), .B0(mai_mai_n422_), .Y(mai_mai_n928_));
  OAI220     m0906(.A0(mai_mai_n928_), .A1(mai_mai_n888_), .B0(mai_mai_n927_), .B1(mai_mai_n926_), .Y(mai_mai_n929_));
  NO2        m0907(.A(mai_mai_n929_), .B(mai_mai_n923_), .Y(mai_mai_n930_));
  NA2        m0908(.A(mai_mai_n677_), .B(mai_mai_n124_), .Y(mai_mai_n931_));
  NO2        m0909(.A(i_6_), .B(mai_mai_n931_), .Y(mai_mai_n932_));
  AOI210     m0910(.A0(mai_mai_n467_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n933_));
  NA2        m0911(.A(mai_mai_n175_), .B(mai_mai_n105_), .Y(mai_mai_n934_));
  NOi32      m0912(.An(mai_mai_n933_), .Bn(mai_mai_n193_), .C(mai_mai_n934_), .Y(mai_mai_n935_));
  NA2        m0913(.A(mai_mai_n623_), .B(mai_mai_n336_), .Y(mai_mai_n936_));
  NO2        m0914(.A(mai_mai_n936_), .B(mai_mai_n877_), .Y(mai_mai_n937_));
  NO3        m0915(.A(mai_mai_n937_), .B(mai_mai_n935_), .C(mai_mai_n932_), .Y(mai_mai_n938_));
  NOi21      m0916(.An(i_7_), .B(i_5_), .Y(mai_mai_n939_));
  OR2        m0917(.A(mai_mai_n934_), .B(mai_mai_n538_), .Y(mai_mai_n940_));
  NO3        m0918(.A(mai_mai_n418_), .B(mai_mai_n372_), .C(mai_mai_n370_), .Y(mai_mai_n941_));
  NO2        m0919(.A(mai_mai_n267_), .B(mai_mai_n325_), .Y(mai_mai_n942_));
  NO2        m0920(.A(mai_mai_n748_), .B(mai_mai_n262_), .Y(mai_mai_n943_));
  AOI210     m0921(.A0(mai_mai_n943_), .A1(mai_mai_n942_), .B0(mai_mai_n941_), .Y(mai_mai_n944_));
  NA4        m0922(.A(mai_mai_n944_), .B(mai_mai_n940_), .C(mai_mai_n938_), .D(mai_mai_n930_), .Y(mai_mai_n945_));
  NO2        m0923(.A(mai_mai_n896_), .B(mai_mai_n242_), .Y(mai_mai_n946_));
  AN2        m0924(.A(mai_mai_n340_), .B(mai_mai_n336_), .Y(mai_mai_n947_));
  AN2        m0925(.A(mai_mai_n947_), .B(mai_mai_n892_), .Y(mai_mai_n948_));
  OAI210     m0926(.A0(mai_mai_n948_), .A1(mai_mai_n946_), .B0(i_10_), .Y(mai_mai_n949_));
  NO2        m0927(.A(mai_mai_n865_), .B(mai_mai_n324_), .Y(mai_mai_n950_));
  OA210      m0928(.A0(mai_mai_n492_), .A1(mai_mai_n226_), .B0(mai_mai_n491_), .Y(mai_mai_n951_));
  NA2        m0929(.A(mai_mai_n950_), .B(mai_mai_n924_), .Y(mai_mai_n952_));
  NO2        m0930(.A(mai_mai_n260_), .B(mai_mai_n47_), .Y(mai_mai_n953_));
  NA2        m0931(.A(mai_mai_n924_), .B(mai_mai_n311_), .Y(mai_mai_n954_));
  OAI210     m0932(.A0(mai_mai_n953_), .A1(mai_mai_n192_), .B0(mai_mai_n954_), .Y(mai_mai_n955_));
  NA2        m0933(.A(mai_mai_n955_), .B(mai_mai_n492_), .Y(mai_mai_n956_));
  NA2        m0934(.A(mai_mai_n94_), .B(mai_mai_n45_), .Y(mai_mai_n957_));
  NO2        m0935(.A(mai_mai_n76_), .B(mai_mai_n771_), .Y(mai_mai_n958_));
  NA2        m0936(.A(mai_mai_n958_), .B(mai_mai_n957_), .Y(mai_mai_n959_));
  NO2        m0937(.A(mai_mai_n959_), .B(mai_mai_n48_), .Y(mai_mai_n960_));
  NA2        m0938(.A(mai_mai_n722_), .B(mai_mai_n569_), .Y(mai_mai_n961_));
  NAi21      m0939(.An(i_9_), .B(i_5_), .Y(mai_mai_n962_));
  NO2        m0940(.A(mai_mai_n962_), .B(mai_mai_n418_), .Y(mai_mai_n963_));
  NO2        m0941(.A(mai_mai_n617_), .B(mai_mai_n107_), .Y(mai_mai_n964_));
  AOI220     m0942(.A0(mai_mai_n964_), .A1(i_0_), .B0(mai_mai_n963_), .B1(mai_mai_n639_), .Y(mai_mai_n965_));
  OAI220     m0943(.A0(mai_mai_n965_), .A1(mai_mai_n87_), .B0(mai_mai_n961_), .B1(mai_mai_n176_), .Y(mai_mai_n966_));
  NO3        m0944(.A(mai_mai_n966_), .B(mai_mai_n960_), .C(mai_mai_n543_), .Y(mai_mai_n967_));
  NA4        m0945(.A(mai_mai_n967_), .B(mai_mai_n956_), .C(mai_mai_n952_), .D(mai_mai_n949_), .Y(mai_mai_n968_));
  NO3        m0946(.A(mai_mai_n968_), .B(mai_mai_n945_), .C(mai_mai_n919_), .Y(mai_mai_n969_));
  NO2        m0947(.A(i_0_), .B(mai_mai_n748_), .Y(mai_mai_n970_));
  NA2        m0948(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n971_));
  NA2        m0949(.A(mai_mai_n910_), .B(mai_mai_n971_), .Y(mai_mai_n972_));
  NO3        m0950(.A(mai_mai_n107_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n973_));
  AO220      m0951(.A0(mai_mai_n973_), .A1(mai_mai_n972_), .B0(mai_mai_n970_), .B1(mai_mai_n178_), .Y(mai_mai_n974_));
  AOI210     m0952(.A0(mai_mai_n820_), .A1(mai_mai_n708_), .B0(mai_mai_n934_), .Y(mai_mai_n975_));
  AOI210     m0953(.A0(mai_mai_n974_), .A1(mai_mai_n358_), .B0(mai_mai_n975_), .Y(mai_mai_n976_));
  NA2        m0954(.A(mai_mai_n757_), .B(mai_mai_n149_), .Y(mai_mai_n977_));
  INV        m0955(.A(mai_mai_n977_), .Y(mai_mai_n978_));
  NA3        m0956(.A(mai_mai_n978_), .B(mai_mai_n695_), .C(mai_mai_n74_), .Y(mai_mai_n979_));
  NO2        m0957(.A(mai_mai_n837_), .B(mai_mai_n418_), .Y(mai_mai_n980_));
  NA3        m0958(.A(mai_mai_n867_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n981_));
  NA2        m0959(.A(mai_mai_n868_), .B(i_9_), .Y(mai_mai_n982_));
  AOI210     m0960(.A0(mai_mai_n981_), .A1(mai_mai_n519_), .B0(mai_mai_n982_), .Y(mai_mai_n983_));
  OAI210     m0961(.A0(mai_mai_n247_), .A1(i_9_), .B0(mai_mai_n232_), .Y(mai_mai_n984_));
  AOI210     m0962(.A0(mai_mai_n984_), .A1(mai_mai_n902_), .B0(mai_mai_n156_), .Y(mai_mai_n985_));
  NO3        m0963(.A(mai_mai_n985_), .B(mai_mai_n983_), .C(mai_mai_n980_), .Y(mai_mai_n986_));
  NA3        m0964(.A(mai_mai_n986_), .B(mai_mai_n979_), .C(mai_mai_n976_), .Y(mai_mai_n987_));
  NA2        m0965(.A(mai_mai_n947_), .B(mai_mai_n385_), .Y(mai_mai_n988_));
  AOI210     m0966(.A0(mai_mai_n306_), .A1(mai_mai_n165_), .B0(mai_mai_n988_), .Y(mai_mai_n989_));
  NA3        m0967(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n990_));
  NA2        m0968(.A(mai_mai_n921_), .B(mai_mai_n508_), .Y(mai_mai_n991_));
  AOI210     m0969(.A0(mai_mai_n990_), .A1(mai_mai_n165_), .B0(mai_mai_n991_), .Y(mai_mai_n992_));
  NO2        m0970(.A(mai_mai_n992_), .B(mai_mai_n989_), .Y(mai_mai_n993_));
  NO3        m0971(.A(mai_mai_n910_), .B(mai_mai_n887_), .C(mai_mai_n195_), .Y(mai_mai_n994_));
  AOI220     m0972(.A0(mai_mai_n994_), .A1(i_11_), .B0(mai_mai_n591_), .B1(mai_mai_n76_), .Y(mai_mai_n995_));
  NO3        m0973(.A(mai_mai_n214_), .B(mai_mai_n396_), .C(i_0_), .Y(mai_mai_n996_));
  OAI210     m0974(.A0(mai_mai_n996_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n997_));
  INV        m0975(.A(mai_mai_n222_), .Y(mai_mai_n998_));
  OAI220     m0976(.A0(mai_mai_n555_), .A1(mai_mai_n142_), .B0(mai_mai_n661_), .B1(mai_mai_n634_), .Y(mai_mai_n999_));
  NA3        m0977(.A(mai_mai_n999_), .B(mai_mai_n410_), .C(mai_mai_n998_), .Y(mai_mai_n1000_));
  NA4        m0978(.A(mai_mai_n1000_), .B(mai_mai_n997_), .C(mai_mai_n995_), .D(mai_mai_n993_), .Y(mai_mai_n1001_));
  INV        m0979(.A(mai_mai_n111_), .Y(mai_mai_n1002_));
  AOI220     m0980(.A0(mai_mai_n939_), .A1(mai_mai_n508_), .B0(mai_mai_n867_), .B1(mai_mai_n166_), .Y(mai_mai_n1003_));
  NA2        m0981(.A(mai_mai_n361_), .B(mai_mai_n180_), .Y(mai_mai_n1004_));
  OA220      m0982(.A0(mai_mai_n1004_), .A1(mai_mai_n1003_), .B0(mai_mai_n1002_), .B1(i_5_), .Y(mai_mai_n1005_));
  AOI210     m0983(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n179_), .Y(mai_mai_n1006_));
  NA2        m0984(.A(mai_mai_n1006_), .B(mai_mai_n951_), .Y(mai_mai_n1007_));
  NA3        m0985(.A(mai_mai_n631_), .B(mai_mai_n190_), .C(mai_mai_n85_), .Y(mai_mai_n1008_));
  INV        m0986(.A(mai_mai_n1008_), .Y(mai_mai_n1009_));
  NO3        m0987(.A(mai_mai_n877_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n1010_));
  NA2        m0988(.A(mai_mai_n513_), .B(mai_mai_n506_), .Y(mai_mai_n1011_));
  NO3        m0989(.A(mai_mai_n1011_), .B(mai_mai_n1010_), .C(mai_mai_n1009_), .Y(mai_mai_n1012_));
  NA3        m0990(.A(mai_mai_n403_), .B(mai_mai_n175_), .C(mai_mai_n174_), .Y(mai_mai_n1013_));
  NA3        m0991(.A(mai_mai_n403_), .B(mai_mai_n342_), .C(mai_mai_n224_), .Y(mai_mai_n1014_));
  INV        m0992(.A(mai_mai_n1014_), .Y(mai_mai_n1015_));
  NOi31      m0993(.An(mai_mai_n402_), .B(mai_mai_n971_), .C(mai_mai_n242_), .Y(mai_mai_n1016_));
  NO3        m0994(.A(mai_mai_n920_), .B(mai_mai_n222_), .C(mai_mai_n195_), .Y(mai_mai_n1017_));
  NO4        m0995(.A(mai_mai_n1017_), .B(mai_mai_n1016_), .C(mai_mai_n1015_), .D(mai_mai_n1080_), .Y(mai_mai_n1018_));
  NA4        m0996(.A(mai_mai_n1018_), .B(mai_mai_n1012_), .C(mai_mai_n1007_), .D(mai_mai_n1005_), .Y(mai_mai_n1019_));
  INV        m0997(.A(mai_mai_n633_), .Y(mai_mai_n1020_));
  NO3        m0998(.A(mai_mai_n1020_), .B(mai_mai_n581_), .C(mai_mai_n355_), .Y(mai_mai_n1021_));
  NO2        m0999(.A(mai_mai_n87_), .B(i_5_), .Y(mai_mai_n1022_));
  NA3        m1000(.A(mai_mai_n868_), .B(mai_mai_n112_), .C(mai_mai_n127_), .Y(mai_mai_n1023_));
  INV        m1001(.A(mai_mai_n1023_), .Y(mai_mai_n1024_));
  AOI210     m1002(.A0(mai_mai_n1024_), .A1(mai_mai_n1022_), .B0(mai_mai_n1021_), .Y(mai_mai_n1025_));
  NAi21      m1003(.An(mai_mai_n244_), .B(mai_mai_n245_), .Y(mai_mai_n1026_));
  NO4        m1004(.A(mai_mai_n242_), .B(mai_mai_n214_), .C(i_0_), .D(i_12_), .Y(mai_mai_n1027_));
  NA2        m1005(.A(mai_mai_n1027_), .B(mai_mai_n1026_), .Y(mai_mai_n1028_));
  AN2        m1006(.A(mai_mai_n910_), .B(mai_mai_n156_), .Y(mai_mai_n1029_));
  NO4        m1007(.A(mai_mai_n1029_), .B(i_12_), .C(mai_mai_n665_), .D(mai_mai_n134_), .Y(mai_mai_n1030_));
  NA2        m1008(.A(mai_mai_n1030_), .B(mai_mai_n222_), .Y(mai_mai_n1031_));
  NA3        m1009(.A(mai_mai_n100_), .B(mai_mai_n595_), .C(i_11_), .Y(mai_mai_n1032_));
  NO2        m1010(.A(mai_mai_n1032_), .B(mai_mai_n158_), .Y(mai_mai_n1033_));
  NA2        m1011(.A(mai_mai_n939_), .B(mai_mai_n490_), .Y(mai_mai_n1034_));
  NO2        m1012(.A(mai_mai_n1034_), .B(mai_mai_n696_), .Y(mai_mai_n1035_));
  AOI210     m1013(.A0(mai_mai_n1035_), .A1(mai_mai_n925_), .B0(mai_mai_n1033_), .Y(mai_mai_n1036_));
  NA4        m1014(.A(mai_mai_n1036_), .B(mai_mai_n1031_), .C(mai_mai_n1028_), .D(mai_mai_n1025_), .Y(mai_mai_n1037_));
  NO4        m1015(.A(mai_mai_n1037_), .B(mai_mai_n1019_), .C(mai_mai_n1001_), .D(mai_mai_n987_), .Y(mai_mai_n1038_));
  OAI210     m1016(.A0(mai_mai_n840_), .A1(mai_mai_n833_), .B0(mai_mai_n37_), .Y(mai_mai_n1039_));
  NA3        m1017(.A(mai_mai_n933_), .B(mai_mai_n380_), .C(i_5_), .Y(mai_mai_n1040_));
  NA3        m1018(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n629_), .Y(mai_mai_n1041_));
  NA2        m1019(.A(mai_mai_n1041_), .B(mai_mai_n211_), .Y(mai_mai_n1042_));
  BUFFER     m1020(.A(mai_mai_n381_), .Y(mai_mai_n1043_));
  NA2        m1021(.A(mai_mai_n191_), .B(mai_mai_n193_), .Y(mai_mai_n1044_));
  AO210      m1022(.A0(mai_mai_n1043_), .A1(mai_mai_n33_), .B0(mai_mai_n1044_), .Y(mai_mai_n1045_));
  OAI210     m1023(.A0(mai_mai_n633_), .A1(mai_mai_n631_), .B0(mai_mai_n324_), .Y(mai_mai_n1046_));
  NAi31      m1024(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n1047_));
  AOI210     m1025(.A0(mai_mai_n120_), .A1(mai_mai_n71_), .B0(mai_mai_n1047_), .Y(mai_mai_n1048_));
  NO2        m1026(.A(mai_mai_n1048_), .B(mai_mai_n662_), .Y(mai_mai_n1049_));
  NA3        m1027(.A(mai_mai_n1049_), .B(mai_mai_n1046_), .C(mai_mai_n1045_), .Y(mai_mai_n1050_));
  NO2        m1028(.A(mai_mai_n481_), .B(mai_mai_n273_), .Y(mai_mai_n1051_));
  NO4        m1029(.A(mai_mai_n235_), .B(mai_mai_n148_), .C(mai_mai_n699_), .D(mai_mai_n37_), .Y(mai_mai_n1052_));
  NO3        m1030(.A(mai_mai_n1052_), .B(mai_mai_n1051_), .C(mai_mai_n903_), .Y(mai_mai_n1053_));
  OAI210     m1031(.A0(mai_mai_n1032_), .A1(mai_mai_n151_), .B0(mai_mai_n1053_), .Y(mai_mai_n1054_));
  AOI210     m1032(.A0(mai_mai_n1050_), .A1(mai_mai_n49_), .B0(mai_mai_n1054_), .Y(mai_mai_n1055_));
  AOI210     m1033(.A0(mai_mai_n1055_), .A1(mai_mai_n1042_), .B0(mai_mai_n74_), .Y(mai_mai_n1056_));
  NO2        m1034(.A(mai_mai_n588_), .B(mai_mai_n392_), .Y(mai_mai_n1057_));
  NO2        m1035(.A(mai_mai_n1057_), .B(mai_mai_n777_), .Y(mai_mai_n1058_));
  NA2        m1036(.A(mai_mai_n267_), .B(mai_mai_n58_), .Y(mai_mai_n1059_));
  AOI220     m1037(.A0(mai_mai_n1059_), .A1(mai_mai_n77_), .B0(mai_mai_n356_), .B1(mai_mai_n259_), .Y(mai_mai_n1060_));
  NO2        m1038(.A(mai_mai_n1060_), .B(mai_mai_n239_), .Y(mai_mai_n1061_));
  NA3        m1039(.A(mai_mai_n98_), .B(mai_mai_n313_), .C(mai_mai_n31_), .Y(mai_mai_n1062_));
  INV        m1040(.A(mai_mai_n1062_), .Y(mai_mai_n1063_));
  NO2        m1041(.A(mai_mai_n1063_), .B(mai_mai_n1061_), .Y(mai_mai_n1064_));
  NA2        m1042(.A(mai_mai_n161_), .B(mai_mai_n88_), .Y(mai_mai_n1065_));
  NO2        m1043(.A(mai_mai_n1065_), .B(i_11_), .Y(mai_mai_n1066_));
  NO4        m1044(.A(mai_mai_n962_), .B(mai_mai_n496_), .C(mai_mai_n256_), .D(mai_mai_n255_), .Y(mai_mai_n1067_));
  NO2        m1045(.A(mai_mai_n1067_), .B(mai_mai_n585_), .Y(mai_mai_n1068_));
  INV        m1046(.A(mai_mai_n373_), .Y(mai_mai_n1069_));
  AOI210     m1047(.A0(mai_mai_n1069_), .A1(mai_mai_n1068_), .B0(mai_mai_n41_), .Y(mai_mai_n1070_));
  NO2        m1048(.A(mai_mai_n1070_), .B(mai_mai_n1066_), .Y(mai_mai_n1071_));
  OAI210     m1049(.A0(mai_mai_n1064_), .A1(i_4_), .B0(mai_mai_n1071_), .Y(mai_mai_n1072_));
  NO3        m1050(.A(mai_mai_n1072_), .B(mai_mai_n1058_), .C(mai_mai_n1056_), .Y(mai_mai_n1073_));
  NA4        m1051(.A(mai_mai_n1073_), .B(mai_mai_n1038_), .C(mai_mai_n969_), .D(mai_mai_n895_), .Y(mai4));
  INV        m1052(.A(mai_mai_n721_), .Y(mai_mai_n1077_));
  INV        m1053(.A(i_2_), .Y(mai_mai_n1078_));
  INV        m1054(.A(mai_mai_n249_), .Y(mai_mai_n1079_));
  INV        m1055(.A(mai_mai_n1013_), .Y(mai_mai_n1080_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u0033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  NA2        u0034(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n57_));
  NA3        u0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n58_));
  NO2        u0036(.A(i_1_), .B(i_6_), .Y(men_men_n59_));
  NA2        u0037(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  OAI210     u0038(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n58_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_12_), .Y(men_men_n62_));
  NAi21      u0040(.An(i_2_), .B(i_7_), .Y(men_men_n63_));
  INV        u0041(.A(i_1_), .Y(men_men_n64_));
  NA2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NA3        u0043(.A(men_men_n65_), .B(men_men_n63_), .C(men_men_n31_), .Y(men_men_n66_));
  NA2        u0044(.A(i_1_), .B(i_10_), .Y(men_men_n67_));
  NO2        u0045(.A(men_men_n67_), .B(i_6_), .Y(men_men_n68_));
  NAi31      u0046(.An(men_men_n68_), .B(men_men_n66_), .C(men_men_n62_), .Y(men_men_n69_));
  NA2        u0047(.A(men_men_n51_), .B(i_2_), .Y(men_men_n70_));
  AOI210     u0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n71_));
  NA2        u0049(.A(i_1_), .B(i_6_), .Y(men_men_n72_));
  NO2        u0050(.A(men_men_n72_), .B(men_men_n25_), .Y(men_men_n73_));
  INV        u0051(.A(i_0_), .Y(men_men_n74_));
  NAi21      u0052(.An(i_5_), .B(i_10_), .Y(men_men_n75_));
  NA2        u0053(.A(i_5_), .B(i_9_), .Y(men_men_n76_));
  AOI210     u0054(.A0(men_men_n76_), .A1(men_men_n75_), .B0(men_men_n74_), .Y(men_men_n77_));
  NO2        u0055(.A(men_men_n77_), .B(men_men_n73_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n78_), .Y(men_men_n79_));
  OAI210     u0057(.A0(men_men_n79_), .A1(men_men_n69_), .B0(i_0_), .Y(men_men_n80_));
  NA2        u0058(.A(i_12_), .B(i_5_), .Y(men_men_n81_));
  NA2        u0059(.A(i_2_), .B(i_8_), .Y(men_men_n82_));
  NO2        u0060(.A(men_men_n82_), .B(men_men_n59_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_9_), .Y(men_men_n84_));
  NO2        u0062(.A(i_3_), .B(i_7_), .Y(men_men_n85_));
  NO3        u0063(.A(men_men_n85_), .B(men_men_n84_), .C(men_men_n64_), .Y(men_men_n86_));
  INV        u0064(.A(i_6_), .Y(men_men_n87_));
  OR4        u0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n88_));
  INV        u0066(.A(men_men_n88_), .Y(men_men_n89_));
  NO2        u0067(.A(i_2_), .B(i_7_), .Y(men_men_n90_));
  NO2        u0068(.A(men_men_n89_), .B(men_men_n90_), .Y(men_men_n91_));
  OAI210     u0069(.A0(men_men_n86_), .A1(men_men_n83_), .B0(men_men_n91_), .Y(men_men_n92_));
  NAi21      u0070(.An(i_6_), .B(i_10_), .Y(men_men_n93_));
  NA2        u0071(.A(i_6_), .B(i_9_), .Y(men_men_n94_));
  AOI210     u0072(.A0(men_men_n94_), .A1(men_men_n93_), .B0(men_men_n64_), .Y(men_men_n95_));
  NA2        u0073(.A(i_2_), .B(i_6_), .Y(men_men_n96_));
  NO3        u0074(.A(men_men_n96_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n97_));
  NO2        u0075(.A(men_men_n97_), .B(men_men_n95_), .Y(men_men_n98_));
  AOI210     u0076(.A0(men_men_n98_), .A1(men_men_n92_), .B0(men_men_n81_), .Y(men_men_n99_));
  AN3        u0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n100_));
  NAi21      u0078(.An(i_6_), .B(i_11_), .Y(men_men_n101_));
  NO2        u0079(.A(i_5_), .B(i_8_), .Y(men_men_n102_));
  NOi21      u0080(.An(men_men_n102_), .B(men_men_n101_), .Y(men_men_n103_));
  AOI220     u0081(.A0(men_men_n103_), .A1(men_men_n63_), .B0(men_men_n100_), .B1(men_men_n32_), .Y(men_men_n104_));
  INV        u0082(.A(i_7_), .Y(men_men_n105_));
  NA2        u0083(.A(men_men_n47_), .B(men_men_n105_), .Y(men_men_n106_));
  NO2        u0084(.A(i_0_), .B(i_5_), .Y(men_men_n107_));
  NO2        u0085(.A(men_men_n107_), .B(men_men_n87_), .Y(men_men_n108_));
  NA2        u0086(.A(i_12_), .B(i_3_), .Y(men_men_n109_));
  INV        u0087(.A(men_men_n109_), .Y(men_men_n110_));
  NA3        u0088(.A(men_men_n110_), .B(men_men_n108_), .C(men_men_n106_), .Y(men_men_n111_));
  NAi21      u0089(.An(i_7_), .B(i_11_), .Y(men_men_n112_));
  AN2        u0090(.A(i_2_), .B(i_10_), .Y(men_men_n113_));
  NO2        u0091(.A(men_men_n113_), .B(i_7_), .Y(men_men_n114_));
  OR2        u0092(.A(men_men_n81_), .B(men_men_n59_), .Y(men_men_n115_));
  NO2        u0093(.A(i_8_), .B(men_men_n105_), .Y(men_men_n116_));
  NO3        u0094(.A(men_men_n116_), .B(men_men_n115_), .C(men_men_n114_), .Y(men_men_n117_));
  NA2        u0095(.A(i_12_), .B(i_7_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n64_), .B(men_men_n26_), .Y(men_men_n119_));
  NA2        u0097(.A(i_11_), .B(i_12_), .Y(men_men_n120_));
  INV        u0098(.A(men_men_n120_), .Y(men_men_n121_));
  NO2        u0099(.A(men_men_n121_), .B(men_men_n117_), .Y(men_men_n122_));
  NA3        u0100(.A(men_men_n122_), .B(men_men_n111_), .C(men_men_n104_), .Y(men_men_n123_));
  NOi21      u0101(.An(i_1_), .B(i_5_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(i_11_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n105_), .B(men_men_n37_), .Y(men_men_n126_));
  NA2        u0104(.A(i_7_), .B(men_men_n25_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO2        u0106(.A(men_men_n128_), .B(men_men_n47_), .Y(men_men_n129_));
  NA2        u0107(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n130_));
  NAi21      u0108(.An(i_3_), .B(i_8_), .Y(men_men_n131_));
  NA2        u0109(.A(men_men_n131_), .B(men_men_n63_), .Y(men_men_n132_));
  NOi31      u0110(.An(men_men_n132_), .B(men_men_n130_), .C(men_men_n129_), .Y(men_men_n133_));
  NO2        u0111(.A(i_1_), .B(men_men_n87_), .Y(men_men_n134_));
  NO2        u0112(.A(i_6_), .B(i_5_), .Y(men_men_n135_));
  NA2        u0113(.A(men_men_n135_), .B(i_3_), .Y(men_men_n136_));
  AO210      u0114(.A0(men_men_n136_), .A1(men_men_n48_), .B0(men_men_n134_), .Y(men_men_n137_));
  OAI220     u0115(.A0(men_men_n137_), .A1(men_men_n112_), .B0(men_men_n133_), .B1(men_men_n125_), .Y(men_men_n138_));
  NO3        u0116(.A(men_men_n138_), .B(men_men_n123_), .C(men_men_n99_), .Y(men_men_n139_));
  NA3        u0117(.A(men_men_n139_), .B(men_men_n80_), .C(men_men_n57_), .Y(men2));
  NO2        u0118(.A(men_men_n64_), .B(men_men_n37_), .Y(men_men_n141_));
  NA2        u0119(.A(i_6_), .B(men_men_n25_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(men_men_n141_), .Y(men_men_n143_));
  NA4        u0121(.A(men_men_n143_), .B(men_men_n78_), .C(men_men_n70_), .D(men_men_n30_), .Y(men0));
  AN2        u0122(.A(i_8_), .B(i_7_), .Y(men_men_n145_));
  NA2        u0123(.A(men_men_n145_), .B(i_6_), .Y(men_men_n146_));
  NO2        u0124(.A(i_12_), .B(i_13_), .Y(men_men_n147_));
  NAi21      u0125(.An(i_5_), .B(i_11_), .Y(men_men_n148_));
  NOi21      u0126(.An(men_men_n147_), .B(men_men_n148_), .Y(men_men_n149_));
  NO2        u0127(.A(i_0_), .B(i_1_), .Y(men_men_n150_));
  NA2        u0128(.A(i_2_), .B(i_3_), .Y(men_men_n151_));
  NO2        u0129(.A(men_men_n151_), .B(i_4_), .Y(men_men_n152_));
  NA3        u0130(.A(men_men_n152_), .B(men_men_n150_), .C(men_men_n149_), .Y(men_men_n153_));
  OR2        u0131(.A(men_men_n153_), .B(men_men_n25_), .Y(men_men_n154_));
  AN2        u0132(.A(men_men_n147_), .B(men_men_n84_), .Y(men_men_n155_));
  NO2        u0133(.A(men_men_n155_), .B(men_men_n27_), .Y(men_men_n156_));
  NA2        u0134(.A(i_1_), .B(i_5_), .Y(men_men_n157_));
  NO2        u0135(.A(men_men_n74_), .B(men_men_n47_), .Y(men_men_n158_));
  NA2        u0136(.A(men_men_n158_), .B(men_men_n36_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n159_), .B(men_men_n157_), .C(men_men_n156_), .Y(men_men_n160_));
  OR2        u0138(.A(i_0_), .B(i_1_), .Y(men_men_n161_));
  NO3        u0139(.A(men_men_n161_), .B(men_men_n81_), .C(i_13_), .Y(men_men_n162_));
  NAi32      u0140(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n163_));
  NAi21      u0141(.An(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0142(.An(i_4_), .B(i_10_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n40_), .Y(men_men_n166_));
  NO2        u0144(.A(i_3_), .B(i_5_), .Y(men_men_n167_));
  NO3        u0145(.A(men_men_n74_), .B(i_2_), .C(i_1_), .Y(men_men_n168_));
  NA2        u0146(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  OAI210     u0147(.A0(men_men_n169_), .A1(men_men_n166_), .B0(men_men_n164_), .Y(men_men_n170_));
  NO2        u0148(.A(men_men_n170_), .B(men_men_n160_), .Y(men_men_n171_));
  AOI210     u0149(.A0(men_men_n171_), .A1(men_men_n154_), .B0(men_men_n146_), .Y(men_men_n172_));
  NA3        u0150(.A(men_men_n74_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n173_));
  NA2        u0151(.A(i_3_), .B(men_men_n49_), .Y(men_men_n174_));
  NOi21      u0152(.An(i_4_), .B(i_9_), .Y(men_men_n175_));
  NOi21      u0153(.An(i_11_), .B(i_13_), .Y(men_men_n176_));
  NA2        u0154(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OR2        u0155(.A(men_men_n177_), .B(men_men_n174_), .Y(men_men_n178_));
  NO2        u0156(.A(i_4_), .B(i_5_), .Y(men_men_n179_));
  NAi21      u0157(.An(i_12_), .B(i_11_), .Y(men_men_n180_));
  NO2        u0158(.A(men_men_n180_), .B(i_13_), .Y(men_men_n181_));
  NA3        u0159(.A(men_men_n181_), .B(men_men_n179_), .C(men_men_n84_), .Y(men_men_n182_));
  AOI210     u0160(.A0(men_men_n182_), .A1(men_men_n178_), .B0(men_men_n173_), .Y(men_men_n183_));
  NO2        u0161(.A(men_men_n74_), .B(men_men_n64_), .Y(men_men_n184_));
  NA2        u0162(.A(men_men_n184_), .B(men_men_n47_), .Y(men_men_n185_));
  NA2        u0163(.A(men_men_n36_), .B(i_5_), .Y(men_men_n186_));
  NAi31      u0164(.An(men_men_n186_), .B(men_men_n155_), .C(i_11_), .Y(men_men_n187_));
  NA2        u0165(.A(i_3_), .B(i_5_), .Y(men_men_n188_));
  OR2        u0166(.A(men_men_n188_), .B(men_men_n177_), .Y(men_men_n189_));
  AOI210     u0167(.A0(men_men_n189_), .A1(men_men_n187_), .B0(men_men_n185_), .Y(men_men_n190_));
  NO2        u0168(.A(men_men_n74_), .B(i_5_), .Y(men_men_n191_));
  NO2        u0169(.A(i_13_), .B(i_10_), .Y(men_men_n192_));
  NA3        u0170(.A(men_men_n192_), .B(men_men_n191_), .C(men_men_n45_), .Y(men_men_n193_));
  NO2        u0171(.A(i_2_), .B(i_1_), .Y(men_men_n194_));
  NA2        u0172(.A(men_men_n194_), .B(i_3_), .Y(men_men_n195_));
  NAi21      u0173(.An(i_4_), .B(i_12_), .Y(men_men_n196_));
  NO4        u0174(.A(men_men_n196_), .B(men_men_n195_), .C(men_men_n193_), .D(men_men_n25_), .Y(men_men_n197_));
  NO3        u0175(.A(men_men_n197_), .B(men_men_n190_), .C(men_men_n183_), .Y(men_men_n198_));
  INV        u0176(.A(i_8_), .Y(men_men_n199_));
  NO2        u0177(.A(men_men_n199_), .B(i_7_), .Y(men_men_n200_));
  NA2        u0178(.A(men_men_n200_), .B(i_6_), .Y(men_men_n201_));
  NO3        u0179(.A(i_3_), .B(men_men_n87_), .C(men_men_n49_), .Y(men_men_n202_));
  NA2        u0180(.A(men_men_n202_), .B(men_men_n116_), .Y(men_men_n203_));
  NO3        u0181(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n204_));
  NA3        u0182(.A(men_men_n204_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n205_));
  NO3        u0183(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n206_));
  OAI210     u0184(.A0(men_men_n100_), .A1(i_12_), .B0(men_men_n206_), .Y(men_men_n207_));
  AOI210     u0185(.A0(men_men_n207_), .A1(men_men_n205_), .B0(men_men_n203_), .Y(men_men_n208_));
  NO2        u0186(.A(i_3_), .B(i_8_), .Y(men_men_n209_));
  NO3        u0187(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n210_));
  NA3        u0188(.A(men_men_n210_), .B(men_men_n209_), .C(men_men_n40_), .Y(men_men_n211_));
  NO2        u0189(.A(men_men_n107_), .B(men_men_n59_), .Y(men_men_n212_));
  INV        u0190(.A(men_men_n212_), .Y(men_men_n213_));
  NO2        u0191(.A(i_13_), .B(i_9_), .Y(men_men_n214_));
  NA3        u0192(.A(men_men_n214_), .B(i_6_), .C(men_men_n199_), .Y(men_men_n215_));
  NAi21      u0193(.An(i_12_), .B(i_3_), .Y(men_men_n216_));
  OR2        u0194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n45_), .B(i_5_), .Y(men_men_n218_));
  NO3        u0196(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n219_));
  NA3        u0197(.A(men_men_n219_), .B(men_men_n218_), .C(i_10_), .Y(men_men_n220_));
  OAI220     u0198(.A0(men_men_n220_), .A1(men_men_n217_), .B0(men_men_n213_), .B1(men_men_n211_), .Y(men_men_n221_));
  AOI210     u0199(.A0(men_men_n221_), .A1(i_7_), .B0(men_men_n208_), .Y(men_men_n222_));
  OAI220     u0200(.A0(men_men_n222_), .A1(i_4_), .B0(men_men_n201_), .B1(men_men_n198_), .Y(men_men_n223_));
  NAi21      u0201(.An(i_12_), .B(i_7_), .Y(men_men_n224_));
  NA3        u0202(.A(i_13_), .B(men_men_n199_), .C(i_10_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NA2        u0204(.A(i_0_), .B(i_5_), .Y(men_men_n227_));
  NA2        u0205(.A(men_men_n227_), .B(men_men_n108_), .Y(men_men_n228_));
  OAI220     u0206(.A0(men_men_n228_), .A1(men_men_n195_), .B0(men_men_n185_), .B1(men_men_n136_), .Y(men_men_n229_));
  NAi31      u0207(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n36_), .B(i_13_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n74_), .B(men_men_n26_), .Y(men_men_n232_));
  NO2        u0210(.A(men_men_n47_), .B(men_men_n64_), .Y(men_men_n233_));
  NA3        u0211(.A(men_men_n233_), .B(men_men_n232_), .C(men_men_n231_), .Y(men_men_n234_));
  INV        u0212(.A(i_13_), .Y(men_men_n235_));
  NO2        u0213(.A(i_12_), .B(men_men_n235_), .Y(men_men_n236_));
  NA3        u0214(.A(men_men_n236_), .B(men_men_n204_), .C(men_men_n202_), .Y(men_men_n237_));
  OAI210     u0215(.A0(men_men_n234_), .A1(men_men_n230_), .B0(men_men_n237_), .Y(men_men_n238_));
  AOI220     u0216(.A0(men_men_n238_), .A1(men_men_n145_), .B0(men_men_n229_), .B1(men_men_n226_), .Y(men_men_n239_));
  NO2        u0217(.A(i_12_), .B(men_men_n37_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n188_), .B(i_4_), .Y(men_men_n241_));
  NA2        u0219(.A(men_men_n241_), .B(men_men_n240_), .Y(men_men_n242_));
  OR2        u0220(.A(i_8_), .B(i_7_), .Y(men_men_n243_));
  NO2        u0221(.A(men_men_n243_), .B(men_men_n87_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n54_), .B(i_1_), .Y(men_men_n245_));
  NA2        u0223(.A(men_men_n245_), .B(men_men_n244_), .Y(men_men_n246_));
  INV        u0224(.A(i_12_), .Y(men_men_n247_));
  NO2        u0225(.A(men_men_n45_), .B(men_men_n247_), .Y(men_men_n248_));
  NO3        u0226(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n249_));
  NA2        u0227(.A(i_2_), .B(i_1_), .Y(men_men_n250_));
  NO2        u0228(.A(men_men_n246_), .B(men_men_n242_), .Y(men_men_n251_));
  NO3        u0229(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n252_));
  NAi21      u0230(.An(i_4_), .B(i_3_), .Y(men_men_n253_));
  NO2        u0231(.A(men_men_n253_), .B(men_men_n76_), .Y(men_men_n254_));
  NO2        u0232(.A(i_0_), .B(i_6_), .Y(men_men_n255_));
  NOi41      u0233(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n256_));
  NA2        u0234(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  NO2        u0235(.A(men_men_n250_), .B(men_men_n188_), .Y(men_men_n258_));
  NAi21      u0236(.An(men_men_n257_), .B(men_men_n258_), .Y(men_men_n259_));
  INV        u0237(.A(men_men_n259_), .Y(men_men_n260_));
  AOI220     u0238(.A0(men_men_n260_), .A1(men_men_n40_), .B0(men_men_n251_), .B1(men_men_n214_), .Y(men_men_n261_));
  NO2        u0239(.A(i_11_), .B(men_men_n235_), .Y(men_men_n262_));
  NOi21      u0240(.An(i_1_), .B(i_6_), .Y(men_men_n263_));
  NAi21      u0241(.An(i_3_), .B(i_7_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n247_), .B(i_9_), .Y(men_men_n265_));
  OR4        u0243(.A(men_men_n265_), .B(men_men_n264_), .C(men_men_n263_), .D(men_men_n191_), .Y(men_men_n266_));
  NO2        u0244(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n267_));
  NO2        u0245(.A(i_12_), .B(i_3_), .Y(men_men_n268_));
  NA2        u0246(.A(men_men_n74_), .B(i_5_), .Y(men_men_n269_));
  NA2        u0247(.A(i_3_), .B(i_9_), .Y(men_men_n270_));
  NAi21      u0248(.An(i_7_), .B(i_10_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n271_), .B(men_men_n270_), .Y(men_men_n272_));
  NA3        u0250(.A(men_men_n272_), .B(men_men_n269_), .C(men_men_n65_), .Y(men_men_n273_));
  NA2        u0251(.A(men_men_n273_), .B(men_men_n266_), .Y(men_men_n274_));
  NA3        u0252(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n275_));
  INV        u0253(.A(men_men_n146_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n247_), .B(i_13_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n277_), .B(men_men_n76_), .Y(men_men_n278_));
  AOI220     u0256(.A0(men_men_n278_), .A1(men_men_n276_), .B0(men_men_n274_), .B1(men_men_n262_), .Y(men_men_n279_));
  NO2        u0257(.A(men_men_n243_), .B(men_men_n37_), .Y(men_men_n280_));
  NA2        u0258(.A(i_12_), .B(i_6_), .Y(men_men_n281_));
  OR2        u0259(.A(i_13_), .B(i_9_), .Y(men_men_n282_));
  NO3        u0260(.A(men_men_n282_), .B(men_men_n281_), .C(men_men_n49_), .Y(men_men_n283_));
  NO2        u0261(.A(men_men_n253_), .B(i_2_), .Y(men_men_n284_));
  NA3        u0262(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n45_), .Y(men_men_n285_));
  NA2        u0263(.A(men_men_n262_), .B(i_9_), .Y(men_men_n286_));
  NA2        u0264(.A(men_men_n269_), .B(men_men_n65_), .Y(men_men_n287_));
  OAI210     u0265(.A0(men_men_n287_), .A1(men_men_n286_), .B0(men_men_n285_), .Y(men_men_n288_));
  NA2        u0266(.A(men_men_n158_), .B(men_men_n64_), .Y(men_men_n289_));
  NO3        u0267(.A(i_11_), .B(men_men_n235_), .C(men_men_n25_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n264_), .B(i_8_), .Y(men_men_n291_));
  NO2        u0269(.A(i_6_), .B(men_men_n49_), .Y(men_men_n292_));
  NA3        u0270(.A(men_men_n292_), .B(men_men_n291_), .C(men_men_n290_), .Y(men_men_n293_));
  NO3        u0271(.A(men_men_n26_), .B(men_men_n87_), .C(i_5_), .Y(men_men_n294_));
  NA3        u0272(.A(men_men_n294_), .B(men_men_n280_), .C(men_men_n236_), .Y(men_men_n295_));
  AOI210     u0273(.A0(men_men_n295_), .A1(men_men_n293_), .B0(men_men_n289_), .Y(men_men_n296_));
  AOI210     u0274(.A0(men_men_n288_), .A1(men_men_n280_), .B0(men_men_n296_), .Y(men_men_n297_));
  NA4        u0275(.A(men_men_n297_), .B(men_men_n279_), .C(men_men_n261_), .D(men_men_n239_), .Y(men_men_n298_));
  NO3        u0276(.A(i_12_), .B(men_men_n235_), .C(men_men_n37_), .Y(men_men_n299_));
  INV        u0277(.A(men_men_n299_), .Y(men_men_n300_));
  NA2        u0278(.A(i_8_), .B(men_men_n105_), .Y(men_men_n301_));
  NOi21      u0279(.An(men_men_n167_), .B(men_men_n87_), .Y(men_men_n302_));
  NO3        u0280(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n303_));
  AOI220     u0281(.A0(men_men_n303_), .A1(men_men_n202_), .B0(men_men_n302_), .B1(men_men_n245_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n304_), .B(men_men_n301_), .Y(men_men_n305_));
  NO3        u0283(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n306_));
  NO2        u0284(.A(men_men_n250_), .B(i_0_), .Y(men_men_n307_));
  AOI220     u0285(.A0(men_men_n307_), .A1(men_men_n200_), .B0(men_men_n306_), .B1(men_men_n145_), .Y(men_men_n308_));
  NA2        u0286(.A(men_men_n292_), .B(men_men_n26_), .Y(men_men_n309_));
  NO2        u0287(.A(men_men_n309_), .B(men_men_n308_), .Y(men_men_n310_));
  NA2        u0288(.A(i_0_), .B(i_1_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n311_), .B(i_2_), .Y(men_men_n312_));
  NO2        u0290(.A(men_men_n60_), .B(i_6_), .Y(men_men_n313_));
  NA3        u0291(.A(men_men_n313_), .B(men_men_n312_), .C(men_men_n167_), .Y(men_men_n314_));
  OAI210     u0292(.A0(men_men_n169_), .A1(men_men_n146_), .B0(men_men_n314_), .Y(men_men_n315_));
  NO3        u0293(.A(men_men_n315_), .B(men_men_n310_), .C(men_men_n305_), .Y(men_men_n316_));
  NO2        u0294(.A(i_3_), .B(i_10_), .Y(men_men_n317_));
  NA3        u0295(.A(men_men_n317_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n318_));
  NO2        u0296(.A(i_2_), .B(men_men_n105_), .Y(men_men_n319_));
  NA2        u0297(.A(i_1_), .B(men_men_n36_), .Y(men_men_n320_));
  NO2        u0298(.A(men_men_n320_), .B(i_8_), .Y(men_men_n321_));
  NOi21      u0299(.An(men_men_n227_), .B(men_men_n107_), .Y(men_men_n322_));
  NA3        u0300(.A(men_men_n322_), .B(men_men_n321_), .C(men_men_n319_), .Y(men_men_n323_));
  AN2        u0301(.A(i_3_), .B(i_10_), .Y(men_men_n324_));
  NA4        u0302(.A(men_men_n324_), .B(men_men_n204_), .C(men_men_n181_), .D(men_men_n179_), .Y(men_men_n325_));
  NO2        u0303(.A(i_5_), .B(men_men_n37_), .Y(men_men_n326_));
  NO2        u0304(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n327_));
  OR2        u0305(.A(men_men_n323_), .B(men_men_n318_), .Y(men_men_n328_));
  OAI220     u0306(.A0(men_men_n328_), .A1(i_6_), .B0(men_men_n316_), .B1(men_men_n300_), .Y(men_men_n329_));
  NO4        u0307(.A(men_men_n329_), .B(men_men_n298_), .C(men_men_n223_), .D(men_men_n172_), .Y(men_men_n330_));
  NO3        u0308(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n331_));
  NO2        u0309(.A(men_men_n60_), .B(men_men_n87_), .Y(men_men_n332_));
  NA2        u0310(.A(men_men_n307_), .B(men_men_n332_), .Y(men_men_n333_));
  NO3        u0311(.A(i_6_), .B(men_men_n199_), .C(i_7_), .Y(men_men_n334_));
  NA2        u0312(.A(men_men_n334_), .B(men_men_n204_), .Y(men_men_n335_));
  AOI210     u0313(.A0(men_men_n335_), .A1(men_men_n333_), .B0(men_men_n174_), .Y(men_men_n336_));
  NO2        u0314(.A(i_2_), .B(i_3_), .Y(men_men_n337_));
  OR2        u0315(.A(i_0_), .B(i_5_), .Y(men_men_n338_));
  NA2        u0316(.A(men_men_n227_), .B(men_men_n338_), .Y(men_men_n339_));
  NA4        u0317(.A(men_men_n339_), .B(men_men_n244_), .C(men_men_n337_), .D(i_1_), .Y(men_men_n340_));
  NA3        u0318(.A(men_men_n307_), .B(men_men_n302_), .C(men_men_n116_), .Y(men_men_n341_));
  NAi21      u0319(.An(i_8_), .B(i_7_), .Y(men_men_n342_));
  NO2        u0320(.A(men_men_n342_), .B(i_6_), .Y(men_men_n343_));
  NO2        u0321(.A(men_men_n161_), .B(men_men_n47_), .Y(men_men_n344_));
  NA3        u0322(.A(men_men_n344_), .B(men_men_n343_), .C(men_men_n167_), .Y(men_men_n345_));
  NA3        u0323(.A(men_men_n345_), .B(men_men_n341_), .C(men_men_n340_), .Y(men_men_n346_));
  OAI210     u0324(.A0(men_men_n346_), .A1(men_men_n336_), .B0(i_4_), .Y(men_men_n347_));
  NO2        u0325(.A(i_12_), .B(i_10_), .Y(men_men_n348_));
  NOi21      u0326(.An(i_5_), .B(i_0_), .Y(men_men_n349_));
  NO3        u0327(.A(men_men_n320_), .B(men_men_n349_), .C(men_men_n131_), .Y(men_men_n350_));
  NA4        u0328(.A(men_men_n85_), .B(men_men_n36_), .C(men_men_n87_), .D(i_8_), .Y(men_men_n351_));
  NA2        u0329(.A(men_men_n350_), .B(men_men_n348_), .Y(men_men_n352_));
  NO2        u0330(.A(i_6_), .B(i_8_), .Y(men_men_n353_));
  NOi21      u0331(.An(i_0_), .B(i_2_), .Y(men_men_n354_));
  AN2        u0332(.A(men_men_n354_), .B(men_men_n353_), .Y(men_men_n355_));
  NO2        u0333(.A(i_1_), .B(i_7_), .Y(men_men_n356_));
  AO220      u0334(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n343_), .B1(men_men_n245_), .Y(men_men_n357_));
  NA3        u0335(.A(men_men_n357_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n358_));
  NA3        u0336(.A(men_men_n358_), .B(men_men_n352_), .C(men_men_n347_), .Y(men_men_n359_));
  NO3        u0337(.A(men_men_n243_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n360_));
  NO3        u0338(.A(men_men_n342_), .B(i_2_), .C(i_1_), .Y(men_men_n361_));
  OAI210     u0339(.A0(men_men_n361_), .A1(men_men_n360_), .B0(i_6_), .Y(men_men_n362_));
  NA3        u0340(.A(men_men_n263_), .B(men_men_n319_), .C(men_men_n199_), .Y(men_men_n363_));
  AOI210     u0341(.A0(men_men_n363_), .A1(men_men_n362_), .B0(men_men_n339_), .Y(men_men_n364_));
  NOi21      u0342(.An(men_men_n157_), .B(men_men_n108_), .Y(men_men_n365_));
  NA2        u0343(.A(men_men_n364_), .B(i_3_), .Y(men_men_n366_));
  INV        u0344(.A(men_men_n85_), .Y(men_men_n367_));
  NO2        u0345(.A(men_men_n311_), .B(men_men_n82_), .Y(men_men_n368_));
  NA2        u0346(.A(men_men_n368_), .B(men_men_n135_), .Y(men_men_n369_));
  NO2        u0347(.A(men_men_n96_), .B(men_men_n199_), .Y(men_men_n370_));
  NA3        u0348(.A(men_men_n322_), .B(men_men_n370_), .C(men_men_n64_), .Y(men_men_n371_));
  AOI210     u0349(.A0(men_men_n371_), .A1(men_men_n369_), .B0(men_men_n367_), .Y(men_men_n372_));
  NO2        u0350(.A(men_men_n199_), .B(i_9_), .Y(men_men_n373_));
  NA2        u0351(.A(men_men_n373_), .B(men_men_n212_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n372_), .B(men_men_n310_), .Y(men_men_n375_));
  AOI210     u0353(.A0(men_men_n375_), .A1(men_men_n366_), .B0(men_men_n166_), .Y(men_men_n376_));
  AOI210     u0354(.A0(men_men_n359_), .A1(men_men_n331_), .B0(men_men_n376_), .Y(men_men_n377_));
  NOi32      u0355(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n378_));
  INV        u0356(.A(men_men_n378_), .Y(men_men_n379_));
  NAi21      u0357(.An(i_0_), .B(i_6_), .Y(men_men_n380_));
  NAi21      u0358(.An(i_1_), .B(i_5_), .Y(men_men_n381_));
  NA2        u0359(.A(men_men_n381_), .B(men_men_n380_), .Y(men_men_n382_));
  NA2        u0360(.A(men_men_n382_), .B(men_men_n25_), .Y(men_men_n383_));
  OAI210     u0361(.A0(men_men_n383_), .A1(men_men_n163_), .B0(men_men_n257_), .Y(men_men_n384_));
  NAi41      u0362(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n385_));
  AOI210     u0363(.A0(men_men_n385_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n386_));
  NOi32      u0364(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n387_));
  NO2        u0365(.A(i_1_), .B(men_men_n105_), .Y(men_men_n388_));
  NAi21      u0366(.An(i_3_), .B(i_4_), .Y(men_men_n389_));
  NO2        u0367(.A(men_men_n389_), .B(i_9_), .Y(men_men_n390_));
  AN2        u0368(.A(i_6_), .B(i_7_), .Y(men_men_n391_));
  OAI210     u0369(.A0(men_men_n391_), .A1(men_men_n388_), .B0(men_men_n390_), .Y(men_men_n392_));
  NA2        u0370(.A(i_2_), .B(i_7_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n389_), .B(i_10_), .Y(men_men_n394_));
  NA3        u0372(.A(men_men_n394_), .B(men_men_n393_), .C(men_men_n255_), .Y(men_men_n395_));
  AOI210     u0373(.A0(men_men_n395_), .A1(men_men_n392_), .B0(men_men_n191_), .Y(men_men_n396_));
  AOI210     u0374(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n397_));
  OAI210     u0375(.A0(men_men_n397_), .A1(men_men_n194_), .B0(men_men_n394_), .Y(men_men_n398_));
  AOI220     u0376(.A0(men_men_n394_), .A1(men_men_n356_), .B0(men_men_n249_), .B1(men_men_n194_), .Y(men_men_n399_));
  AOI210     u0377(.A0(men_men_n399_), .A1(men_men_n398_), .B0(i_5_), .Y(men_men_n400_));
  NO4        u0378(.A(men_men_n400_), .B(men_men_n396_), .C(men_men_n386_), .D(men_men_n384_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n401_), .B(men_men_n379_), .Y(men_men_n402_));
  NO2        u0380(.A(men_men_n60_), .B(men_men_n25_), .Y(men_men_n403_));
  AN2        u0381(.A(i_12_), .B(i_5_), .Y(men_men_n404_));
  NO2        u0382(.A(i_4_), .B(men_men_n26_), .Y(men_men_n405_));
  NA2        u0383(.A(men_men_n405_), .B(men_men_n404_), .Y(men_men_n406_));
  NO2        u0384(.A(i_11_), .B(i_6_), .Y(men_men_n407_));
  NA3        u0385(.A(men_men_n407_), .B(men_men_n344_), .C(men_men_n235_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n408_), .B(men_men_n406_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n253_), .B(i_5_), .Y(men_men_n410_));
  NO2        u0388(.A(i_5_), .B(i_10_), .Y(men_men_n411_));
  AOI220     u0389(.A0(men_men_n411_), .A1(men_men_n284_), .B0(men_men_n410_), .B1(men_men_n204_), .Y(men_men_n412_));
  NA2        u0390(.A(men_men_n147_), .B(men_men_n46_), .Y(men_men_n413_));
  NO2        u0391(.A(men_men_n413_), .B(men_men_n412_), .Y(men_men_n414_));
  OAI210     u0392(.A0(men_men_n414_), .A1(men_men_n409_), .B0(men_men_n403_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n153_), .B(men_men_n87_), .Y(men_men_n417_));
  OAI210     u0395(.A0(men_men_n417_), .A1(men_men_n409_), .B0(men_men_n416_), .Y(men_men_n418_));
  NO3        u0396(.A(men_men_n87_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n419_));
  NO2        u0397(.A(i_11_), .B(i_12_), .Y(men_men_n420_));
  NA2        u0398(.A(men_men_n411_), .B(men_men_n247_), .Y(men_men_n421_));
  NA3        u0399(.A(men_men_n116_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n422_));
  OAI220     u0400(.A0(men_men_n422_), .A1(men_men_n230_), .B0(men_men_n421_), .B1(men_men_n351_), .Y(men_men_n423_));
  NAi21      u0401(.An(i_13_), .B(i_0_), .Y(men_men_n424_));
  NO2        u0402(.A(men_men_n424_), .B(men_men_n250_), .Y(men_men_n425_));
  NA2        u0403(.A(men_men_n423_), .B(men_men_n425_), .Y(men_men_n426_));
  NA3        u0404(.A(men_men_n426_), .B(men_men_n418_), .C(men_men_n415_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n45_), .B(men_men_n235_), .Y(men_men_n428_));
  NO3        u0406(.A(i_1_), .B(i_12_), .C(men_men_n87_), .Y(men_men_n429_));
  NO2        u0407(.A(i_0_), .B(i_11_), .Y(men_men_n430_));
  INV        u0408(.A(i_5_), .Y(men_men_n431_));
  AN2        u0409(.A(i_1_), .B(i_6_), .Y(men_men_n432_));
  NOi21      u0410(.An(i_2_), .B(i_12_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n433_), .B(men_men_n432_), .Y(men_men_n434_));
  NO2        u0412(.A(men_men_n434_), .B(men_men_n431_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n145_), .B(i_9_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(i_4_), .Y(men_men_n437_));
  NA2        u0415(.A(men_men_n435_), .B(men_men_n437_), .Y(men_men_n438_));
  NAi21      u0416(.An(i_9_), .B(i_4_), .Y(men_men_n439_));
  OR2        u0417(.A(i_13_), .B(i_10_), .Y(men_men_n440_));
  NO3        u0418(.A(men_men_n440_), .B(men_men_n120_), .C(men_men_n439_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n177_), .B(men_men_n126_), .Y(men_men_n442_));
  OR2        u0420(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n443_));
  NO2        u0421(.A(men_men_n105_), .B(men_men_n25_), .Y(men_men_n444_));
  NA2        u0422(.A(men_men_n299_), .B(men_men_n444_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n292_), .B(men_men_n219_), .Y(men_men_n446_));
  OAI220     u0424(.A0(men_men_n446_), .A1(men_men_n443_), .B0(men_men_n445_), .B1(men_men_n365_), .Y(men_men_n447_));
  INV        u0425(.A(men_men_n447_), .Y(men_men_n448_));
  AOI210     u0426(.A0(men_men_n448_), .A1(men_men_n438_), .B0(men_men_n26_), .Y(men_men_n449_));
  NA2        u0427(.A(men_men_n341_), .B(men_men_n340_), .Y(men_men_n450_));
  AOI220     u0428(.A0(men_men_n313_), .A1(men_men_n303_), .B0(men_men_n307_), .B1(men_men_n332_), .Y(men_men_n451_));
  NO2        u0429(.A(men_men_n451_), .B(men_men_n174_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n188_), .B(men_men_n87_), .Y(men_men_n453_));
  AOI220     u0431(.A0(men_men_n453_), .A1(men_men_n312_), .B0(men_men_n294_), .B1(men_men_n219_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n454_), .B(men_men_n301_), .Y(men_men_n455_));
  NO3        u0433(.A(men_men_n455_), .B(men_men_n452_), .C(men_men_n450_), .Y(men_men_n456_));
  NA2        u0434(.A(men_men_n202_), .B(men_men_n100_), .Y(men_men_n457_));
  NA3        u0435(.A(men_men_n344_), .B(men_men_n167_), .C(men_men_n87_), .Y(men_men_n458_));
  AOI210     u0436(.A0(men_men_n458_), .A1(men_men_n457_), .B0(men_men_n342_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n313_), .B(men_men_n245_), .Y(men_men_n460_));
  NO2        u0438(.A(men_men_n460_), .B(men_men_n188_), .Y(men_men_n461_));
  NO2        u0439(.A(i_3_), .B(men_men_n49_), .Y(men_men_n462_));
  NA3        u0440(.A(men_men_n356_), .B(men_men_n355_), .C(men_men_n462_), .Y(men_men_n463_));
  NA2        u0441(.A(men_men_n334_), .B(men_men_n339_), .Y(men_men_n464_));
  OAI210     u0442(.A0(men_men_n464_), .A1(men_men_n195_), .B0(men_men_n463_), .Y(men_men_n465_));
  NO3        u0443(.A(men_men_n465_), .B(men_men_n461_), .C(men_men_n459_), .Y(men_men_n466_));
  AOI210     u0444(.A0(men_men_n466_), .A1(men_men_n456_), .B0(men_men_n286_), .Y(men_men_n467_));
  NO4        u0445(.A(men_men_n467_), .B(men_men_n449_), .C(men_men_n427_), .D(men_men_n402_), .Y(men_men_n468_));
  NO2        u0446(.A(men_men_n64_), .B(i_4_), .Y(men_men_n469_));
  NO2        u0447(.A(men_men_n74_), .B(i_13_), .Y(men_men_n470_));
  NO2        u0448(.A(i_10_), .B(i_9_), .Y(men_men_n471_));
  NAi21      u0449(.An(i_12_), .B(i_8_), .Y(men_men_n472_));
  NO2        u0450(.A(men_men_n472_), .B(i_3_), .Y(men_men_n473_));
  NO2        u0451(.A(men_men_n47_), .B(i_4_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n474_), .B(men_men_n108_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n475_), .B(men_men_n211_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n327_), .B(i_0_), .Y(men_men_n477_));
  NO3        u0455(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n281_), .B(men_men_n101_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n479_), .B(men_men_n478_), .Y(men_men_n480_));
  NA2        u0458(.A(i_8_), .B(i_9_), .Y(men_men_n481_));
  AOI210     u0459(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n482_));
  OR2        u0460(.A(men_men_n482_), .B(men_men_n481_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n299_), .B(men_men_n212_), .Y(men_men_n484_));
  OAI220     u0462(.A0(men_men_n484_), .A1(men_men_n483_), .B0(men_men_n480_), .B1(men_men_n477_), .Y(men_men_n485_));
  NA2        u0463(.A(men_men_n262_), .B(men_men_n326_), .Y(men_men_n486_));
  NO3        u0464(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n487_));
  INV        u0465(.A(men_men_n487_), .Y(men_men_n488_));
  NA3        u0466(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n489_));
  NA4        u0467(.A(men_men_n148_), .B(men_men_n119_), .C(men_men_n81_), .D(men_men_n23_), .Y(men_men_n490_));
  OAI220     u0468(.A0(men_men_n490_), .A1(men_men_n489_), .B0(men_men_n488_), .B1(men_men_n486_), .Y(men_men_n491_));
  NO3        u0469(.A(men_men_n491_), .B(men_men_n485_), .C(men_men_n476_), .Y(men_men_n492_));
  NA2        u0470(.A(men_men_n312_), .B(men_men_n112_), .Y(men_men_n493_));
  OR2        u0471(.A(men_men_n493_), .B(men_men_n215_), .Y(men_men_n494_));
  OA210      u0472(.A0(men_men_n374_), .A1(men_men_n105_), .B0(men_men_n314_), .Y(men_men_n495_));
  OA220      u0473(.A0(men_men_n495_), .A1(men_men_n166_), .B0(men_men_n494_), .B1(men_men_n242_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n100_), .B(i_13_), .Y(men_men_n497_));
  NA2        u0475(.A(men_men_n453_), .B(men_men_n403_), .Y(men_men_n498_));
  NO2        u0476(.A(i_2_), .B(i_13_), .Y(men_men_n499_));
  NA3        u0477(.A(men_men_n499_), .B(men_men_n165_), .C(men_men_n103_), .Y(men_men_n500_));
  OAI220     u0478(.A0(men_men_n500_), .A1(men_men_n247_), .B0(men_men_n498_), .B1(men_men_n497_), .Y(men_men_n501_));
  NO3        u0479(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n502_));
  NO2        u0480(.A(i_6_), .B(i_7_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n503_), .B(men_men_n502_), .Y(men_men_n504_));
  NO2        u0482(.A(i_11_), .B(i_1_), .Y(men_men_n505_));
  NO2        u0483(.A(men_men_n74_), .B(i_3_), .Y(men_men_n506_));
  OR2        u0484(.A(i_11_), .B(i_8_), .Y(men_men_n507_));
  NOi21      u0485(.An(i_2_), .B(i_7_), .Y(men_men_n508_));
  NAi31      u0486(.An(men_men_n507_), .B(men_men_n508_), .C(men_men_n506_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n440_), .B(i_6_), .Y(men_men_n510_));
  NA3        u0488(.A(men_men_n510_), .B(men_men_n469_), .C(men_men_n76_), .Y(men_men_n511_));
  NO2        u0489(.A(men_men_n511_), .B(men_men_n509_), .Y(men_men_n512_));
  NO2        u0490(.A(i_3_), .B(men_men_n199_), .Y(men_men_n513_));
  NO2        u0491(.A(i_6_), .B(i_10_), .Y(men_men_n514_));
  NA4        u0492(.A(men_men_n514_), .B(men_men_n331_), .C(men_men_n513_), .D(men_men_n247_), .Y(men_men_n515_));
  NO2        u0493(.A(men_men_n515_), .B(men_men_n159_), .Y(men_men_n516_));
  NA3        u0494(.A(men_men_n256_), .B(men_men_n176_), .C(men_men_n135_), .Y(men_men_n517_));
  NA2        u0495(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n518_));
  NO2        u0496(.A(men_men_n161_), .B(i_3_), .Y(men_men_n519_));
  NAi31      u0497(.An(men_men_n518_), .B(men_men_n519_), .C(men_men_n236_), .Y(men_men_n520_));
  NA3        u0498(.A(men_men_n416_), .B(men_men_n184_), .C(men_men_n152_), .Y(men_men_n521_));
  NA3        u0499(.A(men_men_n521_), .B(men_men_n520_), .C(men_men_n517_), .Y(men_men_n522_));
  NO4        u0500(.A(men_men_n522_), .B(men_men_n516_), .C(men_men_n512_), .D(men_men_n501_), .Y(men_men_n523_));
  NA2        u0501(.A(men_men_n478_), .B(men_men_n404_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n487_), .B(men_men_n411_), .Y(men_men_n525_));
  NO2        u0503(.A(men_men_n525_), .B(men_men_n234_), .Y(men_men_n526_));
  NAi21      u0504(.An(men_men_n225_), .B(men_men_n420_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n356_), .B(men_men_n227_), .Y(men_men_n528_));
  NO2        u0506(.A(men_men_n26_), .B(i_5_), .Y(men_men_n529_));
  NO2        u0507(.A(i_0_), .B(men_men_n87_), .Y(men_men_n530_));
  NA3        u0508(.A(men_men_n530_), .B(men_men_n529_), .C(men_men_n145_), .Y(men_men_n531_));
  OR3        u0509(.A(men_men_n320_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n532_));
  OAI220     u0510(.A0(men_men_n532_), .A1(men_men_n531_), .B0(men_men_n528_), .B1(men_men_n527_), .Y(men_men_n533_));
  NA2        u0511(.A(men_men_n27_), .B(i_10_), .Y(men_men_n534_));
  NO2        u0512(.A(men_men_n534_), .B(men_men_n497_), .Y(men_men_n535_));
  NA4        u0513(.A(men_men_n324_), .B(men_men_n233_), .C(men_men_n74_), .D(men_men_n247_), .Y(men_men_n536_));
  NO2        u0514(.A(men_men_n536_), .B(men_men_n504_), .Y(men_men_n537_));
  NO4        u0515(.A(men_men_n537_), .B(men_men_n535_), .C(men_men_n533_), .D(men_men_n526_), .Y(men_men_n538_));
  NA4        u0516(.A(men_men_n538_), .B(men_men_n523_), .C(men_men_n496_), .D(men_men_n492_), .Y(men_men_n539_));
  NA3        u0517(.A(men_men_n324_), .B(men_men_n181_), .C(men_men_n179_), .Y(men_men_n540_));
  OAI210     u0518(.A0(men_men_n318_), .A1(men_men_n186_), .B0(men_men_n540_), .Y(men_men_n541_));
  AN2        u0519(.A(men_men_n303_), .B(men_men_n244_), .Y(men_men_n542_));
  NA2        u0520(.A(men_men_n542_), .B(men_men_n541_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n125_), .B(men_men_n115_), .Y(men_men_n544_));
  AO220      u0522(.A0(men_men_n544_), .A1(men_men_n478_), .B0(men_men_n441_), .B1(i_6_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n331_), .B(men_men_n168_), .Y(men_men_n546_));
  OAI210     u0524(.A0(men_men_n546_), .A1(men_men_n242_), .B0(men_men_n325_), .Y(men_men_n547_));
  AOI220     u0525(.A0(men_men_n547_), .A1(men_men_n343_), .B0(men_men_n545_), .B1(men_men_n327_), .Y(men_men_n548_));
  NA2        u0526(.A(men_men_n404_), .B(men_men_n235_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n378_), .B(men_men_n74_), .Y(men_men_n550_));
  NA2        u0528(.A(men_men_n391_), .B(men_men_n387_), .Y(men_men_n551_));
  AO210      u0529(.A0(men_men_n550_), .A1(men_men_n549_), .B0(men_men_n551_), .Y(men_men_n552_));
  NO2        u0530(.A(men_men_n36_), .B(i_8_), .Y(men_men_n553_));
  AOI210     u0531(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n441_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n554_), .B(men_men_n552_), .Y(men_men_n555_));
  INV        u0533(.A(men_men_n555_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n269_), .B(men_men_n65_), .Y(men_men_n557_));
  OAI210     u0535(.A0(i_8_), .A1(men_men_n557_), .B0(men_men_n137_), .Y(men_men_n558_));
  NO2        u0536(.A(i_7_), .B(men_men_n205_), .Y(men_men_n559_));
  OR2        u0537(.A(men_men_n188_), .B(i_4_), .Y(men_men_n560_));
  NO2        u0538(.A(men_men_n560_), .B(men_men_n87_), .Y(men_men_n561_));
  AOI220     u0539(.A0(men_men_n561_), .A1(men_men_n559_), .B0(men_men_n558_), .B1(men_men_n442_), .Y(men_men_n562_));
  NA4        u0540(.A(men_men_n562_), .B(men_men_n556_), .C(men_men_n548_), .D(men_men_n543_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n410_), .B(men_men_n312_), .Y(men_men_n564_));
  OAI210     u0542(.A0(men_men_n406_), .A1(men_men_n173_), .B0(men_men_n564_), .Y(men_men_n565_));
  NO2        u0543(.A(i_12_), .B(men_men_n199_), .Y(men_men_n566_));
  NA2        u0544(.A(men_men_n566_), .B(men_men_n235_), .Y(men_men_n567_));
  NO3        u0545(.A(men_men_n1112_), .B(men_men_n567_), .C(men_men_n493_), .Y(men_men_n568_));
  NOi31      u0546(.An(men_men_n334_), .B(men_men_n440_), .C(men_men_n38_), .Y(men_men_n569_));
  OAI210     u0547(.A0(men_men_n569_), .A1(men_men_n568_), .B0(men_men_n565_), .Y(men_men_n570_));
  NO2        u0548(.A(i_8_), .B(i_7_), .Y(men_men_n571_));
  OAI210     u0549(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n572_));
  NA2        u0550(.A(men_men_n572_), .B(men_men_n233_), .Y(men_men_n573_));
  AOI220     u0551(.A0(men_men_n344_), .A1(men_men_n40_), .B0(men_men_n245_), .B1(men_men_n214_), .Y(men_men_n574_));
  OAI220     u0552(.A0(men_men_n574_), .A1(men_men_n560_), .B0(men_men_n573_), .B1(men_men_n253_), .Y(men_men_n575_));
  NA2        u0553(.A(men_men_n45_), .B(i_10_), .Y(men_men_n576_));
  NO2        u0554(.A(men_men_n576_), .B(i_6_), .Y(men_men_n577_));
  NA3        u0555(.A(men_men_n577_), .B(men_men_n575_), .C(men_men_n571_), .Y(men_men_n578_));
  AOI220     u0556(.A0(men_men_n453_), .A1(men_men_n344_), .B0(men_men_n258_), .B1(men_men_n255_), .Y(men_men_n579_));
  OAI220     u0557(.A0(men_men_n579_), .A1(men_men_n277_), .B0(men_men_n497_), .B1(men_men_n136_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n580_), .B(men_men_n280_), .Y(men_men_n581_));
  NOi31      u0559(.An(men_men_n307_), .B(men_men_n318_), .C(men_men_n186_), .Y(men_men_n582_));
  NA3        u0560(.A(men_men_n324_), .B(men_men_n179_), .C(men_men_n100_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n231_), .B(men_men_n45_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n161_), .B(i_5_), .Y(men_men_n585_));
  NA3        u0563(.A(men_men_n585_), .B(men_men_n428_), .C(men_men_n337_), .Y(men_men_n586_));
  OAI210     u0564(.A0(men_men_n586_), .A1(men_men_n584_), .B0(men_men_n583_), .Y(men_men_n587_));
  OAI210     u0565(.A0(men_men_n587_), .A1(men_men_n582_), .B0(men_men_n487_), .Y(men_men_n588_));
  NA4        u0566(.A(men_men_n588_), .B(men_men_n581_), .C(men_men_n578_), .D(men_men_n570_), .Y(men_men_n589_));
  NA3        u0567(.A(men_men_n227_), .B(men_men_n72_), .C(men_men_n45_), .Y(men_men_n590_));
  NA2        u0568(.A(men_men_n299_), .B(men_men_n85_), .Y(men_men_n591_));
  AOI210     u0569(.A0(men_men_n590_), .A1(men_men_n369_), .B0(men_men_n591_), .Y(men_men_n592_));
  NA2        u0570(.A(men_men_n313_), .B(men_men_n303_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n593_), .B(men_men_n178_), .Y(men_men_n594_));
  NA2        u0572(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n595_));
  NA2        u0573(.A(men_men_n471_), .B(men_men_n231_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n595_), .B(men_men_n596_), .Y(men_men_n597_));
  AOI210     u0575(.A0(i_6_), .A1(men_men_n47_), .B0(men_men_n388_), .Y(men_men_n598_));
  NA2        u0576(.A(i_0_), .B(men_men_n49_), .Y(men_men_n599_));
  NA3        u0577(.A(men_men_n566_), .B(men_men_n290_), .C(men_men_n599_), .Y(men_men_n600_));
  NO2        u0578(.A(men_men_n598_), .B(men_men_n600_), .Y(men_men_n601_));
  NO4        u0579(.A(men_men_n601_), .B(men_men_n597_), .C(men_men_n594_), .D(men_men_n592_), .Y(men_men_n602_));
  NO4        u0580(.A(men_men_n263_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n603_));
  NO3        u0581(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n243_), .B(men_men_n36_), .Y(men_men_n605_));
  AN2        u0583(.A(men_men_n605_), .B(men_men_n604_), .Y(men_men_n606_));
  OA210      u0584(.A0(men_men_n606_), .A1(men_men_n603_), .B0(men_men_n378_), .Y(men_men_n607_));
  NO2        u0585(.A(men_men_n440_), .B(i_1_), .Y(men_men_n608_));
  NOi31      u0586(.An(men_men_n608_), .B(men_men_n479_), .C(men_men_n74_), .Y(men_men_n609_));
  AN4        u0587(.A(men_men_n609_), .B(men_men_n437_), .C(men_men_n529_), .D(i_2_), .Y(men_men_n610_));
  NO2        u0588(.A(men_men_n451_), .B(men_men_n182_), .Y(men_men_n611_));
  NO3        u0589(.A(men_men_n611_), .B(men_men_n610_), .C(men_men_n607_), .Y(men_men_n612_));
  NOi21      u0590(.An(i_10_), .B(i_6_), .Y(men_men_n613_));
  NO2        u0591(.A(men_men_n87_), .B(men_men_n25_), .Y(men_men_n614_));
  AOI220     u0592(.A0(men_men_n299_), .A1(men_men_n614_), .B0(men_men_n290_), .B1(men_men_n613_), .Y(men_men_n615_));
  NO2        u0593(.A(men_men_n615_), .B(men_men_n477_), .Y(men_men_n616_));
  NO2        u0594(.A(men_men_n118_), .B(men_men_n23_), .Y(men_men_n617_));
  NA2        u0595(.A(men_men_n334_), .B(men_men_n168_), .Y(men_men_n618_));
  AOI220     u0596(.A0(men_men_n618_), .A1(men_men_n460_), .B0(men_men_n189_), .B1(men_men_n187_), .Y(men_men_n619_));
  NO2        u0597(.A(men_men_n204_), .B(men_men_n37_), .Y(men_men_n620_));
  NOi31      u0598(.An(men_men_n149_), .B(men_men_n620_), .C(men_men_n351_), .Y(men_men_n621_));
  NO3        u0599(.A(men_men_n621_), .B(men_men_n619_), .C(men_men_n616_), .Y(men_men_n622_));
  NO2        u0600(.A(men_men_n550_), .B(men_men_n399_), .Y(men_men_n623_));
  INV        u0601(.A(men_men_n337_), .Y(men_men_n624_));
  NO2        u0602(.A(i_12_), .B(men_men_n87_), .Y(men_men_n625_));
  NA3        u0603(.A(men_men_n625_), .B(men_men_n290_), .C(men_men_n599_), .Y(men_men_n626_));
  NA3        u0604(.A(men_men_n407_), .B(men_men_n299_), .C(men_men_n227_), .Y(men_men_n627_));
  AOI210     u0605(.A0(men_men_n627_), .A1(men_men_n626_), .B0(men_men_n624_), .Y(men_men_n628_));
  NA2        u0606(.A(men_men_n179_), .B(i_0_), .Y(men_men_n629_));
  NO3        u0607(.A(men_men_n629_), .B(men_men_n362_), .C(men_men_n318_), .Y(men_men_n630_));
  OR2        u0608(.A(i_2_), .B(i_5_), .Y(men_men_n631_));
  OR2        u0609(.A(men_men_n631_), .B(men_men_n432_), .Y(men_men_n632_));
  NO2        u0610(.A(men_men_n632_), .B(men_men_n527_), .Y(men_men_n633_));
  NO4        u0611(.A(men_men_n633_), .B(men_men_n630_), .C(men_men_n628_), .D(men_men_n623_), .Y(men_men_n634_));
  NA4        u0612(.A(men_men_n634_), .B(men_men_n622_), .C(men_men_n612_), .D(men_men_n602_), .Y(men_men_n635_));
  NO4        u0613(.A(men_men_n635_), .B(men_men_n589_), .C(men_men_n563_), .D(men_men_n539_), .Y(men_men_n636_));
  NA4        u0614(.A(men_men_n636_), .B(men_men_n468_), .C(men_men_n377_), .D(men_men_n330_), .Y(men7));
  NO2        u0615(.A(men_men_n96_), .B(men_men_n55_), .Y(men_men_n638_));
  NO2        u0616(.A(men_men_n112_), .B(men_men_n93_), .Y(men_men_n639_));
  NA2        u0617(.A(men_men_n405_), .B(men_men_n639_), .Y(men_men_n640_));
  NA2        u0618(.A(men_men_n514_), .B(men_men_n85_), .Y(men_men_n641_));
  NA2        u0619(.A(i_11_), .B(men_men_n199_), .Y(men_men_n642_));
  INV        u0620(.A(men_men_n640_), .Y(men_men_n643_));
  NA3        u0621(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n644_));
  NO2        u0622(.A(men_men_n247_), .B(i_4_), .Y(men_men_n645_));
  NA2        u0623(.A(men_men_n645_), .B(i_8_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n109_), .B(men_men_n644_), .Y(men_men_n647_));
  NA2        u0625(.A(i_2_), .B(men_men_n87_), .Y(men_men_n648_));
  OAI210     u0626(.A0(men_men_n90_), .A1(men_men_n209_), .B0(men_men_n210_), .Y(men_men_n649_));
  NO2        u0627(.A(i_7_), .B(men_men_n37_), .Y(men_men_n650_));
  NA2        u0628(.A(i_4_), .B(i_8_), .Y(men_men_n651_));
  AOI210     u0629(.A0(men_men_n651_), .A1(men_men_n324_), .B0(men_men_n650_), .Y(men_men_n652_));
  OAI220     u0630(.A0(men_men_n652_), .A1(men_men_n648_), .B0(men_men_n649_), .B1(i_13_), .Y(men_men_n653_));
  NO4        u0631(.A(men_men_n653_), .B(men_men_n647_), .C(men_men_n643_), .D(men_men_n638_), .Y(men_men_n654_));
  AOI210     u0632(.A0(men_men_n131_), .A1(men_men_n63_), .B0(i_10_), .Y(men_men_n655_));
  AOI210     u0633(.A0(men_men_n655_), .A1(men_men_n247_), .B0(men_men_n165_), .Y(men_men_n656_));
  OR2        u0634(.A(i_6_), .B(i_10_), .Y(men_men_n657_));
  NO2        u0635(.A(men_men_n657_), .B(men_men_n23_), .Y(men_men_n658_));
  OR3        u0636(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n659_));
  NO3        u0637(.A(men_men_n659_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n660_));
  INV        u0638(.A(men_men_n206_), .Y(men_men_n661_));
  NO2        u0639(.A(men_men_n660_), .B(men_men_n658_), .Y(men_men_n662_));
  OA220      u0640(.A0(men_men_n662_), .A1(men_men_n624_), .B0(men_men_n656_), .B1(men_men_n282_), .Y(men_men_n663_));
  AOI210     u0641(.A0(men_men_n663_), .A1(men_men_n654_), .B0(men_men_n64_), .Y(men_men_n664_));
  NOi21      u0642(.An(i_11_), .B(i_7_), .Y(men_men_n665_));
  AO210      u0643(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n666_));
  NO2        u0644(.A(men_men_n666_), .B(men_men_n665_), .Y(men_men_n667_));
  NA2        u0645(.A(men_men_n667_), .B(men_men_n214_), .Y(men_men_n668_));
  NA3        u0646(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n669_));
  NAi31      u0647(.An(men_men_n669_), .B(men_men_n224_), .C(i_11_), .Y(men_men_n670_));
  AOI210     u0648(.A0(men_men_n670_), .A1(men_men_n668_), .B0(men_men_n64_), .Y(men_men_n671_));
  NA2        u0649(.A(men_men_n89_), .B(men_men_n64_), .Y(men_men_n672_));
  AO210      u0650(.A0(men_men_n672_), .A1(men_men_n399_), .B0(men_men_n41_), .Y(men_men_n673_));
  NO3        u0651(.A(men_men_n271_), .B(men_men_n216_), .C(men_men_n642_), .Y(men_men_n674_));
  OAI210     u0652(.A0(men_men_n674_), .A1(men_men_n236_), .B0(men_men_n64_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n433_), .B(men_men_n31_), .Y(men_men_n676_));
  OR2        u0654(.A(men_men_n216_), .B(men_men_n112_), .Y(men_men_n677_));
  NA2        u0655(.A(men_men_n677_), .B(men_men_n676_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n64_), .B(i_9_), .Y(men_men_n679_));
  NO2        u0657(.A(men_men_n679_), .B(i_4_), .Y(men_men_n680_));
  NA2        u0658(.A(men_men_n680_), .B(men_men_n678_), .Y(men_men_n681_));
  NO2        u0659(.A(i_1_), .B(i_12_), .Y(men_men_n682_));
  NA3        u0660(.A(men_men_n682_), .B(men_men_n113_), .C(men_men_n24_), .Y(men_men_n683_));
  NA4        u0661(.A(men_men_n683_), .B(men_men_n681_), .C(men_men_n675_), .D(men_men_n673_), .Y(men_men_n684_));
  OAI210     u0662(.A0(men_men_n684_), .A1(men_men_n671_), .B0(i_6_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n247_), .B(men_men_n87_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n686_), .B(i_11_), .Y(men_men_n687_));
  INV        u0665(.A(men_men_n480_), .Y(men_men_n688_));
  NO4        u0666(.A(men_men_n224_), .B(men_men_n131_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n689_));
  NA2        u0667(.A(men_men_n689_), .B(men_men_n679_), .Y(men_men_n690_));
  NA2        u0668(.A(men_men_n247_), .B(i_6_), .Y(men_men_n691_));
  NO3        u0669(.A(men_men_n657_), .B(men_men_n243_), .C(men_men_n23_), .Y(men_men_n692_));
  AOI210     u0670(.A0(i_1_), .A1(men_men_n272_), .B0(men_men_n692_), .Y(men_men_n693_));
  OAI210     u0671(.A0(men_men_n693_), .A1(men_men_n45_), .B0(men_men_n690_), .Y(men_men_n694_));
  NA3        u0672(.A(men_men_n571_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n695_));
  NA2        u0673(.A(men_men_n141_), .B(i_9_), .Y(men_men_n696_));
  NA3        u0674(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n47_), .B(i_1_), .Y(men_men_n698_));
  NO2        u0676(.A(men_men_n696_), .B(men_men_n1111_), .Y(men_men_n699_));
  NA3        u0677(.A(men_men_n679_), .B(men_men_n337_), .C(i_6_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n700_), .B(men_men_n23_), .Y(men_men_n701_));
  AOI210     u0679(.A0(men_men_n505_), .A1(men_men_n444_), .B0(men_men_n252_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n702_), .B(men_men_n648_), .Y(men_men_n703_));
  NO2        u0681(.A(i_11_), .B(men_men_n37_), .Y(men_men_n704_));
  NA2        u0682(.A(men_men_n704_), .B(men_men_n24_), .Y(men_men_n705_));
  OR3        u0683(.A(men_men_n703_), .B(men_men_n701_), .C(men_men_n699_), .Y(men_men_n706_));
  NO3        u0684(.A(men_men_n706_), .B(men_men_n694_), .C(men_men_n688_), .Y(men_men_n707_));
  NO2        u0685(.A(men_men_n247_), .B(men_men_n105_), .Y(men_men_n708_));
  NO2        u0686(.A(men_men_n708_), .B(men_men_n665_), .Y(men_men_n709_));
  NA2        u0687(.A(men_men_n709_), .B(i_1_), .Y(men_men_n710_));
  NO2        u0688(.A(men_men_n710_), .B(men_men_n659_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n439_), .B(men_men_n87_), .Y(men_men_n712_));
  NA2        u0690(.A(men_men_n711_), .B(men_men_n47_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n243_), .B(men_men_n45_), .Y(men_men_n714_));
  NO3        u0692(.A(men_men_n714_), .B(men_men_n327_), .C(men_men_n248_), .Y(men_men_n715_));
  NO2        u0693(.A(men_men_n120_), .B(men_men_n37_), .Y(men_men_n716_));
  NO2        u0694(.A(men_men_n716_), .B(i_6_), .Y(men_men_n717_));
  NO2        u0695(.A(men_men_n87_), .B(i_9_), .Y(men_men_n718_));
  NO2        u0696(.A(men_men_n718_), .B(men_men_n64_), .Y(men_men_n719_));
  NO2        u0697(.A(men_men_n719_), .B(men_men_n682_), .Y(men_men_n720_));
  NO4        u0698(.A(men_men_n720_), .B(men_men_n717_), .C(men_men_n715_), .D(i_4_), .Y(men_men_n721_));
  NA2        u0699(.A(i_1_), .B(i_3_), .Y(men_men_n722_));
  INV        u0700(.A(men_men_n721_), .Y(men_men_n723_));
  NA4        u0701(.A(men_men_n723_), .B(men_men_n713_), .C(men_men_n707_), .D(men_men_n685_), .Y(men_men_n724_));
  NO3        u0702(.A(men_men_n507_), .B(i_3_), .C(i_7_), .Y(men_men_n725_));
  NOi21      u0703(.An(men_men_n725_), .B(i_10_), .Y(men_men_n726_));
  OA210      u0704(.A0(men_men_n726_), .A1(men_men_n256_), .B0(men_men_n87_), .Y(men_men_n727_));
  NO3        u0705(.A(men_men_n508_), .B(men_men_n651_), .C(men_men_n87_), .Y(men_men_n728_));
  NA2        u0706(.A(men_men_n728_), .B(men_men_n25_), .Y(men_men_n729_));
  NA3        u0707(.A(men_men_n165_), .B(men_men_n85_), .C(men_men_n87_), .Y(men_men_n730_));
  NA2        u0708(.A(men_men_n730_), .B(men_men_n729_), .Y(men_men_n731_));
  OAI210     u0709(.A0(men_men_n731_), .A1(men_men_n727_), .B0(i_1_), .Y(men_men_n732_));
  AOI210     u0710(.A0(men_men_n281_), .A1(men_men_n101_), .B0(i_1_), .Y(men_men_n733_));
  NO2        u0711(.A(men_men_n389_), .B(i_2_), .Y(men_men_n734_));
  NA2        u0712(.A(men_men_n734_), .B(men_men_n733_), .Y(men_men_n735_));
  OAI210     u0713(.A0(men_men_n700_), .A1(men_men_n472_), .B0(men_men_n735_), .Y(men_men_n736_));
  INV        u0714(.A(men_men_n736_), .Y(men_men_n737_));
  AOI210     u0715(.A0(men_men_n737_), .A1(men_men_n732_), .B0(i_13_), .Y(men_men_n738_));
  OR2        u0716(.A(i_11_), .B(i_7_), .Y(men_men_n739_));
  NA3        u0717(.A(men_men_n739_), .B(men_men_n110_), .C(men_men_n141_), .Y(men_men_n740_));
  AOI220     u0718(.A0(men_men_n499_), .A1(men_men_n165_), .B0(men_men_n474_), .B1(men_men_n141_), .Y(men_men_n741_));
  OAI210     u0719(.A0(men_men_n741_), .A1(men_men_n45_), .B0(men_men_n740_), .Y(men_men_n742_));
  AOI210     u0720(.A0(men_men_n697_), .A1(men_men_n55_), .B0(i_12_), .Y(men_men_n743_));
  NO2        u0721(.A(men_men_n508_), .B(men_men_n24_), .Y(men_men_n744_));
  AOI220     u0722(.A0(men_men_n744_), .A1(men_men_n712_), .B0(men_men_n256_), .B1(men_men_n134_), .Y(men_men_n745_));
  OAI220     u0723(.A0(men_men_n745_), .A1(men_men_n41_), .B0(men_men_n1110_), .B1(men_men_n96_), .Y(men_men_n746_));
  AOI210     u0724(.A0(men_men_n742_), .A1(men_men_n353_), .B0(men_men_n746_), .Y(men_men_n747_));
  NA2        u0725(.A(men_men_n407_), .B(men_men_n698_), .Y(men_men_n748_));
  NO2        u0726(.A(men_men_n748_), .B(men_men_n253_), .Y(men_men_n749_));
  AOI210     u0727(.A0(men_men_n472_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n750_));
  NOi31      u0728(.An(men_men_n750_), .B(men_men_n641_), .C(men_men_n45_), .Y(men_men_n751_));
  NA2        u0729(.A(men_men_n130_), .B(i_13_), .Y(men_men_n752_));
  NO2        u0730(.A(men_men_n697_), .B(men_men_n118_), .Y(men_men_n753_));
  INV        u0731(.A(men_men_n753_), .Y(men_men_n754_));
  OAI220     u0732(.A0(men_men_n754_), .A1(men_men_n72_), .B0(men_men_n752_), .B1(men_men_n733_), .Y(men_men_n755_));
  NO3        u0733(.A(men_men_n72_), .B(men_men_n32_), .C(men_men_n105_), .Y(men_men_n756_));
  NA2        u0734(.A(men_men_n26_), .B(men_men_n199_), .Y(men_men_n757_));
  NA2        u0735(.A(men_men_n757_), .B(i_7_), .Y(men_men_n758_));
  INV        u0736(.A(men_men_n756_), .Y(men_men_n759_));
  AOI220     u0737(.A0(men_men_n407_), .A1(men_men_n698_), .B0(men_men_n95_), .B1(men_men_n106_), .Y(men_men_n760_));
  OAI220     u0738(.A0(men_men_n760_), .A1(men_men_n646_), .B0(men_men_n759_), .B1(men_men_n661_), .Y(men_men_n761_));
  NO4        u0739(.A(men_men_n761_), .B(men_men_n755_), .C(men_men_n751_), .D(men_men_n749_), .Y(men_men_n762_));
  OR2        u0740(.A(i_11_), .B(i_6_), .Y(men_men_n763_));
  NA3        u0741(.A(men_men_n645_), .B(men_men_n757_), .C(i_7_), .Y(men_men_n764_));
  AOI210     u0742(.A0(men_men_n764_), .A1(men_men_n754_), .B0(men_men_n763_), .Y(men_men_n765_));
  NA3        u0743(.A(men_men_n433_), .B(men_men_n650_), .C(men_men_n101_), .Y(men_men_n766_));
  NA2        u0744(.A(men_men_n687_), .B(i_13_), .Y(men_men_n767_));
  NA2        u0745(.A(men_men_n106_), .B(men_men_n757_), .Y(men_men_n768_));
  NAi21      u0746(.An(i_11_), .B(i_12_), .Y(men_men_n769_));
  NOi41      u0747(.An(men_men_n114_), .B(men_men_n769_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n770_));
  NA2        u0748(.A(men_men_n770_), .B(men_men_n768_), .Y(men_men_n771_));
  NA3        u0749(.A(men_men_n771_), .B(men_men_n767_), .C(men_men_n766_), .Y(men_men_n772_));
  OAI210     u0750(.A0(men_men_n772_), .A1(men_men_n765_), .B0(men_men_n64_), .Y(men_men_n773_));
  NO2        u0751(.A(i_2_), .B(i_12_), .Y(men_men_n774_));
  NA2        u0752(.A(men_men_n388_), .B(men_men_n774_), .Y(men_men_n775_));
  NA2        u0753(.A(i_8_), .B(men_men_n25_), .Y(men_men_n776_));
  NO3        u0754(.A(men_men_n776_), .B(men_men_n405_), .C(men_men_n645_), .Y(men_men_n777_));
  OAI210     u0755(.A0(men_men_n777_), .A1(men_men_n390_), .B0(men_men_n388_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n131_), .B(i_2_), .Y(men_men_n779_));
  NA2        u0757(.A(men_men_n779_), .B(men_men_n682_), .Y(men_men_n780_));
  NA3        u0758(.A(men_men_n780_), .B(men_men_n778_), .C(men_men_n775_), .Y(men_men_n781_));
  NA3        u0759(.A(men_men_n781_), .B(men_men_n46_), .C(men_men_n235_), .Y(men_men_n782_));
  NA4        u0760(.A(men_men_n782_), .B(men_men_n773_), .C(men_men_n762_), .D(men_men_n747_), .Y(men_men_n783_));
  OR4        u0761(.A(men_men_n783_), .B(men_men_n738_), .C(men_men_n724_), .D(men_men_n664_), .Y(men5));
  AOI210     u0762(.A0(men_men_n709_), .A1(men_men_n284_), .B0(men_men_n442_), .Y(men_men_n785_));
  AN2        u0763(.A(men_men_n24_), .B(i_10_), .Y(men_men_n786_));
  NA3        u0764(.A(men_men_n786_), .B(men_men_n774_), .C(men_men_n112_), .Y(men_men_n787_));
  NO2        u0765(.A(men_men_n646_), .B(i_11_), .Y(men_men_n788_));
  NA2        u0766(.A(men_men_n90_), .B(men_men_n788_), .Y(men_men_n789_));
  NA3        u0767(.A(men_men_n789_), .B(men_men_n787_), .C(men_men_n785_), .Y(men_men_n790_));
  NO3        u0768(.A(i_11_), .B(men_men_n247_), .C(i_13_), .Y(men_men_n791_));
  NO2        u0769(.A(men_men_n127_), .B(men_men_n23_), .Y(men_men_n792_));
  NA2        u0770(.A(i_12_), .B(i_8_), .Y(men_men_n793_));
  OAI210     u0771(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n793_), .Y(men_men_n794_));
  INV        u0772(.A(men_men_n471_), .Y(men_men_n795_));
  AOI220     u0773(.A0(men_men_n337_), .A1(men_men_n617_), .B0(men_men_n794_), .B1(men_men_n792_), .Y(men_men_n796_));
  INV        u0774(.A(men_men_n796_), .Y(men_men_n797_));
  NO2        u0775(.A(men_men_n797_), .B(men_men_n790_), .Y(men_men_n798_));
  INV        u0776(.A(men_men_n176_), .Y(men_men_n799_));
  INV        u0777(.A(men_men_n256_), .Y(men_men_n800_));
  OAI210     u0778(.A0(men_men_n734_), .A1(men_men_n473_), .B0(men_men_n114_), .Y(men_men_n801_));
  AOI210     u0779(.A0(men_men_n801_), .A1(men_men_n800_), .B0(men_men_n799_), .Y(men_men_n802_));
  NO2        u0780(.A(men_men_n481_), .B(men_men_n26_), .Y(men_men_n803_));
  NO2        u0781(.A(men_men_n803_), .B(men_men_n444_), .Y(men_men_n804_));
  NA2        u0782(.A(men_men_n804_), .B(i_2_), .Y(men_men_n805_));
  INV        u0783(.A(men_men_n805_), .Y(men_men_n806_));
  AOI210     u0784(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n440_), .Y(men_men_n807_));
  AOI210     u0785(.A0(men_men_n807_), .A1(men_men_n806_), .B0(men_men_n802_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n196_), .B(men_men_n128_), .Y(men_men_n809_));
  OAI210     u0787(.A0(men_men_n809_), .A1(men_men_n792_), .B0(i_2_), .Y(men_men_n810_));
  INV        u0788(.A(men_men_n177_), .Y(men_men_n811_));
  NO3        u0789(.A(men_men_n666_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n812_));
  AOI210     u0790(.A0(men_men_n811_), .A1(men_men_n90_), .B0(men_men_n812_), .Y(men_men_n813_));
  AOI210     u0791(.A0(men_men_n813_), .A1(men_men_n810_), .B0(men_men_n199_), .Y(men_men_n814_));
  OA210      u0792(.A0(men_men_n667_), .A1(men_men_n129_), .B0(i_13_), .Y(men_men_n815_));
  NA2        u0793(.A(men_men_n206_), .B(men_men_n209_), .Y(men_men_n816_));
  NA2        u0794(.A(men_men_n155_), .B(men_men_n642_), .Y(men_men_n817_));
  AOI210     u0795(.A0(men_men_n817_), .A1(men_men_n816_), .B0(men_men_n393_), .Y(men_men_n818_));
  AOI210     u0796(.A0(men_men_n216_), .A1(men_men_n151_), .B0(men_men_n553_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n819_), .B(men_men_n444_), .Y(men_men_n820_));
  NO2        u0798(.A(men_men_n106_), .B(men_men_n45_), .Y(men_men_n821_));
  INV        u0799(.A(men_men_n319_), .Y(men_men_n822_));
  NA4        u0800(.A(men_men_n822_), .B(men_men_n324_), .C(men_men_n127_), .D(men_men_n43_), .Y(men_men_n823_));
  OAI210     u0801(.A0(men_men_n823_), .A1(men_men_n821_), .B0(men_men_n820_), .Y(men_men_n824_));
  NO4        u0802(.A(men_men_n824_), .B(men_men_n818_), .C(men_men_n815_), .D(men_men_n814_), .Y(men_men_n825_));
  NA2        u0803(.A(men_men_n617_), .B(men_men_n28_), .Y(men_men_n826_));
  NA2        u0804(.A(men_men_n791_), .B(men_men_n291_), .Y(men_men_n827_));
  NA2        u0805(.A(men_men_n827_), .B(men_men_n826_), .Y(men_men_n828_));
  NO2        u0806(.A(men_men_n63_), .B(i_12_), .Y(men_men_n829_));
  NO2        u0807(.A(men_men_n829_), .B(men_men_n129_), .Y(men_men_n830_));
  NO2        u0808(.A(men_men_n830_), .B(men_men_n642_), .Y(men_men_n831_));
  AOI220     u0809(.A0(men_men_n831_), .A1(men_men_n36_), .B0(men_men_n828_), .B1(men_men_n47_), .Y(men_men_n832_));
  NA4        u0810(.A(men_men_n832_), .B(men_men_n825_), .C(men_men_n808_), .D(men_men_n798_), .Y(men6));
  NO3        u0811(.A(men_men_n267_), .B(men_men_n326_), .C(i_1_), .Y(men_men_n834_));
  NO2        u0812(.A(men_men_n191_), .B(men_men_n142_), .Y(men_men_n835_));
  OAI210     u0813(.A0(men_men_n835_), .A1(men_men_n834_), .B0(men_men_n779_), .Y(men_men_n836_));
  NA4        u0814(.A(men_men_n411_), .B(men_men_n513_), .C(men_men_n72_), .D(men_men_n105_), .Y(men_men_n837_));
  INV        u0815(.A(men_men_n837_), .Y(men_men_n838_));
  NO2        u0816(.A(men_men_n230_), .B(men_men_n518_), .Y(men_men_n839_));
  NO2        u0817(.A(men_men_n838_), .B(men_men_n349_), .Y(men_men_n840_));
  AO210      u0818(.A0(men_men_n840_), .A1(men_men_n836_), .B0(i_12_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n625_), .B(men_men_n64_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n726_), .B(men_men_n72_), .Y(men_men_n843_));
  BUFFER     u0821(.A(men_men_n672_), .Y(men_men_n844_));
  NA3        u0822(.A(men_men_n844_), .B(men_men_n843_), .C(men_men_n842_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n845_), .B(men_men_n74_), .Y(men_men_n846_));
  INV        u0824(.A(men_men_n348_), .Y(men_men_n847_));
  NA2        u0825(.A(men_men_n76_), .B(men_men_n134_), .Y(men_men_n848_));
  INV        u0826(.A(men_men_n127_), .Y(men_men_n849_));
  NA2        u0827(.A(men_men_n849_), .B(men_men_n47_), .Y(men_men_n850_));
  AOI210     u0828(.A0(men_men_n850_), .A1(men_men_n848_), .B0(men_men_n847_), .Y(men_men_n851_));
  NO3        u0829(.A(men_men_n263_), .B(men_men_n135_), .C(i_9_), .Y(men_men_n852_));
  NA2        u0830(.A(men_men_n852_), .B(men_men_n829_), .Y(men_men_n853_));
  AOI210     u0831(.A0(men_men_n853_), .A1(men_men_n551_), .B0(men_men_n191_), .Y(men_men_n854_));
  NO2        u0832(.A(men_men_n32_), .B(i_11_), .Y(men_men_n855_));
  NA3        u0833(.A(men_men_n855_), .B(men_men_n503_), .C(men_men_n411_), .Y(men_men_n856_));
  NAi32      u0834(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n857_));
  AOI210     u0835(.A0(men_men_n763_), .A1(men_men_n88_), .B0(men_men_n857_), .Y(men_men_n858_));
  OAI210     u0836(.A0(men_men_n725_), .A1(men_men_n605_), .B0(men_men_n604_), .Y(men_men_n859_));
  NAi31      u0837(.An(men_men_n858_), .B(men_men_n859_), .C(men_men_n856_), .Y(men_men_n860_));
  OR3        u0838(.A(men_men_n860_), .B(men_men_n854_), .C(men_men_n851_), .Y(men_men_n861_));
  NO2        u0839(.A(men_men_n739_), .B(i_2_), .Y(men_men_n862_));
  NA2        u0840(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n863_));
  OAI210     u0841(.A0(men_men_n863_), .A1(men_men_n432_), .B0(men_men_n383_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n864_), .B(men_men_n862_), .Y(men_men_n865_));
  AO220      u0843(.A0(men_men_n382_), .A1(men_men_n373_), .B0(men_men_n419_), .B1(men_men_n642_), .Y(men_men_n866_));
  NA3        u0844(.A(men_men_n866_), .B(men_men_n268_), .C(i_7_), .Y(men_men_n867_));
  OR2        u0845(.A(men_men_n667_), .B(men_men_n473_), .Y(men_men_n868_));
  NA3        u0846(.A(men_men_n868_), .B(men_men_n150_), .C(men_men_n70_), .Y(men_men_n869_));
  AO210      u0847(.A0(men_men_n525_), .A1(men_men_n795_), .B0(men_men_n36_), .Y(men_men_n870_));
  NA4        u0848(.A(men_men_n870_), .B(men_men_n869_), .C(men_men_n867_), .D(men_men_n865_), .Y(men_men_n871_));
  OAI210     u0849(.A0(men_men_n686_), .A1(i_11_), .B0(men_men_n88_), .Y(men_men_n872_));
  AOI220     u0850(.A0(men_men_n872_), .A1(men_men_n604_), .B0(men_men_n839_), .B1(men_men_n758_), .Y(men_men_n873_));
  NA3        u0851(.A(men_men_n393_), .B(men_men_n249_), .C(men_men_n150_), .Y(men_men_n874_));
  NA2        u0852(.A(men_men_n419_), .B(men_men_n71_), .Y(men_men_n875_));
  NA4        u0853(.A(men_men_n875_), .B(men_men_n874_), .C(men_men_n873_), .D(men_men_n649_), .Y(men_men_n876_));
  AO210      u0854(.A0(men_men_n553_), .A1(men_men_n47_), .B0(men_men_n89_), .Y(men_men_n877_));
  NA3        u0855(.A(men_men_n877_), .B(men_men_n514_), .C(men_men_n227_), .Y(men_men_n878_));
  AOI210     u0856(.A0(men_men_n473_), .A1(men_men_n471_), .B0(men_men_n603_), .Y(men_men_n879_));
  NO2        u0857(.A(men_men_n657_), .B(men_men_n106_), .Y(men_men_n880_));
  OAI210     u0858(.A0(men_men_n880_), .A1(men_men_n115_), .B0(men_men_n430_), .Y(men_men_n881_));
  NA2        u0859(.A(men_men_n255_), .B(men_men_n47_), .Y(men_men_n882_));
  INV        u0860(.A(men_men_n632_), .Y(men_men_n883_));
  NA3        u0861(.A(men_men_n883_), .B(men_men_n348_), .C(i_7_), .Y(men_men_n884_));
  NA4        u0862(.A(men_men_n884_), .B(men_men_n881_), .C(men_men_n879_), .D(men_men_n878_), .Y(men_men_n885_));
  NO4        u0863(.A(men_men_n885_), .B(men_men_n876_), .C(men_men_n871_), .D(men_men_n861_), .Y(men_men_n886_));
  NA4        u0864(.A(men_men_n886_), .B(men_men_n846_), .C(men_men_n841_), .D(men_men_n401_), .Y(men3));
  NA2        u0865(.A(i_6_), .B(i_7_), .Y(men_men_n888_));
  NO2        u0866(.A(men_men_n888_), .B(i_0_), .Y(men_men_n889_));
  NO2        u0867(.A(i_11_), .B(men_men_n247_), .Y(men_men_n890_));
  OAI210     u0868(.A0(men_men_n889_), .A1(men_men_n307_), .B0(men_men_n890_), .Y(men_men_n891_));
  NO2        u0869(.A(men_men_n891_), .B(men_men_n199_), .Y(men_men_n892_));
  NO3        u0870(.A(men_men_n477_), .B(men_men_n93_), .C(men_men_n45_), .Y(men_men_n893_));
  OA210      u0871(.A0(men_men_n893_), .A1(men_men_n892_), .B0(men_men_n179_), .Y(men_men_n894_));
  NA3        u0872(.A(men_men_n874_), .B(men_men_n649_), .C(men_men_n392_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n895_), .B(men_men_n40_), .Y(men_men_n896_));
  NOi21      u0874(.An(men_men_n100_), .B(men_men_n804_), .Y(men_men_n897_));
  NO3        u0875(.A(men_men_n677_), .B(men_men_n481_), .C(men_men_n134_), .Y(men_men_n898_));
  AN2        u0876(.A(men_men_n479_), .B(men_men_n56_), .Y(men_men_n899_));
  NO3        u0877(.A(men_men_n899_), .B(men_men_n898_), .C(men_men_n897_), .Y(men_men_n900_));
  AOI210     u0878(.A0(men_men_n900_), .A1(men_men_n896_), .B0(men_men_n49_), .Y(men_men_n901_));
  NO4        u0879(.A(men_men_n397_), .B(men_men_n404_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n902_));
  NA2        u0880(.A(men_men_n191_), .B(men_men_n613_), .Y(men_men_n903_));
  NOi21      u0881(.An(men_men_n903_), .B(men_men_n902_), .Y(men_men_n904_));
  NA2        u0882(.A(men_men_n750_), .B(men_men_n718_), .Y(men_men_n905_));
  NA2        u0883(.A(men_men_n354_), .B(men_men_n462_), .Y(men_men_n906_));
  OAI220     u0884(.A0(men_men_n906_), .A1(men_men_n905_), .B0(men_men_n904_), .B1(men_men_n64_), .Y(men_men_n907_));
  NOi21      u0885(.An(i_5_), .B(i_9_), .Y(men_men_n908_));
  NA2        u0886(.A(men_men_n908_), .B(men_men_n470_), .Y(men_men_n909_));
  AOI210     u0887(.A0(men_men_n281_), .A1(men_men_n505_), .B0(men_men_n728_), .Y(men_men_n910_));
  NO3        u0888(.A(men_men_n436_), .B(men_men_n281_), .C(men_men_n74_), .Y(men_men_n911_));
  NO2        u0889(.A(men_men_n180_), .B(men_men_n151_), .Y(men_men_n912_));
  AOI210     u0890(.A0(men_men_n912_), .A1(men_men_n255_), .B0(men_men_n911_), .Y(men_men_n913_));
  OAI220     u0891(.A0(men_men_n913_), .A1(men_men_n186_), .B0(men_men_n910_), .B1(men_men_n909_), .Y(men_men_n914_));
  NO4        u0892(.A(men_men_n914_), .B(men_men_n907_), .C(men_men_n901_), .D(men_men_n894_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n191_), .B(men_men_n24_), .Y(men_men_n916_));
  NO2        u0894(.A(men_men_n716_), .B(men_men_n639_), .Y(men_men_n917_));
  NO2        u0895(.A(men_men_n917_), .B(men_men_n916_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n331_), .B(men_men_n132_), .Y(men_men_n919_));
  NAi21      u0897(.An(men_men_n166_), .B(men_men_n462_), .Y(men_men_n920_));
  OAI220     u0898(.A0(men_men_n920_), .A1(men_men_n882_), .B0(men_men_n919_), .B1(men_men_n421_), .Y(men_men_n921_));
  NO2        u0899(.A(men_men_n921_), .B(men_men_n918_), .Y(men_men_n922_));
  NO2        u0900(.A(men_men_n411_), .B(men_men_n311_), .Y(men_men_n923_));
  NA2        u0901(.A(men_men_n923_), .B(men_men_n753_), .Y(men_men_n924_));
  NA2        u0902(.A(men_men_n614_), .B(i_0_), .Y(men_men_n925_));
  NO3        u0903(.A(men_men_n925_), .B(men_men_n406_), .C(men_men_n90_), .Y(men_men_n926_));
  NO4        u0904(.A(men_men_n631_), .B(men_men_n224_), .C(men_men_n440_), .D(men_men_n432_), .Y(men_men_n927_));
  AOI210     u0905(.A0(men_men_n927_), .A1(i_11_), .B0(men_men_n926_), .Y(men_men_n928_));
  INV        u0906(.A(men_men_n503_), .Y(men_men_n929_));
  AN2        u0907(.A(men_men_n100_), .B(men_men_n254_), .Y(men_men_n930_));
  NA2        u0908(.A(men_men_n791_), .B(men_men_n349_), .Y(men_men_n931_));
  AOI210     u0909(.A0(men_men_n514_), .A1(men_men_n90_), .B0(men_men_n59_), .Y(men_men_n932_));
  OAI220     u0910(.A0(men_men_n932_), .A1(men_men_n931_), .B0(men_men_n705_), .B1(men_men_n573_), .Y(men_men_n933_));
  NO2        u0911(.A(men_men_n265_), .B(men_men_n157_), .Y(men_men_n934_));
  NA2        u0912(.A(i_0_), .B(i_10_), .Y(men_men_n935_));
  AN2        u0913(.A(men_men_n934_), .B(i_6_), .Y(men_men_n936_));
  AOI220     u0914(.A0(men_men_n354_), .A1(men_men_n102_), .B0(men_men_n191_), .B1(men_men_n85_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n608_), .B(i_4_), .Y(men_men_n938_));
  NA2        u0916(.A(men_men_n194_), .B(men_men_n209_), .Y(men_men_n939_));
  OAI220     u0917(.A0(men_men_n939_), .A1(men_men_n931_), .B0(men_men_n938_), .B1(men_men_n937_), .Y(men_men_n940_));
  NO4        u0918(.A(men_men_n940_), .B(men_men_n936_), .C(men_men_n933_), .D(men_men_n930_), .Y(men_men_n941_));
  NA4        u0919(.A(men_men_n941_), .B(men_men_n928_), .C(men_men_n924_), .D(men_men_n922_), .Y(men_men_n942_));
  NO2        u0920(.A(men_men_n107_), .B(men_men_n37_), .Y(men_men_n943_));
  NA2        u0921(.A(i_11_), .B(i_9_), .Y(men_men_n944_));
  NO3        u0922(.A(i_12_), .B(men_men_n944_), .C(men_men_n648_), .Y(men_men_n945_));
  AO220      u0923(.A0(men_men_n945_), .A1(men_men_n943_), .B0(men_men_n283_), .B1(men_men_n89_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n49_), .B(i_7_), .Y(men_men_n947_));
  NA2        u0925(.A(men_men_n416_), .B(men_men_n184_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n948_), .B(men_men_n164_), .Y(men_men_n949_));
  NO2        u0927(.A(men_men_n180_), .B(i_0_), .Y(men_men_n950_));
  INV        u0928(.A(men_men_n950_), .Y(men_men_n951_));
  NA2        u0929(.A(men_men_n503_), .B(men_men_n241_), .Y(men_men_n952_));
  AOI210     u0930(.A0(men_men_n391_), .A1(men_men_n42_), .B0(men_men_n429_), .Y(men_men_n953_));
  OAI220     u0931(.A0(men_men_n953_), .A1(men_men_n909_), .B0(men_men_n952_), .B1(men_men_n951_), .Y(men_men_n954_));
  NO3        u0932(.A(men_men_n954_), .B(men_men_n949_), .C(men_men_n946_), .Y(men_men_n955_));
  NA2        u0933(.A(men_men_n704_), .B(men_men_n124_), .Y(men_men_n956_));
  NO2        u0934(.A(i_6_), .B(men_men_n956_), .Y(men_men_n957_));
  AOI210     u0935(.A0(men_men_n472_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n958_));
  NA2        u0936(.A(men_men_n176_), .B(men_men_n107_), .Y(men_men_n959_));
  NOi32      u0937(.An(men_men_n958_), .Bn(men_men_n194_), .C(men_men_n959_), .Y(men_men_n960_));
  NO2        u0938(.A(men_men_n960_), .B(men_men_n957_), .Y(men_men_n961_));
  NOi21      u0939(.An(i_7_), .B(i_5_), .Y(men_men_n962_));
  NOi31      u0940(.An(men_men_n962_), .B(i_0_), .C(men_men_n769_), .Y(men_men_n963_));
  NA3        u0941(.A(men_men_n963_), .B(men_men_n405_), .C(i_6_), .Y(men_men_n964_));
  OA210      u0942(.A0(men_men_n959_), .A1(men_men_n551_), .B0(men_men_n964_), .Y(men_men_n965_));
  NO3        u0943(.A(men_men_n424_), .B(men_men_n385_), .C(men_men_n381_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n275_), .B(men_men_n338_), .Y(men_men_n967_));
  NO2        u0945(.A(men_men_n769_), .B(men_men_n270_), .Y(men_men_n968_));
  AOI210     u0946(.A0(men_men_n968_), .A1(men_men_n967_), .B0(men_men_n966_), .Y(men_men_n969_));
  NA4        u0947(.A(men_men_n969_), .B(men_men_n965_), .C(men_men_n961_), .D(men_men_n955_), .Y(men_men_n970_));
  NO2        u0948(.A(men_men_n916_), .B(men_men_n250_), .Y(men_men_n971_));
  AN2        u0949(.A(men_men_n353_), .B(men_men_n349_), .Y(men_men_n972_));
  AN2        u0950(.A(men_men_n972_), .B(men_men_n912_), .Y(men_men_n973_));
  OAI210     u0951(.A0(men_men_n973_), .A1(men_men_n971_), .B0(i_10_), .Y(men_men_n974_));
  OA210      u0952(.A0(men_men_n503_), .A1(men_men_n233_), .B0(men_men_n502_), .Y(men_men_n975_));
  NA3        u0953(.A(men_men_n502_), .B(men_men_n433_), .C(men_men_n46_), .Y(men_men_n976_));
  OAI210     u0954(.A0(men_men_n920_), .A1(men_men_n929_), .B0(men_men_n976_), .Y(men_men_n977_));
  NO2        u0955(.A(men_men_n268_), .B(men_men_n47_), .Y(men_men_n978_));
  NO2        u0956(.A(men_men_n978_), .B(men_men_n193_), .Y(men_men_n979_));
  AOI220     u0957(.A0(men_men_n979_), .A1(men_men_n503_), .B0(men_men_n977_), .B1(men_men_n74_), .Y(men_men_n980_));
  NA3        u0958(.A(men_men_n863_), .B(men_men_n403_), .C(men_men_n686_), .Y(men_men_n981_));
  NA2        u0959(.A(men_men_n96_), .B(men_men_n45_), .Y(men_men_n982_));
  NO2        u0960(.A(men_men_n76_), .B(men_men_n793_), .Y(men_men_n983_));
  AOI220     u0961(.A0(men_men_n983_), .A1(men_men_n982_), .B0(men_men_n179_), .B1(men_men_n639_), .Y(men_men_n984_));
  AOI210     u0962(.A0(men_men_n984_), .A1(men_men_n981_), .B0(men_men_n48_), .Y(men_men_n985_));
  NO3        u0963(.A(men_men_n631_), .B(men_men_n380_), .C(men_men_n24_), .Y(men_men_n986_));
  AOI210     u0964(.A0(men_men_n744_), .A1(men_men_n585_), .B0(men_men_n986_), .Y(men_men_n987_));
  NO2        u0965(.A(men_men_n644_), .B(men_men_n109_), .Y(men_men_n988_));
  NA2        u0966(.A(men_men_n988_), .B(i_0_), .Y(men_men_n989_));
  OAI220     u0967(.A0(men_men_n989_), .A1(men_men_n87_), .B0(men_men_n987_), .B1(men_men_n177_), .Y(men_men_n990_));
  NO3        u0968(.A(men_men_n990_), .B(men_men_n985_), .C(men_men_n555_), .Y(men_men_n991_));
  NA3        u0969(.A(men_men_n991_), .B(men_men_n980_), .C(men_men_n974_), .Y(men_men_n992_));
  NO3        u0970(.A(men_men_n992_), .B(men_men_n970_), .C(men_men_n942_), .Y(men_men_n993_));
  NO2        u0971(.A(i_0_), .B(men_men_n769_), .Y(men_men_n994_));
  NA2        u0972(.A(men_men_n74_), .B(men_men_n45_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n935_), .B(men_men_n995_), .Y(men_men_n996_));
  NO3        u0974(.A(men_men_n109_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n997_));
  AO220      u0975(.A0(men_men_n997_), .A1(men_men_n996_), .B0(men_men_n994_), .B1(men_men_n179_), .Y(men_men_n998_));
  NO2        u0976(.A(men_men_n842_), .B(men_men_n959_), .Y(men_men_n999_));
  AOI210     u0977(.A0(men_men_n998_), .A1(men_men_n370_), .B0(men_men_n999_), .Y(men_men_n1000_));
  NA2        u0978(.A(men_men_n779_), .B(men_men_n149_), .Y(men_men_n1001_));
  INV        u0979(.A(men_men_n1001_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n1002_), .B(men_men_n718_), .C(men_men_n74_), .Y(men_men_n1003_));
  NO2        u0981(.A(men_men_n859_), .B(men_men_n424_), .Y(men_men_n1004_));
  NA3        u0982(.A(men_men_n889_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n890_), .B(i_9_), .Y(men_men_n1006_));
  AOI210     u0984(.A0(men_men_n1005_), .A1(men_men_n531_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  OAI210     u0985(.A0(men_men_n255_), .A1(i_9_), .B0(men_men_n240_), .Y(men_men_n1008_));
  AOI210     u0986(.A0(men_men_n1008_), .A1(men_men_n925_), .B0(men_men_n157_), .Y(men_men_n1009_));
  NO3        u0987(.A(men_men_n1009_), .B(men_men_n1007_), .C(men_men_n1004_), .Y(men_men_n1010_));
  NA3        u0988(.A(men_men_n1010_), .B(men_men_n1003_), .C(men_men_n1000_), .Y(men_men_n1011_));
  NA2        u0989(.A(men_men_n972_), .B(men_men_n393_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n318_), .A1(men_men_n166_), .B0(men_men_n1012_), .Y(men_men_n1013_));
  NA3        u0991(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n1014_));
  NA2        u0992(.A(men_men_n947_), .B(men_men_n519_), .Y(men_men_n1015_));
  AOI210     u0993(.A0(men_men_n1014_), .A1(men_men_n166_), .B0(men_men_n1015_), .Y(men_men_n1016_));
  NO2        u0994(.A(men_men_n1016_), .B(men_men_n1013_), .Y(men_men_n1017_));
  NO3        u0995(.A(men_men_n935_), .B(men_men_n908_), .C(men_men_n196_), .Y(men_men_n1018_));
  AOI220     u0996(.A0(men_men_n1018_), .A1(i_11_), .B0(men_men_n609_), .B1(men_men_n76_), .Y(men_men_n1019_));
  NO3        u0997(.A(men_men_n218_), .B(men_men_n404_), .C(i_0_), .Y(men_men_n1020_));
  OAI210     u0998(.A0(men_men_n1020_), .A1(men_men_n77_), .B0(i_13_), .Y(men_men_n1021_));
  INV        u0999(.A(men_men_n227_), .Y(men_men_n1022_));
  OAI220     u1000(.A0(men_men_n567_), .A1(men_men_n142_), .B0(men_men_n691_), .B1(men_men_n661_), .Y(men_men_n1023_));
  NA3        u1001(.A(men_men_n1023_), .B(i_7_), .C(men_men_n1022_), .Y(men_men_n1024_));
  NA4        u1002(.A(men_men_n1024_), .B(men_men_n1021_), .C(men_men_n1019_), .D(men_men_n1017_), .Y(men_men_n1025_));
  NO2        u1003(.A(men_men_n253_), .B(men_men_n96_), .Y(men_men_n1026_));
  NA2        u1004(.A(men_men_n1026_), .B(men_men_n994_), .Y(men_men_n1027_));
  AOI220     u1005(.A0(men_men_n962_), .A1(men_men_n519_), .B0(men_men_n889_), .B1(men_men_n167_), .Y(men_men_n1028_));
  NA2        u1006(.A(men_men_n373_), .B(men_men_n181_), .Y(men_men_n1029_));
  OA220      u1007(.A0(men_men_n1029_), .A1(men_men_n1028_), .B0(men_men_n1027_), .B1(i_5_), .Y(men_men_n1030_));
  AOI210     u1008(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n180_), .Y(men_men_n1031_));
  NA2        u1009(.A(men_men_n1031_), .B(men_men_n975_), .Y(men_men_n1032_));
  NA3        u1010(.A(men_men_n658_), .B(men_men_n191_), .C(men_men_n85_), .Y(men_men_n1033_));
  NA2        u1011(.A(men_men_n1033_), .B(men_men_n583_), .Y(men_men_n1034_));
  NA3        u1012(.A(men_men_n524_), .B(men_men_n517_), .C(men_men_n500_), .Y(men_men_n1035_));
  NO2        u1013(.A(men_men_n1035_), .B(men_men_n1034_), .Y(men_men_n1036_));
  NA3        u1014(.A(men_men_n411_), .B(men_men_n176_), .C(men_men_n175_), .Y(men_men_n1037_));
  NA3        u1015(.A(men_men_n947_), .B(men_men_n307_), .C(men_men_n240_), .Y(men_men_n1038_));
  NA2        u1016(.A(men_men_n1038_), .B(men_men_n1037_), .Y(men_men_n1039_));
  NA3        u1017(.A(men_men_n411_), .B(men_men_n355_), .C(men_men_n231_), .Y(men_men_n1040_));
  INV        u1018(.A(men_men_n1040_), .Y(men_men_n1041_));
  NOi31      u1019(.An(men_men_n410_), .B(men_men_n995_), .C(men_men_n250_), .Y(men_men_n1042_));
  NO3        u1020(.A(men_men_n944_), .B(men_men_n227_), .C(men_men_n196_), .Y(men_men_n1043_));
  NO4        u1021(.A(men_men_n1043_), .B(men_men_n1042_), .C(men_men_n1041_), .D(men_men_n1039_), .Y(men_men_n1044_));
  NA4        u1022(.A(men_men_n1044_), .B(men_men_n1036_), .C(men_men_n1032_), .D(men_men_n1030_), .Y(men_men_n1045_));
  INV        u1023(.A(men_men_n660_), .Y(men_men_n1046_));
  NO3        u1024(.A(men_men_n1046_), .B(men_men_n599_), .C(men_men_n367_), .Y(men_men_n1047_));
  INV        u1025(.A(men_men_n1047_), .Y(men_men_n1048_));
  NA3        u1026(.A(men_men_n324_), .B(i_5_), .C(men_men_n199_), .Y(men_men_n1049_));
  NAi31      u1027(.An(men_men_n252_), .B(men_men_n1049_), .C(men_men_n253_), .Y(men_men_n1050_));
  NO4        u1028(.A(men_men_n250_), .B(men_men_n218_), .C(i_0_), .D(i_12_), .Y(men_men_n1051_));
  AOI220     u1029(.A0(men_men_n1051_), .A1(men_men_n1050_), .B0(men_men_n838_), .B1(men_men_n181_), .Y(men_men_n1052_));
  AN2        u1030(.A(men_men_n935_), .B(men_men_n157_), .Y(men_men_n1053_));
  NO4        u1031(.A(men_men_n1053_), .B(i_12_), .C(men_men_n695_), .D(men_men_n134_), .Y(men_men_n1054_));
  NA2        u1032(.A(men_men_n1054_), .B(men_men_n227_), .Y(men_men_n1055_));
  NA3        u1033(.A(men_men_n102_), .B(men_men_n613_), .C(i_11_), .Y(men_men_n1056_));
  NO2        u1034(.A(men_men_n1056_), .B(men_men_n159_), .Y(men_men_n1057_));
  NA2        u1035(.A(men_men_n962_), .B(men_men_n499_), .Y(men_men_n1058_));
  NA2        u1036(.A(men_men_n65_), .B(men_men_n105_), .Y(men_men_n1059_));
  OAI220     u1037(.A0(men_men_n1059_), .A1(men_men_n1049_), .B0(men_men_n1058_), .B1(men_men_n719_), .Y(men_men_n1060_));
  AOI210     u1038(.A0(men_men_n1060_), .A1(men_men_n950_), .B0(men_men_n1057_), .Y(men_men_n1061_));
  NA4        u1039(.A(men_men_n1061_), .B(men_men_n1055_), .C(men_men_n1052_), .D(men_men_n1048_), .Y(men_men_n1062_));
  NO4        u1040(.A(men_men_n1062_), .B(men_men_n1045_), .C(men_men_n1025_), .D(men_men_n1011_), .Y(men_men_n1063_));
  OAI210     u1041(.A0(men_men_n862_), .A1(men_men_n855_), .B0(men_men_n37_), .Y(men_men_n1064_));
  NA3        u1042(.A(men_men_n958_), .B(men_men_n388_), .C(i_5_), .Y(men_men_n1065_));
  NA3        u1043(.A(men_men_n1065_), .B(men_men_n1064_), .C(men_men_n656_), .Y(men_men_n1066_));
  NA2        u1044(.A(men_men_n1066_), .B(men_men_n214_), .Y(men_men_n1067_));
  AN2        u1045(.A(men_men_n739_), .B(men_men_n389_), .Y(men_men_n1068_));
  NA2        u1046(.A(men_men_n192_), .B(men_men_n194_), .Y(men_men_n1069_));
  AO210      u1047(.A0(men_men_n1068_), .A1(men_men_n33_), .B0(men_men_n1069_), .Y(men_men_n1070_));
  OAI210     u1048(.A0(men_men_n660_), .A1(men_men_n658_), .B0(men_men_n337_), .Y(men_men_n1071_));
  NAi31      u1049(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1072_));
  AOI210     u1050(.A0(men_men_n120_), .A1(men_men_n71_), .B0(men_men_n1072_), .Y(men_men_n1073_));
  NO2        u1051(.A(men_men_n1073_), .B(men_men_n692_), .Y(men_men_n1074_));
  NA3        u1052(.A(men_men_n1074_), .B(men_men_n1071_), .C(men_men_n1070_), .Y(men_men_n1075_));
  NO2        u1053(.A(men_men_n489_), .B(men_men_n281_), .Y(men_men_n1076_));
  NO4        u1054(.A(men_men_n243_), .B(men_men_n148_), .C(men_men_n722_), .D(men_men_n37_), .Y(men_men_n1077_));
  NO3        u1055(.A(men_men_n1077_), .B(men_men_n1076_), .C(men_men_n927_), .Y(men_men_n1078_));
  OAI210     u1056(.A0(men_men_n1056_), .A1(men_men_n151_), .B0(men_men_n1078_), .Y(men_men_n1079_));
  AOI210     u1057(.A0(men_men_n1075_), .A1(men_men_n49_), .B0(men_men_n1079_), .Y(men_men_n1080_));
  AOI210     u1058(.A0(men_men_n1080_), .A1(men_men_n1067_), .B0(men_men_n74_), .Y(men_men_n1081_));
  NO2        u1059(.A(men_men_n606_), .B(men_men_n400_), .Y(men_men_n1082_));
  NO2        u1060(.A(men_men_n1082_), .B(men_men_n799_), .Y(men_men_n1083_));
  OAI210     u1061(.A0(men_men_n81_), .A1(men_men_n55_), .B0(men_men_n112_), .Y(men_men_n1084_));
  NA2        u1062(.A(men_men_n1084_), .B(men_men_n77_), .Y(men_men_n1085_));
  AOI210     u1063(.A0(men_men_n1031_), .A1(men_men_n947_), .B0(men_men_n963_), .Y(men_men_n1086_));
  AOI210     u1064(.A0(men_men_n1086_), .A1(men_men_n1085_), .B0(men_men_n722_), .Y(men_men_n1087_));
  NA2        u1065(.A(men_men_n275_), .B(men_men_n58_), .Y(men_men_n1088_));
  AOI220     u1066(.A0(men_men_n1088_), .A1(men_men_n77_), .B0(men_men_n368_), .B1(men_men_n267_), .Y(men_men_n1089_));
  NO2        u1067(.A(men_men_n1089_), .B(men_men_n247_), .Y(men_men_n1090_));
  NA3        u1068(.A(men_men_n100_), .B(men_men_n326_), .C(men_men_n31_), .Y(men_men_n1091_));
  INV        u1069(.A(men_men_n1091_), .Y(men_men_n1092_));
  NO3        u1070(.A(men_men_n1092_), .B(men_men_n1090_), .C(men_men_n1087_), .Y(men_men_n1093_));
  OAI210     u1071(.A0(men_men_n283_), .A1(men_men_n162_), .B0(men_men_n90_), .Y(men_men_n1094_));
  NA3        u1072(.A(men_men_n803_), .B(men_men_n307_), .C(men_men_n81_), .Y(men_men_n1095_));
  AOI210     u1073(.A0(men_men_n1095_), .A1(men_men_n1094_), .B0(i_11_), .Y(men_men_n1096_));
  NA2        u1074(.A(men_men_n651_), .B(men_men_n224_), .Y(men_men_n1097_));
  OAI210     u1075(.A0(men_men_n1097_), .A1(men_men_n958_), .B0(men_men_n214_), .Y(men_men_n1098_));
  NA2        u1076(.A(men_men_n168_), .B(i_5_), .Y(men_men_n1099_));
  NO2        u1077(.A(men_men_n1098_), .B(men_men_n1099_), .Y(men_men_n1100_));
  NO3        u1078(.A(men_men_n60_), .B(men_men_n59_), .C(i_4_), .Y(men_men_n1101_));
  OAI210     u1079(.A0(men_men_n967_), .A1(men_men_n326_), .B0(men_men_n1101_), .Y(men_men_n1102_));
  NO2        u1080(.A(men_men_n1102_), .B(men_men_n769_), .Y(men_men_n1103_));
  NO3        u1081(.A(men_men_n1103_), .B(men_men_n1100_), .C(men_men_n1096_), .Y(men_men_n1104_));
  OAI210     u1082(.A0(men_men_n1093_), .A1(i_4_), .B0(men_men_n1104_), .Y(men_men_n1105_));
  NO3        u1083(.A(men_men_n1105_), .B(men_men_n1083_), .C(men_men_n1081_), .Y(men_men_n1106_));
  NA4        u1084(.A(men_men_n1106_), .B(men_men_n1063_), .C(men_men_n993_), .D(men_men_n915_), .Y(men4));
  INV        u1085(.A(men_men_n743_), .Y(men_men_n1110_));
  INV        u1086(.A(i_2_), .Y(men_men_n1111_));
  INV        u1087(.A(men_men_n514_), .Y(men_men_n1112_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule