// Benchmark "top" written by ABC on Thu Jun 20 14:59:19 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n136_, new_new_n137_, new_new_n138_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n971_,
    new_new_n972_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(mai1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g026(.A(i_5_), .Y(new_new_n49_));
  NO2        g027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g041(.A(i_1_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g064(.A(i_6_), .Y(new_new_n87_));
  NO2        g065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  INV        g066(.A(new_new_n88_), .Y(new_new_n89_));
  OAI210     g067(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n89_), .Y(new_new_n90_));
  NAi21      g068(.An(i_6_), .B(i_10_), .Y(new_new_n91_));
  NA2        g069(.A(i_6_), .B(i_9_), .Y(new_new_n92_));
  AOI210     g070(.A0(new_new_n92_), .A1(new_new_n91_), .B0(new_new_n64_), .Y(new_new_n93_));
  NA2        g071(.A(i_2_), .B(i_6_), .Y(new_new_n94_));
  NO3        g072(.A(new_new_n94_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n93_), .Y(new_new_n96_));
  AOI210     g074(.A0(new_new_n96_), .A1(new_new_n90_), .B0(new_new_n81_), .Y(new_new_n97_));
  AN3        g075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n98_), .B(new_new_n32_), .Y(new_new_n101_));
  INV        g079(.A(i_7_), .Y(new_new_n102_));
  NA2        g080(.A(new_new_n47_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(new_new_n87_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  INV        g084(.A(new_new_n106_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n103_), .Y(new_new_n108_));
  NAi21      g086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n91_), .C(new_new_n54_), .Y(new_new_n110_));
  AN2        g088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g090(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n113_));
  NO2        g091(.A(i_8_), .B(new_new_n102_), .Y(new_new_n114_));
  NA2        g092(.A(i_12_), .B(i_7_), .Y(new_new_n115_));
  NO2        g093(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n116_));
  NA2        g094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  NAi41      g095(.An(new_new_n110_), .B(new_new_n117_), .C(new_new_n108_), .D(new_new_n101_), .Y(new_new_n118_));
  NOi21      g096(.An(i_1_), .B(i_5_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_11_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n121_));
  NA2        g099(.A(i_7_), .B(new_new_n25_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n122_), .B(new_new_n121_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n123_), .B(new_new_n47_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n92_), .B(new_new_n91_), .Y(new_new_n125_));
  NAi21      g103(.An(i_3_), .B(i_8_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n63_), .Y(new_new_n127_));
  NOi31      g105(.An(new_new_n127_), .B(new_new_n125_), .C(new_new_n124_), .Y(new_new_n128_));
  NO2        g106(.A(i_1_), .B(new_new_n87_), .Y(new_new_n129_));
  NO2        g107(.A(i_6_), .B(i_5_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(i_3_), .Y(new_new_n131_));
  AO210      g109(.A0(new_new_n131_), .A1(new_new_n48_), .B0(new_new_n129_), .Y(new_new_n132_));
  OAI220     g110(.A0(new_new_n132_), .A1(new_new_n109_), .B0(new_new_n128_), .B1(new_new_n120_), .Y(new_new_n133_));
  NO3        g111(.A(new_new_n133_), .B(new_new_n118_), .C(new_new_n97_), .Y(new_new_n134_));
  NA3        g112(.A(new_new_n134_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g113(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n136_));
  NA2        g114(.A(i_6_), .B(new_new_n25_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n137_), .B(new_new_n136_), .Y(new_new_n138_));
  NA4        g116(.A(new_new_n138_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g117(.A(i_8_), .B(i_7_), .Y(new_new_n140_));
  NA2        g118(.A(new_new_n140_), .B(i_6_), .Y(new_new_n141_));
  NO2        g119(.A(i_12_), .B(i_13_), .Y(new_new_n142_));
  NAi21      g120(.An(i_5_), .B(i_11_), .Y(new_new_n143_));
  NOi21      g121(.An(new_new_n142_), .B(new_new_n143_), .Y(new_new_n144_));
  NO2        g122(.A(i_0_), .B(i_1_), .Y(new_new_n145_));
  NA2        g123(.A(i_2_), .B(i_3_), .Y(new_new_n146_));
  NO2        g124(.A(new_new_n146_), .B(i_4_), .Y(new_new_n147_));
  NA3        g125(.A(new_new_n147_), .B(new_new_n145_), .C(new_new_n144_), .Y(new_new_n148_));
  OR2        g126(.A(new_new_n148_), .B(new_new_n25_), .Y(new_new_n149_));
  AN2        g127(.A(new_new_n142_), .B(new_new_n84_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n150_), .B(new_new_n27_), .Y(new_new_n151_));
  NA2        g129(.A(i_1_), .B(i_5_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n153_));
  NA2        g131(.A(new_new_n153_), .B(new_new_n36_), .Y(new_new_n154_));
  NO3        g132(.A(new_new_n154_), .B(new_new_n152_), .C(new_new_n151_), .Y(new_new_n155_));
  OR2        g133(.A(i_0_), .B(i_1_), .Y(new_new_n156_));
  NO3        g134(.A(new_new_n156_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n157_));
  NAi32      g135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n158_));
  NOi21      g136(.An(i_4_), .B(i_10_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n159_), .B(new_new_n40_), .Y(new_new_n160_));
  NO2        g138(.A(i_3_), .B(i_5_), .Y(new_new_n161_));
  INV        g139(.A(new_new_n155_), .Y(new_new_n162_));
  AOI210     g140(.A0(new_new_n162_), .A1(new_new_n149_), .B0(new_new_n141_), .Y(new_new_n163_));
  NA3        g141(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n164_));
  NOi21      g142(.An(i_4_), .B(i_9_), .Y(new_new_n165_));
  NOi21      g143(.An(i_11_), .B(i_13_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  BUFFER     g145(.A(new_new_n167_), .Y(new_new_n168_));
  NO2        g146(.A(i_4_), .B(i_5_), .Y(new_new_n169_));
  NAi21      g147(.An(i_12_), .B(i_11_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n170_), .B(i_13_), .Y(new_new_n171_));
  NA3        g149(.A(new_new_n171_), .B(new_new_n169_), .C(new_new_n84_), .Y(new_new_n172_));
  AOI210     g150(.A0(new_new_n172_), .A1(new_new_n168_), .B0(new_new_n164_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n36_), .B(i_5_), .Y(new_new_n175_));
  NA2        g153(.A(i_3_), .B(i_5_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n74_), .B(i_5_), .Y(new_new_n177_));
  NO2        g155(.A(i_13_), .B(i_10_), .Y(new_new_n178_));
  NA3        g156(.A(new_new_n178_), .B(new_new_n177_), .C(new_new_n45_), .Y(new_new_n179_));
  NO2        g157(.A(i_2_), .B(i_1_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(i_3_), .Y(new_new_n181_));
  NAi21      g159(.An(i_4_), .B(i_12_), .Y(new_new_n182_));
  NO4        g160(.A(new_new_n182_), .B(new_new_n181_), .C(new_new_n179_), .D(new_new_n25_), .Y(new_new_n183_));
  NO2        g161(.A(new_new_n183_), .B(new_new_n173_), .Y(new_new_n184_));
  INV        g162(.A(i_8_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(i_7_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n186_), .B(i_6_), .Y(new_new_n187_));
  NO3        g165(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(new_new_n114_), .Y(new_new_n189_));
  NO3        g167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n191_));
  NO3        g169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n192_));
  OAI210     g170(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n192_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n193_), .B(new_new_n189_), .Y(new_new_n194_));
  NO2        g172(.A(i_3_), .B(i_8_), .Y(new_new_n195_));
  NO3        g173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n104_), .B(new_new_n59_), .Y(new_new_n197_));
  NO2        g175(.A(i_13_), .B(i_9_), .Y(new_new_n198_));
  NA3        g176(.A(new_new_n198_), .B(i_6_), .C(new_new_n185_), .Y(new_new_n199_));
  NAi21      g177(.An(i_12_), .B(i_3_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n45_), .B(i_5_), .Y(new_new_n201_));
  NO3        g179(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n202_));
  NA3        g180(.A(new_new_n202_), .B(new_new_n201_), .C(i_10_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n203_), .B(new_new_n199_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n204_), .B(new_new_n194_), .Y(new_new_n205_));
  OAI220     g183(.A0(new_new_n205_), .A1(i_4_), .B0(new_new_n187_), .B1(new_new_n184_), .Y(new_new_n206_));
  NAi21      g184(.An(i_12_), .B(i_7_), .Y(new_new_n207_));
  NA3        g185(.A(i_13_), .B(new_new_n185_), .C(i_10_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n208_), .B(new_new_n207_), .Y(new_new_n209_));
  NA2        g187(.A(i_0_), .B(i_5_), .Y(new_new_n210_));
  NA2        g188(.A(new_new_n210_), .B(new_new_n105_), .Y(new_new_n211_));
  OAI220     g189(.A0(new_new_n211_), .A1(new_new_n181_), .B0(i_2_), .B1(new_new_n131_), .Y(new_new_n212_));
  NAi31      g190(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n36_), .B(i_13_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n216_));
  INV        g194(.A(i_13_), .Y(new_new_n217_));
  NO2        g195(.A(i_12_), .B(new_new_n217_), .Y(new_new_n218_));
  NA3        g196(.A(new_new_n218_), .B(new_new_n190_), .C(new_new_n188_), .Y(new_new_n219_));
  INV        g197(.A(new_new_n219_), .Y(new_new_n220_));
  AOI220     g198(.A0(new_new_n220_), .A1(new_new_n140_), .B0(new_new_n212_), .B1(new_new_n209_), .Y(new_new_n221_));
  NO2        g199(.A(i_12_), .B(new_new_n37_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n176_), .B(i_4_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  OR2        g202(.A(i_8_), .B(i_7_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n225_), .B(new_new_n87_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n54_), .B(i_1_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n228_));
  INV        g206(.A(i_12_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n45_), .B(new_new_n229_), .Y(new_new_n230_));
  NO3        g208(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n231_));
  NA2        g209(.A(i_2_), .B(i_1_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n228_), .B(new_new_n224_), .Y(new_new_n233_));
  NO3        g211(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n234_));
  NAi21      g212(.An(i_4_), .B(i_3_), .Y(new_new_n235_));
  NO2        g213(.A(i_0_), .B(i_6_), .Y(new_new_n236_));
  NOi41      g214(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n232_), .B(new_new_n176_), .Y(new_new_n239_));
  NAi21      g217(.An(new_new_n238_), .B(new_new_n239_), .Y(new_new_n240_));
  INV        g218(.A(new_new_n240_), .Y(new_new_n241_));
  AOI220     g219(.A0(new_new_n241_), .A1(new_new_n40_), .B0(new_new_n233_), .B1(new_new_n198_), .Y(new_new_n242_));
  NO2        g220(.A(i_11_), .B(new_new_n217_), .Y(new_new_n243_));
  NOi21      g221(.An(i_1_), .B(i_6_), .Y(new_new_n244_));
  NAi21      g222(.An(i_3_), .B(i_7_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n246_));
  NO2        g224(.A(i_12_), .B(i_3_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n74_), .B(i_5_), .Y(new_new_n248_));
  NA3        g226(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n225_), .B(new_new_n37_), .Y(new_new_n250_));
  NA2        g228(.A(i_12_), .B(i_6_), .Y(new_new_n251_));
  OR2        g229(.A(i_13_), .B(i_9_), .Y(new_new_n252_));
  NO3        g230(.A(new_new_n252_), .B(new_new_n251_), .C(new_new_n49_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n235_), .B(i_2_), .Y(new_new_n254_));
  NA3        g232(.A(new_new_n254_), .B(new_new_n253_), .C(new_new_n45_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n243_), .B(i_9_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n248_), .B(new_new_n65_), .Y(new_new_n257_));
  OAI210     g235(.A0(new_new_n257_), .A1(new_new_n256_), .B0(new_new_n255_), .Y(new_new_n258_));
  NA2        g236(.A(new_new_n153_), .B(new_new_n64_), .Y(new_new_n259_));
  NO3        g237(.A(i_11_), .B(new_new_n217_), .C(new_new_n25_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n245_), .B(i_8_), .Y(new_new_n261_));
  NA3        g239(.A(i_5_), .B(new_new_n261_), .C(new_new_n260_), .Y(new_new_n262_));
  NO3        g240(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n263_), .B(new_new_n250_), .C(new_new_n218_), .Y(new_new_n264_));
  AOI210     g242(.A0(new_new_n264_), .A1(new_new_n262_), .B0(new_new_n259_), .Y(new_new_n265_));
  AOI210     g243(.A0(new_new_n258_), .A1(new_new_n250_), .B0(new_new_n265_), .Y(new_new_n266_));
  NA3        g244(.A(new_new_n266_), .B(new_new_n242_), .C(new_new_n221_), .Y(new_new_n267_));
  NO3        g245(.A(i_12_), .B(new_new_n217_), .C(new_new_n37_), .Y(new_new_n268_));
  INV        g246(.A(new_new_n268_), .Y(new_new_n269_));
  NA2        g247(.A(i_8_), .B(new_new_n102_), .Y(new_new_n270_));
  NO3        g248(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n232_), .B(i_0_), .Y(new_new_n272_));
  NA2        g250(.A(i_0_), .B(i_1_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(i_2_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n60_), .B(i_6_), .Y(new_new_n275_));
  NA3        g253(.A(new_new_n275_), .B(new_new_n274_), .C(new_new_n161_), .Y(new_new_n276_));
  NO2        g254(.A(i_3_), .B(i_10_), .Y(new_new_n277_));
  NA3        g255(.A(new_new_n277_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n278_));
  NO2        g256(.A(i_2_), .B(new_new_n102_), .Y(new_new_n279_));
  NO2        g257(.A(i_4_), .B(i_8_), .Y(new_new_n280_));
  NOi21      g258(.An(new_new_n210_), .B(new_new_n104_), .Y(new_new_n281_));
  NA3        g259(.A(new_new_n281_), .B(new_new_n280_), .C(new_new_n279_), .Y(new_new_n282_));
  AN2        g260(.A(i_3_), .B(i_10_), .Y(new_new_n283_));
  NA4        g261(.A(new_new_n283_), .B(new_new_n190_), .C(new_new_n171_), .D(new_new_n169_), .Y(new_new_n284_));
  NO2        g262(.A(i_5_), .B(new_new_n37_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n286_));
  OR2        g264(.A(new_new_n282_), .B(new_new_n278_), .Y(new_new_n287_));
  OAI220     g265(.A0(new_new_n287_), .A1(i_6_), .B0(new_new_n276_), .B1(new_new_n269_), .Y(new_new_n288_));
  NO4        g266(.A(new_new_n288_), .B(new_new_n267_), .C(new_new_n206_), .D(new_new_n163_), .Y(new_new_n289_));
  NO3        g267(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n291_));
  NO3        g269(.A(i_6_), .B(new_new_n185_), .C(i_7_), .Y(new_new_n292_));
  NO2        g270(.A(i_2_), .B(i_3_), .Y(new_new_n293_));
  OR2        g271(.A(i_0_), .B(i_5_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n210_), .B(new_new_n294_), .Y(new_new_n295_));
  NA4        g273(.A(new_new_n295_), .B(new_new_n226_), .C(new_new_n293_), .D(i_1_), .Y(new_new_n296_));
  NAi21      g274(.An(i_8_), .B(i_7_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n297_), .B(i_6_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n156_), .B(new_new_n47_), .Y(new_new_n299_));
  NA3        g277(.A(new_new_n299_), .B(new_new_n298_), .C(new_new_n161_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n300_), .B(new_new_n296_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n301_), .B(i_4_), .Y(new_new_n302_));
  NO2        g280(.A(i_12_), .B(i_10_), .Y(new_new_n303_));
  NOi21      g281(.An(i_5_), .B(i_0_), .Y(new_new_n304_));
  NO2        g282(.A(i_6_), .B(i_8_), .Y(new_new_n305_));
  NOi21      g283(.An(i_0_), .B(i_2_), .Y(new_new_n306_));
  AN2        g284(.A(new_new_n306_), .B(new_new_n305_), .Y(new_new_n307_));
  NO2        g285(.A(i_1_), .B(i_7_), .Y(new_new_n308_));
  AO220      g286(.A0(new_new_n308_), .A1(new_new_n307_), .B0(new_new_n298_), .B1(new_new_n227_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n309_), .B(new_new_n42_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n310_), .B(new_new_n302_), .Y(new_new_n311_));
  NO3        g289(.A(new_new_n225_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n312_));
  NO3        g290(.A(new_new_n297_), .B(i_2_), .C(i_1_), .Y(new_new_n313_));
  OAI210     g291(.A0(new_new_n313_), .A1(new_new_n312_), .B0(i_6_), .Y(new_new_n314_));
  INV        g292(.A(new_new_n314_), .Y(new_new_n315_));
  NOi21      g293(.An(new_new_n152_), .B(new_new_n105_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n316_), .B(new_new_n122_), .Y(new_new_n317_));
  OAI210     g295(.A0(new_new_n317_), .A1(new_new_n315_), .B0(i_3_), .Y(new_new_n318_));
  NO2        g296(.A(new_new_n273_), .B(new_new_n82_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n319_), .B(new_new_n130_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n94_), .B(new_new_n185_), .Y(new_new_n321_));
  NA3        g299(.A(new_new_n281_), .B(new_new_n321_), .C(new_new_n64_), .Y(new_new_n322_));
  AOI210     g300(.A0(new_new_n322_), .A1(new_new_n320_), .B0(i_7_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n185_), .B(i_9_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n324_), .B(new_new_n197_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n325_), .B(new_new_n47_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n326_), .B(new_new_n323_), .Y(new_new_n327_));
  AOI210     g305(.A0(new_new_n327_), .A1(new_new_n318_), .B0(new_new_n160_), .Y(new_new_n328_));
  AOI210     g306(.A0(new_new_n311_), .A1(new_new_n290_), .B0(new_new_n328_), .Y(new_new_n329_));
  NOi32      g307(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n330_));
  INV        g308(.A(new_new_n330_), .Y(new_new_n331_));
  NAi21      g309(.An(i_0_), .B(i_6_), .Y(new_new_n332_));
  NAi21      g310(.An(i_1_), .B(i_5_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n333_), .B(new_new_n332_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n25_), .Y(new_new_n335_));
  OAI210     g313(.A0(new_new_n335_), .A1(new_new_n158_), .B0(new_new_n238_), .Y(new_new_n336_));
  NAi41      g314(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n337_));
  OAI220     g315(.A0(new_new_n337_), .A1(new_new_n333_), .B0(new_new_n213_), .B1(new_new_n158_), .Y(new_new_n338_));
  AOI210     g316(.A0(new_new_n337_), .A1(new_new_n158_), .B0(new_new_n156_), .Y(new_new_n339_));
  NOi32      g317(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n340_));
  NAi21      g318(.An(i_6_), .B(i_1_), .Y(new_new_n341_));
  NA3        g319(.A(new_new_n341_), .B(new_new_n340_), .C(new_new_n47_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n342_), .B(i_0_), .Y(new_new_n343_));
  OR3        g321(.A(new_new_n343_), .B(new_new_n339_), .C(new_new_n338_), .Y(new_new_n344_));
  NO2        g322(.A(i_1_), .B(new_new_n102_), .Y(new_new_n345_));
  NAi21      g323(.An(i_3_), .B(i_4_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n346_), .B(i_9_), .Y(new_new_n347_));
  AN2        g325(.A(i_6_), .B(i_7_), .Y(new_new_n348_));
  OAI210     g326(.A0(new_new_n348_), .A1(new_new_n345_), .B0(new_new_n347_), .Y(new_new_n349_));
  NA2        g327(.A(i_2_), .B(i_7_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n346_), .B(i_10_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n349_), .B(new_new_n177_), .Y(new_new_n352_));
  AOI210     g330(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n353_));
  OAI210     g331(.A0(new_new_n353_), .A1(new_new_n180_), .B0(new_new_n351_), .Y(new_new_n354_));
  AOI220     g332(.A0(new_new_n351_), .A1(new_new_n308_), .B0(new_new_n231_), .B1(new_new_n180_), .Y(new_new_n355_));
  AOI210     g333(.A0(new_new_n355_), .A1(new_new_n354_), .B0(i_5_), .Y(new_new_n356_));
  NO4        g334(.A(new_new_n356_), .B(new_new_n352_), .C(new_new_n344_), .D(new_new_n336_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(new_new_n331_), .Y(new_new_n358_));
  AN2        g336(.A(i_12_), .B(i_5_), .Y(new_new_n359_));
  NO2        g337(.A(i_11_), .B(i_6_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n235_), .B(i_5_), .Y(new_new_n361_));
  NO2        g339(.A(i_5_), .B(i_10_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n363_));
  NO3        g341(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n364_));
  NO2        g342(.A(i_11_), .B(i_12_), .Y(new_new_n365_));
  NA3        g343(.A(new_new_n114_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n366_), .B(new_new_n213_), .Y(new_new_n367_));
  NAi21      g345(.An(i_13_), .B(i_0_), .Y(new_new_n368_));
  INV        g346(.A(new_new_n368_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n367_), .B(new_new_n369_), .Y(new_new_n370_));
  INV        g348(.A(new_new_n370_), .Y(new_new_n371_));
  NO3        g349(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n372_));
  NO2        g350(.A(i_0_), .B(i_11_), .Y(new_new_n373_));
  INV        g351(.A(i_5_), .Y(new_new_n374_));
  AN2        g352(.A(i_1_), .B(i_6_), .Y(new_new_n375_));
  NOi21      g353(.An(i_2_), .B(i_12_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n377_), .B(new_new_n374_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n140_), .B(i_9_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(i_4_), .Y(new_new_n380_));
  NA2        g358(.A(new_new_n378_), .B(new_new_n380_), .Y(new_new_n381_));
  NAi21      g359(.An(i_9_), .B(i_4_), .Y(new_new_n382_));
  OR2        g360(.A(i_13_), .B(i_10_), .Y(new_new_n383_));
  NO3        g361(.A(new_new_n383_), .B(new_new_n117_), .C(new_new_n382_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n167_), .B(new_new_n121_), .Y(new_new_n385_));
  OR2        g363(.A(new_new_n208_), .B(new_new_n207_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n268_), .B(new_new_n387_), .Y(new_new_n388_));
  NA2        g366(.A(i_5_), .B(new_new_n202_), .Y(new_new_n389_));
  OAI220     g367(.A0(new_new_n389_), .A1(new_new_n386_), .B0(new_new_n388_), .B1(new_new_n316_), .Y(new_new_n390_));
  INV        g368(.A(new_new_n390_), .Y(new_new_n391_));
  AOI210     g369(.A0(new_new_n391_), .A1(new_new_n381_), .B0(new_new_n26_), .Y(new_new_n392_));
  INV        g370(.A(new_new_n296_), .Y(new_new_n393_));
  AOI220     g371(.A0(new_new_n275_), .A1(new_new_n271_), .B0(new_new_n272_), .B1(new_new_n291_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n394_), .B(i_5_), .Y(new_new_n395_));
  AOI220     g373(.A0(i_3_), .A1(new_new_n274_), .B0(new_new_n263_), .B1(new_new_n202_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n396_), .B(new_new_n270_), .Y(new_new_n397_));
  NO3        g375(.A(new_new_n397_), .B(new_new_n395_), .C(new_new_n393_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n188_), .B(new_new_n98_), .Y(new_new_n399_));
  NA3        g377(.A(new_new_n299_), .B(new_new_n161_), .C(new_new_n87_), .Y(new_new_n400_));
  AOI210     g378(.A0(new_new_n400_), .A1(new_new_n399_), .B0(new_new_n297_), .Y(new_new_n401_));
  NA3        g379(.A(new_new_n308_), .B(new_new_n307_), .C(i_5_), .Y(new_new_n402_));
  INV        g380(.A(new_new_n292_), .Y(new_new_n403_));
  OAI210     g381(.A0(new_new_n403_), .A1(new_new_n181_), .B0(new_new_n402_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n404_), .B(new_new_n401_), .Y(new_new_n405_));
  AOI210     g383(.A0(new_new_n405_), .A1(new_new_n398_), .B0(new_new_n256_), .Y(new_new_n406_));
  NO4        g384(.A(new_new_n406_), .B(new_new_n392_), .C(new_new_n371_), .D(new_new_n358_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n64_), .B(i_4_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n74_), .B(i_13_), .Y(new_new_n409_));
  NO2        g387(.A(i_10_), .B(i_9_), .Y(new_new_n410_));
  NAi21      g388(.An(i_12_), .B(i_8_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(i_3_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n286_), .B(i_0_), .Y(new_new_n413_));
  NO3        g391(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n251_), .B(new_new_n99_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(new_new_n414_), .Y(new_new_n416_));
  NA2        g394(.A(i_8_), .B(i_9_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n268_), .B(new_new_n197_), .Y(new_new_n418_));
  OAI220     g396(.A0(new_new_n418_), .A1(new_new_n417_), .B0(new_new_n416_), .B1(new_new_n413_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n243_), .B(new_new_n285_), .Y(new_new_n420_));
  NO3        g398(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n421_));
  INV        g399(.A(new_new_n421_), .Y(new_new_n422_));
  NA3        g400(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n423_));
  NA4        g401(.A(new_new_n143_), .B(new_new_n116_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n424_));
  OAI220     g402(.A0(new_new_n424_), .A1(new_new_n423_), .B0(new_new_n422_), .B1(new_new_n420_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(new_new_n419_), .Y(new_new_n426_));
  OR2        g404(.A(new_new_n273_), .B(new_new_n199_), .Y(new_new_n427_));
  OA210      g405(.A0(new_new_n325_), .A1(new_new_n102_), .B0(new_new_n276_), .Y(new_new_n428_));
  OA220      g406(.A0(new_new_n428_), .A1(new_new_n160_), .B0(new_new_n427_), .B1(new_new_n224_), .Y(new_new_n429_));
  NO2        g407(.A(i_2_), .B(i_13_), .Y(new_new_n430_));
  NO3        g408(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n431_));
  NO2        g409(.A(i_6_), .B(i_7_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n433_));
  NO2        g411(.A(i_11_), .B(i_1_), .Y(new_new_n434_));
  OR2        g412(.A(i_11_), .B(i_8_), .Y(new_new_n435_));
  NOi21      g413(.An(i_2_), .B(i_7_), .Y(new_new_n436_));
  NAi31      g414(.An(new_new_n435_), .B(new_new_n436_), .C(i_0_), .Y(new_new_n437_));
  INV        g415(.A(new_new_n383_), .Y(new_new_n438_));
  NA3        g416(.A(new_new_n438_), .B(new_new_n408_), .C(new_new_n76_), .Y(new_new_n439_));
  NO2        g417(.A(new_new_n439_), .B(new_new_n437_), .Y(new_new_n440_));
  NO2        g418(.A(i_3_), .B(new_new_n185_), .Y(new_new_n441_));
  NO2        g419(.A(i_6_), .B(i_10_), .Y(new_new_n442_));
  NA4        g420(.A(new_new_n442_), .B(new_new_n290_), .C(new_new_n441_), .D(new_new_n229_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n443_), .B(new_new_n154_), .Y(new_new_n444_));
  NA3        g422(.A(new_new_n237_), .B(new_new_n166_), .C(new_new_n130_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n156_), .B(i_3_), .Y(new_new_n447_));
  NAi31      g425(.An(new_new_n446_), .B(new_new_n447_), .C(new_new_n218_), .Y(new_new_n448_));
  NA3        g426(.A(new_new_n363_), .B(new_new_n174_), .C(new_new_n147_), .Y(new_new_n449_));
  NA3        g427(.A(new_new_n449_), .B(new_new_n448_), .C(new_new_n445_), .Y(new_new_n450_));
  NO3        g428(.A(new_new_n450_), .B(new_new_n444_), .C(new_new_n440_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n414_), .B(new_new_n359_), .Y(new_new_n452_));
  NAi21      g430(.An(new_new_n208_), .B(new_new_n365_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n308_), .B(new_new_n210_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n26_), .B(i_5_), .Y(new_new_n455_));
  NO2        g433(.A(i_0_), .B(new_new_n87_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n456_), .B(new_new_n455_), .C(new_new_n140_), .Y(new_new_n457_));
  OR3        g435(.A(i_4_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n458_));
  OAI220     g436(.A0(new_new_n458_), .A1(new_new_n457_), .B0(new_new_n454_), .B1(new_new_n453_), .Y(new_new_n459_));
  NA4        g437(.A(new_new_n283_), .B(new_new_n216_), .C(new_new_n74_), .D(new_new_n229_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n460_), .B(new_new_n433_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n461_), .B(new_new_n459_), .Y(new_new_n462_));
  NA4        g440(.A(new_new_n462_), .B(new_new_n451_), .C(new_new_n429_), .D(new_new_n426_), .Y(new_new_n463_));
  NA3        g441(.A(new_new_n283_), .B(new_new_n171_), .C(new_new_n169_), .Y(new_new_n464_));
  INV        g442(.A(new_new_n464_), .Y(new_new_n465_));
  BUFFER     g443(.A(new_new_n226_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n466_), .B(new_new_n465_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n290_), .B(i_0_), .Y(new_new_n468_));
  OAI210     g446(.A0(new_new_n468_), .A1(new_new_n224_), .B0(new_new_n284_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n469_), .B(new_new_n298_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n359_), .B(new_new_n217_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n330_), .B(new_new_n74_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n348_), .B(new_new_n340_), .Y(new_new_n473_));
  OR2        g451(.A(new_new_n471_), .B(new_new_n473_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n36_), .B(i_8_), .Y(new_new_n475_));
  NAi41      g453(.An(new_new_n472_), .B(new_new_n442_), .C(new_new_n475_), .D(new_new_n47_), .Y(new_new_n476_));
  AOI210     g454(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n384_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n477_), .B(new_new_n476_), .C(new_new_n474_), .Y(new_new_n478_));
  INV        g456(.A(new_new_n478_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n248_), .B(new_new_n65_), .Y(new_new_n480_));
  OAI210     g458(.A0(i_8_), .A1(new_new_n480_), .B0(new_new_n132_), .Y(new_new_n481_));
  AOI210     g459(.A0(new_new_n186_), .A1(i_9_), .B0(new_new_n250_), .Y(new_new_n482_));
  NO2        g460(.A(new_new_n482_), .B(new_new_n191_), .Y(new_new_n483_));
  OR2        g461(.A(new_new_n176_), .B(i_4_), .Y(new_new_n484_));
  INV        g462(.A(new_new_n484_), .Y(new_new_n485_));
  AOI220     g463(.A0(new_new_n485_), .A1(new_new_n483_), .B0(new_new_n481_), .B1(new_new_n385_), .Y(new_new_n486_));
  NA4        g464(.A(new_new_n486_), .B(new_new_n479_), .C(new_new_n470_), .D(new_new_n467_), .Y(new_new_n487_));
  NA2        g465(.A(new_new_n361_), .B(new_new_n274_), .Y(new_new_n488_));
  OAI210     g466(.A0(new_new_n972_), .A1(new_new_n164_), .B0(new_new_n488_), .Y(new_new_n489_));
  NO2        g467(.A(i_12_), .B(new_new_n185_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(new_new_n217_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n442_), .B(new_new_n27_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n492_), .B(new_new_n491_), .Y(new_new_n493_));
  NOi31      g471(.An(new_new_n292_), .B(new_new_n383_), .C(new_new_n38_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n494_), .A1(new_new_n493_), .B0(new_new_n489_), .Y(new_new_n495_));
  AOI220     g473(.A0(new_new_n299_), .A1(new_new_n40_), .B0(new_new_n227_), .B1(new_new_n198_), .Y(new_new_n496_));
  NO2        g474(.A(new_new_n496_), .B(new_new_n484_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n45_), .B(i_10_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(i_6_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n499_), .B(new_new_n497_), .Y(new_new_n500_));
  NOi31      g478(.An(new_new_n272_), .B(new_new_n278_), .C(new_new_n175_), .Y(new_new_n501_));
  NA3        g479(.A(new_new_n283_), .B(new_new_n169_), .C(new_new_n98_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n156_), .B(i_5_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n503_), .B(new_new_n293_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n504_), .B(new_new_n502_), .Y(new_new_n505_));
  OAI210     g483(.A0(new_new_n505_), .A1(new_new_n501_), .B0(new_new_n421_), .Y(new_new_n506_));
  NA3        g484(.A(new_new_n506_), .B(new_new_n500_), .C(new_new_n495_), .Y(new_new_n507_));
  NA3        g485(.A(new_new_n210_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n268_), .B(new_new_n85_), .Y(new_new_n509_));
  AOI210     g487(.A0(new_new_n508_), .A1(new_new_n320_), .B0(new_new_n509_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n275_), .B(new_new_n271_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n511_), .B(new_new_n168_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n410_), .B(new_new_n214_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n513_), .B(new_new_n514_), .Y(new_new_n515_));
  AOI210     g493(.A0(new_new_n341_), .A1(new_new_n47_), .B0(new_new_n345_), .Y(new_new_n516_));
  NA2        g494(.A(i_0_), .B(new_new_n49_), .Y(new_new_n517_));
  NA3        g495(.A(new_new_n490_), .B(new_new_n260_), .C(new_new_n517_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n516_), .B(new_new_n518_), .Y(new_new_n519_));
  NO4        g497(.A(new_new_n519_), .B(new_new_n515_), .C(new_new_n512_), .D(new_new_n510_), .Y(new_new_n520_));
  NO4        g498(.A(new_new_n244_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n521_));
  NO3        g499(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n225_), .B(new_new_n36_), .Y(new_new_n523_));
  AN2        g501(.A(new_new_n523_), .B(new_new_n522_), .Y(new_new_n524_));
  OA210      g502(.A0(new_new_n524_), .A1(new_new_n521_), .B0(new_new_n330_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n383_), .B(i_1_), .Y(new_new_n526_));
  NOi31      g504(.An(new_new_n526_), .B(new_new_n415_), .C(new_new_n74_), .Y(new_new_n527_));
  AN4        g505(.A(new_new_n527_), .B(new_new_n380_), .C(new_new_n455_), .D(i_2_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n394_), .B(new_new_n172_), .Y(new_new_n529_));
  NO3        g507(.A(new_new_n529_), .B(new_new_n528_), .C(new_new_n525_), .Y(new_new_n530_));
  NOi21      g508(.An(i_10_), .B(i_6_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n532_));
  AOI220     g510(.A0(new_new_n268_), .A1(new_new_n532_), .B0(new_new_n260_), .B1(new_new_n531_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n533_), .B(new_new_n413_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n535_));
  INV        g513(.A(new_new_n534_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n472_), .B(new_new_n355_), .Y(new_new_n537_));
  INV        g515(.A(new_new_n293_), .Y(new_new_n538_));
  NO2        g516(.A(i_12_), .B(new_new_n87_), .Y(new_new_n539_));
  NA3        g517(.A(new_new_n539_), .B(new_new_n260_), .C(new_new_n517_), .Y(new_new_n540_));
  NA3        g518(.A(new_new_n360_), .B(new_new_n268_), .C(new_new_n210_), .Y(new_new_n541_));
  AOI210     g519(.A0(new_new_n541_), .A1(new_new_n540_), .B0(new_new_n538_), .Y(new_new_n542_));
  NO3        g520(.A(i_4_), .B(new_new_n314_), .C(new_new_n278_), .Y(new_new_n543_));
  OR2        g521(.A(i_2_), .B(i_5_), .Y(new_new_n544_));
  OR2        g522(.A(new_new_n544_), .B(new_new_n375_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n545_), .B(new_new_n453_), .Y(new_new_n546_));
  NO4        g524(.A(new_new_n546_), .B(new_new_n543_), .C(new_new_n542_), .D(new_new_n537_), .Y(new_new_n547_));
  NA4        g525(.A(new_new_n547_), .B(new_new_n536_), .C(new_new_n530_), .D(new_new_n520_), .Y(new_new_n548_));
  NO4        g526(.A(new_new_n548_), .B(new_new_n507_), .C(new_new_n487_), .D(new_new_n463_), .Y(new_new_n549_));
  NA4        g527(.A(new_new_n549_), .B(new_new_n407_), .C(new_new_n329_), .D(new_new_n289_), .Y(mai7));
  NO2        g528(.A(new_new_n94_), .B(new_new_n55_), .Y(new_new_n551_));
  NA2        g529(.A(i_11_), .B(new_new_n185_), .Y(new_new_n552_));
  NA3        g530(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n229_), .B(i_4_), .Y(new_new_n554_));
  NA2        g532(.A(new_new_n554_), .B(i_8_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n106_), .B(new_new_n553_), .Y(new_new_n556_));
  NA2        g534(.A(i_2_), .B(new_new_n87_), .Y(new_new_n557_));
  OAI210     g535(.A0(new_new_n88_), .A1(new_new_n195_), .B0(new_new_n196_), .Y(new_new_n558_));
  NO2        g536(.A(i_7_), .B(new_new_n37_), .Y(new_new_n559_));
  NA2        g537(.A(i_4_), .B(i_8_), .Y(new_new_n560_));
  AOI210     g538(.A0(new_new_n560_), .A1(new_new_n283_), .B0(new_new_n559_), .Y(new_new_n561_));
  OAI220     g539(.A0(new_new_n561_), .A1(new_new_n557_), .B0(new_new_n558_), .B1(i_13_), .Y(new_new_n562_));
  NO3        g540(.A(new_new_n562_), .B(new_new_n556_), .C(new_new_n551_), .Y(new_new_n563_));
  INV        g541(.A(new_new_n159_), .Y(new_new_n564_));
  OR2        g542(.A(i_6_), .B(i_10_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n565_), .B(new_new_n23_), .Y(new_new_n566_));
  OR3        g544(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n567_));
  NO3        g545(.A(new_new_n567_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n568_));
  INV        g546(.A(new_new_n192_), .Y(new_new_n569_));
  NO2        g547(.A(new_new_n568_), .B(new_new_n566_), .Y(new_new_n570_));
  OA220      g548(.A0(new_new_n570_), .A1(new_new_n538_), .B0(new_new_n564_), .B1(new_new_n252_), .Y(new_new_n571_));
  AOI210     g549(.A0(new_new_n571_), .A1(new_new_n563_), .B0(new_new_n64_), .Y(new_new_n572_));
  NOi21      g550(.An(i_11_), .B(i_7_), .Y(new_new_n573_));
  AO210      g551(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n574_), .B(new_new_n573_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n575_), .B(new_new_n198_), .Y(new_new_n576_));
  NA3        g554(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n577_));
  NAi31      g555(.An(new_new_n577_), .B(new_new_n207_), .C(i_11_), .Y(new_new_n578_));
  AOI210     g556(.A0(new_new_n578_), .A1(new_new_n576_), .B0(new_new_n64_), .Y(new_new_n579_));
  NO3        g557(.A(i_7_), .B(new_new_n200_), .C(new_new_n552_), .Y(new_new_n580_));
  OAI210     g558(.A0(new_new_n580_), .A1(new_new_n218_), .B0(new_new_n64_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n64_), .B(i_9_), .Y(new_new_n582_));
  NO2        g560(.A(i_1_), .B(i_12_), .Y(new_new_n583_));
  NA3        g561(.A(new_new_n583_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n584_));
  BUFFER     g562(.A(new_new_n584_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n585_), .B(new_new_n581_), .Y(new_new_n586_));
  OAI210     g564(.A0(new_new_n586_), .A1(new_new_n579_), .B0(i_6_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n577_), .B(new_new_n109_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(new_new_n539_), .Y(new_new_n589_));
  NO2        g567(.A(i_6_), .B(i_11_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n589_), .B(new_new_n416_), .Y(new_new_n591_));
  NO4        g569(.A(new_new_n207_), .B(new_new_n126_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n592_), .B(new_new_n582_), .Y(new_new_n593_));
  NA2        g571(.A(new_new_n229_), .B(i_6_), .Y(new_new_n594_));
  INV        g572(.A(new_new_n593_), .Y(new_new_n595_));
  INV        g573(.A(i_2_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n136_), .B(i_9_), .Y(new_new_n597_));
  NA3        g575(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n47_), .B(i_1_), .Y(new_new_n599_));
  NA3        g577(.A(new_new_n599_), .B(new_new_n251_), .C(new_new_n45_), .Y(new_new_n600_));
  OAI220     g578(.A0(new_new_n600_), .A1(new_new_n598_), .B0(new_new_n597_), .B1(new_new_n596_), .Y(new_new_n601_));
  NA3        g579(.A(new_new_n582_), .B(new_new_n293_), .C(i_6_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n602_), .B(new_new_n23_), .Y(new_new_n603_));
  AOI210     g581(.A0(new_new_n434_), .A1(new_new_n387_), .B0(new_new_n234_), .Y(new_new_n604_));
  NO2        g582(.A(new_new_n604_), .B(new_new_n557_), .Y(new_new_n605_));
  NO2        g583(.A(i_11_), .B(new_new_n37_), .Y(new_new_n606_));
  OR3        g584(.A(new_new_n605_), .B(new_new_n603_), .C(new_new_n601_), .Y(new_new_n607_));
  NO3        g585(.A(new_new_n607_), .B(new_new_n595_), .C(new_new_n591_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n229_), .B(new_new_n102_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n609_), .B(new_new_n573_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(i_1_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n611_), .B(new_new_n567_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n382_), .B(new_new_n87_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n612_), .B(new_new_n47_), .Y(new_new_n614_));
  NA2        g592(.A(i_3_), .B(new_new_n185_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(new_new_n115_), .Y(new_new_n616_));
  AN2        g594(.A(new_new_n616_), .B(new_new_n499_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n225_), .B(new_new_n45_), .Y(new_new_n618_));
  NO3        g596(.A(new_new_n618_), .B(new_new_n286_), .C(new_new_n230_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n620_), .B(i_6_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n87_), .B(i_9_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n622_), .B(new_new_n64_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n623_), .B(new_new_n583_), .Y(new_new_n624_));
  NO4        g602(.A(new_new_n624_), .B(new_new_n621_), .C(new_new_n619_), .D(i_4_), .Y(new_new_n625_));
  NA2        g603(.A(i_1_), .B(i_3_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n417_), .B(new_new_n94_), .Y(new_new_n627_));
  AOI210     g605(.A0(new_new_n618_), .A1(new_new_n531_), .B0(new_new_n627_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n626_), .Y(new_new_n629_));
  NO3        g607(.A(new_new_n629_), .B(new_new_n625_), .C(new_new_n617_), .Y(new_new_n630_));
  NA4        g608(.A(new_new_n630_), .B(new_new_n614_), .C(new_new_n608_), .D(new_new_n587_), .Y(new_new_n631_));
  NO3        g609(.A(new_new_n435_), .B(i_3_), .C(i_7_), .Y(new_new_n632_));
  NOi21      g610(.An(new_new_n632_), .B(i_10_), .Y(new_new_n633_));
  OA210      g611(.A0(new_new_n633_), .A1(new_new_n237_), .B0(new_new_n87_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n348_), .B(new_new_n347_), .Y(new_new_n635_));
  NA3        g613(.A(new_new_n159_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n636_), .B(new_new_n635_), .Y(new_new_n637_));
  OAI210     g615(.A0(new_new_n637_), .A1(new_new_n634_), .B0(i_1_), .Y(new_new_n638_));
  AOI210     g616(.A0(new_new_n251_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n346_), .B(i_2_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n640_), .B(new_new_n639_), .Y(new_new_n641_));
  OAI210     g619(.A0(new_new_n602_), .A1(new_new_n411_), .B0(new_new_n641_), .Y(new_new_n642_));
  INV        g620(.A(new_new_n642_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n643_), .A1(new_new_n638_), .B0(i_13_), .Y(new_new_n644_));
  OR2        g622(.A(i_11_), .B(i_7_), .Y(new_new_n645_));
  NA3        g623(.A(new_new_n645_), .B(new_new_n107_), .C(new_new_n136_), .Y(new_new_n646_));
  AOI220     g624(.A0(new_new_n430_), .A1(new_new_n159_), .B0(i_2_), .B1(new_new_n136_), .Y(new_new_n647_));
  OAI210     g625(.A0(new_new_n647_), .A1(new_new_n45_), .B0(new_new_n646_), .Y(new_new_n648_));
  NO2        g626(.A(new_new_n55_), .B(i_12_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n436_), .B(new_new_n24_), .Y(new_new_n650_));
  AOI220     g628(.A0(new_new_n650_), .A1(new_new_n613_), .B0(new_new_n237_), .B1(new_new_n129_), .Y(new_new_n651_));
  OAI220     g629(.A0(new_new_n651_), .A1(new_new_n41_), .B0(new_new_n971_), .B1(new_new_n94_), .Y(new_new_n652_));
  AOI210     g630(.A0(new_new_n648_), .A1(new_new_n305_), .B0(new_new_n652_), .Y(new_new_n653_));
  INV        g631(.A(new_new_n115_), .Y(new_new_n654_));
  AOI220     g632(.A0(new_new_n654_), .A1(new_new_n73_), .B0(new_new_n360_), .B1(new_new_n599_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n655_), .B(new_new_n235_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n125_), .B(i_13_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n598_), .B(new_new_n115_), .Y(new_new_n658_));
  INV        g636(.A(new_new_n658_), .Y(new_new_n659_));
  OAI220     g637(.A0(new_new_n659_), .A1(new_new_n72_), .B0(new_new_n657_), .B1(new_new_n639_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n26_), .B(new_new_n185_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n661_), .B(i_7_), .Y(new_new_n662_));
  NO3        g640(.A(new_new_n436_), .B(new_new_n229_), .C(new_new_n87_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n663_), .B(new_new_n662_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n93_), .B(new_new_n103_), .Y(new_new_n665_));
  OAI220     g643(.A0(new_new_n665_), .A1(new_new_n555_), .B0(new_new_n664_), .B1(new_new_n569_), .Y(new_new_n666_));
  NO3        g644(.A(new_new_n666_), .B(new_new_n660_), .C(new_new_n656_), .Y(new_new_n667_));
  OR2        g645(.A(i_11_), .B(i_6_), .Y(new_new_n668_));
  NA3        g646(.A(new_new_n554_), .B(new_new_n661_), .C(i_7_), .Y(new_new_n669_));
  AOI210     g647(.A0(new_new_n669_), .A1(new_new_n659_), .B0(new_new_n668_), .Y(new_new_n670_));
  NA3        g648(.A(new_new_n376_), .B(new_new_n559_), .C(new_new_n99_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n590_), .B(i_13_), .Y(new_new_n672_));
  NAi21      g650(.An(i_11_), .B(i_12_), .Y(new_new_n673_));
  NOi41      g651(.An(new_new_n112_), .B(new_new_n673_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n674_));
  NO3        g652(.A(new_new_n436_), .B(new_new_n539_), .C(new_new_n560_), .Y(new_new_n675_));
  AOI210     g653(.A0(new_new_n675_), .A1(new_new_n290_), .B0(new_new_n674_), .Y(new_new_n676_));
  NA3        g654(.A(new_new_n676_), .B(new_new_n672_), .C(new_new_n671_), .Y(new_new_n677_));
  OAI210     g655(.A0(new_new_n677_), .A1(new_new_n670_), .B0(new_new_n64_), .Y(new_new_n678_));
  NO2        g656(.A(i_2_), .B(i_12_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n345_), .B(new_new_n679_), .Y(new_new_n680_));
  NO3        g658(.A(i_9_), .B(i_3_), .C(new_new_n554_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n681_), .B(new_new_n345_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n682_), .B(new_new_n680_), .Y(new_new_n683_));
  NA3        g661(.A(new_new_n683_), .B(new_new_n46_), .C(new_new_n217_), .Y(new_new_n684_));
  NA4        g662(.A(new_new_n684_), .B(new_new_n678_), .C(new_new_n667_), .D(new_new_n653_), .Y(new_new_n685_));
  OR4        g663(.A(new_new_n685_), .B(new_new_n644_), .C(new_new_n631_), .D(new_new_n572_), .Y(mai5));
  NA2        g664(.A(new_new_n610_), .B(new_new_n254_), .Y(new_new_n687_));
  AN2        g665(.A(new_new_n24_), .B(i_10_), .Y(new_new_n688_));
  NA3        g666(.A(new_new_n688_), .B(new_new_n679_), .C(new_new_n109_), .Y(new_new_n689_));
  NO2        g667(.A(new_new_n555_), .B(i_11_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n88_), .B(new_new_n690_), .Y(new_new_n691_));
  NA3        g669(.A(new_new_n691_), .B(new_new_n689_), .C(new_new_n687_), .Y(new_new_n692_));
  NO3        g670(.A(i_11_), .B(new_new_n229_), .C(i_13_), .Y(new_new_n693_));
  NO2        g671(.A(new_new_n122_), .B(new_new_n23_), .Y(new_new_n694_));
  NA2        g672(.A(i_12_), .B(i_8_), .Y(new_new_n695_));
  OAI210     g673(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n695_), .Y(new_new_n696_));
  INV        g674(.A(new_new_n410_), .Y(new_new_n697_));
  AOI220     g675(.A0(new_new_n293_), .A1(new_new_n535_), .B0(new_new_n696_), .B1(new_new_n694_), .Y(new_new_n698_));
  INV        g676(.A(new_new_n698_), .Y(new_new_n699_));
  NO2        g677(.A(new_new_n699_), .B(new_new_n692_), .Y(new_new_n700_));
  INV        g678(.A(new_new_n166_), .Y(new_new_n701_));
  INV        g679(.A(new_new_n237_), .Y(new_new_n702_));
  OAI210     g680(.A0(new_new_n640_), .A1(new_new_n412_), .B0(new_new_n112_), .Y(new_new_n703_));
  AOI210     g681(.A0(new_new_n703_), .A1(new_new_n702_), .B0(new_new_n701_), .Y(new_new_n704_));
  NO2        g682(.A(new_new_n417_), .B(new_new_n26_), .Y(new_new_n705_));
  NO2        g683(.A(new_new_n705_), .B(new_new_n387_), .Y(new_new_n706_));
  NA2        g684(.A(new_new_n706_), .B(i_2_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n707_), .Y(new_new_n708_));
  AOI210     g686(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n383_), .Y(new_new_n709_));
  AOI210     g687(.A0(new_new_n709_), .A1(new_new_n708_), .B0(new_new_n704_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n182_), .B(new_new_n123_), .Y(new_new_n711_));
  OAI210     g689(.A0(new_new_n711_), .A1(new_new_n694_), .B0(i_2_), .Y(new_new_n712_));
  INV        g690(.A(new_new_n167_), .Y(new_new_n713_));
  NO3        g691(.A(new_new_n574_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n714_));
  AOI210     g692(.A0(new_new_n713_), .A1(new_new_n88_), .B0(new_new_n714_), .Y(new_new_n715_));
  AOI210     g693(.A0(new_new_n715_), .A1(new_new_n712_), .B0(new_new_n185_), .Y(new_new_n716_));
  OA210      g694(.A0(new_new_n575_), .A1(new_new_n124_), .B0(i_13_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n192_), .B(new_new_n195_), .Y(new_new_n718_));
  NA2        g696(.A(new_new_n150_), .B(new_new_n552_), .Y(new_new_n719_));
  AOI210     g697(.A0(new_new_n719_), .A1(new_new_n718_), .B0(new_new_n350_), .Y(new_new_n720_));
  AOI210     g698(.A0(new_new_n200_), .A1(new_new_n146_), .B0(new_new_n475_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n721_), .B(new_new_n387_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n103_), .B(new_new_n45_), .Y(new_new_n723_));
  INV        g701(.A(new_new_n279_), .Y(new_new_n724_));
  NA4        g702(.A(new_new_n724_), .B(new_new_n283_), .C(new_new_n122_), .D(new_new_n43_), .Y(new_new_n725_));
  OAI210     g703(.A0(new_new_n725_), .A1(new_new_n723_), .B0(new_new_n722_), .Y(new_new_n726_));
  NO4        g704(.A(new_new_n726_), .B(new_new_n720_), .C(new_new_n717_), .D(new_new_n716_), .Y(new_new_n727_));
  NA2        g705(.A(new_new_n535_), .B(new_new_n28_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n693_), .B(new_new_n261_), .Y(new_new_n729_));
  NA2        g707(.A(new_new_n729_), .B(new_new_n728_), .Y(new_new_n730_));
  NO2        g708(.A(new_new_n63_), .B(i_12_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n731_), .B(new_new_n124_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n732_), .B(new_new_n552_), .Y(new_new_n733_));
  AOI220     g711(.A0(new_new_n733_), .A1(new_new_n36_), .B0(new_new_n730_), .B1(new_new_n47_), .Y(new_new_n734_));
  NA4        g712(.A(new_new_n734_), .B(new_new_n727_), .C(new_new_n710_), .D(new_new_n700_), .Y(mai6));
  NA4        g713(.A(new_new_n362_), .B(new_new_n441_), .C(new_new_n72_), .D(new_new_n102_), .Y(new_new_n736_));
  INV        g714(.A(new_new_n736_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n213_), .B(new_new_n446_), .Y(new_new_n738_));
  NO2        g716(.A(i_11_), .B(i_9_), .Y(new_new_n739_));
  NO2        g717(.A(new_new_n737_), .B(new_new_n304_), .Y(new_new_n740_));
  OR2        g718(.A(new_new_n740_), .B(i_12_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n351_), .B(new_new_n308_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n539_), .B(new_new_n64_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n633_), .B(new_new_n72_), .Y(new_new_n744_));
  NA3        g722(.A(new_new_n744_), .B(new_new_n743_), .C(new_new_n742_), .Y(new_new_n745_));
  INV        g723(.A(new_new_n189_), .Y(new_new_n746_));
  AOI220     g724(.A0(new_new_n746_), .A1(new_new_n739_), .B0(new_new_n745_), .B1(new_new_n74_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n303_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n76_), .B(new_new_n129_), .Y(new_new_n749_));
  INV        g727(.A(new_new_n122_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n750_), .B(new_new_n47_), .Y(new_new_n751_));
  AOI210     g729(.A0(new_new_n751_), .A1(new_new_n749_), .B0(new_new_n748_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n32_), .B(i_11_), .Y(new_new_n753_));
  NA3        g731(.A(new_new_n753_), .B(new_new_n432_), .C(new_new_n362_), .Y(new_new_n754_));
  NAi32      g732(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n668_), .B(new_new_n755_), .Y(new_new_n756_));
  OAI210     g734(.A0(new_new_n632_), .A1(new_new_n523_), .B0(new_new_n522_), .Y(new_new_n757_));
  NAi31      g735(.An(new_new_n756_), .B(new_new_n757_), .C(new_new_n754_), .Y(new_new_n758_));
  OR2        g736(.A(new_new_n758_), .B(new_new_n752_), .Y(new_new_n759_));
  NO2        g737(.A(new_new_n645_), .B(i_2_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n761_), .B(new_new_n375_), .Y(new_new_n762_));
  NA2        g740(.A(new_new_n762_), .B(new_new_n760_), .Y(new_new_n763_));
  AO210      g741(.A0(new_new_n334_), .A1(new_new_n324_), .B0(new_new_n364_), .Y(new_new_n764_));
  NA3        g742(.A(new_new_n764_), .B(new_new_n247_), .C(i_7_), .Y(new_new_n765_));
  BUFFER     g743(.A(new_new_n575_), .Y(new_new_n766_));
  NA3        g744(.A(new_new_n766_), .B(new_new_n145_), .C(new_new_n70_), .Y(new_new_n767_));
  OR2        g745(.A(new_new_n697_), .B(new_new_n36_), .Y(new_new_n768_));
  NA4        g746(.A(new_new_n768_), .B(new_new_n767_), .C(new_new_n765_), .D(new_new_n763_), .Y(new_new_n769_));
  NO2        g747(.A(i_6_), .B(i_11_), .Y(new_new_n770_));
  AOI220     g748(.A0(new_new_n770_), .A1(new_new_n522_), .B0(new_new_n738_), .B1(new_new_n662_), .Y(new_new_n771_));
  NA3        g749(.A(new_new_n350_), .B(new_new_n231_), .C(new_new_n145_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n364_), .B(new_new_n71_), .Y(new_new_n773_));
  NA4        g751(.A(new_new_n773_), .B(new_new_n772_), .C(new_new_n771_), .D(new_new_n558_), .Y(new_new_n774_));
  AOI210     g752(.A0(new_new_n412_), .A1(new_new_n410_), .B0(new_new_n521_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n565_), .B(new_new_n103_), .Y(new_new_n776_));
  OAI210     g754(.A0(new_new_n776_), .A1(new_new_n113_), .B0(new_new_n373_), .Y(new_new_n777_));
  INV        g755(.A(new_new_n545_), .Y(new_new_n778_));
  NA3        g756(.A(new_new_n778_), .B(new_new_n303_), .C(i_7_), .Y(new_new_n779_));
  NA3        g757(.A(new_new_n779_), .B(new_new_n777_), .C(new_new_n775_), .Y(new_new_n780_));
  NO4        g758(.A(new_new_n780_), .B(new_new_n774_), .C(new_new_n769_), .D(new_new_n759_), .Y(new_new_n781_));
  NA4        g759(.A(new_new_n781_), .B(new_new_n747_), .C(new_new_n741_), .D(new_new_n357_), .Y(mai3));
  NA2        g760(.A(i_12_), .B(i_10_), .Y(new_new_n783_));
  NA2        g761(.A(i_6_), .B(i_7_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n784_), .B(i_0_), .Y(new_new_n785_));
  NO2        g763(.A(i_11_), .B(new_new_n229_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n272_), .B(new_new_n786_), .Y(new_new_n787_));
  NO2        g765(.A(new_new_n787_), .B(new_new_n185_), .Y(new_new_n788_));
  NO3        g766(.A(new_new_n413_), .B(new_new_n91_), .C(new_new_n45_), .Y(new_new_n789_));
  OA210      g767(.A0(new_new_n789_), .A1(new_new_n788_), .B0(new_new_n169_), .Y(new_new_n790_));
  NA2        g768(.A(new_new_n772_), .B(new_new_n349_), .Y(new_new_n791_));
  NA2        g769(.A(new_new_n791_), .B(new_new_n40_), .Y(new_new_n792_));
  NOi21      g770(.An(new_new_n98_), .B(new_new_n706_), .Y(new_new_n793_));
  NA2        g771(.A(new_new_n376_), .B(new_new_n46_), .Y(new_new_n794_));
  AN2        g772(.A(new_new_n415_), .B(new_new_n56_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n795_), .B(new_new_n793_), .Y(new_new_n796_));
  AOI210     g774(.A0(new_new_n796_), .A1(new_new_n792_), .B0(new_new_n49_), .Y(new_new_n797_));
  NO4        g775(.A(new_new_n353_), .B(new_new_n359_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n177_), .B(new_new_n531_), .Y(new_new_n799_));
  NOi21      g777(.An(new_new_n799_), .B(new_new_n798_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n64_), .Y(new_new_n801_));
  NOi21      g779(.An(i_5_), .B(i_9_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n802_), .B(new_new_n409_), .Y(new_new_n803_));
  BUFFER     g781(.A(new_new_n251_), .Y(new_new_n804_));
  NA2        g782(.A(new_new_n804_), .B(new_new_n434_), .Y(new_new_n805_));
  NO3        g783(.A(new_new_n379_), .B(new_new_n251_), .C(new_new_n74_), .Y(new_new_n806_));
  NO2        g784(.A(new_new_n170_), .B(new_new_n146_), .Y(new_new_n807_));
  AOI210     g785(.A0(new_new_n807_), .A1(new_new_n236_), .B0(new_new_n806_), .Y(new_new_n808_));
  OAI220     g786(.A0(new_new_n808_), .A1(new_new_n175_), .B0(new_new_n805_), .B1(new_new_n803_), .Y(new_new_n809_));
  NO4        g787(.A(new_new_n809_), .B(new_new_n801_), .C(new_new_n797_), .D(new_new_n790_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n177_), .B(new_new_n24_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n362_), .B(new_new_n273_), .Y(new_new_n812_));
  NA2        g790(.A(new_new_n812_), .B(new_new_n658_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n532_), .B(i_0_), .Y(new_new_n814_));
  NO4        g792(.A(new_new_n544_), .B(new_new_n207_), .C(new_new_n383_), .D(new_new_n375_), .Y(new_new_n815_));
  NA2        g793(.A(new_new_n815_), .B(i_11_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n693_), .B(new_new_n304_), .Y(new_new_n817_));
  AOI210     g795(.A0(new_new_n442_), .A1(new_new_n88_), .B0(new_new_n59_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n818_), .B(new_new_n817_), .Y(new_new_n819_));
  INV        g797(.A(new_new_n498_), .Y(new_new_n820_));
  NO4        g798(.A(new_new_n115_), .B(new_new_n59_), .C(new_new_n615_), .D(i_5_), .Y(new_new_n821_));
  AN2        g799(.A(new_new_n821_), .B(new_new_n820_), .Y(new_new_n822_));
  AOI220     g800(.A0(new_new_n306_), .A1(new_new_n100_), .B0(new_new_n177_), .B1(new_new_n85_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n526_), .B(i_4_), .Y(new_new_n824_));
  NO2        g802(.A(new_new_n824_), .B(new_new_n823_), .Y(new_new_n825_));
  NO3        g803(.A(new_new_n825_), .B(new_new_n822_), .C(new_new_n819_), .Y(new_new_n826_));
  NA3        g804(.A(new_new_n826_), .B(new_new_n816_), .C(new_new_n813_), .Y(new_new_n827_));
  NO2        g805(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n828_));
  NA2        g806(.A(i_11_), .B(i_9_), .Y(new_new_n829_));
  NO3        g807(.A(i_12_), .B(new_new_n829_), .C(new_new_n557_), .Y(new_new_n830_));
  AN2        g808(.A(new_new_n830_), .B(new_new_n828_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n49_), .B(i_7_), .Y(new_new_n832_));
  NA2        g810(.A(new_new_n363_), .B(new_new_n174_), .Y(new_new_n833_));
  INV        g811(.A(new_new_n833_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n829_), .B(new_new_n74_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n170_), .B(i_0_), .Y(new_new_n836_));
  INV        g814(.A(new_new_n836_), .Y(new_new_n837_));
  NA2        g815(.A(new_new_n432_), .B(new_new_n223_), .Y(new_new_n838_));
  AOI210     g816(.A0(new_new_n348_), .A1(new_new_n42_), .B0(new_new_n372_), .Y(new_new_n839_));
  OAI220     g817(.A0(new_new_n839_), .A1(new_new_n803_), .B0(new_new_n838_), .B1(new_new_n837_), .Y(new_new_n840_));
  NO3        g818(.A(new_new_n840_), .B(new_new_n834_), .C(new_new_n831_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n606_), .B(new_new_n119_), .Y(new_new_n842_));
  NO2        g820(.A(i_6_), .B(new_new_n842_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n166_), .B(new_new_n104_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n559_), .B(new_new_n304_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n845_), .B(new_new_n794_), .Y(new_new_n846_));
  NO2        g824(.A(new_new_n846_), .B(new_new_n843_), .Y(new_new_n847_));
  NOi21      g825(.An(i_7_), .B(i_5_), .Y(new_new_n848_));
  NO3        g826(.A(new_new_n368_), .B(new_new_n337_), .C(new_new_n333_), .Y(new_new_n849_));
  NO2        g827(.A(new_new_n249_), .B(new_new_n294_), .Y(new_new_n850_));
  INV        g828(.A(new_new_n673_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n851_), .A1(new_new_n850_), .B0(new_new_n849_), .Y(new_new_n852_));
  NA3        g830(.A(new_new_n852_), .B(new_new_n847_), .C(new_new_n841_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n811_), .B(new_new_n232_), .Y(new_new_n854_));
  AN2        g832(.A(new_new_n305_), .B(new_new_n304_), .Y(new_new_n855_));
  AN2        g833(.A(new_new_n855_), .B(new_new_n807_), .Y(new_new_n856_));
  OAI210     g834(.A0(new_new_n856_), .A1(new_new_n854_), .B0(i_10_), .Y(new_new_n857_));
  NO2        g835(.A(new_new_n783_), .B(new_new_n293_), .Y(new_new_n858_));
  OA210      g836(.A0(new_new_n432_), .A1(new_new_n216_), .B0(new_new_n431_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n858_), .B(new_new_n835_), .Y(new_new_n860_));
  NA2        g838(.A(new_new_n835_), .B(new_new_n283_), .Y(new_new_n861_));
  OAI210     g839(.A0(i_2_), .A1(new_new_n179_), .B0(new_new_n861_), .Y(new_new_n862_));
  NA2        g840(.A(new_new_n862_), .B(new_new_n432_), .Y(new_new_n863_));
  NO3        g841(.A(new_new_n544_), .B(new_new_n332_), .C(new_new_n24_), .Y(new_new_n864_));
  AOI210     g842(.A0(new_new_n650_), .A1(new_new_n503_), .B0(new_new_n864_), .Y(new_new_n865_));
  NAi21      g843(.An(i_9_), .B(i_5_), .Y(new_new_n866_));
  NO2        g844(.A(new_new_n866_), .B(new_new_n368_), .Y(new_new_n867_));
  NO2        g845(.A(new_new_n553_), .B(new_new_n106_), .Y(new_new_n868_));
  AOI220     g846(.A0(new_new_n868_), .A1(i_0_), .B0(new_new_n867_), .B1(new_new_n575_), .Y(new_new_n869_));
  OAI220     g847(.A0(new_new_n869_), .A1(new_new_n87_), .B0(new_new_n865_), .B1(new_new_n167_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n870_), .B(new_new_n478_), .Y(new_new_n871_));
  NA4        g849(.A(new_new_n871_), .B(new_new_n863_), .C(new_new_n860_), .D(new_new_n857_), .Y(new_new_n872_));
  NO3        g850(.A(new_new_n872_), .B(new_new_n853_), .C(new_new_n827_), .Y(new_new_n873_));
  NO2        g851(.A(i_0_), .B(new_new_n673_), .Y(new_new_n874_));
  NO3        g852(.A(new_new_n106_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n875_));
  AO220      g853(.A0(new_new_n875_), .A1(new_new_n45_), .B0(new_new_n874_), .B1(new_new_n169_), .Y(new_new_n876_));
  AOI210     g854(.A0(new_new_n743_), .A1(new_new_n635_), .B0(new_new_n844_), .Y(new_new_n877_));
  AOI210     g855(.A0(new_new_n876_), .A1(new_new_n321_), .B0(new_new_n877_), .Y(new_new_n878_));
  NA2        g856(.A(i_8_), .B(new_new_n144_), .Y(new_new_n879_));
  INV        g857(.A(new_new_n879_), .Y(new_new_n880_));
  NA3        g858(.A(new_new_n880_), .B(new_new_n622_), .C(new_new_n74_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n757_), .B(new_new_n368_), .Y(new_new_n882_));
  NA3        g860(.A(new_new_n785_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n883_));
  NA2        g861(.A(new_new_n786_), .B(i_9_), .Y(new_new_n884_));
  AOI210     g862(.A0(new_new_n883_), .A1(new_new_n457_), .B0(new_new_n884_), .Y(new_new_n885_));
  OAI210     g863(.A0(new_new_n236_), .A1(i_9_), .B0(new_new_n222_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n886_), .A1(new_new_n814_), .B0(new_new_n152_), .Y(new_new_n887_));
  NO3        g865(.A(new_new_n887_), .B(new_new_n885_), .C(new_new_n882_), .Y(new_new_n888_));
  NA3        g866(.A(new_new_n888_), .B(new_new_n881_), .C(new_new_n878_), .Y(new_new_n889_));
  NA2        g867(.A(new_new_n855_), .B(new_new_n350_), .Y(new_new_n890_));
  AOI210     g868(.A0(new_new_n278_), .A1(new_new_n160_), .B0(new_new_n890_), .Y(new_new_n891_));
  NA3        g869(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n892_));
  NA2        g870(.A(new_new_n832_), .B(new_new_n447_), .Y(new_new_n893_));
  AOI210     g871(.A0(new_new_n892_), .A1(new_new_n160_), .B0(new_new_n893_), .Y(new_new_n894_));
  NO2        g872(.A(new_new_n894_), .B(new_new_n891_), .Y(new_new_n895_));
  NA2        g873(.A(new_new_n527_), .B(new_new_n76_), .Y(new_new_n896_));
  NO3        g874(.A(new_new_n201_), .B(new_new_n359_), .C(i_0_), .Y(new_new_n897_));
  OAI210     g875(.A0(new_new_n897_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n898_));
  INV        g876(.A(new_new_n210_), .Y(new_new_n899_));
  OAI220     g877(.A0(new_new_n491_), .A1(new_new_n137_), .B0(new_new_n594_), .B1(new_new_n569_), .Y(new_new_n900_));
  NA3        g878(.A(new_new_n900_), .B(i_7_), .C(new_new_n899_), .Y(new_new_n901_));
  NA4        g879(.A(new_new_n901_), .B(new_new_n898_), .C(new_new_n896_), .D(new_new_n895_), .Y(new_new_n902_));
  NO2        g880(.A(new_new_n235_), .B(new_new_n94_), .Y(new_new_n903_));
  AOI210     g881(.A0(new_new_n903_), .A1(new_new_n874_), .B0(new_new_n110_), .Y(new_new_n904_));
  NA2        g882(.A(new_new_n848_), .B(new_new_n447_), .Y(new_new_n905_));
  NA2        g883(.A(new_new_n324_), .B(new_new_n171_), .Y(new_new_n906_));
  OA220      g884(.A0(new_new_n906_), .A1(new_new_n905_), .B0(new_new_n904_), .B1(i_5_), .Y(new_new_n907_));
  AOI210     g885(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n170_), .Y(new_new_n908_));
  NA2        g886(.A(new_new_n908_), .B(new_new_n859_), .Y(new_new_n909_));
  NA3        g887(.A(new_new_n566_), .B(new_new_n177_), .C(new_new_n85_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n910_), .B(new_new_n502_), .Y(new_new_n911_));
  NO3        g889(.A(new_new_n794_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n452_), .B(new_new_n445_), .Y(new_new_n913_));
  NO3        g891(.A(new_new_n913_), .B(new_new_n912_), .C(new_new_n911_), .Y(new_new_n914_));
  NA3        g892(.A(new_new_n832_), .B(new_new_n272_), .C(new_new_n222_), .Y(new_new_n915_));
  INV        g893(.A(new_new_n915_), .Y(new_new_n916_));
  NO3        g894(.A(new_new_n829_), .B(new_new_n210_), .C(new_new_n182_), .Y(new_new_n917_));
  NO2        g895(.A(new_new_n917_), .B(new_new_n916_), .Y(new_new_n918_));
  NA4        g896(.A(new_new_n918_), .B(new_new_n914_), .C(new_new_n909_), .D(new_new_n907_), .Y(new_new_n919_));
  INV        g897(.A(new_new_n568_), .Y(new_new_n920_));
  NO3        g898(.A(new_new_n920_), .B(new_new_n517_), .C(i_7_), .Y(new_new_n921_));
  INV        g899(.A(new_new_n921_), .Y(new_new_n922_));
  NA3        g900(.A(new_new_n283_), .B(i_5_), .C(new_new_n185_), .Y(new_new_n923_));
  NAi31      g901(.An(new_new_n234_), .B(new_new_n923_), .C(new_new_n235_), .Y(new_new_n924_));
  NO4        g902(.A(new_new_n232_), .B(new_new_n201_), .C(i_0_), .D(i_12_), .Y(new_new_n925_));
  AOI220     g903(.A0(new_new_n925_), .A1(new_new_n924_), .B0(new_new_n737_), .B1(new_new_n171_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n848_), .B(new_new_n430_), .Y(new_new_n927_));
  OAI220     g905(.A0(i_7_), .A1(new_new_n923_), .B0(new_new_n927_), .B1(new_new_n623_), .Y(new_new_n928_));
  NA2        g906(.A(new_new_n928_), .B(new_new_n836_), .Y(new_new_n929_));
  NA3        g907(.A(new_new_n929_), .B(new_new_n926_), .C(new_new_n922_), .Y(new_new_n930_));
  NO4        g908(.A(new_new_n930_), .B(new_new_n919_), .C(new_new_n902_), .D(new_new_n889_), .Y(new_new_n931_));
  OAI210     g909(.A0(new_new_n760_), .A1(new_new_n753_), .B0(new_new_n37_), .Y(new_new_n932_));
  NA2        g910(.A(new_new_n932_), .B(new_new_n564_), .Y(new_new_n933_));
  NA2        g911(.A(new_new_n933_), .B(new_new_n198_), .Y(new_new_n934_));
  NA2        g912(.A(new_new_n178_), .B(new_new_n180_), .Y(new_new_n935_));
  AO210      g913(.A0(new_new_n645_), .A1(new_new_n33_), .B0(new_new_n935_), .Y(new_new_n936_));
  OAI210     g914(.A0(new_new_n568_), .A1(new_new_n566_), .B0(new_new_n293_), .Y(new_new_n937_));
  NAi31      g915(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n938_));
  NO2        g916(.A(new_new_n71_), .B(new_new_n938_), .Y(new_new_n939_));
  INV        g917(.A(new_new_n939_), .Y(new_new_n940_));
  NA3        g918(.A(new_new_n940_), .B(new_new_n937_), .C(new_new_n936_), .Y(new_new_n941_));
  NO2        g919(.A(new_new_n423_), .B(new_new_n251_), .Y(new_new_n942_));
  NO4        g920(.A(new_new_n225_), .B(new_new_n143_), .C(new_new_n626_), .D(new_new_n37_), .Y(new_new_n943_));
  NO3        g921(.A(new_new_n943_), .B(new_new_n942_), .C(new_new_n815_), .Y(new_new_n944_));
  INV        g922(.A(new_new_n944_), .Y(new_new_n945_));
  AOI210     g923(.A0(new_new_n941_), .A1(new_new_n49_), .B0(new_new_n945_), .Y(new_new_n946_));
  AOI210     g924(.A0(new_new_n946_), .A1(new_new_n934_), .B0(new_new_n74_), .Y(new_new_n947_));
  NO2        g925(.A(new_new_n524_), .B(new_new_n356_), .Y(new_new_n948_));
  NO2        g926(.A(new_new_n948_), .B(new_new_n701_), .Y(new_new_n949_));
  NA2        g927(.A(new_new_n908_), .B(new_new_n832_), .Y(new_new_n950_));
  NO2        g928(.A(new_new_n950_), .B(new_new_n626_), .Y(new_new_n951_));
  NA2        g929(.A(new_new_n249_), .B(new_new_n58_), .Y(new_new_n952_));
  AOI220     g930(.A0(new_new_n952_), .A1(new_new_n77_), .B0(new_new_n319_), .B1(new_new_n246_), .Y(new_new_n953_));
  NO2        g931(.A(new_new_n953_), .B(new_new_n229_), .Y(new_new_n954_));
  NA3        g932(.A(new_new_n98_), .B(new_new_n285_), .C(new_new_n31_), .Y(new_new_n955_));
  INV        g933(.A(new_new_n955_), .Y(new_new_n956_));
  NO3        g934(.A(new_new_n956_), .B(new_new_n954_), .C(new_new_n951_), .Y(new_new_n957_));
  OAI210     g935(.A0(new_new_n253_), .A1(new_new_n157_), .B0(new_new_n88_), .Y(new_new_n958_));
  NA3        g936(.A(new_new_n705_), .B(new_new_n272_), .C(new_new_n81_), .Y(new_new_n959_));
  AOI210     g937(.A0(new_new_n959_), .A1(new_new_n958_), .B0(i_11_), .Y(new_new_n960_));
  NO4        g938(.A(new_new_n866_), .B(new_new_n435_), .C(new_new_n245_), .D(new_new_n244_), .Y(new_new_n961_));
  NO2        g939(.A(new_new_n961_), .B(new_new_n521_), .Y(new_new_n962_));
  INV        g940(.A(new_new_n338_), .Y(new_new_n963_));
  AOI210     g941(.A0(new_new_n963_), .A1(new_new_n962_), .B0(new_new_n41_), .Y(new_new_n964_));
  NO2        g942(.A(new_new_n964_), .B(new_new_n960_), .Y(new_new_n965_));
  OAI210     g943(.A0(new_new_n957_), .A1(i_4_), .B0(new_new_n965_), .Y(new_new_n966_));
  NO3        g944(.A(new_new_n966_), .B(new_new_n949_), .C(new_new_n947_), .Y(new_new_n967_));
  NA4        g945(.A(new_new_n967_), .B(new_new_n931_), .C(new_new_n873_), .D(new_new_n810_), .Y(mai4));
  INV        g946(.A(new_new_n649_), .Y(new_new_n971_));
  INV        g947(.A(i_12_), .Y(new_new_n972_));
endmodule


