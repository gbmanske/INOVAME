//Benchmark atmr_intb_466_0.0156

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n349_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n411_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n390_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n393_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n466_, men_men_n467_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n53_));
  NOi21      o031(.An(x01), .B(x09), .Y(ori_ori_n54_));
  INV        o032(.A(x00), .Y(ori_ori_n55_));
  NO2        o033(.A(ori_ori_n51_), .B(ori_ori_n55_), .Y(ori_ori_n56_));
  NO2        o034(.A(ori_ori_n56_), .B(ori_ori_n54_), .Y(ori_ori_n57_));
  NA2        o035(.A(x09), .B(ori_ori_n55_), .Y(ori_ori_n58_));
  INV        o036(.A(x07), .Y(ori_ori_n59_));
  AOI220     o037(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n59_), .Y(ori_ori_n60_));
  INV        o038(.A(ori_ori_n57_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n62_), .B(ori_ori_n24_), .Y(ori_ori_n63_));
  OAI220     o041(.A0(ori_ori_n63_), .A1(ori_ori_n61_), .B0(ori_ori_n60_), .B1(ori_ori_n58_), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n59_), .B(ori_ori_n48_), .Y(ori_ori_n65_));
  OAI210     o043(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n65_), .Y(ori_ori_n66_));
  AOI220     o044(.A0(ori_ori_n66_), .A1(ori_ori_n57_), .B0(ori_ori_n64_), .B1(ori_ori_n31_), .Y(ori_ori_n67_));
  AOI210     o045(.A0(ori_ori_n67_), .A1(ori_ori_n53_), .B0(x05), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n59_), .B(ori_ori_n23_), .Y(ori_ori_n69_));
  NA2        o047(.A(x09), .B(x05), .Y(ori_ori_n70_));
  NA2        o048(.A(x10), .B(x06), .Y(ori_ori_n71_));
  NA3        o049(.A(ori_ori_n71_), .B(ori_ori_n70_), .C(ori_ori_n28_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n59_), .B(ori_ori_n41_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n72_), .A1(ori_ori_n69_), .B0(x03), .Y(ori_ori_n74_));
  NOi31      o052(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n75_));
  INV        o053(.A(x07), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n24_), .Y(ori_ori_n77_));
  NO2        o055(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n36_), .Y(ori_ori_n79_));
  OAI210     o057(.A0(ori_ori_n78_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n80_));
  AOI210     o058(.A0(ori_ori_n79_), .A1(ori_ori_n48_), .B0(ori_ori_n80_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n82_));
  NO2        o060(.A(x08), .B(x01), .Y(ori_ori_n83_));
  OAI210     o061(.A0(ori_ori_n83_), .A1(ori_ori_n82_), .B0(ori_ori_n35_), .Y(ori_ori_n84_));
  NA2        o062(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n85_));
  NO3        o063(.A(ori_ori_n84_), .B(ori_ori_n81_), .C(ori_ori_n77_), .Y(ori_ori_n86_));
  AN2        o064(.A(ori_ori_n86_), .B(ori_ori_n74_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n84_), .Y(ori_ori_n88_));
  NO2        o066(.A(x06), .B(x05), .Y(ori_ori_n89_));
  NA2        o067(.A(x11), .B(x00), .Y(ori_ori_n90_));
  NO2        o068(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n91_));
  NOi21      o069(.An(ori_ori_n90_), .B(ori_ori_n91_), .Y(ori_ori_n92_));
  AOI210     o070(.A0(ori_ori_n89_), .A1(ori_ori_n88_), .B0(ori_ori_n92_), .Y(ori_ori_n93_));
  NOi21      o071(.An(x01), .B(x10), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n29_), .B(ori_ori_n55_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n94_), .C(x06), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n96_), .B(ori_ori_n27_), .Y(ori_ori_n97_));
  OAI210     o075(.A0(ori_ori_n93_), .A1(x07), .B0(ori_ori_n97_), .Y(ori_ori_n98_));
  NO3        o076(.A(ori_ori_n98_), .B(ori_ori_n87_), .C(ori_ori_n68_), .Y(ori01));
  INV        o077(.A(x12), .Y(ori_ori_n100_));
  INV        o078(.A(x13), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n94_), .B(ori_ori_n28_), .Y(ori_ori_n102_));
  NO2        o080(.A(x10), .B(x01), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(ori_ori_n103_), .Y(ori_ori_n105_));
  NA2        o083(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n107_));
  NOi21      o085(.An(ori_ori_n107_), .B(ori_ori_n56_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n83_), .B(x13), .Y(ori_ori_n110_));
  NA2        o088(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n111_));
  NA2        o089(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n112_), .B(x05), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n35_), .B(ori_ori_n55_), .Y(ori_ori_n114_));
  AOI210     o092(.A0(x13), .A1(ori_ori_n79_), .B0(ori_ori_n108_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n115_), .B(ori_ori_n71_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n117_));
  NA2        o095(.A(x10), .B(ori_ori_n55_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(ori_ori_n117_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n121_));
  NA3        o099(.A(ori_ori_n121_), .B(ori_ori_n120_), .C(x13), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n123_));
  NOi31      o101(.An(ori_ori_n122_), .B(ori_ori_n123_), .C(ori_ori_n119_), .Y(ori_ori_n124_));
  NO3        o102(.A(ori_ori_n124_), .B(x06), .C(x03), .Y(ori_ori_n125_));
  NO2        o103(.A(ori_ori_n125_), .B(ori_ori_n116_), .Y(ori_ori_n126_));
  NA2        o104(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n127_));
  OAI210     o105(.A0(ori_ori_n83_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n131_));
  AOI210     o109(.A0(ori_ori_n131_), .A1(ori_ori_n49_), .B0(ori_ori_n130_), .Y(ori_ori_n132_));
  AN2        o110(.A(ori_ori_n132_), .B(ori_ori_n129_), .Y(ori_ori_n133_));
  NO2        o111(.A(x09), .B(x05), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n134_), .B(ori_ori_n47_), .Y(ori_ori_n135_));
  AOI210     o113(.A0(ori_ori_n135_), .A1(ori_ori_n105_), .B0(ori_ori_n49_), .Y(ori_ori_n136_));
  NA2        o114(.A(x09), .B(x00), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n107_), .B(ori_ori_n137_), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n138_), .B(ori_ori_n131_), .Y(ori_ori_n139_));
  NO3        o117(.A(ori_ori_n139_), .B(ori_ori_n136_), .C(ori_ori_n133_), .Y(ori_ori_n140_));
  NO2        o118(.A(x03), .B(x02), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n84_), .B(ori_ori_n101_), .Y(ori_ori_n142_));
  OAI210     o120(.A0(ori_ori_n142_), .A1(ori_ori_n108_), .B0(ori_ori_n141_), .Y(ori_ori_n143_));
  OA210      o121(.A0(ori_ori_n140_), .A1(x11), .B0(ori_ori_n143_), .Y(ori_ori_n144_));
  OAI210     o122(.A0(ori_ori_n126_), .A1(ori_ori_n23_), .B0(ori_ori_n144_), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n105_), .B(ori_ori_n40_), .Y(ori_ori_n146_));
  NAi21      o124(.An(x06), .B(x10), .Y(ori_ori_n147_));
  NOi21      o125(.An(x01), .B(x13), .Y(ori_ori_n148_));
  NA2        o126(.A(ori_ori_n148_), .B(ori_ori_n147_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n146_), .B(ori_ori_n41_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n101_), .B(x01), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n152_), .B(x08), .Y(ori_ori_n153_));
  NO2        o131(.A(ori_ori_n151_), .B(ori_ori_n48_), .Y(ori_ori_n154_));
  AOI210     o132(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n155_));
  OAI210     o133(.A0(ori_ori_n154_), .A1(ori_ori_n150_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o134(.A(x04), .B(x02), .Y(ori_ori_n157_));
  NA2        o135(.A(x10), .B(x05), .Y(ori_ori_n158_));
  NO2        o136(.A(x09), .B(x01), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n107_), .B(x08), .Y(ori_ori_n160_));
  INV        o138(.A(ori_ori_n25_), .Y(ori_ori_n161_));
  NAi21      o139(.An(x13), .B(x00), .Y(ori_ori_n162_));
  AOI210     o140(.A0(ori_ori_n29_), .A1(ori_ori_n48_), .B0(ori_ori_n162_), .Y(ori_ori_n163_));
  AN2        o141(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n164_));
  NO2        o142(.A(ori_ori_n95_), .B(x06), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n162_), .B(ori_ori_n36_), .Y(ori_ori_n166_));
  INV        o144(.A(ori_ori_n166_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n165_), .B(ori_ori_n164_), .Y(ori_ori_n168_));
  NA2        o146(.A(ori_ori_n168_), .B(ori_ori_n161_), .Y(ori_ori_n169_));
  NOi21      o147(.An(x09), .B(x00), .Y(ori_ori_n170_));
  NO3        o148(.A(ori_ori_n82_), .B(ori_ori_n170_), .C(ori_ori_n47_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(ori_ori_n118_), .Y(ori_ori_n172_));
  NA2        o150(.A(x06), .B(x05), .Y(ori_ori_n173_));
  OAI210     o151(.A0(ori_ori_n173_), .A1(ori_ori_n35_), .B0(ori_ori_n100_), .Y(ori_ori_n174_));
  AOI210     o152(.A0(x10), .A1(ori_ori_n56_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n172_), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n101_), .B(x12), .Y(ori_ori_n177_));
  AOI210     o155(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n177_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n179_), .B(x02), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n178_), .B(ori_ori_n176_), .Y(ori_ori_n181_));
  NA3        o159(.A(ori_ori_n181_), .B(ori_ori_n169_), .C(ori_ori_n156_), .Y(ori_ori_n182_));
  AOI210     o160(.A0(ori_ori_n145_), .A1(ori_ori_n100_), .B0(ori_ori_n182_), .Y(ori_ori_n183_));
  INV        o161(.A(ori_ori_n72_), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n184_), .B(ori_ori_n129_), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n186_), .B(ori_ori_n128_), .Y(ori_ori_n187_));
  AOI210     o165(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n117_), .B(x06), .Y(ori_ori_n189_));
  AOI210     o167(.A0(ori_ori_n188_), .A1(ori_ori_n187_), .B0(ori_ori_n189_), .Y(ori_ori_n190_));
  AOI210     o168(.A0(ori_ori_n190_), .A1(ori_ori_n185_), .B0(x12), .Y(ori_ori_n191_));
  INV        o169(.A(ori_ori_n75_), .Y(ori_ori_n192_));
  NO2        o170(.A(x05), .B(ori_ori_n51_), .Y(ori_ori_n193_));
  OAI210     o171(.A0(ori_ori_n193_), .A1(ori_ori_n149_), .B0(ori_ori_n55_), .Y(ori_ori_n194_));
  NA2        o172(.A(ori_ori_n194_), .B(ori_ori_n192_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n94_), .B(x06), .Y(ori_ori_n196_));
  AOI210     o174(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n197_));
  NO3        o175(.A(ori_ori_n197_), .B(ori_ori_n196_), .C(ori_ori_n41_), .Y(ori_ori_n198_));
  INV        o176(.A(ori_ori_n131_), .Y(ori_ori_n199_));
  OAI210     o177(.A0(ori_ori_n199_), .A1(ori_ori_n198_), .B0(x02), .Y(ori_ori_n200_));
  AOI210     o178(.A0(ori_ori_n200_), .A1(ori_ori_n195_), .B0(ori_ori_n23_), .Y(ori_ori_n201_));
  OAI210     o179(.A0(ori_ori_n191_), .A1(ori_ori_n55_), .B0(ori_ori_n201_), .Y(ori_ori_n202_));
  INV        o180(.A(ori_ori_n131_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n204_));
  OAI210     o182(.A0(ori_ori_n78_), .A1(ori_ori_n36_), .B0(ori_ori_n111_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n101_), .B(x03), .Y(ori_ori_n206_));
  AOI220     o184(.A0(ori_ori_n206_), .A1(ori_ori_n205_), .B0(ori_ori_n75_), .B1(ori_ori_n204_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n208_));
  INV        o186(.A(ori_ori_n147_), .Y(ori_ori_n209_));
  NOi21      o187(.An(x13), .B(x04), .Y(ori_ori_n210_));
  NO3        o188(.A(ori_ori_n210_), .B(ori_ori_n75_), .C(ori_ori_n170_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(x05), .Y(ori_ori_n212_));
  AOI220     o190(.A0(ori_ori_n212_), .A1(ori_ori_n208_), .B0(ori_ori_n209_), .B1(ori_ori_n55_), .Y(ori_ori_n213_));
  OAI210     o191(.A0(ori_ori_n207_), .A1(ori_ori_n203_), .B0(ori_ori_n213_), .Y(ori_ori_n214_));
  INV        o192(.A(ori_ori_n91_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n215_), .B(x12), .Y(ori_ori_n216_));
  NA2        o194(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n163_), .Y(ori_ori_n219_));
  AOI210     o197(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n220_));
  NO2        o198(.A(x06), .B(x00), .Y(ori_ori_n221_));
  NO3        o199(.A(ori_ori_n221_), .B(ori_ori_n220_), .C(ori_ori_n41_), .Y(ori_ori_n222_));
  INV        o200(.A(ori_ori_n71_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n225_));
  NA2        o203(.A(ori_ori_n225_), .B(x03), .Y(ori_ori_n226_));
  OA210      o204(.A0(ori_ori_n226_), .A1(ori_ori_n224_), .B0(ori_ori_n219_), .Y(ori_ori_n227_));
  NA2        o205(.A(x13), .B(ori_ori_n100_), .Y(ori_ori_n228_));
  NA3        o206(.A(ori_ori_n228_), .B(ori_ori_n174_), .C(ori_ori_n92_), .Y(ori_ori_n229_));
  OAI210     o207(.A0(ori_ori_n227_), .A1(ori_ori_n217_), .B0(ori_ori_n229_), .Y(ori_ori_n230_));
  AOI210     o208(.A0(ori_ori_n216_), .A1(ori_ori_n214_), .B0(ori_ori_n230_), .Y(ori_ori_n231_));
  AOI210     o209(.A0(ori_ori_n231_), .A1(ori_ori_n202_), .B0(x07), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n70_), .B(ori_ori_n29_), .Y(ori_ori_n233_));
  NOi31      o211(.An(ori_ori_n127_), .B(ori_ori_n210_), .C(ori_ori_n170_), .Y(ori_ori_n234_));
  NO2        o212(.A(ori_ori_n234_), .B(ori_ori_n233_), .Y(ori_ori_n235_));
  NO2        o213(.A(x08), .B(x05), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n220_), .Y(ori_ori_n237_));
  OAI210     o215(.A0(ori_ori_n75_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n238_));
  INV        o216(.A(ori_ori_n238_), .Y(ori_ori_n239_));
  NO2        o217(.A(x12), .B(x02), .Y(ori_ori_n240_));
  INV        o218(.A(ori_ori_n240_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n241_), .B(ori_ori_n215_), .Y(ori_ori_n242_));
  OA210      o220(.A0(ori_ori_n239_), .A1(ori_ori_n235_), .B0(ori_ori_n242_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(x01), .Y(ori_ori_n245_));
  INV        o223(.A(ori_ori_n245_), .Y(ori_ori_n246_));
  AOI210     o224(.A0(ori_ori_n246_), .A1(ori_ori_n122_), .B0(ori_ori_n29_), .Y(ori_ori_n247_));
  NA2        o225(.A(ori_ori_n101_), .B(x04), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n248_), .B(ori_ori_n28_), .Y(ori_ori_n249_));
  NO2        o227(.A(ori_ori_n249_), .B(ori_ori_n110_), .Y(ori_ori_n250_));
  NO3        o228(.A(ori_ori_n90_), .B(x12), .C(x03), .Y(ori_ori_n251_));
  OAI210     o229(.A0(ori_ori_n250_), .A1(ori_ori_n247_), .B0(ori_ori_n251_), .Y(ori_ori_n252_));
  NOi21      o230(.An(ori_ori_n233_), .B(ori_ori_n196_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n254_));
  NA2        o232(.A(ori_ori_n253_), .B(ori_ori_n254_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n256_));
  NO3        o234(.A(ori_ori_n256_), .B(ori_ori_n197_), .C(ori_ori_n165_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n217_), .B(ori_ori_n28_), .Y(ori_ori_n258_));
  OAI210     o236(.A0(ori_ori_n257_), .A1(ori_ori_n203_), .B0(ori_ori_n258_), .Y(ori_ori_n259_));
  NA3        o237(.A(ori_ori_n259_), .B(ori_ori_n255_), .C(ori_ori_n252_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n260_), .B(ori_ori_n243_), .C(ori_ori_n232_), .Y(ori_ori_n261_));
  OAI210     o239(.A0(ori_ori_n183_), .A1(ori_ori_n59_), .B0(ori_ori_n261_), .Y(ori02));
  AOI210     o240(.A0(ori_ori_n127_), .A1(ori_ori_n84_), .B0(ori_ori_n120_), .Y(ori_ori_n263_));
  NOi21      o241(.An(ori_ori_n211_), .B(ori_ori_n159_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n101_), .B(ori_ori_n35_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n264_), .B(ori_ori_n32_), .Y(ori_ori_n266_));
  OAI210     o244(.A0(ori_ori_n266_), .A1(ori_ori_n263_), .B0(ori_ori_n158_), .Y(ori_ori_n267_));
  INV        o245(.A(ori_ori_n158_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n109_), .A1(ori_ori_n85_), .B0(ori_ori_n197_), .Y(ori_ori_n269_));
  OAI220     o247(.A0(ori_ori_n269_), .A1(ori_ori_n101_), .B0(ori_ori_n84_), .B1(ori_ori_n51_), .Y(ori_ori_n270_));
  AOI220     o248(.A0(ori_ori_n270_), .A1(ori_ori_n268_), .B0(ori_ori_n142_), .B1(ori_ori_n141_), .Y(ori_ori_n271_));
  AOI210     o249(.A0(ori_ori_n271_), .A1(ori_ori_n267_), .B0(ori_ori_n48_), .Y(ori_ori_n272_));
  NO2        o250(.A(x05), .B(x02), .Y(ori_ori_n273_));
  OAI210     o251(.A0(ori_ori_n187_), .A1(ori_ori_n170_), .B0(ori_ori_n273_), .Y(ori_ori_n274_));
  AOI220     o252(.A0(ori_ori_n236_), .A1(ori_ori_n56_), .B0(ori_ori_n54_), .B1(ori_ori_n36_), .Y(ori_ori_n275_));
  NOi21      o253(.An(ori_ori_n265_), .B(ori_ori_n275_), .Y(ori_ori_n276_));
  AOI210     o254(.A0(ori_ori_n210_), .A1(ori_ori_n78_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  AOI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n274_), .B0(ori_ori_n131_), .Y(ori_ori_n278_));
  NAi21      o256(.An(ori_ori_n212_), .B(ori_ori_n207_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n225_), .B(ori_ori_n47_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n279_), .Y(ori_ori_n281_));
  AN2        o259(.A(ori_ori_n206_), .B(ori_ori_n205_), .Y(ori_ori_n282_));
  OAI210     o260(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n283_));
  NA2        o261(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n284_));
  OA210      o262(.A0(ori_ori_n284_), .A1(x08), .B0(ori_ori_n135_), .Y(ori_ori_n285_));
  AOI210     o263(.A0(ori_ori_n285_), .A1(ori_ori_n128_), .B0(ori_ori_n283_), .Y(ori_ori_n286_));
  OAI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n282_), .B0(ori_ori_n95_), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n141_), .Y(ori_ori_n288_));
  OAI220     o266(.A0(ori_ori_n237_), .A1(ori_ori_n102_), .B0(ori_ori_n288_), .B1(ori_ori_n119_), .Y(ori_ori_n289_));
  NA2        o267(.A(ori_ori_n289_), .B(x13), .Y(ori_ori_n290_));
  NA3        o268(.A(ori_ori_n290_), .B(ori_ori_n287_), .C(ori_ori_n281_), .Y(ori_ori_n291_));
  NO3        o269(.A(ori_ori_n291_), .B(ori_ori_n278_), .C(ori_ori_n272_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n130_), .B(x03), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n162_), .Y(ori_ori_n294_));
  OAI210     o272(.A0(ori_ori_n51_), .A1(ori_ori_n35_), .B0(ori_ori_n36_), .Y(ori_ori_n295_));
  AOI220     o273(.A0(ori_ori_n295_), .A1(ori_ori_n294_), .B0(ori_ori_n179_), .B1(x08), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n296_), .A1(ori_ori_n256_), .B0(ori_ori_n293_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n297_), .B(ori_ori_n103_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n157_), .B(ori_ori_n152_), .Y(ori_ori_n299_));
  AN2        o277(.A(ori_ori_n299_), .B(ori_ori_n160_), .Y(ori_ori_n300_));
  INV        o278(.A(ori_ori_n54_), .Y(ori_ori_n301_));
  OAI220     o279(.A0(ori_ori_n248_), .A1(ori_ori_n301_), .B0(ori_ori_n120_), .B1(ori_ori_n28_), .Y(ori_ori_n302_));
  OAI210     o280(.A0(ori_ori_n302_), .A1(ori_ori_n300_), .B0(ori_ori_n104_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n248_), .B(ori_ori_n100_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n100_), .B(ori_ori_n41_), .Y(ori_ori_n305_));
  NA3        o283(.A(ori_ori_n305_), .B(ori_ori_n304_), .C(ori_ori_n119_), .Y(ori_ori_n306_));
  NA4        o284(.A(ori_ori_n306_), .B(ori_ori_n303_), .C(ori_ori_n298_), .D(ori_ori_n48_), .Y(ori_ori_n307_));
  INV        o285(.A(ori_ori_n179_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n309_));
  OAI220     o287(.A0(ori_ori_n309_), .A1(ori_ori_n411_), .B0(ori_ori_n308_), .B1(ori_ori_n57_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n310_), .B(x02), .Y(ori_ori_n311_));
  INV        o289(.A(ori_ori_n218_), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n177_), .B(x04), .Y(ori_ori_n313_));
  NO3        o291(.A(ori_ori_n177_), .B(ori_ori_n151_), .C(ori_ori_n52_), .Y(ori_ori_n314_));
  OAI210     o292(.A0(ori_ori_n137_), .A1(ori_ori_n36_), .B0(ori_ori_n100_), .Y(ori_ori_n315_));
  OAI210     o293(.A0(ori_ori_n315_), .A1(ori_ori_n171_), .B0(ori_ori_n314_), .Y(ori_ori_n316_));
  NA3        o294(.A(ori_ori_n316_), .B(ori_ori_n311_), .C(x06), .Y(ori_ori_n317_));
  NA2        o295(.A(x09), .B(x03), .Y(ori_ori_n318_));
  OAI220     o296(.A0(ori_ori_n318_), .A1(ori_ori_n118_), .B0(ori_ori_n186_), .B1(ori_ori_n62_), .Y(ori_ori_n319_));
  NO3        o297(.A(ori_ori_n256_), .B(ori_ori_n117_), .C(x08), .Y(ori_ori_n320_));
  INV        o298(.A(ori_ori_n320_), .Y(ori_ori_n321_));
  NO2        o299(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n322_));
  NO3        o300(.A(ori_ori_n107_), .B(ori_ori_n118_), .C(ori_ori_n38_), .Y(ori_ori_n323_));
  AOI210     o301(.A0(ori_ori_n314_), .A1(ori_ori_n322_), .B0(ori_ori_n323_), .Y(ori_ori_n324_));
  OAI210     o302(.A0(ori_ori_n321_), .A1(ori_ori_n28_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  AO220      o303(.A0(ori_ori_n325_), .A1(x04), .B0(ori_ori_n319_), .B1(x05), .Y(ori_ori_n326_));
  AOI210     o304(.A0(ori_ori_n317_), .A1(ori_ori_n307_), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  OAI210     o305(.A0(ori_ori_n292_), .A1(x12), .B0(ori_ori_n327_), .Y(ori03));
  OR2        o306(.A(ori_ori_n42_), .B(ori_ori_n204_), .Y(ori_ori_n329_));
  AOI210     o307(.A0(ori_ori_n142_), .A1(ori_ori_n100_), .B0(ori_ori_n329_), .Y(ori_ori_n330_));
  AO210      o308(.A0(ori_ori_n312_), .A1(ori_ori_n85_), .B0(ori_ori_n313_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n177_), .B(ori_ori_n141_), .Y(ori_ori_n332_));
  NA3        o310(.A(ori_ori_n332_), .B(ori_ori_n331_), .C(ori_ori_n180_), .Y(ori_ori_n333_));
  OAI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n330_), .B0(x05), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n329_), .B(x05), .Y(ori_ori_n335_));
  AOI210     o313(.A0(ori_ori_n128_), .A1(ori_ori_n192_), .B0(ori_ori_n335_), .Y(ori_ori_n336_));
  AOI210     o314(.A0(ori_ori_n206_), .A1(ori_ori_n79_), .B0(ori_ori_n113_), .Y(ori_ori_n337_));
  OAI220     o315(.A0(ori_ori_n337_), .A1(ori_ori_n57_), .B0(ori_ori_n284_), .B1(ori_ori_n275_), .Y(ori_ori_n338_));
  OAI210     o316(.A0(ori_ori_n338_), .A1(ori_ori_n336_), .B0(ori_ori_n100_), .Y(ori_ori_n339_));
  AOI210     o317(.A0(ori_ori_n135_), .A1(ori_ori_n58_), .B0(ori_ori_n38_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n159_), .B(ori_ori_n123_), .Y(ori_ori_n341_));
  OAI220     o319(.A0(ori_ori_n341_), .A1(ori_ori_n37_), .B0(ori_ori_n138_), .B1(x13), .Y(ori_ori_n342_));
  OAI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n340_), .B0(x04), .Y(ori_ori_n343_));
  NO3        o321(.A(ori_ori_n305_), .B(ori_ori_n84_), .C(ori_ori_n57_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n167_), .A1(ori_ori_n100_), .B0(ori_ori_n135_), .Y(ori_ori_n345_));
  OA210      o323(.A0(ori_ori_n153_), .A1(x12), .B0(ori_ori_n123_), .Y(ori_ori_n346_));
  NO3        o324(.A(ori_ori_n346_), .B(ori_ori_n345_), .C(ori_ori_n344_), .Y(ori_ori_n347_));
  NA4        o325(.A(ori_ori_n347_), .B(ori_ori_n343_), .C(ori_ori_n339_), .D(ori_ori_n334_), .Y(ori04));
  NO2        o326(.A(ori_ori_n88_), .B(ori_ori_n39_), .Y(ori_ori_n349_));
  XO2        o327(.A(ori_ori_n349_), .B(ori_ori_n228_), .Y(ori05));
  AOI210     o328(.A0(ori_ori_n70_), .A1(ori_ori_n52_), .B0(ori_ori_n189_), .Y(ori_ori_n351_));
  AOI210     o329(.A0(ori_ori_n351_), .A1(ori_ori_n283_), .B0(ori_ori_n25_), .Y(ori_ori_n352_));
  NA3        o330(.A(ori_ori_n131_), .B(ori_ori_n120_), .C(ori_ori_n31_), .Y(ori_ori_n353_));
  AOI210     o331(.A0(ori_ori_n209_), .A1(ori_ori_n55_), .B0(ori_ori_n89_), .Y(ori_ori_n354_));
  AOI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n353_), .B0(ori_ori_n24_), .Y(ori_ori_n355_));
  OAI210     o333(.A0(ori_ori_n355_), .A1(ori_ori_n352_), .B0(ori_ori_n100_), .Y(ori_ori_n356_));
  NA2        o334(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n233_), .B(x03), .Y(ori_ori_n359_));
  OAI220     o337(.A0(ori_ori_n359_), .A1(ori_ori_n358_), .B0(ori_ori_n357_), .B1(ori_ori_n80_), .Y(ori_ori_n360_));
  OAI210     o338(.A0(ori_ori_n26_), .A1(ori_ori_n100_), .B0(x07), .Y(ori_ori_n361_));
  AOI210     o339(.A0(ori_ori_n360_), .A1(x06), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  AOI220     o340(.A0(ori_ori_n80_), .A1(ori_ori_n31_), .B0(ori_ori_n52_), .B1(ori_ori_n51_), .Y(ori_ori_n363_));
  NO3        o341(.A(ori_ori_n363_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n364_));
  OR2        o342(.A(x02), .B(ori_ori_n217_), .Y(ori_ori_n365_));
  NA2        o343(.A(ori_ori_n221_), .B(ori_ori_n215_), .Y(ori_ori_n366_));
  NA2        o344(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n367_));
  OAI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n364_), .B0(ori_ori_n100_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n33_), .B(ori_ori_n100_), .Y(ori_ori_n369_));
  AOI210     o347(.A0(ori_ori_n369_), .A1(ori_ori_n91_), .B0(x07), .Y(ori_ori_n370_));
  AOI220     o348(.A0(ori_ori_n370_), .A1(ori_ori_n368_), .B0(ori_ori_n362_), .B1(ori_ori_n356_), .Y(ori_ori_n371_));
  OR2        o349(.A(ori_ori_n244_), .B(ori_ori_n241_), .Y(ori_ori_n372_));
  NO2        o350(.A(ori_ori_n134_), .B(ori_ori_n28_), .Y(ori_ori_n373_));
  AOI210     o351(.A0(ori_ori_n372_), .A1(ori_ori_n47_), .B0(ori_ori_n373_), .Y(ori_ori_n374_));
  NA2        o352(.A(ori_ori_n374_), .B(ori_ori_n101_), .Y(ori_ori_n375_));
  AOI210     o353(.A0(ori_ori_n313_), .A1(ori_ori_n106_), .B0(ori_ori_n240_), .Y(ori_ori_n376_));
  NOi21      o354(.An(ori_ori_n293_), .B(ori_ori_n123_), .Y(ori_ori_n377_));
  NO2        o355(.A(ori_ori_n377_), .B(ori_ori_n241_), .Y(ori_ori_n378_));
  OAI210     o356(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n379_));
  AOI210     o357(.A0(ori_ori_n228_), .A1(ori_ori_n47_), .B0(ori_ori_n379_), .Y(ori_ori_n380_));
  NO4        o358(.A(ori_ori_n380_), .B(ori_ori_n378_), .C(ori_ori_n376_), .D(x08), .Y(ori_ori_n381_));
  NA2        o359(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n382_));
  NO2        o360(.A(ori_ori_n382_), .B(x03), .Y(ori_ori_n383_));
  NO2        o361(.A(x13), .B(x12), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n120_), .B(ori_ori_n28_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n385_), .B(ori_ori_n245_), .Y(ori_ori_n386_));
  OR3        o364(.A(ori_ori_n386_), .B(x12), .C(x03), .Y(ori_ori_n387_));
  NA3        o365(.A(ori_ori_n308_), .B(ori_ori_n114_), .C(x12), .Y(ori_ori_n388_));
  AO210      o366(.A0(ori_ori_n308_), .A1(ori_ori_n114_), .B0(ori_ori_n228_), .Y(ori_ori_n389_));
  NA4        o367(.A(ori_ori_n389_), .B(ori_ori_n388_), .C(ori_ori_n387_), .D(x08), .Y(ori_ori_n390_));
  AOI210     o368(.A0(ori_ori_n384_), .A1(ori_ori_n383_), .B0(ori_ori_n390_), .Y(ori_ori_n391_));
  AOI210     o369(.A0(ori_ori_n381_), .A1(ori_ori_n375_), .B0(ori_ori_n391_), .Y(ori_ori_n392_));
  INV        o370(.A(x03), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n134_), .B(ori_ori_n43_), .Y(ori_ori_n394_));
  OAI210     o372(.A0(ori_ori_n394_), .A1(ori_ori_n393_), .B0(ori_ori_n166_), .Y(ori_ori_n395_));
  NA3        o373(.A(ori_ori_n386_), .B(ori_ori_n377_), .C(ori_ori_n304_), .Y(ori_ori_n396_));
  INV        o374(.A(x14), .Y(ori_ori_n397_));
  NO3        o375(.A(ori_ori_n152_), .B(ori_ori_n73_), .C(ori_ori_n55_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n397_), .Y(ori_ori_n399_));
  NA3        o377(.A(ori_ori_n399_), .B(ori_ori_n396_), .C(ori_ori_n395_), .Y(ori_ori_n400_));
  AOI220     o378(.A0(ori_ori_n369_), .A1(ori_ori_n59_), .B0(ori_ori_n385_), .B1(ori_ori_n151_), .Y(ori_ori_n401_));
  NOi21      o379(.An(ori_ori_n248_), .B(ori_ori_n138_), .Y(ori_ori_n402_));
  NO3        o380(.A(ori_ori_n117_), .B(ori_ori_n24_), .C(x06), .Y(ori_ori_n403_));
  AOI210     o381(.A0(ori_ori_n254_), .A1(ori_ori_n209_), .B0(ori_ori_n403_), .Y(ori_ori_n404_));
  OAI210     o382(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n404_), .Y(ori_ori_n405_));
  OAI210     o383(.A0(ori_ori_n405_), .A1(ori_ori_n402_), .B0(ori_ori_n100_), .Y(ori_ori_n406_));
  OAI210     o384(.A0(ori_ori_n401_), .A1(ori_ori_n90_), .B0(ori_ori_n406_), .Y(ori_ori_n407_));
  NO4        o385(.A(ori_ori_n407_), .B(ori_ori_n400_), .C(ori_ori_n392_), .D(ori_ori_n371_), .Y(ori06));
  INV        o386(.A(ori_ori_n40_), .Y(ori_ori_n411_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NA2        m029(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(x07), .Y(mai_mai_n53_));
  NA2        m031(.A(mai_mai_n53_), .B(mai_mai_n47_), .Y(mai_mai_n54_));
  NOi21      m032(.An(x01), .B(x09), .Y(mai_mai_n55_));
  INV        m033(.A(x00), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n56_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(x09), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m037(.A(x07), .Y(mai_mai_n60_));
  AOI220     m038(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n60_), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n58_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n63_), .B(mai_mai_n24_), .Y(mai_mai_n64_));
  OAI220     m042(.A0(mai_mai_n64_), .A1(mai_mai_n62_), .B0(mai_mai_n61_), .B1(mai_mai_n59_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n60_), .B(mai_mai_n48_), .Y(mai_mai_n66_));
  OAI210     m044(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  AOI220     m045(.A0(mai_mai_n67_), .A1(mai_mai_n58_), .B0(mai_mai_n65_), .B1(mai_mai_n31_), .Y(mai_mai_n68_));
  AOI210     m046(.A0(mai_mai_n68_), .A1(mai_mai_n54_), .B0(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x10), .B(x09), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA3        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n28_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(x11), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n456_), .B(mai_mai_n24_), .Y(mai_mai_n76_));
  NO2        m054(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n36_), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n77_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n79_));
  AOI210     m057(.A0(mai_mai_n78_), .A1(mai_mai_n48_), .B0(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m058(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n81_));
  NO2        m059(.A(x08), .B(x01), .Y(mai_mai_n82_));
  OAI210     m060(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n35_), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n84_));
  NO3        m062(.A(mai_mai_n83_), .B(mai_mai_n80_), .C(mai_mai_n76_), .Y(mai_mai_n85_));
  AN2        m063(.A(mai_mai_n85_), .B(mai_mai_n74_), .Y(mai_mai_n86_));
  INV        m064(.A(mai_mai_n83_), .Y(mai_mai_n87_));
  NO2        m065(.A(x06), .B(x05), .Y(mai_mai_n88_));
  NA2        m066(.A(x11), .B(x00), .Y(mai_mai_n89_));
  NO2        m067(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  AOI210     m069(.A0(mai_mai_n88_), .A1(mai_mai_n87_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NOi21      m070(.An(x01), .B(x10), .Y(mai_mai_n93_));
  NO2        m071(.A(mai_mai_n29_), .B(mai_mai_n56_), .Y(mai_mai_n94_));
  NO3        m072(.A(mai_mai_n94_), .B(mai_mai_n93_), .C(x06), .Y(mai_mai_n95_));
  NA2        m073(.A(mai_mai_n95_), .B(mai_mai_n27_), .Y(mai_mai_n96_));
  OAI210     m074(.A0(mai_mai_n92_), .A1(x07), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  NO3        m075(.A(mai_mai_n97_), .B(mai_mai_n86_), .C(mai_mai_n69_), .Y(mai01));
  INV        m076(.A(x12), .Y(mai_mai_n99_));
  INV        m077(.A(x13), .Y(mai_mai_n100_));
  NA2        m078(.A(x08), .B(x04), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n101_), .B(mai_mai_n56_), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n102_), .B(mai_mai_n88_), .Y(mai_mai_n103_));
  NA2        m081(.A(mai_mai_n93_), .B(mai_mai_n28_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n104_), .B(mai_mai_n71_), .Y(mai_mai_n105_));
  NO2        m083(.A(x10), .B(x01), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(mai_mai_n106_), .Y(mai_mai_n108_));
  NA2        m086(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n109_));
  NO3        m087(.A(mai_mai_n109_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n110_));
  AOI210     m088(.A0(mai_mai_n110_), .A1(mai_mai_n108_), .B0(mai_mai_n105_), .Y(mai_mai_n111_));
  AOI210     m089(.A0(mai_mai_n111_), .A1(mai_mai_n103_), .B0(mai_mai_n100_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n55_), .B(x05), .Y(mai_mai_n113_));
  NOi21      m091(.An(mai_mai_n113_), .B(mai_mai_n57_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n100_), .B(mai_mai_n36_), .Y(mai_mai_n116_));
  NA3        m094(.A(mai_mai_n116_), .B(mai_mai_n115_), .C(x06), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n117_), .B(mai_mai_n114_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n82_), .B(x13), .Y(mai_mai_n119_));
  NA2        m097(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(mai_mai_n119_), .Y(mai_mai_n121_));
  NA2        m099(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n122_), .B(x05), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n123_), .B(mai_mai_n121_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n35_), .B(mai_mai_n56_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(mai_mai_n100_), .Y(mai_mai_n126_));
  AOI210     m104(.A0(mai_mai_n126_), .A1(mai_mai_n78_), .B0(mai_mai_n114_), .Y(mai_mai_n127_));
  AOI210     m105(.A0(mai_mai_n127_), .A1(mai_mai_n124_), .B0(mai_mai_n72_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n129_));
  NA2        m107(.A(x10), .B(mai_mai_n56_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n129_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n132_));
  NO3        m110(.A(mai_mai_n125_), .B(mai_mai_n77_), .C(mai_mai_n36_), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n59_), .B(x05), .Y(mai_mai_n134_));
  NO3        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n131_), .Y(mai_mai_n135_));
  NO3        m113(.A(mai_mai_n135_), .B(x06), .C(x03), .Y(mai_mai_n136_));
  NO4        m114(.A(mai_mai_n136_), .B(mai_mai_n128_), .C(mai_mai_n118_), .D(mai_mai_n112_), .Y(mai_mai_n137_));
  NA2        m115(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n138_));
  OAI210     m116(.A0(mai_mai_n82_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n139_));
  NA2        m117(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NO2        m118(.A(mai_mai_n35_), .B(mai_mai_n47_), .Y(mai_mai_n141_));
  NO2        m119(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n143_));
  AOI210     m121(.A0(mai_mai_n143_), .A1(mai_mai_n49_), .B0(mai_mai_n142_), .Y(mai_mai_n144_));
  OA210      m122(.A0(mai_mai_n144_), .A1(mai_mai_n141_), .B0(mai_mai_n140_), .Y(mai_mai_n145_));
  NO2        m123(.A(x09), .B(x05), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n146_), .B(mai_mai_n47_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n108_), .B(mai_mai_n49_), .Y(mai_mai_n148_));
  NA2        m126(.A(x09), .B(x00), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n113_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n75_), .B(mai_mai_n50_), .Y(mai_mai_n151_));
  AOI210     m129(.A0(mai_mai_n151_), .A1(mai_mai_n150_), .B0(mai_mai_n143_), .Y(mai_mai_n152_));
  NO3        m130(.A(mai_mai_n152_), .B(mai_mai_n148_), .C(mai_mai_n145_), .Y(mai_mai_n153_));
  NO2        m131(.A(x03), .B(x02), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n83_), .B(mai_mai_n100_), .Y(mai_mai_n155_));
  OAI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n114_), .B0(mai_mai_n154_), .Y(mai_mai_n156_));
  OA210      m134(.A0(mai_mai_n153_), .A1(x11), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  OAI210     m135(.A0(mai_mai_n137_), .A1(mai_mai_n23_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n108_), .B(mai_mai_n40_), .Y(mai_mai_n159_));
  NAi21      m137(.An(x06), .B(x10), .Y(mai_mai_n160_));
  NOi21      m138(.An(x01), .B(x13), .Y(mai_mai_n161_));
  NA2        m139(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  BUFFER     m140(.A(mai_mai_n162_), .Y(mai_mai_n163_));
  AOI210     m141(.A0(mai_mai_n163_), .A1(mai_mai_n159_), .B0(mai_mai_n41_), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n100_), .B(x01), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n166_), .B(x08), .Y(mai_mai_n167_));
  OAI210     m145(.A0(x05), .A1(mai_mai_n167_), .B0(mai_mai_n50_), .Y(mai_mai_n168_));
  AOI210     m146(.A0(mai_mai_n168_), .A1(mai_mai_n165_), .B0(mai_mai_n48_), .Y(mai_mai_n169_));
  AOI210     m147(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n170_));
  OAI210     m148(.A0(mai_mai_n169_), .A1(mai_mai_n164_), .B0(mai_mai_n170_), .Y(mai_mai_n171_));
  NA2        m149(.A(x04), .B(x02), .Y(mai_mai_n172_));
  NA2        m150(.A(x10), .B(x05), .Y(mai_mai_n173_));
  NA2        m151(.A(x09), .B(x06), .Y(mai_mai_n174_));
  AOI210     m152(.A0(mai_mai_n174_), .A1(mai_mai_n173_), .B0(x11), .Y(mai_mai_n175_));
  NO2        m153(.A(x09), .B(x01), .Y(mai_mai_n176_));
  NO3        m154(.A(mai_mai_n176_), .B(mai_mai_n106_), .C(mai_mai_n31_), .Y(mai_mai_n177_));
  OAI210     m155(.A0(mai_mai_n177_), .A1(mai_mai_n175_), .B0(x00), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n113_), .B(x08), .Y(mai_mai_n179_));
  NA3        m157(.A(mai_mai_n161_), .B(mai_mai_n160_), .C(mai_mai_n50_), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n93_), .B(x05), .Y(mai_mai_n181_));
  NA2        m159(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  AOI210     m160(.A0(mai_mai_n179_), .A1(x06), .B0(mai_mai_n182_), .Y(mai_mai_n183_));
  OAI210     m161(.A0(mai_mai_n183_), .A1(x11), .B0(mai_mai_n178_), .Y(mai_mai_n184_));
  NAi21      m162(.An(mai_mai_n172_), .B(mai_mai_n184_), .Y(mai_mai_n185_));
  INV        m163(.A(mai_mai_n25_), .Y(mai_mai_n186_));
  NAi21      m164(.An(x13), .B(x00), .Y(mai_mai_n187_));
  AOI210     m165(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  AOI220     m166(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n189_));
  OAI210     m167(.A0(mai_mai_n173_), .A1(mai_mai_n35_), .B0(mai_mai_n189_), .Y(mai_mai_n190_));
  AN2        m168(.A(mai_mai_n190_), .B(mai_mai_n188_), .Y(mai_mai_n191_));
  BUFFER     m169(.A(mai_mai_n71_), .Y(mai_mai_n192_));
  NO2        m170(.A(mai_mai_n94_), .B(x06), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n187_), .B(mai_mai_n36_), .Y(mai_mai_n194_));
  INV        m172(.A(mai_mai_n194_), .Y(mai_mai_n195_));
  OAI220     m173(.A0(mai_mai_n195_), .A1(mai_mai_n174_), .B0(mai_mai_n193_), .B1(mai_mai_n192_), .Y(mai_mai_n196_));
  OAI210     m174(.A0(mai_mai_n196_), .A1(mai_mai_n191_), .B0(mai_mai_n186_), .Y(mai_mai_n197_));
  NOi21      m175(.An(x09), .B(x00), .Y(mai_mai_n198_));
  NO3        m176(.A(mai_mai_n81_), .B(mai_mai_n198_), .C(mai_mai_n47_), .Y(mai_mai_n199_));
  NA2        m177(.A(mai_mai_n199_), .B(mai_mai_n130_), .Y(mai_mai_n200_));
  NA2        m178(.A(x10), .B(x08), .Y(mai_mai_n201_));
  INV        m179(.A(mai_mai_n201_), .Y(mai_mai_n202_));
  NA2        m180(.A(x06), .B(x05), .Y(mai_mai_n203_));
  OAI210     m181(.A0(mai_mai_n203_), .A1(mai_mai_n35_), .B0(mai_mai_n99_), .Y(mai_mai_n204_));
  NA2        m182(.A(mai_mai_n99_), .B(mai_mai_n200_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n100_), .B(x12), .Y(mai_mai_n206_));
  AOI210     m184(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n206_), .Y(mai_mai_n207_));
  NA2        m185(.A(mai_mai_n93_), .B(mai_mai_n50_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n209_));
  NA2        m187(.A(mai_mai_n209_), .B(x02), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n210_), .B(mai_mai_n208_), .Y(mai_mai_n211_));
  AOI210     m189(.A0(mai_mai_n207_), .A1(mai_mai_n205_), .B0(mai_mai_n211_), .Y(mai_mai_n212_));
  NA4        m190(.A(mai_mai_n212_), .B(mai_mai_n197_), .C(mai_mai_n185_), .D(mai_mai_n171_), .Y(mai_mai_n213_));
  AOI210     m191(.A0(mai_mai_n158_), .A1(mai_mai_n99_), .B0(mai_mai_n213_), .Y(mai_mai_n214_));
  INV        m192(.A(mai_mai_n73_), .Y(mai_mai_n215_));
  NA2        m193(.A(mai_mai_n215_), .B(mai_mai_n140_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n217_), .B(mai_mai_n139_), .Y(mai_mai_n218_));
  AOI210     m196(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n129_), .B(x06), .Y(mai_mai_n220_));
  AOI210     m198(.A0(mai_mai_n219_), .A1(mai_mai_n218_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  AOI210     m199(.A0(mai_mai_n221_), .A1(mai_mai_n216_), .B0(x12), .Y(mai_mai_n222_));
  INV        m200(.A(mai_mai_n75_), .Y(mai_mai_n223_));
  OAI210     m201(.A0(x09), .A1(mai_mai_n162_), .B0(mai_mai_n56_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n226_));
  AOI210     m204(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n227_));
  NO3        m205(.A(mai_mai_n227_), .B(mai_mai_n226_), .C(mai_mai_n41_), .Y(mai_mai_n228_));
  NA4        m206(.A(mai_mai_n160_), .B(mai_mai_n55_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n229_));
  NA2        m207(.A(mai_mai_n229_), .B(mai_mai_n143_), .Y(mai_mai_n230_));
  OAI210     m208(.A0(mai_mai_n230_), .A1(mai_mai_n228_), .B0(x02), .Y(mai_mai_n231_));
  AOI210     m209(.A0(mai_mai_n231_), .A1(mai_mai_n225_), .B0(mai_mai_n23_), .Y(mai_mai_n232_));
  OAI210     m210(.A0(mai_mai_n222_), .A1(mai_mai_n56_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  INV        m211(.A(mai_mai_n143_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n235_));
  OAI210     m213(.A0(mai_mai_n77_), .A1(mai_mai_n36_), .B0(mai_mai_n120_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n100_), .B(x03), .Y(mai_mai_n237_));
  AOI220     m215(.A0(mai_mai_n237_), .A1(mai_mai_n236_), .B0(mai_mai_n75_), .B1(mai_mai_n235_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n239_));
  INV        m217(.A(mai_mai_n160_), .Y(mai_mai_n240_));
  NOi21      m218(.An(x13), .B(x04), .Y(mai_mai_n241_));
  NO3        m219(.A(mai_mai_n241_), .B(mai_mai_n75_), .C(mai_mai_n198_), .Y(mai_mai_n242_));
  NO2        m220(.A(mai_mai_n242_), .B(x05), .Y(mai_mai_n243_));
  AOI220     m221(.A0(mai_mai_n243_), .A1(mai_mai_n239_), .B0(mai_mai_n240_), .B1(mai_mai_n56_), .Y(mai_mai_n244_));
  OAI210     m222(.A0(mai_mai_n238_), .A1(mai_mai_n234_), .B0(mai_mai_n244_), .Y(mai_mai_n245_));
  INV        m223(.A(mai_mai_n90_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n246_), .B(x12), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n249_));
  OAI210     m227(.A0(mai_mai_n249_), .A1(mai_mai_n190_), .B0(mai_mai_n188_), .Y(mai_mai_n250_));
  AOI210     m228(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n251_));
  NO2        m229(.A(x06), .B(x00), .Y(mai_mai_n252_));
  NO3        m230(.A(mai_mai_n252_), .B(mai_mai_n251_), .C(mai_mai_n41_), .Y(mai_mai_n253_));
  OAI210     m231(.A0(mai_mai_n101_), .A1(mai_mai_n149_), .B0(mai_mai_n72_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n254_), .B(mai_mai_n253_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n256_), .B(x03), .Y(mai_mai_n257_));
  OA210      m235(.A0(mai_mai_n257_), .A1(mai_mai_n255_), .B0(mai_mai_n250_), .Y(mai_mai_n258_));
  NA2        m236(.A(x13), .B(mai_mai_n99_), .Y(mai_mai_n259_));
  NA3        m237(.A(mai_mai_n259_), .B(mai_mai_n204_), .C(mai_mai_n91_), .Y(mai_mai_n260_));
  OAI210     m238(.A0(mai_mai_n258_), .A1(mai_mai_n248_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  AOI210     m239(.A0(mai_mai_n247_), .A1(mai_mai_n245_), .B0(mai_mai_n261_), .Y(mai_mai_n262_));
  AOI210     m240(.A0(mai_mai_n262_), .A1(mai_mai_n233_), .B0(x07), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n264_));
  NOi31      m242(.An(mai_mai_n138_), .B(mai_mai_n241_), .C(mai_mai_n198_), .Y(mai_mai_n265_));
  AOI210     m243(.A0(mai_mai_n265_), .A1(mai_mai_n151_), .B0(mai_mai_n264_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n100_), .B(x06), .Y(mai_mai_n267_));
  INV        m245(.A(mai_mai_n267_), .Y(mai_mai_n268_));
  NO2        m246(.A(x08), .B(x05), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n269_), .B(mai_mai_n251_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n271_));
  OAI210     m249(.A0(mai_mai_n270_), .A1(mai_mai_n268_), .B0(mai_mai_n271_), .Y(mai_mai_n272_));
  NO2        m250(.A(x12), .B(x02), .Y(mai_mai_n273_));
  INV        m251(.A(mai_mai_n273_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n274_), .B(mai_mai_n246_), .Y(mai_mai_n275_));
  OA210      m253(.A0(mai_mai_n272_), .A1(mai_mai_n266_), .B0(mai_mai_n275_), .Y(mai_mai_n276_));
  NA2        m254(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n277_), .B(x01), .Y(mai_mai_n278_));
  NOi21      m256(.An(mai_mai_n82_), .B(mai_mai_n120_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n279_), .B(mai_mai_n278_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n280_), .B(mai_mai_n29_), .Y(mai_mai_n281_));
  NA2        m259(.A(mai_mai_n267_), .B(mai_mai_n236_), .Y(mai_mai_n282_));
  NA2        m260(.A(mai_mai_n100_), .B(x04), .Y(mai_mai_n283_));
  NA2        m261(.A(mai_mai_n283_), .B(mai_mai_n28_), .Y(mai_mai_n284_));
  OAI210     m262(.A0(mai_mai_n284_), .A1(mai_mai_n119_), .B0(mai_mai_n282_), .Y(mai_mai_n285_));
  NO3        m263(.A(mai_mai_n89_), .B(x12), .C(x03), .Y(mai_mai_n286_));
  OAI210     m264(.A0(mai_mai_n285_), .A1(mai_mai_n281_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  AOI210     m265(.A0(mai_mai_n208_), .A1(mai_mai_n203_), .B0(mai_mai_n101_), .Y(mai_mai_n288_));
  NOi21      m266(.An(mai_mai_n264_), .B(mai_mai_n226_), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n290_));
  OAI210     m268(.A0(mai_mai_n289_), .A1(mai_mai_n288_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n57_), .B(x05), .Y(mai_mai_n292_));
  NO3        m270(.A(mai_mai_n292_), .B(mai_mai_n227_), .C(mai_mai_n193_), .Y(mai_mai_n293_));
  NO2        m271(.A(mai_mai_n248_), .B(mai_mai_n28_), .Y(mai_mai_n294_));
  OAI210     m272(.A0(mai_mai_n293_), .A1(mai_mai_n234_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  NA3        m273(.A(mai_mai_n295_), .B(mai_mai_n291_), .C(mai_mai_n287_), .Y(mai_mai_n296_));
  NO3        m274(.A(mai_mai_n296_), .B(mai_mai_n276_), .C(mai_mai_n263_), .Y(mai_mai_n297_));
  OAI210     m275(.A0(mai_mai_n214_), .A1(mai_mai_n60_), .B0(mai_mai_n297_), .Y(mai02));
  AOI210     m276(.A0(mai_mai_n138_), .A1(mai_mai_n83_), .B0(mai_mai_n132_), .Y(mai_mai_n299_));
  NOi21      m277(.An(mai_mai_n242_), .B(mai_mai_n176_), .Y(mai_mai_n300_));
  NO2        m278(.A(mai_mai_n100_), .B(mai_mai_n35_), .Y(mai_mai_n301_));
  NA3        m279(.A(mai_mai_n301_), .B(mai_mai_n202_), .C(mai_mai_n55_), .Y(mai_mai_n302_));
  OAI210     m280(.A0(mai_mai_n300_), .A1(mai_mai_n32_), .B0(mai_mai_n302_), .Y(mai_mai_n303_));
  OAI210     m281(.A0(mai_mai_n303_), .A1(mai_mai_n299_), .B0(mai_mai_n173_), .Y(mai_mai_n304_));
  INV        m282(.A(mai_mai_n173_), .Y(mai_mai_n305_));
  AOI210     m283(.A0(mai_mai_n115_), .A1(mai_mai_n84_), .B0(mai_mai_n227_), .Y(mai_mai_n306_));
  OAI220     m284(.A0(mai_mai_n306_), .A1(mai_mai_n100_), .B0(mai_mai_n83_), .B1(mai_mai_n50_), .Y(mai_mai_n307_));
  AOI220     m285(.A0(mai_mai_n307_), .A1(mai_mai_n305_), .B0(mai_mai_n155_), .B1(mai_mai_n154_), .Y(mai_mai_n308_));
  AOI210     m286(.A0(mai_mai_n308_), .A1(mai_mai_n304_), .B0(mai_mai_n48_), .Y(mai_mai_n309_));
  NO2        m287(.A(x05), .B(x02), .Y(mai_mai_n310_));
  OAI210     m288(.A0(mai_mai_n218_), .A1(mai_mai_n198_), .B0(mai_mai_n310_), .Y(mai_mai_n311_));
  AOI220     m289(.A0(mai_mai_n269_), .A1(mai_mai_n57_), .B0(mai_mai_n55_), .B1(mai_mai_n36_), .Y(mai_mai_n312_));
  NO2        m290(.A(mai_mai_n311_), .B(mai_mai_n143_), .Y(mai_mai_n313_));
  NAi21      m291(.An(mai_mai_n243_), .B(mai_mai_n238_), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n256_), .B(mai_mai_n47_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n315_), .B(mai_mai_n314_), .Y(mai_mai_n316_));
  AN2        m294(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n317_));
  OAI210     m295(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n318_));
  NA2        m296(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n319_));
  OA210      m297(.A0(mai_mai_n319_), .A1(x08), .B0(mai_mai_n147_), .Y(mai_mai_n320_));
  AOI210     m298(.A0(mai_mai_n320_), .A1(mai_mai_n139_), .B0(mai_mai_n318_), .Y(mai_mai_n321_));
  OAI210     m299(.A0(mai_mai_n321_), .A1(mai_mai_n317_), .B0(mai_mai_n94_), .Y(mai_mai_n322_));
  NA3        m300(.A(mai_mai_n94_), .B(mai_mai_n82_), .C(mai_mai_n235_), .Y(mai_mai_n323_));
  NA3        m301(.A(mai_mai_n93_), .B(mai_mai_n81_), .C(mai_mai_n42_), .Y(mai_mai_n324_));
  AOI210     m302(.A0(mai_mai_n324_), .A1(mai_mai_n323_), .B0(x04), .Y(mai_mai_n325_));
  INV        m303(.A(mai_mai_n154_), .Y(mai_mai_n326_));
  OAI220     m304(.A0(mai_mai_n270_), .A1(mai_mai_n104_), .B0(mai_mai_n326_), .B1(mai_mai_n131_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n327_), .A1(x13), .B0(mai_mai_n325_), .Y(mai_mai_n328_));
  NA3        m306(.A(mai_mai_n328_), .B(mai_mai_n322_), .C(mai_mai_n316_), .Y(mai_mai_n329_));
  NO3        m307(.A(mai_mai_n329_), .B(mai_mai_n313_), .C(mai_mai_n309_), .Y(mai_mai_n330_));
  NA2        m308(.A(mai_mai_n142_), .B(x03), .Y(mai_mai_n331_));
  INV        m309(.A(mai_mai_n187_), .Y(mai_mai_n332_));
  AOI220     m310(.A0(x08), .A1(mai_mai_n332_), .B0(mai_mai_n209_), .B1(x08), .Y(mai_mai_n333_));
  OAI210     m311(.A0(mai_mai_n333_), .A1(mai_mai_n292_), .B0(mai_mai_n331_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n334_), .B(mai_mai_n106_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n172_), .B(mai_mai_n166_), .Y(mai_mai_n336_));
  AN2        m314(.A(mai_mai_n336_), .B(mai_mai_n179_), .Y(mai_mai_n337_));
  NO2        m315(.A(mai_mai_n132_), .B(mai_mai_n28_), .Y(mai_mai_n338_));
  OAI210     m316(.A0(mai_mai_n338_), .A1(mai_mai_n337_), .B0(mai_mai_n107_), .Y(mai_mai_n339_));
  NA2        m317(.A(mai_mai_n283_), .B(mai_mai_n99_), .Y(mai_mai_n340_));
  NA2        m318(.A(mai_mai_n99_), .B(mai_mai_n41_), .Y(mai_mai_n341_));
  NA3        m319(.A(mai_mai_n341_), .B(mai_mai_n340_), .C(mai_mai_n131_), .Y(mai_mai_n342_));
  NA4        m320(.A(mai_mai_n342_), .B(mai_mai_n339_), .C(mai_mai_n335_), .D(mai_mai_n48_), .Y(mai_mai_n343_));
  INV        m321(.A(mai_mai_n209_), .Y(mai_mai_n344_));
  NO2        m322(.A(mai_mai_n167_), .B(mai_mai_n40_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n346_));
  OAI220     m324(.A0(mai_mai_n346_), .A1(mai_mai_n345_), .B0(mai_mai_n344_), .B1(mai_mai_n58_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n347_), .B(x02), .Y(mai_mai_n348_));
  INV        m326(.A(mai_mai_n249_), .Y(mai_mai_n349_));
  NA2        m327(.A(mai_mai_n206_), .B(x04), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n351_));
  NO3        m329(.A(mai_mai_n189_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n352_));
  OAI210     m330(.A0(mai_mai_n352_), .A1(mai_mai_n351_), .B0(mai_mai_n94_), .Y(mai_mai_n353_));
  NO3        m331(.A(mai_mai_n206_), .B(mai_mai_n165_), .C(mai_mai_n51_), .Y(mai_mai_n354_));
  OAI210     m332(.A0(mai_mai_n149_), .A1(mai_mai_n36_), .B0(mai_mai_n99_), .Y(mai_mai_n355_));
  OAI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n199_), .B0(mai_mai_n354_), .Y(mai_mai_n356_));
  NA4        m334(.A(mai_mai_n356_), .B(mai_mai_n353_), .C(mai_mai_n348_), .D(x06), .Y(mai_mai_n357_));
  NA2        m335(.A(x09), .B(x03), .Y(mai_mai_n358_));
  OAI220     m336(.A0(mai_mai_n358_), .A1(mai_mai_n130_), .B0(mai_mai_n217_), .B1(mai_mai_n63_), .Y(mai_mai_n359_));
  OAI220     m337(.A0(mai_mai_n166_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n360_));
  NO3        m338(.A(mai_mai_n292_), .B(mai_mai_n129_), .C(x08), .Y(mai_mai_n361_));
  AOI210     m339(.A0(mai_mai_n360_), .A1(mai_mai_n234_), .B0(mai_mai_n361_), .Y(mai_mai_n362_));
  NO2        m340(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n363_));
  NO3        m341(.A(mai_mai_n113_), .B(mai_mai_n130_), .C(mai_mai_n38_), .Y(mai_mai_n364_));
  AOI210     m342(.A0(mai_mai_n354_), .A1(mai_mai_n363_), .B0(mai_mai_n364_), .Y(mai_mai_n365_));
  OAI210     m343(.A0(mai_mai_n362_), .A1(mai_mai_n28_), .B0(mai_mai_n365_), .Y(mai_mai_n366_));
  AO220      m344(.A0(mai_mai_n366_), .A1(x04), .B0(mai_mai_n359_), .B1(x05), .Y(mai_mai_n367_));
  AOI210     m345(.A0(mai_mai_n357_), .A1(mai_mai_n343_), .B0(mai_mai_n367_), .Y(mai_mai_n368_));
  OAI210     m346(.A0(mai_mai_n330_), .A1(x12), .B0(mai_mai_n368_), .Y(mai03));
  OR2        m347(.A(mai_mai_n42_), .B(mai_mai_n235_), .Y(mai_mai_n370_));
  AOI210     m348(.A0(mai_mai_n155_), .A1(mai_mai_n99_), .B0(mai_mai_n370_), .Y(mai_mai_n371_));
  AO210      m349(.A0(mai_mai_n349_), .A1(mai_mai_n84_), .B0(mai_mai_n350_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n206_), .B(mai_mai_n154_), .Y(mai_mai_n373_));
  NA3        m351(.A(mai_mai_n373_), .B(mai_mai_n372_), .C(mai_mai_n210_), .Y(mai_mai_n374_));
  OAI210     m352(.A0(mai_mai_n374_), .A1(mai_mai_n371_), .B0(x05), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n370_), .B(x05), .Y(mai_mai_n376_));
  AOI210     m354(.A0(mai_mai_n139_), .A1(mai_mai_n223_), .B0(mai_mai_n376_), .Y(mai_mai_n377_));
  AOI210     m355(.A0(mai_mai_n237_), .A1(mai_mai_n78_), .B0(mai_mai_n123_), .Y(mai_mai_n378_));
  OAI220     m356(.A0(mai_mai_n378_), .A1(mai_mai_n58_), .B0(mai_mai_n319_), .B1(mai_mai_n312_), .Y(mai_mai_n379_));
  OAI210     m357(.A0(mai_mai_n379_), .A1(mai_mai_n377_), .B0(mai_mai_n99_), .Y(mai_mai_n380_));
  AOI210     m358(.A0(mai_mai_n147_), .A1(mai_mai_n59_), .B0(mai_mai_n38_), .Y(mai_mai_n381_));
  NO2        m359(.A(mai_mai_n176_), .B(mai_mai_n134_), .Y(mai_mai_n382_));
  OAI220     m360(.A0(mai_mai_n382_), .A1(mai_mai_n37_), .B0(mai_mai_n150_), .B1(x13), .Y(mai_mai_n383_));
  OAI210     m361(.A0(mai_mai_n383_), .A1(mai_mai_n381_), .B0(x04), .Y(mai_mai_n384_));
  NO3        m362(.A(mai_mai_n341_), .B(mai_mai_n83_), .C(mai_mai_n58_), .Y(mai_mai_n385_));
  AOI210     m363(.A0(mai_mai_n195_), .A1(mai_mai_n99_), .B0(mai_mai_n147_), .Y(mai_mai_n386_));
  OA210      m364(.A0(mai_mai_n167_), .A1(x12), .B0(mai_mai_n134_), .Y(mai_mai_n387_));
  NO3        m365(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(mai_mai_n385_), .Y(mai_mai_n388_));
  NA4        m366(.A(mai_mai_n388_), .B(mai_mai_n384_), .C(mai_mai_n380_), .D(mai_mai_n375_), .Y(mai04));
  NO2        m367(.A(mai_mai_n87_), .B(mai_mai_n39_), .Y(mai_mai_n390_));
  XO2        m368(.A(mai_mai_n390_), .B(mai_mai_n259_), .Y(mai05));
  AOI210     m369(.A0(mai_mai_n458_), .A1(mai_mai_n318_), .B0(mai_mai_n25_), .Y(mai_mai_n392_));
  NO2        m370(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n393_));
  OAI210     m371(.A0(mai_mai_n393_), .A1(mai_mai_n392_), .B0(mai_mai_n99_), .Y(mai_mai_n394_));
  NA2        m372(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n395_));
  NA2        m373(.A(mai_mai_n264_), .B(x03), .Y(mai_mai_n396_));
  OAI210     m374(.A0(mai_mai_n26_), .A1(mai_mai_n99_), .B0(x07), .Y(mai_mai_n397_));
  INV        m375(.A(mai_mai_n397_), .Y(mai_mai_n398_));
  AOI220     m376(.A0(mai_mai_n79_), .A1(mai_mai_n31_), .B0(mai_mai_n51_), .B1(mai_mai_n50_), .Y(mai_mai_n399_));
  NO3        m377(.A(mai_mai_n399_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n70_), .B(x02), .Y(mai_mai_n401_));
  AOI210     m379(.A0(mai_mai_n401_), .A1(mai_mai_n396_), .B0(mai_mai_n267_), .Y(mai_mai_n402_));
  OR2        m380(.A(mai_mai_n402_), .B(mai_mai_n248_), .Y(mai_mai_n403_));
  NA2        m381(.A(mai_mai_n161_), .B(x05), .Y(mai_mai_n404_));
  NA3        m382(.A(mai_mai_n404_), .B(mai_mai_n252_), .C(mai_mai_n246_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n406_));
  OAI210     m384(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n407_));
  OR3        m385(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(mai_mai_n44_), .Y(mai_mai_n408_));
  NA3        m386(.A(mai_mai_n408_), .B(mai_mai_n405_), .C(mai_mai_n403_), .Y(mai_mai_n409_));
  OAI210     m387(.A0(mai_mai_n409_), .A1(mai_mai_n400_), .B0(mai_mai_n99_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n33_), .B(mai_mai_n99_), .Y(mai_mai_n411_));
  AOI210     m389(.A0(mai_mai_n411_), .A1(mai_mai_n90_), .B0(x07), .Y(mai_mai_n412_));
  AOI220     m390(.A0(mai_mai_n412_), .A1(mai_mai_n410_), .B0(mai_mai_n398_), .B1(mai_mai_n394_), .Y(mai_mai_n413_));
  AOI210     m391(.A0(mai_mai_n406_), .A1(x07), .B0(mai_mai_n142_), .Y(mai_mai_n414_));
  OR2        m392(.A(mai_mai_n414_), .B(x03), .Y(mai_mai_n415_));
  NO2        m393(.A(x07), .B(x11), .Y(mai_mai_n416_));
  NO3        m394(.A(mai_mai_n416_), .B(mai_mai_n146_), .C(mai_mai_n28_), .Y(mai_mai_n417_));
  AOI210     m395(.A0(mai_mai_n417_), .A1(mai_mai_n415_), .B0(mai_mai_n47_), .Y(mai_mai_n418_));
  NO4        m396(.A(mai_mai_n341_), .B(mai_mai_n32_), .C(x11), .D(x09), .Y(mai_mai_n419_));
  OAI210     m397(.A0(mai_mai_n419_), .A1(mai_mai_n418_), .B0(mai_mai_n100_), .Y(mai_mai_n420_));
  AOI210     m398(.A0(mai_mai_n350_), .A1(mai_mai_n109_), .B0(mai_mai_n273_), .Y(mai_mai_n421_));
  NOi21      m399(.An(mai_mai_n331_), .B(mai_mai_n134_), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n422_), .B(mai_mai_n274_), .Y(mai_mai_n423_));
  OAI210     m401(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n424_));
  AOI210     m402(.A0(mai_mai_n259_), .A1(mai_mai_n47_), .B0(mai_mai_n424_), .Y(mai_mai_n425_));
  NO4        m403(.A(mai_mai_n425_), .B(mai_mai_n423_), .C(mai_mai_n421_), .D(x08), .Y(mai_mai_n426_));
  AOI210     m404(.A0(mai_mai_n406_), .A1(mai_mai_n28_), .B0(mai_mai_n31_), .Y(mai_mai_n427_));
  NA2        m405(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n428_));
  NO2        m406(.A(mai_mai_n428_), .B(mai_mai_n427_), .Y(mai_mai_n429_));
  NO2        m407(.A(x13), .B(x12), .Y(mai_mai_n430_));
  NO2        m408(.A(mai_mai_n132_), .B(mai_mai_n28_), .Y(mai_mai_n431_));
  NO2        m409(.A(mai_mai_n431_), .B(mai_mai_n278_), .Y(mai_mai_n432_));
  OR3        m410(.A(mai_mai_n432_), .B(x12), .C(x03), .Y(mai_mai_n433_));
  NA3        m411(.A(mai_mai_n344_), .B(mai_mai_n125_), .C(x12), .Y(mai_mai_n434_));
  AO210      m412(.A0(mai_mai_n344_), .A1(mai_mai_n125_), .B0(mai_mai_n259_), .Y(mai_mai_n435_));
  NA4        m413(.A(mai_mai_n435_), .B(mai_mai_n434_), .C(mai_mai_n433_), .D(x08), .Y(mai_mai_n436_));
  AOI210     m414(.A0(mai_mai_n430_), .A1(mai_mai_n429_), .B0(mai_mai_n436_), .Y(mai_mai_n437_));
  AOI210     m415(.A0(mai_mai_n426_), .A1(mai_mai_n420_), .B0(mai_mai_n437_), .Y(mai_mai_n438_));
  OAI210     m416(.A0(x07), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n439_));
  OAI220     m417(.A0(mai_mai_n457_), .A1(mai_mai_n395_), .B0(mai_mai_n146_), .B1(mai_mai_n43_), .Y(mai_mai_n440_));
  OAI210     m418(.A0(mai_mai_n440_), .A1(mai_mai_n439_), .B0(mai_mai_n194_), .Y(mai_mai_n441_));
  NA3        m419(.A(mai_mai_n432_), .B(mai_mai_n422_), .C(mai_mai_n340_), .Y(mai_mai_n442_));
  INV        m420(.A(x14), .Y(mai_mai_n443_));
  NO3        m421(.A(mai_mai_n331_), .B(mai_mai_n104_), .C(x11), .Y(mai_mai_n444_));
  NO3        m422(.A(x06), .B(mai_mai_n341_), .C(mai_mai_n187_), .Y(mai_mai_n445_));
  NO3        m423(.A(mai_mai_n445_), .B(mai_mai_n444_), .C(mai_mai_n443_), .Y(mai_mai_n446_));
  NA3        m424(.A(mai_mai_n446_), .B(mai_mai_n442_), .C(mai_mai_n441_), .Y(mai_mai_n447_));
  AOI220     m425(.A0(mai_mai_n411_), .A1(mai_mai_n60_), .B0(mai_mai_n431_), .B1(mai_mai_n165_), .Y(mai_mai_n448_));
  NOi21      m426(.An(mai_mai_n283_), .B(mai_mai_n150_), .Y(mai_mai_n449_));
  NO2        m427(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n450_));
  OAI210     m428(.A0(mai_mai_n450_), .A1(mai_mai_n449_), .B0(mai_mai_n99_), .Y(mai_mai_n451_));
  OAI210     m429(.A0(mai_mai_n448_), .A1(mai_mai_n89_), .B0(mai_mai_n451_), .Y(mai_mai_n452_));
  NO4        m430(.A(mai_mai_n452_), .B(mai_mai_n447_), .C(mai_mai_n438_), .D(mai_mai_n413_), .Y(mai06));
  INV        m431(.A(x07), .Y(mai_mai_n456_));
  INV        m432(.A(x07), .Y(mai_mai_n457_));
  INV        m433(.A(mai_mai_n51_), .Y(mai_mai_n458_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  INV        u039(.A(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  NO2        u042(.A(men_men_n64_), .B(men_men_n62_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  AOI210     u048(.A0(men_men_n70_), .A1(men_men_n61_), .B0(men_men_n23_), .Y(men_men_n71_));
  NA2        u049(.A(x09), .B(x05), .Y(men_men_n72_));
  NA2        u050(.A(x10), .B(x06), .Y(men_men_n73_));
  NA3        u051(.A(men_men_n73_), .B(men_men_n72_), .C(men_men_n28_), .Y(men_men_n74_));
  NO2        u052(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n75_));
  OAI210     u053(.A0(men_men_n74_), .A1(men_men_n71_), .B0(x03), .Y(men_men_n76_));
  NOi31      u054(.An(x08), .B(x04), .C(x00), .Y(men_men_n77_));
  NO2        u055(.A(x10), .B(x09), .Y(men_men_n78_));
  AOI210     u056(.A0(men_men_n466_), .A1(men_men_n77_), .B0(men_men_n24_), .Y(men_men_n79_));
  NO2        u057(.A(x09), .B(men_men_n41_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n80_), .B(men_men_n36_), .Y(men_men_n81_));
  OAI210     u059(.A0(men_men_n80_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n82_));
  AOI210     u060(.A0(men_men_n81_), .A1(men_men_n48_), .B0(men_men_n82_), .Y(men_men_n83_));
  NO2        u061(.A(men_men_n36_), .B(x00), .Y(men_men_n84_));
  NO2        u062(.A(x08), .B(x01), .Y(men_men_n85_));
  OAI210     u063(.A0(men_men_n85_), .A1(men_men_n84_), .B0(men_men_n35_), .Y(men_men_n86_));
  NA2        u064(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n87_));
  NO3        u065(.A(men_men_n86_), .B(men_men_n83_), .C(men_men_n79_), .Y(men_men_n88_));
  AN2        u066(.A(men_men_n88_), .B(men_men_n76_), .Y(men_men_n89_));
  INV        u067(.A(men_men_n86_), .Y(men_men_n90_));
  NO2        u068(.A(x06), .B(x05), .Y(men_men_n91_));
  NA2        u069(.A(x11), .B(x00), .Y(men_men_n92_));
  NO2        u070(.A(x11), .B(men_men_n47_), .Y(men_men_n93_));
  NOi21      u071(.An(men_men_n92_), .B(men_men_n93_), .Y(men_men_n94_));
  AOI210     u072(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n94_), .Y(men_men_n95_));
  NOi21      u073(.An(x01), .B(x10), .Y(men_men_n96_));
  NO2        u074(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n97_));
  NO3        u075(.A(men_men_n97_), .B(men_men_n96_), .C(x06), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n98_), .B(men_men_n27_), .Y(men_men_n99_));
  OAI210     u077(.A0(men_men_n95_), .A1(x07), .B0(men_men_n99_), .Y(men_men_n100_));
  NO3        u078(.A(men_men_n100_), .B(men_men_n89_), .C(men_men_n69_), .Y(men01));
  INV        u079(.A(x12), .Y(men_men_n102_));
  INV        u080(.A(x13), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n91_), .B(x01), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n104_), .B(men_men_n70_), .Y(men_men_n105_));
  NA2        u083(.A(x08), .B(x04), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n57_), .Y(men_men_n107_));
  NA2        u085(.A(men_men_n107_), .B(men_men_n105_), .Y(men_men_n108_));
  NA2        u086(.A(men_men_n96_), .B(men_men_n28_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n72_), .Y(men_men_n110_));
  NO2        u088(.A(x10), .B(x01), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n29_), .B(x00), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NA2        u091(.A(x04), .B(men_men_n28_), .Y(men_men_n114_));
  NO3        u092(.A(men_men_n114_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n115_));
  AOI210     u093(.A0(men_men_n115_), .A1(men_men_n113_), .B0(men_men_n110_), .Y(men_men_n116_));
  AOI210     u094(.A0(men_men_n116_), .A1(men_men_n108_), .B0(men_men_n103_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n56_), .B(x05), .Y(men_men_n118_));
  NOi21      u096(.An(men_men_n118_), .B(men_men_n58_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n35_), .B(x02), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n103_), .B(men_men_n36_), .Y(men_men_n121_));
  NA3        u099(.A(men_men_n121_), .B(men_men_n120_), .C(x06), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(men_men_n119_), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n85_), .B(x13), .Y(men_men_n124_));
  NA2        u102(.A(x09), .B(men_men_n35_), .Y(men_men_n125_));
  NO2        u103(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n126_));
  NA2        u104(.A(x13), .B(men_men_n35_), .Y(men_men_n127_));
  NO2        u105(.A(men_men_n127_), .B(x05), .Y(men_men_n128_));
  NO2        u106(.A(men_men_n128_), .B(men_men_n126_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n130_));
  AOI210     u108(.A0(men_men_n57_), .A1(men_men_n81_), .B0(men_men_n119_), .Y(men_men_n131_));
  AOI210     u109(.A0(men_men_n131_), .A1(men_men_n129_), .B0(men_men_n73_), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n133_));
  NA2        u111(.A(x10), .B(men_men_n57_), .Y(men_men_n134_));
  NA2        u112(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n51_), .B(x05), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n36_), .B(x04), .Y(men_men_n137_));
  NA3        u115(.A(men_men_n137_), .B(men_men_n136_), .C(x13), .Y(men_men_n138_));
  NO3        u116(.A(men_men_n130_), .B(men_men_n80_), .C(men_men_n36_), .Y(men_men_n139_));
  NO2        u117(.A(men_men_n60_), .B(x05), .Y(men_men_n140_));
  NOi41      u118(.An(men_men_n138_), .B(men_men_n140_), .C(men_men_n139_), .D(men_men_n135_), .Y(men_men_n141_));
  NO3        u119(.A(men_men_n141_), .B(x06), .C(x03), .Y(men_men_n142_));
  NO4        u120(.A(men_men_n142_), .B(men_men_n132_), .C(men_men_n123_), .D(men_men_n117_), .Y(men_men_n143_));
  NA2        u121(.A(x13), .B(men_men_n36_), .Y(men_men_n144_));
  OAI210     u122(.A0(men_men_n85_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n145_));
  NA2        u123(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n146_));
  NOi21      u124(.An(men_men_n91_), .B(men_men_n57_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n148_));
  OA210      u126(.A0(men_men_n147_), .A1(men_men_n78_), .B0(men_men_n148_), .Y(men_men_n149_));
  NO2        u127(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n29_), .B(x06), .Y(men_men_n151_));
  AN2        u129(.A(men_men_n149_), .B(men_men_n146_), .Y(men_men_n152_));
  NO2        u130(.A(x09), .B(x05), .Y(men_men_n153_));
  NA2        u131(.A(men_men_n153_), .B(men_men_n47_), .Y(men_men_n154_));
  AOI210     u132(.A0(men_men_n154_), .A1(men_men_n113_), .B0(men_men_n49_), .Y(men_men_n155_));
  NA2        u133(.A(x09), .B(x00), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n118_), .B(men_men_n156_), .Y(men_men_n157_));
  NA2        u135(.A(men_men_n77_), .B(men_men_n51_), .Y(men_men_n158_));
  AOI210     u136(.A0(men_men_n158_), .A1(men_men_n157_), .B0(men_men_n151_), .Y(men_men_n159_));
  NO3        u137(.A(men_men_n159_), .B(men_men_n155_), .C(men_men_n152_), .Y(men_men_n160_));
  NO2        u138(.A(x03), .B(x02), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n86_), .B(men_men_n103_), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n162_), .A1(men_men_n119_), .B0(men_men_n161_), .Y(men_men_n163_));
  OA210      u141(.A0(men_men_n160_), .A1(x11), .B0(men_men_n163_), .Y(men_men_n164_));
  OAI210     u142(.A0(men_men_n143_), .A1(men_men_n23_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u143(.A(men_men_n113_), .B(men_men_n40_), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n167_));
  NAi21      u145(.An(x06), .B(x10), .Y(men_men_n168_));
  NOi21      u146(.An(x01), .B(x13), .Y(men_men_n169_));
  NA2        u147(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  OR2        u148(.A(men_men_n170_), .B(men_men_n167_), .Y(men_men_n171_));
  AOI210     u149(.A0(men_men_n171_), .A1(men_men_n166_), .B0(men_men_n41_), .Y(men_men_n172_));
  NO2        u150(.A(men_men_n29_), .B(x03), .Y(men_men_n173_));
  NA2        u151(.A(men_men_n103_), .B(x01), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n174_), .B(x08), .Y(men_men_n175_));
  OAI210     u153(.A0(x05), .A1(men_men_n175_), .B0(men_men_n51_), .Y(men_men_n176_));
  AOI210     u154(.A0(men_men_n176_), .A1(men_men_n173_), .B0(men_men_n48_), .Y(men_men_n177_));
  AOI210     u155(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n177_), .A1(men_men_n172_), .B0(men_men_n178_), .Y(men_men_n179_));
  NA2        u157(.A(x04), .B(x02), .Y(men_men_n180_));
  NA2        u158(.A(x10), .B(x05), .Y(men_men_n181_));
  NA2        u159(.A(x09), .B(x06), .Y(men_men_n182_));
  AOI210     u160(.A0(men_men_n182_), .A1(men_men_n181_), .B0(men_men_n167_), .Y(men_men_n183_));
  NO2        u161(.A(x09), .B(x01), .Y(men_men_n184_));
  NO3        u162(.A(men_men_n184_), .B(men_men_n111_), .C(men_men_n31_), .Y(men_men_n185_));
  OAI210     u163(.A0(men_men_n185_), .A1(men_men_n183_), .B0(x00), .Y(men_men_n186_));
  NO2        u164(.A(men_men_n118_), .B(x08), .Y(men_men_n187_));
  NA3        u165(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n51_), .Y(men_men_n188_));
  NA2        u166(.A(men_men_n96_), .B(x05), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n121_), .B0(men_men_n188_), .Y(men_men_n190_));
  AOI210     u168(.A0(men_men_n187_), .A1(x06), .B0(men_men_n190_), .Y(men_men_n191_));
  OAI210     u169(.A0(men_men_n191_), .A1(x11), .B0(men_men_n186_), .Y(men_men_n192_));
  NAi21      u170(.An(men_men_n180_), .B(men_men_n192_), .Y(men_men_n193_));
  INV        u171(.A(men_men_n25_), .Y(men_men_n194_));
  NAi21      u172(.An(x13), .B(x00), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n195_), .Y(men_men_n196_));
  AOI220     u174(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n197_));
  OAI210     u175(.A0(men_men_n181_), .A1(men_men_n35_), .B0(men_men_n197_), .Y(men_men_n198_));
  AN2        u176(.A(men_men_n198_), .B(men_men_n196_), .Y(men_men_n199_));
  NO2        u177(.A(men_men_n195_), .B(men_men_n36_), .Y(men_men_n200_));
  INV        u178(.A(men_men_n200_), .Y(men_men_n201_));
  OAI210     u179(.A0(men_men_n201_), .A1(men_men_n182_), .B0(men_men_n73_), .Y(men_men_n202_));
  OAI210     u180(.A0(men_men_n202_), .A1(men_men_n199_), .B0(men_men_n194_), .Y(men_men_n203_));
  NOi21      u181(.An(x09), .B(x00), .Y(men_men_n204_));
  NO3        u182(.A(men_men_n84_), .B(men_men_n204_), .C(men_men_n47_), .Y(men_men_n205_));
  NA2        u183(.A(men_men_n205_), .B(men_men_n134_), .Y(men_men_n206_));
  NA2        u184(.A(x10), .B(x08), .Y(men_men_n207_));
  INV        u185(.A(men_men_n207_), .Y(men_men_n208_));
  NA2        u186(.A(x06), .B(x05), .Y(men_men_n209_));
  OAI210     u187(.A0(men_men_n209_), .A1(men_men_n35_), .B0(men_men_n102_), .Y(men_men_n210_));
  AOI210     u188(.A0(men_men_n208_), .A1(men_men_n58_), .B0(men_men_n210_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n211_), .B(men_men_n206_), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n103_), .B(x12), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n213_), .Y(men_men_n214_));
  NA2        u192(.A(men_men_n96_), .B(men_men_n51_), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n216_), .B(x02), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n217_), .B(men_men_n215_), .Y(men_men_n218_));
  AOI210     u196(.A0(men_men_n214_), .A1(men_men_n212_), .B0(men_men_n218_), .Y(men_men_n219_));
  NA4        u197(.A(men_men_n219_), .B(men_men_n203_), .C(men_men_n193_), .D(men_men_n179_), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n165_), .A1(men_men_n102_), .B0(men_men_n220_), .Y(men_men_n221_));
  NA2        u199(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n222_), .B(men_men_n145_), .Y(men_men_n223_));
  AOI210     u201(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n133_), .B(x06), .Y(men_men_n225_));
  AOI210     u203(.A0(men_men_n224_), .A1(men_men_n223_), .B0(men_men_n225_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n226_), .B(x12), .Y(men_men_n227_));
  INV        u205(.A(men_men_n77_), .Y(men_men_n228_));
  AOI210     u206(.A0(men_men_n207_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n229_), .A1(men_men_n170_), .B0(men_men_n57_), .Y(men_men_n230_));
  NA2        u208(.A(men_men_n230_), .B(men_men_n228_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n96_), .B(x06), .Y(men_men_n232_));
  AOI210     u210(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n233_));
  NO3        u211(.A(men_men_n233_), .B(men_men_n232_), .C(men_men_n41_), .Y(men_men_n234_));
  NA4        u212(.A(men_men_n168_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n235_));
  NA2        u213(.A(men_men_n235_), .B(men_men_n151_), .Y(men_men_n236_));
  OAI210     u214(.A0(men_men_n236_), .A1(men_men_n234_), .B0(x02), .Y(men_men_n237_));
  AOI210     u215(.A0(men_men_n237_), .A1(men_men_n231_), .B0(men_men_n23_), .Y(men_men_n238_));
  OAI210     u216(.A0(men_men_n227_), .A1(men_men_n57_), .B0(men_men_n238_), .Y(men_men_n239_));
  INV        u217(.A(men_men_n151_), .Y(men_men_n240_));
  NO2        u218(.A(men_men_n51_), .B(x03), .Y(men_men_n241_));
  OAI210     u219(.A0(men_men_n80_), .A1(men_men_n36_), .B0(men_men_n125_), .Y(men_men_n242_));
  NO2        u220(.A(men_men_n103_), .B(x03), .Y(men_men_n243_));
  AOI220     u221(.A0(men_men_n243_), .A1(men_men_n242_), .B0(men_men_n77_), .B1(men_men_n241_), .Y(men_men_n244_));
  NA2        u222(.A(men_men_n32_), .B(x06), .Y(men_men_n245_));
  INV        u223(.A(men_men_n168_), .Y(men_men_n246_));
  NOi21      u224(.An(x13), .B(x04), .Y(men_men_n247_));
  NO3        u225(.A(men_men_n247_), .B(men_men_n77_), .C(men_men_n204_), .Y(men_men_n248_));
  NO2        u226(.A(men_men_n248_), .B(x05), .Y(men_men_n249_));
  AOI220     u227(.A0(men_men_n249_), .A1(men_men_n245_), .B0(men_men_n246_), .B1(men_men_n57_), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n240_), .B0(men_men_n250_), .Y(men_men_n251_));
  INV        u229(.A(men_men_n93_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(x12), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n255_));
  OAI210     u233(.A0(men_men_n255_), .A1(men_men_n198_), .B0(men_men_n196_), .Y(men_men_n256_));
  AOI210     u234(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n257_));
  NA2        u235(.A(men_men_n156_), .B(men_men_n73_), .Y(men_men_n258_));
  INV        u236(.A(men_men_n258_), .Y(men_men_n259_));
  NA2        u237(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n260_), .B(x03), .Y(men_men_n261_));
  OA210      u239(.A0(men_men_n261_), .A1(men_men_n259_), .B0(men_men_n256_), .Y(men_men_n262_));
  NA2        u240(.A(x13), .B(men_men_n102_), .Y(men_men_n263_));
  NA3        u241(.A(men_men_n263_), .B(men_men_n210_), .C(men_men_n94_), .Y(men_men_n264_));
  OAI210     u242(.A0(men_men_n262_), .A1(men_men_n254_), .B0(men_men_n264_), .Y(men_men_n265_));
  AOI210     u243(.A0(men_men_n253_), .A1(men_men_n251_), .B0(men_men_n265_), .Y(men_men_n266_));
  AOI210     u244(.A0(men_men_n266_), .A1(men_men_n239_), .B0(x07), .Y(men_men_n267_));
  NA2        u245(.A(men_men_n72_), .B(men_men_n29_), .Y(men_men_n268_));
  AOI210     u246(.A0(men_men_n144_), .A1(men_men_n158_), .B0(men_men_n268_), .Y(men_men_n269_));
  NO2        u247(.A(men_men_n103_), .B(x06), .Y(men_men_n270_));
  INV        u248(.A(men_men_n270_), .Y(men_men_n271_));
  NO2        u249(.A(x08), .B(x05), .Y(men_men_n272_));
  NO2        u250(.A(men_men_n272_), .B(men_men_n257_), .Y(men_men_n273_));
  OAI210     u251(.A0(men_men_n77_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n273_), .A1(men_men_n271_), .B0(men_men_n274_), .Y(men_men_n275_));
  NO2        u253(.A(x12), .B(x02), .Y(men_men_n276_));
  INV        u254(.A(men_men_n276_), .Y(men_men_n277_));
  NO2        u255(.A(men_men_n277_), .B(men_men_n252_), .Y(men_men_n278_));
  OA210      u256(.A0(men_men_n275_), .A1(men_men_n269_), .B0(men_men_n278_), .Y(men_men_n279_));
  NA2        u257(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n280_));
  NO2        u258(.A(men_men_n280_), .B(x01), .Y(men_men_n281_));
  NOi21      u259(.An(men_men_n85_), .B(men_men_n125_), .Y(men_men_n282_));
  NO2        u260(.A(men_men_n282_), .B(men_men_n281_), .Y(men_men_n283_));
  AOI210     u261(.A0(men_men_n283_), .A1(men_men_n138_), .B0(men_men_n29_), .Y(men_men_n284_));
  NA2        u262(.A(men_men_n270_), .B(men_men_n242_), .Y(men_men_n285_));
  NA2        u263(.A(men_men_n103_), .B(x04), .Y(men_men_n286_));
  NA2        u264(.A(men_men_n286_), .B(men_men_n28_), .Y(men_men_n287_));
  OAI210     u265(.A0(men_men_n287_), .A1(men_men_n124_), .B0(men_men_n285_), .Y(men_men_n288_));
  NO3        u266(.A(men_men_n92_), .B(x12), .C(x03), .Y(men_men_n289_));
  OAI210     u267(.A0(men_men_n288_), .A1(men_men_n284_), .B0(men_men_n289_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n215_), .A1(men_men_n209_), .B0(men_men_n106_), .Y(men_men_n291_));
  NOi21      u269(.An(men_men_n268_), .B(men_men_n232_), .Y(men_men_n292_));
  NO2        u270(.A(men_men_n25_), .B(x00), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n292_), .A1(men_men_n291_), .B0(men_men_n293_), .Y(men_men_n294_));
  NO2        u272(.A(men_men_n58_), .B(x05), .Y(men_men_n295_));
  NO2        u273(.A(men_men_n254_), .B(men_men_n28_), .Y(men_men_n296_));
  NA2        u274(.A(men_men_n240_), .B(men_men_n296_), .Y(men_men_n297_));
  NA3        u275(.A(men_men_n297_), .B(men_men_n294_), .C(men_men_n290_), .Y(men_men_n298_));
  NO3        u276(.A(men_men_n298_), .B(men_men_n279_), .C(men_men_n267_), .Y(men_men_n299_));
  OAI210     u277(.A0(men_men_n221_), .A1(men_men_n61_), .B0(men_men_n299_), .Y(men02));
  NOi21      u278(.An(men_men_n248_), .B(men_men_n184_), .Y(men_men_n301_));
  NO2        u279(.A(men_men_n103_), .B(men_men_n35_), .Y(men_men_n302_));
  NA3        u280(.A(men_men_n302_), .B(men_men_n208_), .C(men_men_n56_), .Y(men_men_n303_));
  OAI210     u281(.A0(men_men_n301_), .A1(men_men_n32_), .B0(men_men_n303_), .Y(men_men_n304_));
  NA2        u282(.A(men_men_n304_), .B(men_men_n181_), .Y(men_men_n305_));
  INV        u283(.A(men_men_n181_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n120_), .A1(men_men_n87_), .B0(men_men_n233_), .Y(men_men_n307_));
  OAI220     u285(.A0(men_men_n307_), .A1(men_men_n103_), .B0(men_men_n86_), .B1(men_men_n51_), .Y(men_men_n308_));
  AOI220     u286(.A0(men_men_n308_), .A1(men_men_n306_), .B0(men_men_n162_), .B1(men_men_n161_), .Y(men_men_n309_));
  AOI210     u287(.A0(men_men_n309_), .A1(men_men_n305_), .B0(men_men_n48_), .Y(men_men_n310_));
  NO2        u288(.A(x05), .B(x02), .Y(men_men_n311_));
  OAI210     u289(.A0(men_men_n223_), .A1(men_men_n204_), .B0(men_men_n311_), .Y(men_men_n312_));
  AOI220     u290(.A0(men_men_n272_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n313_));
  NOi21      u291(.An(men_men_n302_), .B(men_men_n313_), .Y(men_men_n314_));
  AOI210     u292(.A0(men_men_n247_), .A1(men_men_n80_), .B0(men_men_n314_), .Y(men_men_n315_));
  AOI210     u293(.A0(men_men_n315_), .A1(men_men_n312_), .B0(men_men_n151_), .Y(men_men_n316_));
  NAi21      u294(.An(men_men_n249_), .B(men_men_n244_), .Y(men_men_n317_));
  NO2        u295(.A(men_men_n260_), .B(men_men_n47_), .Y(men_men_n318_));
  NA2        u296(.A(men_men_n318_), .B(men_men_n317_), .Y(men_men_n319_));
  AN2        u297(.A(men_men_n243_), .B(men_men_n242_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n321_));
  NA2        u299(.A(x13), .B(men_men_n28_), .Y(men_men_n322_));
  AOI210     u300(.A0(men_men_n154_), .A1(men_men_n145_), .B0(men_men_n321_), .Y(men_men_n323_));
  OAI210     u301(.A0(men_men_n323_), .A1(men_men_n320_), .B0(men_men_n97_), .Y(men_men_n324_));
  NA3        u302(.A(men_men_n97_), .B(men_men_n85_), .C(men_men_n241_), .Y(men_men_n325_));
  NA3        u303(.A(men_men_n96_), .B(men_men_n84_), .C(men_men_n42_), .Y(men_men_n326_));
  AOI210     u304(.A0(men_men_n326_), .A1(men_men_n325_), .B0(x04), .Y(men_men_n327_));
  INV        u305(.A(men_men_n161_), .Y(men_men_n328_));
  OAI220     u306(.A0(men_men_n273_), .A1(men_men_n109_), .B0(men_men_n328_), .B1(men_men_n135_), .Y(men_men_n329_));
  AOI210     u307(.A0(men_men_n329_), .A1(x13), .B0(men_men_n327_), .Y(men_men_n330_));
  NA3        u308(.A(men_men_n330_), .B(men_men_n324_), .C(men_men_n319_), .Y(men_men_n331_));
  NO3        u309(.A(men_men_n331_), .B(men_men_n316_), .C(men_men_n310_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n150_), .B(x03), .Y(men_men_n333_));
  INV        u311(.A(men_men_n195_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n335_));
  AOI220     u313(.A0(men_men_n335_), .A1(men_men_n334_), .B0(men_men_n216_), .B1(x08), .Y(men_men_n336_));
  OAI210     u314(.A0(men_men_n336_), .A1(men_men_n295_), .B0(men_men_n333_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n337_), .B(men_men_n111_), .Y(men_men_n338_));
  NA2        u316(.A(men_men_n180_), .B(men_men_n174_), .Y(men_men_n339_));
  AN2        u317(.A(men_men_n339_), .B(men_men_n187_), .Y(men_men_n340_));
  INV        u318(.A(men_men_n56_), .Y(men_men_n341_));
  OAI220     u319(.A0(men_men_n286_), .A1(men_men_n341_), .B0(men_men_n136_), .B1(men_men_n28_), .Y(men_men_n342_));
  OAI210     u320(.A0(men_men_n342_), .A1(men_men_n340_), .B0(men_men_n112_), .Y(men_men_n343_));
  NA2        u321(.A(men_men_n286_), .B(men_men_n102_), .Y(men_men_n344_));
  NA2        u322(.A(men_men_n102_), .B(men_men_n41_), .Y(men_men_n345_));
  NA3        u323(.A(men_men_n345_), .B(men_men_n344_), .C(men_men_n135_), .Y(men_men_n346_));
  NA4        u324(.A(men_men_n346_), .B(men_men_n343_), .C(men_men_n338_), .D(men_men_n48_), .Y(men_men_n347_));
  INV        u325(.A(men_men_n216_), .Y(men_men_n348_));
  NO2        u326(.A(men_men_n175_), .B(men_men_n40_), .Y(men_men_n349_));
  NA2        u327(.A(men_men_n32_), .B(x05), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n350_), .A1(men_men_n349_), .B0(men_men_n348_), .B1(men_men_n59_), .Y(men_men_n351_));
  NA2        u329(.A(men_men_n351_), .B(x02), .Y(men_men_n352_));
  INV        u330(.A(men_men_n255_), .Y(men_men_n353_));
  NA2        u331(.A(men_men_n213_), .B(x04), .Y(men_men_n354_));
  NO2        u332(.A(men_men_n354_), .B(men_men_n353_), .Y(men_men_n355_));
  NO3        u333(.A(men_men_n197_), .B(x13), .C(men_men_n31_), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n97_), .Y(men_men_n357_));
  NO3        u335(.A(men_men_n213_), .B(men_men_n173_), .C(men_men_n52_), .Y(men_men_n358_));
  OAI210     u336(.A0(men_men_n156_), .A1(men_men_n36_), .B0(men_men_n102_), .Y(men_men_n359_));
  OAI210     u337(.A0(men_men_n359_), .A1(men_men_n205_), .B0(men_men_n358_), .Y(men_men_n360_));
  NA4        u338(.A(men_men_n360_), .B(men_men_n357_), .C(men_men_n352_), .D(x06), .Y(men_men_n361_));
  NA2        u339(.A(x09), .B(x03), .Y(men_men_n362_));
  OAI220     u340(.A0(men_men_n362_), .A1(men_men_n134_), .B0(men_men_n222_), .B1(men_men_n63_), .Y(men_men_n363_));
  OAI220     u341(.A0(men_men_n174_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n364_));
  NO3        u342(.A(men_men_n295_), .B(men_men_n133_), .C(x08), .Y(men_men_n365_));
  AOI210     u343(.A0(men_men_n364_), .A1(men_men_n240_), .B0(men_men_n365_), .Y(men_men_n366_));
  NO2        u344(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n367_));
  NA2        u345(.A(men_men_n358_), .B(men_men_n367_), .Y(men_men_n368_));
  OAI210     u346(.A0(men_men_n366_), .A1(men_men_n28_), .B0(men_men_n368_), .Y(men_men_n369_));
  AO220      u347(.A0(men_men_n369_), .A1(x04), .B0(men_men_n363_), .B1(x05), .Y(men_men_n370_));
  AOI210     u348(.A0(men_men_n361_), .A1(men_men_n347_), .B0(men_men_n370_), .Y(men_men_n371_));
  OAI210     u349(.A0(men_men_n332_), .A1(x12), .B0(men_men_n371_), .Y(men03));
  OR2        u350(.A(men_men_n42_), .B(men_men_n241_), .Y(men_men_n373_));
  AOI210     u351(.A0(men_men_n162_), .A1(men_men_n102_), .B0(men_men_n373_), .Y(men_men_n374_));
  AO210      u352(.A0(men_men_n353_), .A1(men_men_n87_), .B0(men_men_n354_), .Y(men_men_n375_));
  NA2        u353(.A(men_men_n213_), .B(men_men_n161_), .Y(men_men_n376_));
  NA3        u354(.A(men_men_n376_), .B(men_men_n375_), .C(men_men_n217_), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n377_), .A1(men_men_n374_), .B0(x05), .Y(men_men_n378_));
  NA2        u356(.A(men_men_n373_), .B(x05), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n145_), .A1(men_men_n228_), .B0(men_men_n379_), .Y(men_men_n380_));
  AOI210     u358(.A0(men_men_n243_), .A1(men_men_n81_), .B0(men_men_n128_), .Y(men_men_n381_));
  OAI220     u359(.A0(men_men_n381_), .A1(men_men_n59_), .B0(men_men_n322_), .B1(men_men_n313_), .Y(men_men_n382_));
  OAI210     u360(.A0(men_men_n382_), .A1(men_men_n380_), .B0(men_men_n102_), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n154_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n384_));
  NO2        u362(.A(men_men_n184_), .B(men_men_n140_), .Y(men_men_n385_));
  OAI220     u363(.A0(men_men_n385_), .A1(men_men_n37_), .B0(men_men_n157_), .B1(x13), .Y(men_men_n386_));
  OAI210     u364(.A0(men_men_n386_), .A1(men_men_n384_), .B0(x04), .Y(men_men_n387_));
  NO3        u365(.A(men_men_n345_), .B(men_men_n86_), .C(men_men_n59_), .Y(men_men_n388_));
  AOI210     u366(.A0(men_men_n201_), .A1(men_men_n102_), .B0(men_men_n154_), .Y(men_men_n389_));
  OA210      u367(.A0(men_men_n175_), .A1(x12), .B0(men_men_n140_), .Y(men_men_n390_));
  NO3        u368(.A(men_men_n390_), .B(men_men_n389_), .C(men_men_n388_), .Y(men_men_n391_));
  NA4        u369(.A(men_men_n391_), .B(men_men_n387_), .C(men_men_n383_), .D(men_men_n378_), .Y(men04));
  NO2        u370(.A(men_men_n90_), .B(men_men_n39_), .Y(men_men_n393_));
  XO2        u371(.A(men_men_n393_), .B(men_men_n263_), .Y(men05));
  AOI210     u372(.A0(men_men_n72_), .A1(men_men_n52_), .B0(men_men_n225_), .Y(men_men_n395_));
  AOI210     u373(.A0(men_men_n395_), .A1(men_men_n321_), .B0(men_men_n25_), .Y(men_men_n396_));
  NAi41      u374(.An(men_men_n78_), .B(men_men_n151_), .C(men_men_n136_), .D(men_men_n31_), .Y(men_men_n397_));
  AOI210     u375(.A0(men_men_n467_), .A1(men_men_n397_), .B0(men_men_n24_), .Y(men_men_n398_));
  OAI210     u376(.A0(men_men_n398_), .A1(men_men_n396_), .B0(men_men_n102_), .Y(men_men_n399_));
  NA2        u377(.A(x11), .B(men_men_n31_), .Y(men_men_n400_));
  NA2        u378(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n268_), .B(x03), .Y(men_men_n402_));
  OAI220     u380(.A0(men_men_n402_), .A1(men_men_n401_), .B0(men_men_n400_), .B1(men_men_n82_), .Y(men_men_n403_));
  OAI210     u381(.A0(men_men_n26_), .A1(men_men_n102_), .B0(x07), .Y(men_men_n404_));
  AOI210     u382(.A0(men_men_n403_), .A1(x06), .B0(men_men_n404_), .Y(men_men_n405_));
  AOI220     u383(.A0(men_men_n82_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n406_));
  NO3        u384(.A(men_men_n406_), .B(men_men_n23_), .C(x00), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n402_), .B(men_men_n270_), .Y(men_men_n408_));
  OR2        u386(.A(men_men_n408_), .B(men_men_n254_), .Y(men_men_n409_));
  NO2        u387(.A(men_men_n23_), .B(x10), .Y(men_men_n410_));
  OAI210     u388(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n411_));
  OR3        u389(.A(men_men_n411_), .B(men_men_n410_), .C(men_men_n44_), .Y(men_men_n412_));
  NA2        u390(.A(men_men_n412_), .B(men_men_n409_), .Y(men_men_n413_));
  OAI210     u391(.A0(men_men_n413_), .A1(men_men_n407_), .B0(men_men_n102_), .Y(men_men_n414_));
  NA2        u392(.A(men_men_n33_), .B(men_men_n102_), .Y(men_men_n415_));
  AOI210     u393(.A0(men_men_n415_), .A1(men_men_n93_), .B0(x07), .Y(men_men_n416_));
  AOI220     u394(.A0(men_men_n416_), .A1(men_men_n414_), .B0(men_men_n405_), .B1(men_men_n399_), .Y(men_men_n417_));
  NA3        u395(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n418_));
  AO210      u396(.A0(men_men_n418_), .A1(men_men_n280_), .B0(men_men_n277_), .Y(men_men_n419_));
  AOI210     u397(.A0(men_men_n410_), .A1(men_men_n75_), .B0(men_men_n150_), .Y(men_men_n420_));
  OR2        u398(.A(men_men_n420_), .B(x03), .Y(men_men_n421_));
  NA2        u399(.A(men_men_n367_), .B(men_men_n61_), .Y(men_men_n422_));
  NO2        u400(.A(men_men_n422_), .B(x11), .Y(men_men_n423_));
  NO3        u401(.A(men_men_n423_), .B(men_men_n153_), .C(men_men_n28_), .Y(men_men_n424_));
  AOI220     u402(.A0(men_men_n424_), .A1(men_men_n421_), .B0(men_men_n419_), .B1(men_men_n47_), .Y(men_men_n425_));
  NO4        u403(.A(men_men_n345_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n426_));
  OAI210     u404(.A0(men_men_n426_), .A1(men_men_n425_), .B0(men_men_n103_), .Y(men_men_n427_));
  AOI210     u405(.A0(men_men_n354_), .A1(men_men_n114_), .B0(men_men_n276_), .Y(men_men_n428_));
  NOi21      u406(.An(men_men_n333_), .B(men_men_n140_), .Y(men_men_n429_));
  NO2        u407(.A(men_men_n429_), .B(men_men_n277_), .Y(men_men_n430_));
  OAI210     u408(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n263_), .A1(men_men_n47_), .B0(men_men_n431_), .Y(men_men_n432_));
  NO4        u410(.A(men_men_n432_), .B(men_men_n430_), .C(men_men_n428_), .D(x08), .Y(men_men_n433_));
  NA2        u411(.A(x09), .B(men_men_n41_), .Y(men_men_n434_));
  OAI220     u412(.A0(men_men_n434_), .A1(x10), .B0(men_men_n400_), .B1(men_men_n66_), .Y(men_men_n435_));
  NO2        u413(.A(x13), .B(x12), .Y(men_men_n436_));
  NO2        u414(.A(men_men_n136_), .B(men_men_n28_), .Y(men_men_n437_));
  NO2        u415(.A(men_men_n437_), .B(men_men_n281_), .Y(men_men_n438_));
  OR3        u416(.A(men_men_n438_), .B(x12), .C(x03), .Y(men_men_n439_));
  NA3        u417(.A(men_men_n348_), .B(men_men_n130_), .C(x12), .Y(men_men_n440_));
  AO210      u418(.A0(men_men_n348_), .A1(men_men_n130_), .B0(men_men_n263_), .Y(men_men_n441_));
  NA4        u419(.A(men_men_n441_), .B(men_men_n440_), .C(men_men_n439_), .D(x08), .Y(men_men_n442_));
  AOI210     u420(.A0(men_men_n436_), .A1(men_men_n435_), .B0(men_men_n442_), .Y(men_men_n443_));
  AOI210     u421(.A0(men_men_n433_), .A1(men_men_n427_), .B0(men_men_n443_), .Y(men_men_n444_));
  OAI210     u422(.A0(men_men_n422_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n445_));
  NA2        u423(.A(men_men_n306_), .B(x07), .Y(men_men_n446_));
  OAI220     u424(.A0(men_men_n446_), .A1(men_men_n401_), .B0(men_men_n153_), .B1(men_men_n43_), .Y(men_men_n447_));
  OAI210     u425(.A0(men_men_n447_), .A1(men_men_n445_), .B0(men_men_n200_), .Y(men_men_n448_));
  NA3        u426(.A(men_men_n438_), .B(men_men_n429_), .C(men_men_n344_), .Y(men_men_n449_));
  INV        u427(.A(x14), .Y(men_men_n450_));
  NO3        u428(.A(men_men_n333_), .B(men_men_n109_), .C(x11), .Y(men_men_n451_));
  NO3        u429(.A(men_men_n174_), .B(men_men_n75_), .C(men_men_n57_), .Y(men_men_n452_));
  NO3        u430(.A(men_men_n418_), .B(men_men_n345_), .C(men_men_n195_), .Y(men_men_n453_));
  NO4        u431(.A(men_men_n453_), .B(men_men_n452_), .C(men_men_n451_), .D(men_men_n450_), .Y(men_men_n454_));
  NA3        u432(.A(men_men_n454_), .B(men_men_n449_), .C(men_men_n448_), .Y(men_men_n455_));
  AOI220     u433(.A0(men_men_n415_), .A1(men_men_n61_), .B0(men_men_n437_), .B1(men_men_n173_), .Y(men_men_n456_));
  NOi21      u434(.An(men_men_n286_), .B(men_men_n157_), .Y(men_men_n457_));
  NO3        u435(.A(men_men_n133_), .B(men_men_n24_), .C(x06), .Y(men_men_n458_));
  AOI210     u436(.A0(men_men_n293_), .A1(men_men_n246_), .B0(men_men_n458_), .Y(men_men_n459_));
  OAI210     u437(.A0(men_men_n44_), .A1(x04), .B0(men_men_n459_), .Y(men_men_n460_));
  OAI210     u438(.A0(men_men_n460_), .A1(men_men_n457_), .B0(men_men_n102_), .Y(men_men_n461_));
  OAI210     u439(.A0(men_men_n456_), .A1(men_men_n92_), .B0(men_men_n461_), .Y(men_men_n462_));
  NO4        u440(.A(men_men_n462_), .B(men_men_n455_), .C(men_men_n444_), .D(men_men_n417_), .Y(men06));
  INV        u441(.A(x07), .Y(men_men_n466_));
  INV        u442(.A(men_men_n91_), .Y(men_men_n467_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule