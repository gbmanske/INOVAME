// Benchmark "top" written by ABC on Thu Jun 20 14:00:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n42_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n120_, new_new_n121_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n355_, new_new_n356_, new_new_n357_,
    new_new_n358_, new_new_n359_, new_new_n360_, new_new_n361_,
    new_new_n362_, new_new_n363_, new_new_n364_, new_new_n365_,
    new_new_n366_, new_new_n367_, new_new_n368_, new_new_n369_,
    new_new_n370_, new_new_n371_, new_new_n372_, new_new_n373_,
    new_new_n374_, new_new_n375_, new_new_n376_, new_new_n377_,
    new_new_n378_, new_new_n379_, new_new_n380_, new_new_n381_,
    new_new_n382_, new_new_n383_, new_new_n384_, new_new_n385_,
    new_new_n386_, new_new_n387_, new_new_n388_, new_new_n389_,
    new_new_n390_, new_new_n391_, new_new_n392_, new_new_n393_,
    new_new_n394_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n472_, new_new_n473_, new_new_n474_,
    new_new_n475_, new_new_n476_, new_new_n477_, new_new_n478_,
    new_new_n479_, new_new_n480_, new_new_n481_, new_new_n482_,
    new_new_n483_, new_new_n484_, new_new_n485_, new_new_n486_,
    new_new_n487_, new_new_n488_, new_new_n489_, new_new_n490_,
    new_new_n491_, new_new_n492_, new_new_n493_, new_new_n494_,
    new_new_n495_, new_new_n496_, new_new_n497_, new_new_n498_,
    new_new_n499_, new_new_n500_, new_new_n501_, new_new_n502_,
    new_new_n503_, new_new_n504_, new_new_n505_, new_new_n507_,
    new_new_n508_, new_new_n509_, new_new_n510_, new_new_n511_,
    new_new_n512_, new_new_n513_, new_new_n514_, new_new_n515_,
    new_new_n516_, new_new_n517_, new_new_n518_, new_new_n519_,
    new_new_n520_, new_new_n521_, new_new_n522_, new_new_n523_,
    new_new_n524_, new_new_n525_, new_new_n526_, new_new_n527_,
    new_new_n528_, new_new_n529_, new_new_n530_, new_new_n531_,
    new_new_n532_, new_new_n533_, new_new_n534_, new_new_n535_,
    new_new_n536_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n656_, new_new_n657_, new_new_n658_, new_new_n659_,
    new_new_n660_, new_new_n661_, new_new_n662_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NOi21      g015(.An(i_12_), .B(i_13_), .Y(new_new_n38_));
  INV        g016(.A(new_new_n38_), .Y(new_new_n39_));
  NAi31      g017(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n35_), .Y(ori1));
  INV        g019(.A(i_11_), .Y(new_new_n42_));
  NO2        g020(.A(new_new_n42_), .B(i_6_), .Y(new_new_n43_));
  INV        g021(.A(i_2_), .Y(new_new_n44_));
  NA2        g022(.A(i_0_), .B(i_3_), .Y(new_new_n45_));
  INV        g023(.A(i_5_), .Y(new_new_n46_));
  NO2        g024(.A(i_7_), .B(i_10_), .Y(new_new_n47_));
  AOI210     g025(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n47_), .Y(new_new_n48_));
  NO2        g026(.A(i_5_), .B(new_new_n44_), .Y(new_new_n49_));
  NA2        g027(.A(i_0_), .B(i_2_), .Y(new_new_n50_));
  NA2        g028(.A(i_7_), .B(i_9_), .Y(new_new_n51_));
  NO2        g029(.A(new_new_n51_), .B(new_new_n50_), .Y(new_new_n52_));
  NA2        g030(.A(new_new_n49_), .B(new_new_n43_), .Y(new_new_n53_));
  NA3        g031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  OAI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n59_), .B(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi31      g042(.An(new_new_n64_), .B(new_new_n62_), .C(new_new_n58_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n48_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  INV        g055(.A(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(new_new_n78_), .B(new_new_n55_), .Y(new_new_n79_));
  INV        g057(.A(i_3_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n80_), .B(new_new_n60_), .Y(new_new_n82_));
  INV        g060(.A(i_6_), .Y(new_new_n83_));
  NO2        g061(.A(i_2_), .B(i_7_), .Y(new_new_n84_));
  NO2        g062(.A(new_new_n82_), .B(new_new_n79_), .Y(new_new_n85_));
  NAi21      g063(.An(i_6_), .B(i_10_), .Y(new_new_n86_));
  NA2        g064(.A(i_6_), .B(i_9_), .Y(new_new_n87_));
  NA2        g065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n87_), .A1(new_new_n85_), .B0(new_new_n77_), .Y(new_new_n89_));
  AN3        g067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  NA2        g069(.A(new_new_n90_), .B(new_new_n32_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n44_), .B(new_new_n93_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n83_), .Y(new_new_n96_));
  NAi21      g074(.An(i_7_), .B(i_11_), .Y(new_new_n97_));
  NO3        g075(.A(new_new_n97_), .B(new_new_n86_), .C(new_new_n50_), .Y(new_new_n98_));
  AN2        g076(.A(i_2_), .B(i_10_), .Y(new_new_n99_));
  NA2        g077(.A(i_12_), .B(i_7_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n60_), .B(new_new_n26_), .Y(new_new_n101_));
  NA2        g079(.A(new_new_n101_), .B(i_0_), .Y(new_new_n102_));
  NA2        g080(.A(i_11_), .B(i_12_), .Y(new_new_n103_));
  OAI210     g081(.A0(new_new_n102_), .A1(new_new_n100_), .B0(new_new_n103_), .Y(new_new_n104_));
  INV        g082(.A(new_new_n104_), .Y(new_new_n105_));
  NAi31      g083(.An(new_new_n98_), .B(new_new_n105_), .C(new_new_n92_), .Y(new_new_n106_));
  NA2        g084(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n107_));
  NA2        g085(.A(i_7_), .B(new_new_n25_), .Y(new_new_n108_));
  NA2        g086(.A(new_new_n108_), .B(new_new_n107_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n109_), .B(new_new_n44_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n87_), .B(new_new_n86_), .Y(new_new_n111_));
  NAi21      g089(.An(i_3_), .B(i_8_), .Y(new_new_n112_));
  NO2        g090(.A(i_1_), .B(new_new_n83_), .Y(new_new_n113_));
  NO2        g091(.A(i_6_), .B(i_5_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(i_3_), .Y(new_new_n115_));
  AO210      g093(.A0(new_new_n115_), .A1(new_new_n45_), .B0(new_new_n113_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n116_), .B(new_new_n97_), .Y(new_new_n117_));
  NO3        g095(.A(new_new_n117_), .B(new_new_n106_), .C(new_new_n89_), .Y(new_new_n118_));
  NA3        g096(.A(new_new_n118_), .B(new_new_n76_), .C(new_new_n53_), .Y(ori2));
  NO2        g097(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n657_), .B(new_new_n120_), .Y(new_new_n121_));
  NA4        g099(.A(new_new_n121_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(ori0));
  NO2        g100(.A(i_12_), .B(i_13_), .Y(new_new_n123_));
  NAi21      g101(.An(i_5_), .B(i_11_), .Y(new_new_n124_));
  NOi21      g102(.An(new_new_n123_), .B(new_new_n124_), .Y(new_new_n125_));
  NO2        g103(.A(i_0_), .B(i_1_), .Y(new_new_n126_));
  NA2        g104(.A(i_1_), .B(i_5_), .Y(new_new_n127_));
  OR2        g105(.A(i_0_), .B(i_1_), .Y(new_new_n128_));
  NAi32      g106(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n129_));
  NOi21      g107(.An(i_4_), .B(i_10_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n38_), .Y(new_new_n131_));
  NOi21      g109(.An(i_4_), .B(i_9_), .Y(new_new_n132_));
  NOi21      g110(.An(i_11_), .B(i_13_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n132_), .Y(new_new_n134_));
  NO2        g112(.A(i_4_), .B(i_5_), .Y(new_new_n135_));
  NAi21      g113(.An(i_12_), .B(i_11_), .Y(new_new_n136_));
  NO2        g114(.A(new_new_n136_), .B(i_13_), .Y(new_new_n137_));
  NO2        g115(.A(new_new_n70_), .B(i_5_), .Y(new_new_n138_));
  NO2        g116(.A(i_13_), .B(i_10_), .Y(new_new_n139_));
  NO2        g117(.A(i_2_), .B(i_1_), .Y(new_new_n140_));
  NAi21      g118(.An(i_4_), .B(i_12_), .Y(new_new_n141_));
  INV        g119(.A(i_8_), .Y(new_new_n142_));
  NO3        g120(.A(i_3_), .B(new_new_n83_), .C(new_new_n46_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(i_7_), .Y(new_new_n144_));
  NO3        g122(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n145_));
  NO2        g123(.A(i_3_), .B(i_8_), .Y(new_new_n146_));
  NO3        g124(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n147_));
  NA3        g125(.A(new_new_n147_), .B(new_new_n146_), .C(new_new_n38_), .Y(new_new_n148_));
  NO2        g126(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n149_));
  INV        g127(.A(new_new_n149_), .Y(new_new_n150_));
  NO2        g128(.A(i_13_), .B(i_9_), .Y(new_new_n151_));
  NAi21      g129(.An(i_12_), .B(i_3_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n42_), .B(i_5_), .Y(new_new_n153_));
  NO2        g131(.A(new_new_n150_), .B(new_new_n148_), .Y(new_new_n154_));
  INV        g132(.A(new_new_n154_), .Y(new_new_n155_));
  NO2        g133(.A(new_new_n155_), .B(i_4_), .Y(new_new_n156_));
  NA3        g134(.A(i_13_), .B(new_new_n142_), .C(i_10_), .Y(new_new_n157_));
  NA2        g135(.A(i_0_), .B(i_5_), .Y(new_new_n158_));
  NAi31      g136(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n36_), .B(i_13_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n161_));
  NO2        g139(.A(new_new_n44_), .B(new_new_n60_), .Y(new_new_n162_));
  INV        g140(.A(i_13_), .Y(new_new_n163_));
  NO2        g141(.A(i_12_), .B(new_new_n163_), .Y(new_new_n164_));
  NO2        g142(.A(i_12_), .B(new_new_n37_), .Y(new_new_n165_));
  OR2        g143(.A(i_8_), .B(i_7_), .Y(new_new_n166_));
  INV        g144(.A(i_12_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n42_), .B(new_new_n167_), .Y(new_new_n168_));
  NO3        g146(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n169_));
  NA2        g147(.A(i_2_), .B(i_1_), .Y(new_new_n170_));
  NO3        g148(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n171_));
  NAi21      g149(.An(i_4_), .B(i_3_), .Y(new_new_n172_));
  NO2        g150(.A(i_0_), .B(i_6_), .Y(new_new_n173_));
  NOi41      g151(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  NO2        g153(.A(i_11_), .B(new_new_n163_), .Y(new_new_n176_));
  NOi21      g154(.An(i_1_), .B(i_6_), .Y(new_new_n177_));
  NAi21      g155(.An(i_3_), .B(i_7_), .Y(new_new_n178_));
  NA2        g156(.A(new_new_n167_), .B(i_9_), .Y(new_new_n179_));
  OR4        g157(.A(new_new_n179_), .B(new_new_n178_), .C(new_new_n177_), .D(new_new_n138_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n70_), .B(i_5_), .Y(new_new_n181_));
  NA2        g159(.A(i_3_), .B(i_9_), .Y(new_new_n182_));
  NAi21      g160(.An(i_7_), .B(i_10_), .Y(new_new_n183_));
  NO2        g161(.A(new_new_n183_), .B(new_new_n182_), .Y(new_new_n184_));
  NA3        g162(.A(new_new_n184_), .B(new_new_n181_), .C(new_new_n61_), .Y(new_new_n185_));
  NA2        g163(.A(new_new_n185_), .B(new_new_n180_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n186_), .B(new_new_n176_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n166_), .B(new_new_n37_), .Y(new_new_n188_));
  NA2        g166(.A(i_12_), .B(i_6_), .Y(new_new_n189_));
  OR2        g167(.A(i_13_), .B(i_9_), .Y(new_new_n190_));
  NO2        g168(.A(new_new_n190_), .B(new_new_n46_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n172_), .B(i_2_), .Y(new_new_n192_));
  NA3        g170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n42_), .Y(new_new_n193_));
  NA2        g171(.A(new_new_n176_), .B(i_9_), .Y(new_new_n194_));
  OAI210     g172(.A0(new_new_n70_), .A1(new_new_n194_), .B0(new_new_n193_), .Y(new_new_n195_));
  NO3        g173(.A(i_11_), .B(new_new_n163_), .C(new_new_n25_), .Y(new_new_n196_));
  NA2        g174(.A(new_new_n195_), .B(new_new_n188_), .Y(new_new_n197_));
  NA2        g175(.A(new_new_n197_), .B(new_new_n187_), .Y(new_new_n198_));
  NO3        g176(.A(i_12_), .B(new_new_n163_), .C(new_new_n37_), .Y(new_new_n199_));
  AN2        g177(.A(i_3_), .B(i_10_), .Y(new_new_n200_));
  NO2        g178(.A(i_5_), .B(new_new_n37_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n44_), .B(new_new_n26_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n198_), .B(new_new_n156_), .Y(new_new_n203_));
  NO3        g181(.A(new_new_n42_), .B(i_13_), .C(i_9_), .Y(new_new_n204_));
  NO2        g182(.A(i_2_), .B(i_3_), .Y(new_new_n205_));
  NO2        g183(.A(i_12_), .B(i_10_), .Y(new_new_n206_));
  NOi21      g184(.An(i_5_), .B(i_0_), .Y(new_new_n207_));
  NA4        g185(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n208_));
  INV        g186(.A(i_6_), .Y(new_new_n209_));
  NO2        g187(.A(i_1_), .B(i_7_), .Y(new_new_n210_));
  NOi21      g188(.An(new_new_n127_), .B(new_new_n96_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(new_new_n108_), .Y(new_new_n212_));
  NA2        g190(.A(new_new_n212_), .B(i_3_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n142_), .B(i_9_), .Y(new_new_n214_));
  NA2        g192(.A(new_new_n214_), .B(new_new_n149_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n215_), .B(new_new_n44_), .Y(new_new_n216_));
  INV        g194(.A(new_new_n216_), .Y(new_new_n217_));
  AOI210     g195(.A0(new_new_n217_), .A1(new_new_n213_), .B0(new_new_n131_), .Y(new_new_n218_));
  INV        g196(.A(new_new_n218_), .Y(new_new_n219_));
  NOi32      g197(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n220_));
  INV        g198(.A(new_new_n220_), .Y(new_new_n221_));
  NAi21      g199(.An(i_0_), .B(i_6_), .Y(new_new_n222_));
  NAi21      g200(.An(i_1_), .B(i_5_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n224_), .B(new_new_n25_), .Y(new_new_n225_));
  OAI210     g203(.A0(new_new_n225_), .A1(new_new_n129_), .B0(new_new_n175_), .Y(new_new_n226_));
  NAi41      g204(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n227_));
  OAI220     g205(.A0(new_new_n227_), .A1(new_new_n223_), .B0(new_new_n159_), .B1(new_new_n129_), .Y(new_new_n228_));
  NOi32      g206(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n229_));
  NAi21      g207(.An(i_6_), .B(i_1_), .Y(new_new_n230_));
  NA3        g208(.A(new_new_n230_), .B(new_new_n229_), .C(new_new_n44_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n231_), .B(i_0_), .Y(new_new_n232_));
  OR2        g210(.A(new_new_n232_), .B(new_new_n228_), .Y(new_new_n233_));
  NO2        g211(.A(i_1_), .B(new_new_n93_), .Y(new_new_n234_));
  NAi21      g212(.An(i_3_), .B(i_4_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n235_), .B(i_9_), .Y(new_new_n236_));
  AN2        g214(.A(i_6_), .B(i_7_), .Y(new_new_n237_));
  OAI210     g215(.A0(new_new_n237_), .A1(new_new_n234_), .B0(new_new_n236_), .Y(new_new_n238_));
  NA2        g216(.A(i_2_), .B(i_7_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n233_), .B(new_new_n226_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n240_), .B(new_new_n221_), .Y(new_new_n241_));
  AN2        g219(.A(i_12_), .B(i_5_), .Y(new_new_n242_));
  INV        g220(.A(new_new_n242_), .Y(new_new_n243_));
  NO2        g221(.A(i_11_), .B(i_6_), .Y(new_new_n244_));
  NO2        g222(.A(i_5_), .B(i_10_), .Y(new_new_n245_));
  NO2        g223(.A(i_11_), .B(i_12_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n246_), .B(new_new_n36_), .Y(new_new_n247_));
  NO2        g225(.A(i_3_), .B(new_new_n247_), .Y(new_new_n248_));
  NAi21      g226(.An(i_13_), .B(i_0_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n249_), .B(new_new_n170_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n248_), .B(new_new_n250_), .Y(new_new_n251_));
  INV        g229(.A(new_new_n251_), .Y(new_new_n252_));
  NO2        g230(.A(i_0_), .B(i_11_), .Y(new_new_n253_));
  AN2        g231(.A(i_1_), .B(i_6_), .Y(new_new_n254_));
  NOi21      g232(.An(i_2_), .B(i_12_), .Y(new_new_n255_));
  NAi21      g233(.An(i_9_), .B(i_4_), .Y(new_new_n256_));
  OR2        g234(.A(i_13_), .B(i_10_), .Y(new_new_n257_));
  NO3        g235(.A(new_new_n257_), .B(new_new_n103_), .C(new_new_n256_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n134_), .B(new_new_n107_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n260_));
  NA2        g238(.A(new_new_n199_), .B(new_new_n260_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n261_), .B(new_new_n211_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n142_), .B(i_10_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n181_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n264_), .B(new_new_n263_), .Y(new_new_n265_));
  INV        g243(.A(new_new_n265_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n266_), .B(new_new_n194_), .Y(new_new_n267_));
  NO4        g245(.A(new_new_n267_), .B(new_new_n262_), .C(new_new_n252_), .D(new_new_n241_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n70_), .B(i_13_), .Y(new_new_n269_));
  NO2        g247(.A(i_10_), .B(i_9_), .Y(new_new_n270_));
  NAi21      g248(.An(i_12_), .B(i_8_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n271_), .B(i_3_), .Y(new_new_n272_));
  NA2        g250(.A(new_new_n202_), .B(i_0_), .Y(new_new_n273_));
  NO3        g251(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n189_), .B(new_new_n91_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n275_), .B(new_new_n274_), .Y(new_new_n276_));
  NA2        g254(.A(i_8_), .B(i_9_), .Y(new_new_n277_));
  NO2        g255(.A(i_7_), .B(i_2_), .Y(new_new_n278_));
  OR2        g256(.A(new_new_n278_), .B(new_new_n277_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n199_), .B(new_new_n149_), .Y(new_new_n280_));
  OAI220     g258(.A0(new_new_n280_), .A1(new_new_n279_), .B0(new_new_n276_), .B1(new_new_n273_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n176_), .B(new_new_n201_), .Y(new_new_n282_));
  NO3        g260(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n283_));
  INV        g261(.A(new_new_n283_), .Y(new_new_n284_));
  NA3        g262(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n285_));
  NA4        g263(.A(new_new_n124_), .B(new_new_n101_), .C(new_new_n77_), .D(new_new_n23_), .Y(new_new_n286_));
  OAI220     g264(.A0(new_new_n286_), .A1(new_new_n285_), .B0(new_new_n284_), .B1(new_new_n282_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(new_new_n281_), .Y(new_new_n288_));
  OR2        g266(.A(new_new_n215_), .B(new_new_n93_), .Y(new_new_n289_));
  OR2        g267(.A(new_new_n289_), .B(new_new_n131_), .Y(new_new_n290_));
  NO2        g268(.A(i_2_), .B(i_13_), .Y(new_new_n291_));
  NO3        g269(.A(i_4_), .B(new_new_n46_), .C(i_8_), .Y(new_new_n292_));
  NO2        g270(.A(i_6_), .B(i_7_), .Y(new_new_n293_));
  NO2        g271(.A(i_11_), .B(i_1_), .Y(new_new_n294_));
  NOi21      g272(.An(i_2_), .B(i_7_), .Y(new_new_n295_));
  NO2        g273(.A(i_3_), .B(new_new_n142_), .Y(new_new_n296_));
  NO2        g274(.A(i_6_), .B(i_10_), .Y(new_new_n297_));
  NA3        g275(.A(new_new_n174_), .B(new_new_n133_), .C(new_new_n114_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n44_), .B(new_new_n42_), .Y(new_new_n299_));
  NA2        g277(.A(new_new_n283_), .B(new_new_n245_), .Y(new_new_n300_));
  NAi21      g278(.An(new_new_n157_), .B(new_new_n246_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n210_), .B(new_new_n158_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n302_), .B(new_new_n301_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n204_), .B(new_new_n169_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n304_), .B(new_new_n264_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n305_), .B(new_new_n303_), .Y(new_new_n306_));
  NA4        g284(.A(new_new_n306_), .B(new_new_n298_), .C(new_new_n290_), .D(new_new_n288_), .Y(new_new_n307_));
  NA2        g285(.A(new_new_n242_), .B(new_new_n163_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n237_), .B(new_new_n229_), .Y(new_new_n309_));
  OR2        g287(.A(new_new_n308_), .B(new_new_n309_), .Y(new_new_n310_));
  INV        g288(.A(new_new_n258_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n311_), .B(new_new_n310_), .Y(new_new_n312_));
  INV        g290(.A(new_new_n312_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n181_), .B(new_new_n61_), .Y(new_new_n314_));
  OAI210     g292(.A0(i_8_), .A1(new_new_n314_), .B0(new_new_n116_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n315_), .B(new_new_n259_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n313_), .Y(new_new_n317_));
  NO2        g295(.A(i_12_), .B(new_new_n142_), .Y(new_new_n318_));
  NA3        g296(.A(new_new_n200_), .B(new_new_n135_), .C(new_new_n90_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n128_), .B(i_5_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n658_), .B(new_new_n283_), .Y(new_new_n321_));
  INV        g299(.A(new_new_n321_), .Y(new_new_n322_));
  NA3        g300(.A(new_new_n158_), .B(new_new_n68_), .C(new_new_n42_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n199_), .B(new_new_n81_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n323_), .B(new_new_n324_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n270_), .B(new_new_n160_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n326_), .B(new_new_n327_), .Y(new_new_n328_));
  AOI210     g306(.A0(new_new_n230_), .A1(new_new_n44_), .B0(new_new_n234_), .Y(new_new_n329_));
  NA2        g307(.A(i_0_), .B(new_new_n46_), .Y(new_new_n330_));
  NA3        g308(.A(new_new_n318_), .B(new_new_n196_), .C(new_new_n330_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n329_), .B(new_new_n331_), .Y(new_new_n332_));
  NO3        g310(.A(new_new_n332_), .B(new_new_n328_), .C(new_new_n325_), .Y(new_new_n333_));
  NO4        g311(.A(new_new_n177_), .B(new_new_n40_), .C(i_2_), .D(new_new_n46_), .Y(new_new_n334_));
  NOi21      g312(.An(i_10_), .B(i_6_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n336_));
  AOI220     g314(.A0(new_new_n199_), .A1(new_new_n336_), .B0(new_new_n196_), .B1(new_new_n335_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n337_), .B(new_new_n273_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n100_), .B(new_new_n23_), .Y(new_new_n339_));
  NOi31      g317(.An(new_new_n125_), .B(i_10_), .C(new_new_n208_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n340_), .B(new_new_n338_), .Y(new_new_n341_));
  INV        g319(.A(new_new_n205_), .Y(new_new_n342_));
  NO2        g320(.A(i_12_), .B(new_new_n83_), .Y(new_new_n343_));
  NA3        g321(.A(new_new_n343_), .B(new_new_n196_), .C(new_new_n330_), .Y(new_new_n344_));
  NA3        g322(.A(new_new_n244_), .B(new_new_n199_), .C(new_new_n158_), .Y(new_new_n345_));
  AOI210     g323(.A0(new_new_n345_), .A1(new_new_n344_), .B0(new_new_n342_), .Y(new_new_n346_));
  OR2        g324(.A(i_2_), .B(i_5_), .Y(new_new_n347_));
  OR2        g325(.A(new_new_n347_), .B(new_new_n254_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n239_), .B(new_new_n173_), .Y(new_new_n349_));
  AOI210     g327(.A0(new_new_n349_), .A1(new_new_n348_), .B0(new_new_n301_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n350_), .B(new_new_n346_), .Y(new_new_n351_));
  NA3        g329(.A(new_new_n351_), .B(new_new_n341_), .C(new_new_n333_), .Y(new_new_n352_));
  NO4        g330(.A(new_new_n352_), .B(new_new_n322_), .C(new_new_n317_), .D(new_new_n307_), .Y(new_new_n353_));
  NA4        g331(.A(new_new_n353_), .B(new_new_n268_), .C(new_new_n219_), .D(new_new_n203_), .Y(ori7));
  NO2        g332(.A(new_new_n88_), .B(new_new_n51_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n97_), .B(new_new_n86_), .Y(new_new_n356_));
  INV        g334(.A(new_new_n356_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n297_), .B(new_new_n81_), .Y(new_new_n358_));
  NA2        g336(.A(i_11_), .B(new_new_n142_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n123_), .B(new_new_n359_), .Y(new_new_n360_));
  OAI210     g338(.A0(new_new_n360_), .A1(new_new_n358_), .B0(new_new_n357_), .Y(new_new_n361_));
  NA2        g339(.A(i_2_), .B(new_new_n83_), .Y(new_new_n362_));
  OAI210     g340(.A0(new_new_n84_), .A1(new_new_n146_), .B0(new_new_n147_), .Y(new_new_n363_));
  NO2        g341(.A(i_7_), .B(new_new_n37_), .Y(new_new_n364_));
  NA2        g342(.A(i_4_), .B(i_8_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n361_), .B(new_new_n355_), .Y(new_new_n366_));
  AOI210     g344(.A0(new_new_n112_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n367_));
  AOI210     g345(.A0(new_new_n367_), .A1(new_new_n167_), .B0(new_new_n130_), .Y(new_new_n368_));
  OR2        g346(.A(i_6_), .B(i_10_), .Y(new_new_n369_));
  OR3        g347(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n370_));
  INV        g348(.A(new_new_n145_), .Y(new_new_n371_));
  OR2        g349(.A(new_new_n368_), .B(new_new_n190_), .Y(new_new_n372_));
  AOI210     g350(.A0(new_new_n372_), .A1(new_new_n366_), .B0(new_new_n60_), .Y(new_new_n373_));
  NOi21      g351(.An(i_11_), .B(i_7_), .Y(new_new_n374_));
  AO210      g352(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n375_), .B(new_new_n374_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n376_), .B(new_new_n151_), .Y(new_new_n377_));
  NA3        g355(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n378_));
  NAi31      g356(.An(new_new_n378_), .B(i_12_), .C(i_11_), .Y(new_new_n379_));
  AOI210     g357(.A0(new_new_n379_), .A1(new_new_n377_), .B0(new_new_n60_), .Y(new_new_n380_));
  NO3        g358(.A(new_new_n183_), .B(new_new_n152_), .C(new_new_n359_), .Y(new_new_n381_));
  OAI210     g359(.A0(new_new_n381_), .A1(new_new_n164_), .B0(new_new_n60_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n255_), .B(new_new_n31_), .Y(new_new_n383_));
  OR2        g361(.A(new_new_n152_), .B(new_new_n97_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n384_), .B(new_new_n383_), .Y(new_new_n385_));
  NO2        g363(.A(i_1_), .B(i_4_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  NO2        g365(.A(i_1_), .B(i_12_), .Y(new_new_n388_));
  NA3        g366(.A(new_new_n388_), .B(new_new_n99_), .C(new_new_n24_), .Y(new_new_n389_));
  BUFFER     g367(.A(new_new_n389_), .Y(new_new_n390_));
  NA3        g368(.A(new_new_n390_), .B(new_new_n387_), .C(new_new_n382_), .Y(new_new_n391_));
  OAI210     g369(.A0(new_new_n391_), .A1(new_new_n380_), .B0(i_6_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n378_), .B(new_new_n97_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n393_), .B(new_new_n343_), .Y(new_new_n394_));
  NO2        g372(.A(i_6_), .B(i_11_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n394_), .B(new_new_n276_), .Y(new_new_n396_));
  NO3        g374(.A(new_new_n369_), .B(new_new_n166_), .C(new_new_n23_), .Y(new_new_n397_));
  AOI210     g375(.A0(i_1_), .A1(new_new_n184_), .B0(new_new_n397_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n42_), .Y(new_new_n399_));
  NA3        g377(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n44_), .B(i_1_), .Y(new_new_n401_));
  NA3        g379(.A(new_new_n401_), .B(new_new_n189_), .C(new_new_n42_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(new_new_n400_), .Y(new_new_n403_));
  AOI210     g381(.A0(new_new_n294_), .A1(new_new_n260_), .B0(new_new_n171_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n404_), .B(new_new_n362_), .Y(new_new_n405_));
  OR2        g383(.A(new_new_n405_), .B(new_new_n403_), .Y(new_new_n406_));
  NO3        g384(.A(new_new_n406_), .B(new_new_n399_), .C(new_new_n396_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n167_), .B(new_new_n93_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n408_), .B(new_new_n374_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n409_), .B(i_1_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n410_), .B(new_new_n370_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n256_), .B(new_new_n83_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n411_), .B(new_new_n44_), .Y(new_new_n413_));
  NA2        g391(.A(i_3_), .B(new_new_n142_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n166_), .B(new_new_n42_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n202_), .C(new_new_n168_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n417_));
  INV        g395(.A(i_6_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n83_), .B(i_9_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n419_), .B(new_new_n60_), .Y(new_new_n420_));
  NO2        g398(.A(new_new_n420_), .B(new_new_n388_), .Y(new_new_n421_));
  NO4        g399(.A(new_new_n421_), .B(new_new_n418_), .C(new_new_n416_), .D(i_4_), .Y(new_new_n422_));
  NA2        g400(.A(i_1_), .B(i_3_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n277_), .B(new_new_n88_), .Y(new_new_n424_));
  INV        g402(.A(new_new_n424_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(new_new_n423_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n426_), .B(new_new_n422_), .Y(new_new_n427_));
  NA4        g405(.A(new_new_n427_), .B(new_new_n413_), .C(new_new_n407_), .D(new_new_n392_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n295_), .B(new_new_n365_), .C(new_new_n83_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n430_), .B(new_new_n25_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n431_), .B(new_new_n429_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n432_), .B(i_1_), .Y(new_new_n433_));
  INV        g411(.A(i_1_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n433_), .B(i_13_), .Y(new_new_n435_));
  NA3        g413(.A(i_7_), .B(i_12_), .C(new_new_n120_), .Y(new_new_n436_));
  AOI220     g414(.A0(new_new_n291_), .A1(new_new_n130_), .B0(i_2_), .B1(new_new_n120_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n437_), .B(new_new_n436_), .Y(new_new_n438_));
  NO2        g416(.A(new_new_n295_), .B(new_new_n24_), .Y(new_new_n439_));
  AOI220     g417(.A0(new_new_n439_), .A1(new_new_n412_), .B0(new_new_n174_), .B1(new_new_n113_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n440_), .B(new_new_n39_), .Y(new_new_n441_));
  AOI210     g419(.A0(new_new_n438_), .A1(new_new_n209_), .B0(new_new_n441_), .Y(new_new_n442_));
  INV        g420(.A(new_new_n100_), .Y(new_new_n443_));
  AOI220     g421(.A0(new_new_n443_), .A1(new_new_n69_), .B0(new_new_n244_), .B1(new_new_n401_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n444_), .B(new_new_n172_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n111_), .B(i_13_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n400_), .B(new_new_n100_), .Y(new_new_n447_));
  INV        g425(.A(new_new_n447_), .Y(new_new_n448_));
  OAI220     g426(.A0(new_new_n448_), .A1(new_new_n68_), .B0(new_new_n446_), .B1(new_new_n434_), .Y(new_new_n449_));
  NO3        g427(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n93_), .Y(new_new_n450_));
  NA2        g428(.A(new_new_n26_), .B(new_new_n142_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n660_), .B(new_new_n371_), .Y(new_new_n452_));
  NO3        g430(.A(new_new_n452_), .B(new_new_n449_), .C(new_new_n445_), .Y(new_new_n453_));
  OR2        g431(.A(i_11_), .B(i_6_), .Y(new_new_n454_));
  NA3        g432(.A(i_12_), .B(new_new_n451_), .C(i_7_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n395_), .B(i_13_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n94_), .B(new_new_n451_), .Y(new_new_n458_));
  NAi21      g436(.An(i_11_), .B(i_12_), .Y(new_new_n459_));
  NO3        g437(.A(new_new_n459_), .B(i_13_), .C(new_new_n83_), .Y(new_new_n460_));
  NO3        g438(.A(new_new_n295_), .B(new_new_n343_), .C(new_new_n365_), .Y(new_new_n461_));
  AOI220     g439(.A0(new_new_n461_), .A1(new_new_n204_), .B0(new_new_n460_), .B1(new_new_n458_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n462_), .B(new_new_n457_), .Y(new_new_n463_));
  OAI210     g441(.A0(new_new_n463_), .A1(new_new_n456_), .B0(new_new_n60_), .Y(new_new_n464_));
  NO2        g442(.A(i_2_), .B(i_12_), .Y(new_new_n465_));
  INV        g443(.A(i_2_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n466_), .B(new_new_n388_), .Y(new_new_n467_));
  INV        g445(.A(new_new_n467_), .Y(new_new_n468_));
  NA3        g446(.A(new_new_n468_), .B(new_new_n43_), .C(new_new_n163_), .Y(new_new_n469_));
  NA4        g447(.A(new_new_n469_), .B(new_new_n464_), .C(new_new_n453_), .D(new_new_n442_), .Y(new_new_n470_));
  OR4        g448(.A(new_new_n470_), .B(new_new_n435_), .C(new_new_n428_), .D(new_new_n373_), .Y(ori5));
  NA2        g449(.A(new_new_n409_), .B(new_new_n192_), .Y(new_new_n472_));
  AN2        g450(.A(new_new_n24_), .B(i_10_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n465_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n474_), .B(new_new_n472_), .Y(new_new_n475_));
  NO3        g453(.A(i_11_), .B(new_new_n167_), .C(i_13_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n108_), .B(new_new_n23_), .Y(new_new_n477_));
  INV        g455(.A(new_new_n270_), .Y(new_new_n478_));
  INV        g456(.A(new_new_n475_), .Y(new_new_n479_));
  INV        g457(.A(new_new_n133_), .Y(new_new_n480_));
  INV        g458(.A(new_new_n174_), .Y(new_new_n481_));
  NO2        g459(.A(new_new_n481_), .B(new_new_n480_), .Y(new_new_n482_));
  NO2        g460(.A(new_new_n277_), .B(new_new_n26_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n260_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n484_), .B(i_2_), .Y(new_new_n485_));
  INV        g463(.A(new_new_n485_), .Y(new_new_n486_));
  AOI210     g464(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n257_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n487_), .A1(new_new_n486_), .B0(new_new_n482_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n141_), .B(new_new_n109_), .Y(new_new_n489_));
  OAI210     g467(.A0(new_new_n489_), .A1(new_new_n477_), .B0(i_2_), .Y(new_new_n490_));
  AOI210     g468(.A0(new_new_n134_), .A1(new_new_n490_), .B0(new_new_n142_), .Y(new_new_n491_));
  OA210      g469(.A0(new_new_n376_), .A1(new_new_n110_), .B0(i_13_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n145_), .B(new_new_n146_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n493_), .B(new_new_n239_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n152_), .B(new_new_n661_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n260_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n93_), .B(new_new_n200_), .Y(new_new_n497_));
  OAI210     g475(.A0(new_new_n497_), .A1(i_11_), .B0(new_new_n496_), .Y(new_new_n498_));
  NO4        g476(.A(new_new_n498_), .B(new_new_n494_), .C(new_new_n492_), .D(new_new_n491_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n339_), .B(new_new_n28_), .Y(new_new_n500_));
  INV        g478(.A(new_new_n500_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n59_), .B(i_12_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n502_), .B(new_new_n110_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(new_new_n359_), .Y(new_new_n504_));
  AOI220     g482(.A0(new_new_n504_), .A1(new_new_n36_), .B0(new_new_n501_), .B1(new_new_n44_), .Y(new_new_n505_));
  NA4        g483(.A(new_new_n505_), .B(new_new_n499_), .C(new_new_n488_), .D(new_new_n479_), .Y(ori6));
  NA4        g484(.A(new_new_n245_), .B(new_new_n296_), .C(new_new_n68_), .D(new_new_n93_), .Y(new_new_n507_));
  INV        g485(.A(new_new_n507_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n159_), .B(new_new_n299_), .Y(new_new_n509_));
  NO2        g487(.A(i_11_), .B(i_9_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n508_), .B(new_new_n207_), .Y(new_new_n511_));
  OR2        g489(.A(new_new_n511_), .B(i_12_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n343_), .B(new_new_n60_), .Y(new_new_n513_));
  INV        g491(.A(new_new_n513_), .Y(new_new_n514_));
  INV        g492(.A(new_new_n144_), .Y(new_new_n515_));
  AOI220     g493(.A0(new_new_n515_), .A1(new_new_n510_), .B0(new_new_n514_), .B1(new_new_n70_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n177_), .B(i_9_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n517_), .B(new_new_n502_), .Y(new_new_n518_));
  AOI210     g496(.A0(new_new_n518_), .A1(new_new_n309_), .B0(new_new_n138_), .Y(new_new_n519_));
  NAi32      g497(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n454_), .B(new_new_n520_), .Y(new_new_n521_));
  OR2        g499(.A(new_new_n521_), .B(new_new_n519_), .Y(new_new_n522_));
  BUFFER     g500(.A(new_new_n272_), .Y(new_new_n523_));
  NA3        g501(.A(new_new_n523_), .B(new_new_n126_), .C(new_new_n66_), .Y(new_new_n524_));
  AO210      g502(.A0(new_new_n300_), .A1(new_new_n478_), .B0(new_new_n36_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n525_), .B(new_new_n524_), .Y(new_new_n526_));
  INV        g504(.A(new_new_n509_), .Y(new_new_n527_));
  NA3        g505(.A(new_new_n239_), .B(new_new_n169_), .C(new_new_n126_), .Y(new_new_n528_));
  NA3        g506(.A(new_new_n528_), .B(new_new_n527_), .C(new_new_n363_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n272_), .B(new_new_n270_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n369_), .B(new_new_n94_), .Y(new_new_n531_));
  OAI210     g509(.A0(new_new_n531_), .A1(new_new_n77_), .B0(new_new_n253_), .Y(new_new_n532_));
  INV        g510(.A(new_new_n348_), .Y(new_new_n533_));
  NA3        g511(.A(new_new_n533_), .B(new_new_n206_), .C(i_7_), .Y(new_new_n534_));
  NA3        g512(.A(new_new_n534_), .B(new_new_n532_), .C(new_new_n530_), .Y(new_new_n535_));
  NO4        g513(.A(new_new_n535_), .B(new_new_n529_), .C(new_new_n526_), .D(new_new_n522_), .Y(new_new_n536_));
  NA4        g514(.A(new_new_n536_), .B(new_new_n516_), .C(new_new_n512_), .D(new_new_n240_), .Y(ori3));
  NA2        g515(.A(i_12_), .B(i_10_), .Y(new_new_n538_));
  NO2        g516(.A(i_11_), .B(new_new_n167_), .Y(new_new_n539_));
  NA3        g517(.A(new_new_n528_), .B(new_new_n363_), .C(new_new_n238_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n540_), .B(new_new_n38_), .Y(new_new_n541_));
  NOi21      g519(.An(new_new_n90_), .B(new_new_n484_), .Y(new_new_n542_));
  NO3        g520(.A(new_new_n384_), .B(new_new_n277_), .C(new_new_n113_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n255_), .B(new_new_n43_), .Y(new_new_n544_));
  AN2        g522(.A(new_new_n275_), .B(new_new_n52_), .Y(new_new_n545_));
  NO3        g523(.A(new_new_n545_), .B(new_new_n543_), .C(new_new_n542_), .Y(new_new_n546_));
  AOI210     g524(.A0(new_new_n546_), .A1(new_new_n541_), .B0(new_new_n46_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n138_), .B(new_new_n335_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n548_), .B(new_new_n60_), .Y(new_new_n549_));
  NOi21      g527(.An(i_5_), .B(i_9_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n550_), .B(new_new_n269_), .Y(new_new_n551_));
  BUFFER     g529(.A(new_new_n189_), .Y(new_new_n552_));
  AOI210     g530(.A0(new_new_n552_), .A1(new_new_n294_), .B0(new_new_n430_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n553_), .B(new_new_n551_), .Y(new_new_n554_));
  NO3        g532(.A(new_new_n554_), .B(new_new_n549_), .C(new_new_n547_), .Y(new_new_n555_));
  BUFFER     g533(.A(i_0_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n138_), .B(new_new_n24_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n417_), .B(new_new_n356_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n558_), .B(new_new_n557_), .Y(new_new_n559_));
  INV        g537(.A(new_new_n559_), .Y(new_new_n560_));
  NA2        g538(.A(new_new_n336_), .B(i_0_), .Y(new_new_n561_));
  NO3        g539(.A(new_new_n561_), .B(new_new_n243_), .C(new_new_n84_), .Y(new_new_n562_));
  NO4        g540(.A(new_new_n347_), .B(i_12_), .C(new_new_n257_), .D(new_new_n254_), .Y(new_new_n563_));
  AOI210     g541(.A0(new_new_n563_), .A1(i_11_), .B0(new_new_n562_), .Y(new_new_n564_));
  NA2        g542(.A(new_new_n476_), .B(new_new_n207_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n297_), .A1(new_new_n84_), .B0(new_new_n55_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n566_), .B(new_new_n565_), .Y(new_new_n567_));
  NO2        g545(.A(new_new_n179_), .B(new_new_n127_), .Y(new_new_n568_));
  NO4        g546(.A(new_new_n100_), .B(new_new_n55_), .C(new_new_n414_), .D(i_5_), .Y(new_new_n569_));
  AO220      g547(.A0(new_new_n569_), .A1(i_10_), .B0(new_new_n568_), .B1(i_6_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n570_), .B(new_new_n567_), .Y(new_new_n571_));
  NA3        g549(.A(new_new_n571_), .B(new_new_n564_), .C(new_new_n560_), .Y(new_new_n572_));
  NA2        g550(.A(i_11_), .B(i_9_), .Y(new_new_n573_));
  NO3        g551(.A(i_12_), .B(new_new_n573_), .C(new_new_n362_), .Y(new_new_n574_));
  AN2        g552(.A(new_new_n574_), .B(i_10_), .Y(new_new_n575_));
  NO2        g553(.A(new_new_n573_), .B(new_new_n70_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n136_), .B(i_0_), .Y(new_new_n577_));
  INV        g555(.A(new_new_n575_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n133_), .B(new_new_n95_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n364_), .B(new_new_n207_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n580_), .B(new_new_n544_), .Y(new_new_n581_));
  INV        g559(.A(new_new_n581_), .Y(new_new_n582_));
  NOi21      g560(.An(i_7_), .B(i_5_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n582_), .B(new_new_n578_), .Y(new_new_n584_));
  INV        g562(.A(new_new_n538_), .Y(new_new_n585_));
  OA210      g563(.A0(new_new_n293_), .A1(new_new_n162_), .B0(new_new_n292_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n585_), .B(new_new_n576_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n576_), .B(new_new_n200_), .Y(new_new_n588_));
  INV        g566(.A(new_new_n588_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n589_), .B(new_new_n293_), .Y(new_new_n590_));
  NO3        g568(.A(new_new_n347_), .B(new_new_n222_), .C(new_new_n24_), .Y(new_new_n591_));
  AOI210     g569(.A0(new_new_n439_), .A1(new_new_n320_), .B0(new_new_n591_), .Y(new_new_n592_));
  NAi21      g570(.An(i_9_), .B(i_5_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n593_), .B(new_new_n249_), .Y(new_new_n594_));
  NA2        g572(.A(new_new_n594_), .B(new_new_n376_), .Y(new_new_n595_));
  OAI220     g573(.A0(new_new_n595_), .A1(new_new_n83_), .B0(new_new_n592_), .B1(new_new_n134_), .Y(new_new_n596_));
  NO2        g574(.A(new_new_n596_), .B(new_new_n312_), .Y(new_new_n597_));
  NA3        g575(.A(new_new_n597_), .B(new_new_n590_), .C(new_new_n587_), .Y(new_new_n598_));
  NO3        g576(.A(new_new_n598_), .B(new_new_n584_), .C(new_new_n572_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n556_), .B(new_new_n459_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n513_), .A1(new_new_n429_), .B0(new_new_n579_), .Y(new_new_n601_));
  INV        g579(.A(new_new_n601_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n173_), .B(new_new_n165_), .Y(new_new_n603_));
  AOI210     g581(.A0(new_new_n603_), .A1(new_new_n561_), .B0(new_new_n127_), .Y(new_new_n604_));
  INV        g582(.A(new_new_n604_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n605_), .B(new_new_n602_), .Y(new_new_n606_));
  NO3        g584(.A(new_new_n153_), .B(new_new_n242_), .C(i_0_), .Y(new_new_n607_));
  OAI210     g585(.A0(new_new_n607_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n608_));
  INV        g586(.A(new_new_n608_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n172_), .B(new_new_n88_), .Y(new_new_n610_));
  AOI210     g588(.A0(new_new_n610_), .A1(new_new_n600_), .B0(new_new_n98_), .Y(new_new_n611_));
  OR2        g589(.A(new_new_n611_), .B(i_5_), .Y(new_new_n612_));
  AOI210     g590(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n136_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n586_), .Y(new_new_n614_));
  NO3        g592(.A(new_new_n544_), .B(new_new_n51_), .C(new_new_n46_), .Y(new_new_n615_));
  NO3        g593(.A(new_new_n659_), .B(new_new_n615_), .C(new_new_n656_), .Y(new_new_n616_));
  NO3        g594(.A(new_new_n573_), .B(new_new_n158_), .C(new_new_n141_), .Y(new_new_n617_));
  INV        g595(.A(new_new_n617_), .Y(new_new_n618_));
  NA4        g596(.A(new_new_n618_), .B(new_new_n616_), .C(new_new_n614_), .D(new_new_n612_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n83_), .B(i_5_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n539_), .B(new_new_n99_), .C(new_new_n108_), .Y(new_new_n621_));
  INV        g599(.A(new_new_n621_), .Y(new_new_n622_));
  NA2        g600(.A(new_new_n622_), .B(new_new_n620_), .Y(new_new_n623_));
  NAi21      g601(.An(new_new_n171_), .B(new_new_n172_), .Y(new_new_n624_));
  NO4        g602(.A(new_new_n170_), .B(new_new_n153_), .C(i_0_), .D(i_12_), .Y(new_new_n625_));
  AOI220     g603(.A0(new_new_n625_), .A1(new_new_n624_), .B0(new_new_n508_), .B1(new_new_n137_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n583_), .B(new_new_n291_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n627_), .B(new_new_n420_), .Y(new_new_n628_));
  NA2        g606(.A(new_new_n628_), .B(new_new_n577_), .Y(new_new_n629_));
  NA3        g607(.A(new_new_n629_), .B(new_new_n626_), .C(new_new_n623_), .Y(new_new_n630_));
  NO4        g608(.A(new_new_n630_), .B(new_new_n619_), .C(new_new_n609_), .D(new_new_n606_), .Y(new_new_n631_));
  INV        g609(.A(new_new_n368_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n632_), .B(new_new_n151_), .Y(new_new_n633_));
  BUFFER     g611(.A(i_7_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n139_), .B(new_new_n140_), .Y(new_new_n635_));
  AO210      g613(.A0(new_new_n634_), .A1(new_new_n33_), .B0(new_new_n635_), .Y(new_new_n636_));
  NAi31      g614(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n637_));
  NO2        g615(.A(new_new_n67_), .B(new_new_n637_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n397_), .Y(new_new_n639_));
  NA2        g617(.A(new_new_n639_), .B(new_new_n636_), .Y(new_new_n640_));
  AOI210     g618(.A0(new_new_n640_), .A1(new_new_n46_), .B0(new_new_n563_), .Y(new_new_n641_));
  AOI210     g619(.A0(new_new_n641_), .A1(new_new_n633_), .B0(new_new_n70_), .Y(new_new_n642_));
  NO3        g620(.A(new_new_n56_), .B(new_new_n55_), .C(i_4_), .Y(new_new_n643_));
  OAI210     g621(.A0(new_new_n662_), .A1(new_new_n201_), .B0(new_new_n643_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n459_), .Y(new_new_n645_));
  NO4        g623(.A(new_new_n593_), .B(i_11_), .C(new_new_n178_), .D(new_new_n177_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n646_), .B(new_new_n334_), .Y(new_new_n647_));
  INV        g625(.A(new_new_n228_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n648_), .A1(new_new_n647_), .B0(new_new_n39_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n649_), .B(new_new_n645_), .Y(new_new_n650_));
  INV        g628(.A(new_new_n650_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n651_), .B(new_new_n642_), .Y(new_new_n652_));
  NA4        g630(.A(new_new_n652_), .B(new_new_n631_), .C(new_new_n599_), .D(new_new_n555_), .Y(ori4));
  INV        g631(.A(new_new_n319_), .Y(new_new_n656_));
  INV        g632(.A(i_6_), .Y(new_new_n657_));
  INV        g633(.A(new_new_n319_), .Y(new_new_n658_));
  INV        g634(.A(new_new_n298_), .Y(new_new_n659_));
  INV        g635(.A(new_new_n450_), .Y(new_new_n660_));
  INV        g636(.A(i_8_), .Y(new_new_n661_));
  INV        g637(.A(i_0_), .Y(new_new_n662_));
endmodule


