library verilog;
use verilog.vl_types.all;
entity dffrs_vlg_vec_tst is
end dffrs_vlg_vec_tst;
