//Benchmark atmr_misex3_1774_0.25

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n534_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  NOi21      o000(.An(i), .B(h), .Y(ori_ori_n29_));
  NOi32      o001(.An(j), .Bn(g), .C(k), .Y(ori_ori_n30_));
  NA2        o002(.A(ori_ori_n30_), .B(m), .Y(ori_ori_n31_));
  INV        o003(.A(h), .Y(ori_ori_n32_));
  INV        o004(.A(i), .Y(ori_ori_n33_));
  AN2        o005(.A(h), .B(g), .Y(ori_ori_n34_));
  NAi21      o006(.An(n), .B(m), .Y(ori_ori_n35_));
  NOi32      o007(.An(k), .Bn(h), .C(l), .Y(ori_ori_n36_));
  NOi32      o008(.An(k), .Bn(h), .C(g), .Y(ori_ori_n37_));
  INV        o009(.A(c), .Y(ori_ori_n38_));
  INV        o010(.A(d), .Y(ori_ori_n39_));
  INV        o011(.A(n), .Y(ori_ori_n40_));
  INV        o012(.A(j), .Y(ori_ori_n41_));
  NOi32      o013(.An(m), .Bn(j), .C(k), .Y(ori_ori_n42_));
  NAi41      o014(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n43_));
  AN2        o015(.A(e), .B(b), .Y(ori_ori_n44_));
  INV        o016(.A(a), .Y(ori_ori_n45_));
  NOi21      o017(.An(m), .B(n), .Y(ori_ori_n46_));
  AN2        o018(.A(k), .B(h), .Y(ori_ori_n47_));
  INV        o019(.A(b), .Y(ori_ori_n48_));
  NOi31      o020(.An(k), .B(m), .C(j), .Y(ori_ori_n49_));
  NA3        o021(.A(ori_ori_n49_), .B(h), .C(n), .Y(ori_ori_n50_));
  NOi31      o022(.An(k), .B(m), .C(i), .Y(ori_ori_n51_));
  INV        o023(.A(ori_ori_n50_), .Y(ori_ori_n52_));
  NOi32      o024(.An(f), .Bn(b), .C(e), .Y(ori_ori_n53_));
  NAi21      o025(.An(m), .B(n), .Y(ori_ori_n54_));
  NAi31      o026(.An(j), .B(k), .C(h), .Y(ori_ori_n55_));
  NAi21      o027(.An(c), .B(b), .Y(ori_ori_n56_));
  NA2        o028(.A(d), .B(b), .Y(ori_ori_n57_));
  NAi21      o029(.An(c), .B(d), .Y(ori_ori_n58_));
  NAi31      o030(.An(l), .B(k), .C(h), .Y(ori_ori_n59_));
  NO2        o031(.A(ori_ori_n54_), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NAi31      o032(.An(e), .B(f), .C(b), .Y(ori_ori_n61_));
  NOi21      o033(.An(h), .B(i), .Y(ori_ori_n62_));
  NOi21      o034(.An(k), .B(m), .Y(ori_ori_n63_));
  NOi21      o035(.An(h), .B(g), .Y(ori_ori_n64_));
  NAi31      o036(.An(d), .B(f), .C(c), .Y(ori_ori_n65_));
  NAi31      o037(.An(e), .B(f), .C(c), .Y(ori_ori_n66_));
  NA2        o038(.A(j), .B(h), .Y(ori_ori_n67_));
  OR3        o039(.A(n), .B(m), .C(k), .Y(ori_ori_n68_));
  NO2        o040(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  NAi21      o041(.An(m), .B(n), .Y(ori_ori_n70_));
  NO2        o042(.A(n), .B(m), .Y(ori_ori_n71_));
  NA2        o043(.A(ori_ori_n71_), .B(ori_ori_n36_), .Y(ori_ori_n72_));
  NAi21      o044(.An(f), .B(e), .Y(ori_ori_n73_));
  NA2        o045(.A(d), .B(c), .Y(ori_ori_n74_));
  NO2        o046(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  NOi21      o047(.An(ori_ori_n75_), .B(ori_ori_n72_), .Y(ori_ori_n76_));
  NAi31      o048(.An(m), .B(n), .C(b), .Y(ori_ori_n77_));
  NAi21      o049(.An(h), .B(f), .Y(ori_ori_n78_));
  NO2        o050(.A(ori_ori_n77_), .B(ori_ori_n58_), .Y(ori_ori_n79_));
  NA2        o051(.A(ori_ori_n79_), .B(k), .Y(ori_ori_n80_));
  NOi32      o052(.An(f), .Bn(c), .C(d), .Y(ori_ori_n81_));
  NOi32      o053(.An(f), .Bn(c), .C(e), .Y(ori_ori_n82_));
  NO2        o054(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n83_));
  NO3        o055(.A(n), .B(m), .C(j), .Y(ori_ori_n84_));
  NA2        o056(.A(ori_ori_n84_), .B(ori_ori_n47_), .Y(ori_ori_n85_));
  AO210      o057(.A0(ori_ori_n85_), .A1(ori_ori_n72_), .B0(ori_ori_n83_), .Y(ori_ori_n86_));
  NAi31      o058(.An(ori_ori_n76_), .B(ori_ori_n86_), .C(ori_ori_n80_), .Y(ori_ori_n87_));
  OR2        o059(.A(ori_ori_n87_), .B(ori_ori_n52_), .Y(ori_ori_n88_));
  INV        o060(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  NA2        o061(.A(m), .B(j), .Y(ori_ori_n90_));
  NAi31      o062(.An(n), .B(h), .C(g), .Y(ori_ori_n91_));
  BUFFER     o063(.A(k), .Y(ori_ori_n92_));
  NAi41      o064(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n93_));
  INV        o065(.A(f), .Y(ori_ori_n94_));
  INV        o066(.A(g), .Y(ori_ori_n95_));
  NOi31      o067(.An(i), .B(j), .C(h), .Y(ori_ori_n96_));
  NOi21      o068(.An(l), .B(m), .Y(ori_ori_n97_));
  NA2        o069(.A(ori_ori_n97_), .B(ori_ori_n96_), .Y(ori_ori_n98_));
  NOi21      o070(.An(n), .B(m), .Y(ori_ori_n99_));
  NAi21      o071(.An(j), .B(h), .Y(ori_ori_n100_));
  XN2        o072(.A(i), .B(h), .Y(ori_ori_n101_));
  NA2        o073(.A(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NOi31      o074(.An(k), .B(n), .C(m), .Y(ori_ori_n103_));
  NOi31      o075(.An(ori_ori_n103_), .B(ori_ori_n74_), .C(ori_ori_n73_), .Y(ori_ori_n104_));
  INV        o076(.A(ori_ori_n104_), .Y(ori_ori_n105_));
  NAi31      o077(.An(f), .B(e), .C(c), .Y(ori_ori_n106_));
  NO3        o078(.A(ori_ori_n106_), .B(ori_ori_n68_), .C(ori_ori_n67_), .Y(ori_ori_n107_));
  NA3        o079(.A(e), .B(c), .C(b), .Y(ori_ori_n108_));
  NAi32      o080(.An(m), .Bn(i), .C(k), .Y(ori_ori_n109_));
  INV        o081(.A(k), .Y(ori_ori_n110_));
  INV        o082(.A(ori_ori_n107_), .Y(ori_ori_n111_));
  BUFFER     o083(.A(n), .Y(ori_ori_n112_));
  NAi41      o084(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n113_));
  NO2        o085(.A(ori_ori_n113_), .B(e), .Y(ori_ori_n114_));
  AN2        o086(.A(ori_ori_n111_), .B(ori_ori_n105_), .Y(ori_ori_n115_));
  BUFFER     o087(.A(g), .Y(ori_ori_n116_));
  NO2        o088(.A(ori_ori_n116_), .B(ori_ori_n43_), .Y(ori_ori_n117_));
  NA2        o089(.A(ori_ori_n117_), .B(ori_ori_n53_), .Y(ori_ori_n118_));
  NA2        o090(.A(ori_ori_n63_), .B(i), .Y(ori_ori_n119_));
  NO2        o091(.A(n), .B(a), .Y(ori_ori_n120_));
  NAi31      o092(.An(ori_ori_n113_), .B(ori_ori_n120_), .C(ori_ori_n44_), .Y(ori_ori_n121_));
  NAi21      o093(.An(h), .B(i), .Y(ori_ori_n122_));
  NA2        o094(.A(ori_ori_n71_), .B(k), .Y(ori_ori_n123_));
  NO2        o095(.A(ori_ori_n123_), .B(ori_ori_n122_), .Y(ori_ori_n124_));
  NA2        o096(.A(ori_ori_n124_), .B(ori_ori_n81_), .Y(ori_ori_n125_));
  NA3        o097(.A(ori_ori_n125_), .B(ori_ori_n121_), .C(ori_ori_n118_), .Y(ori_ori_n126_));
  INV        o098(.A(e), .Y(ori_ori_n127_));
  NOi21      o099(.An(ori_ori_n115_), .B(ori_ori_n126_), .Y(ori_ori_n128_));
  NA3        o100(.A(ori_ori_n39_), .B(c), .C(b), .Y(ori_ori_n129_));
  NA2        o101(.A(k), .B(h), .Y(ori_ori_n130_));
  NA2        o102(.A(ori_ori_n63_), .B(ori_ori_n62_), .Y(ori_ori_n131_));
  NO2        o103(.A(ori_ori_n131_), .B(ori_ori_n83_), .Y(ori_ori_n132_));
  NA2        o104(.A(e), .B(b), .Y(ori_ori_n133_));
  NAi32      o105(.An(j), .Bn(h), .C(i), .Y(ori_ori_n134_));
  NAi21      o106(.An(m), .B(l), .Y(ori_ori_n135_));
  NO3        o107(.A(ori_ori_n135_), .B(ori_ori_n134_), .C(ori_ori_n40_), .Y(ori_ori_n136_));
  INV        o108(.A(h), .Y(ori_ori_n137_));
  NAi32      o109(.An(n), .Bn(m), .C(l), .Y(ori_ori_n138_));
  NO2        o110(.A(ori_ori_n138_), .B(ori_ori_n134_), .Y(ori_ori_n139_));
  NA2        o111(.A(ori_ori_n139_), .B(ori_ori_n75_), .Y(ori_ori_n140_));
  INV        o112(.A(ori_ori_n140_), .Y(ori_ori_n141_));
  NO2        o113(.A(ori_ori_n141_), .B(ori_ori_n132_), .Y(ori_ori_n142_));
  NA2        o114(.A(ori_ori_n124_), .B(ori_ori_n82_), .Y(ori_ori_n143_));
  NAi21      o115(.An(m), .B(k), .Y(ori_ori_n144_));
  NO2        o116(.A(ori_ori_n101_), .B(ori_ori_n144_), .Y(ori_ori_n145_));
  NAi41      o117(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n146_));
  INV        o118(.A(ori_ori_n146_), .Y(ori_ori_n147_));
  NA2        o119(.A(ori_ori_n147_), .B(ori_ori_n145_), .Y(ori_ori_n148_));
  NA2        o120(.A(e), .B(c), .Y(ori_ori_n149_));
  NO3        o121(.A(ori_ori_n149_), .B(n), .C(d), .Y(ori_ori_n150_));
  NOi21      o122(.An(f), .B(h), .Y(ori_ori_n151_));
  NAi31      o123(.An(d), .B(e), .C(b), .Y(ori_ori_n152_));
  NA2        o124(.A(ori_ori_n148_), .B(ori_ori_n143_), .Y(ori_ori_n153_));
  NA2        o125(.A(ori_ori_n120_), .B(ori_ori_n44_), .Y(ori_ori_n154_));
  NOi31      o126(.An(l), .B(n), .C(m), .Y(ori_ori_n155_));
  NA2        o127(.A(ori_ori_n155_), .B(ori_ori_n96_), .Y(ori_ori_n156_));
  NO2        o128(.A(ori_ori_n156_), .B(ori_ori_n83_), .Y(ori_ori_n157_));
  NAi32      o129(.An(m), .Bn(j), .C(k), .Y(ori_ori_n158_));
  NAi41      o130(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n159_));
  NA2        o131(.A(ori_ori_n93_), .B(ori_ori_n159_), .Y(ori_ori_n160_));
  NOi31      o132(.An(j), .B(m), .C(k), .Y(ori_ori_n161_));
  NO2        o133(.A(ori_ori_n49_), .B(ori_ori_n161_), .Y(ori_ori_n162_));
  NAi31      o134(.An(ori_ori_n162_), .B(h), .C(ori_ori_n160_), .Y(ori_ori_n163_));
  NO2        o135(.A(ori_ori_n135_), .B(ori_ori_n134_), .Y(ori_ori_n164_));
  INV        o136(.A(ori_ori_n163_), .Y(ori_ori_n165_));
  NOi32      o137(.An(e), .Bn(b), .C(a), .Y(ori_ori_n166_));
  NA2        o138(.A(ori_ori_n37_), .B(ori_ori_n46_), .Y(ori_ori_n167_));
  NO3        o139(.A(ori_ori_n165_), .B(ori_ori_n157_), .C(ori_ori_n153_), .Y(ori_ori_n168_));
  NA4        o140(.A(ori_ori_n168_), .B(ori_ori_n142_), .C(ori_ori_n128_), .D(ori_ori_n89_), .Y(ori10));
  NO3        o141(.A(ori_ori_n58_), .B(n), .C(ori_ori_n45_), .Y(ori_ori_n170_));
  NAi31      o142(.An(b), .B(f), .C(c), .Y(ori_ori_n171_));
  INV        o143(.A(ori_ori_n171_), .Y(ori_ori_n172_));
  NOi32      o144(.An(k), .Bn(h), .C(j), .Y(ori_ori_n173_));
  NA2        o145(.A(ori_ori_n173_), .B(ori_ori_n99_), .Y(ori_ori_n174_));
  AN2        o146(.A(j), .B(h), .Y(ori_ori_n175_));
  NO3        o147(.A(n), .B(m), .C(k), .Y(ori_ori_n176_));
  NA2        o148(.A(ori_ori_n176_), .B(ori_ori_n175_), .Y(ori_ori_n177_));
  NO3        o149(.A(ori_ori_n177_), .B(ori_ori_n58_), .C(ori_ori_n94_), .Y(ori_ori_n178_));
  OR2        o150(.A(m), .B(k), .Y(ori_ori_n179_));
  NO2        o151(.A(ori_ori_n67_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NA4        o152(.A(n), .B(f), .C(c), .D(ori_ori_n48_), .Y(ori_ori_n181_));
  NOi21      o153(.An(ori_ori_n180_), .B(ori_ori_n181_), .Y(ori_ori_n182_));
  NO2        o154(.A(ori_ori_n182_), .B(ori_ori_n178_), .Y(ori_ori_n183_));
  NO2        o155(.A(ori_ori_n181_), .B(ori_ori_n135_), .Y(ori_ori_n184_));
  NOi32      o156(.An(f), .Bn(d), .C(c), .Y(ori_ori_n185_));
  AOI220     o157(.A0(ori_ori_n185_), .A1(ori_ori_n139_), .B0(ori_ori_n184_), .B1(ori_ori_n96_), .Y(ori_ori_n186_));
  NA2        o158(.A(ori_ori_n186_), .B(ori_ori_n183_), .Y(ori_ori_n187_));
  NA2        o159(.A(ori_ori_n120_), .B(b), .Y(ori_ori_n188_));
  INV        o160(.A(e), .Y(ori_ori_n189_));
  NA2        o161(.A(ori_ori_n34_), .B(e), .Y(ori_ori_n190_));
  NO2        o162(.A(ori_ori_n190_), .B(ori_ori_n90_), .Y(ori_ori_n191_));
  INV        o163(.A(ori_ori_n191_), .Y(ori_ori_n192_));
  NO2        o164(.A(ori_ori_n192_), .B(ori_ori_n188_), .Y(ori_ori_n193_));
  NO2        o165(.A(ori_ori_n193_), .B(ori_ori_n187_), .Y(ori_ori_n194_));
  NOi21      o166(.An(d), .B(c), .Y(ori_ori_n195_));
  OR2        o167(.A(n), .B(m), .Y(ori_ori_n196_));
  NO2        o168(.A(ori_ori_n196_), .B(ori_ori_n59_), .Y(ori_ori_n197_));
  INV        o169(.A(ori_ori_n167_), .Y(ori_ori_n198_));
  NA2        o170(.A(ori_ori_n198_), .B(ori_ori_n166_), .Y(ori_ori_n199_));
  NAi21      o171(.An(k), .B(j), .Y(ori_ori_n200_));
  NAi21      o172(.An(e), .B(d), .Y(ori_ori_n201_));
  INV        o173(.A(ori_ori_n201_), .Y(ori_ori_n202_));
  NO2        o174(.A(ori_ori_n123_), .B(ori_ori_n94_), .Y(ori_ori_n203_));
  NA3        o175(.A(ori_ori_n203_), .B(ori_ori_n202_), .C(ori_ori_n102_), .Y(ori_ori_n204_));
  NA2        o176(.A(ori_ori_n204_), .B(ori_ori_n199_), .Y(ori_ori_n205_));
  NO2        o177(.A(ori_ori_n156_), .B(ori_ori_n94_), .Y(ori_ori_n206_));
  NA2        o178(.A(ori_ori_n206_), .B(ori_ori_n202_), .Y(ori_ori_n207_));
  NOi31      o179(.An(n), .B(m), .C(k), .Y(ori_ori_n208_));
  AOI220     o180(.A0(ori_ori_n208_), .A1(ori_ori_n175_), .B0(ori_ori_n99_), .B1(ori_ori_n36_), .Y(ori_ori_n209_));
  NAi31      o181(.An(g), .B(f), .C(c), .Y(ori_ori_n210_));
  NA2        o182(.A(ori_ori_n207_), .B(ori_ori_n140_), .Y(ori_ori_n211_));
  NO2        o183(.A(ori_ori_n211_), .B(ori_ori_n205_), .Y(ori_ori_n212_));
  AN2        o184(.A(e), .B(d), .Y(ori_ori_n213_));
  NO4        o185(.A(ori_ori_n78_), .B(ori_ori_n43_), .C(ori_ori_n38_), .D(b), .Y(ori_ori_n214_));
  NA2        o186(.A(ori_ori_n172_), .B(ori_ori_n60_), .Y(ori_ori_n215_));
  AOI210     o187(.A0(ori_ori_n109_), .A1(ori_ori_n158_), .B0(ori_ori_n40_), .Y(ori_ori_n216_));
  INV        o188(.A(ori_ori_n50_), .Y(ori_ori_n217_));
  NA2        o189(.A(ori_ori_n50_), .B(ori_ori_n215_), .Y(ori_ori_n218_));
  NO2        o190(.A(ori_ori_n218_), .B(ori_ori_n214_), .Y(ori_ori_n219_));
  INV        o191(.A(ori_ori_n76_), .Y(ori_ori_n220_));
  NA2        o192(.A(ori_ori_n220_), .B(ori_ori_n115_), .Y(ori_ori_n221_));
  OAI210     o193(.A0(ori_ori_n51_), .A1(ori_ori_n49_), .B0(n), .Y(ori_ori_n222_));
  XO2        o194(.A(i), .B(h), .Y(ori_ori_n223_));
  NA3        o195(.A(ori_ori_n223_), .B(ori_ori_n63_), .C(n), .Y(ori_ori_n224_));
  NAi41      o196(.An(ori_ori_n136_), .B(ori_ori_n224_), .C(ori_ori_n209_), .D(ori_ori_n174_), .Y(ori_ori_n225_));
  NOi21      o197(.An(ori_ori_n225_), .B(ori_ori_n129_), .Y(ori_ori_n226_));
  NAi31      o198(.An(c), .B(f), .C(d), .Y(ori_ori_n227_));
  AOI210     o199(.A0(ori_ori_n131_), .A1(ori_ori_n85_), .B0(ori_ori_n227_), .Y(ori_ori_n228_));
  NA2        o200(.A(ori_ori_n103_), .B(i), .Y(ori_ori_n229_));
  NO3        o201(.A(ori_ori_n228_), .B(ori_ori_n226_), .C(ori_ori_n221_), .Y(ori_ori_n230_));
  NA4        o202(.A(ori_ori_n230_), .B(ori_ori_n219_), .C(ori_ori_n212_), .D(ori_ori_n194_), .Y(ori11));
  INV        o203(.A(k), .Y(ori_ori_n232_));
  INV        o204(.A(j), .Y(ori_ori_n233_));
  NAi31      o205(.An(n), .B(m), .C(k), .Y(ori_ori_n234_));
  NO2        o206(.A(ori_ori_n130_), .B(ori_ori_n35_), .Y(ori_ori_n235_));
  NA2        o207(.A(k), .B(ori_ori_n29_), .Y(ori_ori_n236_));
  OAI220     o208(.A0(ori_ori_n236_), .A1(m), .B0(ori_ori_n534_), .B1(ori_ori_n109_), .Y(ori_ori_n237_));
  NOi41      o209(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n238_));
  NAi32      o210(.An(e), .Bn(b), .C(c), .Y(ori_ori_n239_));
  OR2        o211(.A(ori_ori_n239_), .B(ori_ori_n40_), .Y(ori_ori_n240_));
  AN2        o212(.A(ori_ori_n159_), .B(ori_ori_n146_), .Y(ori_ori_n241_));
  NA2        o213(.A(ori_ori_n241_), .B(ori_ori_n240_), .Y(ori_ori_n242_));
  OA210      o214(.A0(ori_ori_n242_), .A1(ori_ori_n238_), .B0(ori_ori_n237_), .Y(ori_ori_n243_));
  AN2        o215(.A(j), .B(h), .Y(ori_ori_n244_));
  NO2        o216(.A(ori_ori_n57_), .B(c), .Y(ori_ori_n245_));
  NA3        o217(.A(ori_ori_n245_), .B(ori_ori_n244_), .C(ori_ori_n208_), .Y(ori_ori_n246_));
  NA3        o218(.A(f), .B(d), .C(b), .Y(ori_ori_n247_));
  NO4        o219(.A(ori_ori_n247_), .B(ori_ori_n70_), .C(ori_ori_n67_), .D(g), .Y(ori_ori_n248_));
  INV        o220(.A(ori_ori_n246_), .Y(ori_ori_n249_));
  NO2        o221(.A(ori_ori_n249_), .B(ori_ori_n243_), .Y(ori_ori_n250_));
  INV        o222(.A(k), .Y(ori_ori_n251_));
  NO2        o223(.A(ori_ori_n144_), .B(n), .Y(ori_ori_n252_));
  NA3        o224(.A(ori_ori_n227_), .B(ori_ori_n66_), .C(ori_ori_n65_), .Y(ori_ori_n253_));
  NA2        o225(.A(ori_ori_n210_), .B(ori_ori_n106_), .Y(ori_ori_n254_));
  OR2        o226(.A(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n255_));
  NA2        o227(.A(ori_ori_n255_), .B(ori_ori_n252_), .Y(ori_ori_n256_));
  NO2        o228(.A(ori_ori_n256_), .B(ori_ori_n41_), .Y(ori_ori_n257_));
  NA3        o229(.A(ori_ori_n238_), .B(ori_ori_n161_), .C(ori_ori_n34_), .Y(ori_ori_n258_));
  NOi32      o230(.An(e), .Bn(c), .C(f), .Y(ori_ori_n259_));
  NOi21      o231(.An(f), .B(g), .Y(ori_ori_n260_));
  NO2        o232(.A(ori_ori_n260_), .B(ori_ori_n93_), .Y(ori_ori_n261_));
  INV        o233(.A(ori_ori_n258_), .Y(ori_ori_n262_));
  NA2        o234(.A(ori_ori_n223_), .B(ori_ori_n63_), .Y(ori_ori_n263_));
  AN3        o235(.A(f), .B(d), .C(b), .Y(ori_ori_n264_));
  OAI210     o236(.A0(ori_ori_n264_), .A1(ori_ori_n53_), .B0(n), .Y(ori_ori_n265_));
  NA3        o237(.A(ori_ori_n223_), .B(ori_ori_n63_), .C(ori_ori_n95_), .Y(ori_ori_n266_));
  AOI210     o238(.A0(ori_ori_n265_), .A1(ori_ori_n108_), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  NAi31      o239(.An(m), .B(n), .C(k), .Y(ori_ori_n268_));
  INV        o240(.A(ori_ori_n121_), .Y(ori_ori_n269_));
  NO2        o241(.A(ori_ori_n269_), .B(ori_ori_n267_), .Y(ori_ori_n270_));
  INV        o242(.A(ori_ori_n270_), .Y(ori_ori_n271_));
  NO3        o243(.A(ori_ori_n271_), .B(ori_ori_n262_), .C(ori_ori_n257_), .Y(ori_ori_n272_));
  NA2        o244(.A(ori_ori_n170_), .B(ori_ori_n64_), .Y(ori_ori_n273_));
  NA2        o245(.A(h), .B(f), .Y(ori_ori_n274_));
  NO2        o246(.A(ori_ori_n273_), .B(ori_ori_n232_), .Y(ori_ori_n275_));
  NO3        o247(.A(g), .B(ori_ori_n94_), .C(ori_ori_n38_), .Y(ori_ori_n276_));
  NA2        o248(.A(ori_ori_n180_), .B(ori_ori_n276_), .Y(ori_ori_n277_));
  NA2        o249(.A(h), .B(ori_ori_n30_), .Y(ori_ori_n278_));
  NA2        o250(.A(ori_ori_n42_), .B(ori_ori_n34_), .Y(ori_ori_n279_));
  NO2        o251(.A(ori_ori_n279_), .B(ori_ori_n154_), .Y(ori_ori_n280_));
  INV        o252(.A(ori_ori_n280_), .Y(ori_ori_n281_));
  NA2        o253(.A(ori_ori_n281_), .B(ori_ori_n277_), .Y(ori_ori_n282_));
  NO3        o254(.A(ori_ori_n185_), .B(ori_ori_n82_), .C(ori_ori_n81_), .Y(ori_ori_n283_));
  NA2        o255(.A(ori_ori_n283_), .B(ori_ori_n106_), .Y(ori_ori_n284_));
  NO3        o256(.A(ori_ori_n210_), .B(ori_ori_n67_), .C(i), .Y(ori_ori_n285_));
  INV        o257(.A(ori_ori_n183_), .Y(ori_ori_n286_));
  NO3        o258(.A(ori_ori_n286_), .B(ori_ori_n282_), .C(ori_ori_n275_), .Y(ori_ori_n287_));
  NA3        o259(.A(ori_ori_n287_), .B(ori_ori_n272_), .C(ori_ori_n250_), .Y(ori08));
  NO2        o260(.A(k), .B(h), .Y(ori_ori_n289_));
  AO210      o261(.A0(ori_ori_n122_), .A1(ori_ori_n200_), .B0(ori_ori_n289_), .Y(ori_ori_n290_));
  NO2        o262(.A(ori_ori_n290_), .B(ori_ori_n135_), .Y(ori_ori_n291_));
  NA2        o263(.A(ori_ori_n259_), .B(ori_ori_n40_), .Y(ori_ori_n292_));
  NA2        o264(.A(ori_ori_n292_), .B(ori_ori_n210_), .Y(ori_ori_n293_));
  NA2        o265(.A(ori_ori_n293_), .B(ori_ori_n291_), .Y(ori_ori_n294_));
  AOI210     o266(.A0(ori_ori_n247_), .A1(ori_ori_n61_), .B0(ori_ori_n40_), .Y(ori_ori_n295_));
  NA3        o267(.A(ori_ori_n97_), .B(k), .C(h), .Y(ori_ori_n296_));
  INV        o268(.A(ori_ori_n294_), .Y(ori_ori_n297_));
  NO2        o269(.A(ori_ori_n144_), .B(g), .Y(ori_ori_n298_));
  NA2        o270(.A(ori_ori_n290_), .B(ori_ori_n55_), .Y(ori_ori_n299_));
  NA2        o271(.A(ori_ori_n299_), .B(ori_ori_n184_), .Y(ori_ori_n300_));
  INV        o272(.A(ori_ori_n300_), .Y(ori_ori_n301_));
  NA3        o273(.A(ori_ori_n284_), .B(ori_ori_n155_), .C(ori_ori_n173_), .Y(ori_ori_n302_));
  INV        o274(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  NO3        o275(.A(ori_ori_n303_), .B(ori_ori_n301_), .C(ori_ori_n297_), .Y(ori_ori_n304_));
  NA2        o276(.A(ori_ori_n261_), .B(ori_ori_n180_), .Y(ori_ori_n305_));
  NA3        o277(.A(ori_ori_n167_), .B(ori_ori_n305_), .C(ori_ori_n121_), .Y(ori_ori_n306_));
  NO4        o278(.A(ori_ori_n283_), .B(ori_ori_n67_), .C(n), .D(i), .Y(ori_ori_n307_));
  NO2        o279(.A(ori_ori_n307_), .B(ori_ori_n285_), .Y(ori_ori_n308_));
  NO2        o280(.A(ori_ori_n308_), .B(m), .Y(ori_ori_n309_));
  AOI210     o281(.A0(ori_ori_n306_), .A1(l), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  NA2        o282(.A(ori_ori_n254_), .B(ori_ori_n139_), .Y(ori_ori_n311_));
  INV        o283(.A(ori_ori_n311_), .Y(ori_ori_n312_));
  NO2        o284(.A(ori_ori_n135_), .B(ori_ori_n55_), .Y(ori_ori_n313_));
  AOI220     o285(.A0(ori_ori_n313_), .A1(ori_ori_n261_), .B0(ori_ori_n298_), .B1(ori_ori_n295_), .Y(ori_ori_n314_));
  INV        o286(.A(ori_ori_n314_), .Y(ori_ori_n315_));
  OR2        o287(.A(ori_ori_n315_), .B(ori_ori_n312_), .Y(ori_ori_n316_));
  INV        o288(.A(ori_ori_n240_), .Y(ori_ori_n317_));
  NA4        o289(.A(ori_ori_n317_), .B(ori_ori_n97_), .C(ori_ori_n200_), .D(ori_ori_n29_), .Y(ori_ori_n318_));
  NO2        o290(.A(ori_ori_n154_), .B(ori_ori_n31_), .Y(ori_ori_n319_));
  INV        o291(.A(ori_ori_n319_), .Y(ori_ori_n320_));
  NA2        o292(.A(ori_ori_n320_), .B(ori_ori_n318_), .Y(ori_ori_n321_));
  NO3        o293(.A(ori_ori_n157_), .B(ori_ori_n321_), .C(ori_ori_n316_), .Y(ori_ori_n322_));
  NO2        o294(.A(ori_ori_n162_), .B(ori_ori_n137_), .Y(ori_ori_n323_));
  INV        o295(.A(ori_ori_n186_), .Y(ori_ori_n324_));
  NO2        o296(.A(ori_ori_n239_), .B(ori_ori_n40_), .Y(ori_ori_n325_));
  NA2        o297(.A(ori_ori_n323_), .B(ori_ori_n325_), .Y(ori_ori_n326_));
  OAI210     o298(.A0(ori_ori_n296_), .A1(ori_ori_n181_), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  NO2        o299(.A(ori_ori_n283_), .B(n), .Y(ori_ori_n328_));
  BUFFER     o300(.A(ori_ori_n313_), .Y(ori_ori_n329_));
  AOI220     o301(.A0(ori_ori_n329_), .A1(ori_ori_n276_), .B0(ori_ori_n328_), .B1(ori_ori_n291_), .Y(ori_ori_n330_));
  INV        o302(.A(ori_ori_n330_), .Y(ori_ori_n331_));
  NO3        o303(.A(ori_ori_n331_), .B(ori_ori_n327_), .C(ori_ori_n324_), .Y(ori_ori_n332_));
  NA4        o304(.A(ori_ori_n332_), .B(ori_ori_n322_), .C(ori_ori_n310_), .D(ori_ori_n304_), .Y(ori09));
  INV        o305(.A(ori_ori_n159_), .Y(ori_ori_n334_));
  NO2        o306(.A(ori_ori_n51_), .B(ori_ori_n49_), .Y(ori_ori_n335_));
  NO2        o307(.A(ori_ori_n335_), .B(f), .Y(ori_ori_n336_));
  NA2        o308(.A(ori_ori_n336_), .B(ori_ori_n334_), .Y(ori_ori_n337_));
  NA2        o309(.A(ori_ori_n290_), .B(ori_ori_n55_), .Y(ori_ori_n338_));
  NA2        o310(.A(ori_ori_n338_), .B(ori_ori_n79_), .Y(ori_ori_n339_));
  NA2        o311(.A(ori_ori_n339_), .B(ori_ori_n337_), .Y(ori_ori_n340_));
  NO2        o312(.A(ori_ori_n268_), .B(ori_ori_n152_), .Y(ori_ori_n341_));
  NA3        o313(.A(c), .B(ori_ori_n225_), .C(f), .Y(ori_ori_n342_));
  OR2        o314(.A(ori_ori_n274_), .B(ori_ori_n234_), .Y(ori_ori_n343_));
  INV        o315(.A(ori_ori_n343_), .Y(ori_ori_n344_));
  NA2        o316(.A(ori_ori_n44_), .B(ori_ori_n344_), .Y(ori_ori_n345_));
  NA2        o317(.A(ori_ori_n345_), .B(ori_ori_n342_), .Y(ori_ori_n346_));
  NO3        o318(.A(ori_ori_n346_), .B(ori_ori_n217_), .C(ori_ori_n340_), .Y(ori_ori_n347_));
  NO2        o319(.A(ori_ori_n106_), .B(ori_ori_n100_), .Y(ori_ori_n348_));
  NA2        o320(.A(ori_ori_n348_), .B(ori_ori_n103_), .Y(ori_ori_n349_));
  NA2        o321(.A(e), .B(d), .Y(ori_ori_n350_));
  OAI220     o322(.A0(ori_ori_n350_), .A1(c), .B0(ori_ori_n149_), .B1(d), .Y(ori_ori_n351_));
  NA2        o323(.A(ori_ori_n351_), .B(ori_ori_n203_), .Y(ori_ori_n352_));
  AOI210     o324(.A0(ori_ori_n229_), .A1(ori_ori_n72_), .B0(ori_ori_n106_), .Y(ori_ori_n353_));
  INV        o325(.A(ori_ori_n353_), .Y(ori_ori_n354_));
  NA2        o326(.A(ori_ori_n354_), .B(ori_ori_n352_), .Y(ori_ori_n355_));
  INV        o327(.A(ori_ori_n355_), .Y(ori_ori_n356_));
  OR2        o328(.A(ori_ori_n292_), .B(ori_ori_n98_), .Y(ori_ori_n357_));
  NA2        o329(.A(h), .B(ori_ori_n341_), .Y(ori_ori_n358_));
  BUFFER     o330(.A(ori_ori_n69_), .Y(ori_ori_n359_));
  OAI210     o331(.A0(ori_ori_n359_), .A1(ori_ori_n206_), .B0(ori_ori_n351_), .Y(ori_ori_n360_));
  AN3        o332(.A(ori_ori_n360_), .B(ori_ori_n358_), .C(ori_ori_n357_), .Y(ori_ori_n361_));
  NA3        o333(.A(ori_ori_n361_), .B(ori_ori_n356_), .C(ori_ori_n347_), .Y(ori12));
  NO2        o334(.A(ori_ori_n201_), .B(c), .Y(ori_ori_n363_));
  NO4        o335(.A(ori_ori_n196_), .B(ori_ori_n122_), .C(ori_ori_n251_), .D(ori_ori_n95_), .Y(ori_ori_n364_));
  NA2        o336(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NO2        o337(.A(ori_ori_n201_), .B(ori_ori_n48_), .Y(ori_ori_n366_));
  NA2        o338(.A(ori_ori_n51_), .B(ori_ori_n366_), .Y(ori_ori_n367_));
  NA2        o339(.A(ori_ori_n367_), .B(ori_ori_n365_), .Y(ori_ori_n368_));
  AOI210     o340(.A0(ori_ori_n109_), .A1(ori_ori_n158_), .B0(ori_ori_n91_), .Y(ori_ori_n369_));
  OR2        o341(.A(ori_ori_n369_), .B(ori_ori_n364_), .Y(ori_ori_n370_));
  AOI210     o342(.A0(ori_ori_n156_), .A1(ori_ori_n177_), .B0(ori_ori_n95_), .Y(ori_ori_n371_));
  OAI210     o343(.A0(ori_ori_n371_), .A1(ori_ori_n370_), .B0(ori_ori_n185_), .Y(ori_ori_n372_));
  NO2        o344(.A(ori_ori_n58_), .B(ori_ori_n112_), .Y(ori_ori_n373_));
  NA2        o345(.A(ori_ori_n373_), .B(ori_ori_n114_), .Y(ori_ori_n374_));
  NA2        o346(.A(ori_ori_n374_), .B(ori_ori_n372_), .Y(ori_ori_n375_));
  NA3        o347(.A(ori_ori_n197_), .B(ori_ori_n195_), .C(ori_ori_n73_), .Y(ori_ori_n376_));
  INV        o348(.A(ori_ori_n376_), .Y(ori_ori_n377_));
  NO3        o349(.A(ori_ori_n377_), .B(ori_ori_n375_), .C(ori_ori_n368_), .Y(ori_ori_n378_));
  NOi21      o350(.An(ori_ori_n29_), .B(ori_ori_n268_), .Y(ori_ori_n379_));
  INV        o351(.A(ori_ori_n121_), .Y(ori_ori_n380_));
  INV        o352(.A(ori_ori_n148_), .Y(ori_ori_n381_));
  NO2        o353(.A(ori_ori_n222_), .B(ori_ori_n137_), .Y(ori_ori_n382_));
  NO3        o354(.A(ori_ori_n382_), .B(ori_ori_n381_), .C(ori_ori_n380_), .Y(ori_ori_n383_));
  INV        o355(.A(ori_ori_n164_), .Y(ori_ori_n384_));
  NA2        o356(.A(ori_ori_n64_), .B(i), .Y(ori_ori_n385_));
  NA2        o357(.A(ori_ori_n34_), .B(i), .Y(ori_ori_n386_));
  NO2        o358(.A(ori_ori_n386_), .B(ori_ori_n90_), .Y(ori_ori_n387_));
  INV        o359(.A(ori_ori_n387_), .Y(ori_ori_n388_));
  NA2        o360(.A(ori_ori_n239_), .B(ori_ori_n171_), .Y(ori_ori_n389_));
  AOI210     o361(.A0(ori_ori_n389_), .A1(n), .B0(ori_ori_n238_), .Y(ori_ori_n390_));
  OAI220     o362(.A0(ori_ori_n390_), .A1(ori_ori_n384_), .B0(ori_ori_n388_), .B1(ori_ori_n154_), .Y(ori_ori_n391_));
  NA3        o363(.A(ori_ori_n151_), .B(i), .C(g), .Y(ori_ori_n392_));
  AOI210     o364(.A0(ori_ori_n278_), .A1(ori_ori_n392_), .B0(m), .Y(ori_ori_n393_));
  OAI210     o365(.A0(ori_ori_n393_), .A1(ori_ori_n51_), .B0(ori_ori_n150_), .Y(ori_ori_n394_));
  INV        o366(.A(ori_ori_n394_), .Y(ori_ori_n395_));
  NO2        o367(.A(ori_ori_n209_), .B(ori_ori_n95_), .Y(ori_ori_n396_));
  NA2        o368(.A(ori_ori_n396_), .B(ori_ori_n172_), .Y(ori_ori_n397_));
  INV        o369(.A(ori_ori_n397_), .Y(ori_ori_n398_));
  NA2        o370(.A(ori_ori_n393_), .B(ori_ori_n366_), .Y(ori_ori_n399_));
  INV        o371(.A(ori_ori_n399_), .Y(ori_ori_n400_));
  NO4        o372(.A(ori_ori_n400_), .B(ori_ori_n398_), .C(ori_ori_n395_), .D(ori_ori_n391_), .Y(ori_ori_n401_));
  NAi31      o373(.An(ori_ori_n56_), .B(h), .C(n), .Y(ori_ori_n402_));
  NO2        o374(.A(ori_ori_n49_), .B(ori_ori_n161_), .Y(ori_ori_n403_));
  NO2        o375(.A(ori_ori_n403_), .B(ori_ori_n402_), .Y(ori_ori_n404_));
  NA2        o376(.A(ori_ori_n106_), .B(ori_ori_n66_), .Y(ori_ori_n405_));
  NO3        o377(.A(ori_ori_n139_), .B(ori_ori_n197_), .C(ori_ori_n69_), .Y(ori_ori_n406_));
  NOi31      o378(.An(ori_ori_n405_), .B(ori_ori_n406_), .C(ori_ori_n95_), .Y(ori_ori_n407_));
  NAi21      o379(.An(ori_ori_n239_), .B(ori_ori_n396_), .Y(ori_ori_n408_));
  INV        o380(.A(ori_ori_n214_), .Y(ori_ori_n409_));
  NA2        o381(.A(ori_ori_n409_), .B(ori_ori_n408_), .Y(ori_ori_n410_));
  NA2        o382(.A(ori_ori_n369_), .B(ori_ori_n363_), .Y(ori_ori_n411_));
  NA2        o383(.A(ori_ori_n411_), .B(ori_ori_n258_), .Y(ori_ori_n412_));
  OAI210     o384(.A0(ori_ori_n369_), .A1(ori_ori_n364_), .B0(ori_ori_n405_), .Y(ori_ori_n413_));
  NA3        o385(.A(ori_ori_n389_), .B(ori_ori_n216_), .C(ori_ori_n34_), .Y(ori_ori_n414_));
  NA2        o386(.A(ori_ori_n414_), .B(ori_ori_n413_), .Y(ori_ori_n415_));
  OR2        o387(.A(ori_ori_n415_), .B(ori_ori_n412_), .Y(ori_ori_n416_));
  NO4        o388(.A(ori_ori_n416_), .B(ori_ori_n410_), .C(ori_ori_n407_), .D(ori_ori_n404_), .Y(ori_ori_n417_));
  NA4        o389(.A(ori_ori_n417_), .B(ori_ori_n401_), .C(ori_ori_n383_), .D(ori_ori_n378_), .Y(ori13));
  NA2        o390(.A(c), .B(ori_ori_n48_), .Y(ori_ori_n419_));
  NA3        o391(.A(k), .B(j), .C(i), .Y(ori_ori_n420_));
  NO2        o392(.A(f), .B(c), .Y(ori_ori_n421_));
  NOi21      o393(.An(ori_ori_n421_), .B(ori_ori_n196_), .Y(ori_ori_n422_));
  OR2        o394(.A(m), .B(i), .Y(ori_ori_n423_));
  AN3        o395(.A(g), .B(f), .C(c), .Y(ori_ori_n424_));
  NA2        o396(.A(i), .B(h), .Y(ori_ori_n425_));
  NO2        o397(.A(n), .B(f), .Y(ori_ori_n426_));
  NO2        o398(.A(ori_ori_n133_), .B(a), .Y(ori_ori_n427_));
  INV        o399(.A(b), .Y(ori_ori_n428_));
  NO2        o400(.A(a), .B(ori_ori_n428_), .Y(ori_ori_n429_));
  NA2        o401(.A(ori_ori_n191_), .B(ori_ori_n429_), .Y(ori_ori_n430_));
  NA2        o402(.A(ori_ori_n235_), .B(ori_ori_n427_), .Y(ori_ori_n431_));
  NA2        o403(.A(ori_ori_n431_), .B(ori_ori_n430_), .Y(ori00));
  NA2        o404(.A(ori_ori_n225_), .B(f), .Y(ori_ori_n433_));
  OAI210     o405(.A0(ori_ori_n403_), .A1(ori_ori_n32_), .B0(ori_ori_n263_), .Y(ori_ori_n434_));
  NA3        o406(.A(ori_ori_n434_), .B(ori_ori_n127_), .C(n), .Y(ori_ori_n435_));
  AOI210     o407(.A0(ori_ori_n435_), .A1(ori_ori_n433_), .B0(ori_ori_n419_), .Y(ori_ori_n436_));
  INV        o408(.A(ori_ori_n436_), .Y(ori_ori_n437_));
  NA2        o409(.A(ori_ori_n173_), .B(ori_ori_n99_), .Y(ori_ori_n438_));
  OR2        o410(.A(ori_ori_n438_), .B(c), .Y(ori_ori_n439_));
  INV        o411(.A(ori_ori_n248_), .Y(ori_ori_n440_));
  AN3        o412(.A(ori_ori_n440_), .B(ori_ori_n439_), .C(ori_ori_n246_), .Y(ori_ori_n441_));
  NA4        o413(.A(ori_ori_n264_), .B(ori_ori_n92_), .C(ori_ori_n99_), .D(ori_ori_n64_), .Y(ori_ori_n442_));
  INV        o414(.A(ori_ori_n442_), .Y(ori_ori_n443_));
  AOI220     o415(.A0(ori_ori_n379_), .A1(ori_ori_n245_), .B0(ori_ori_n264_), .B1(ori_ori_n117_), .Y(ori_ori_n444_));
  INV        o416(.A(ori_ori_n444_), .Y(ori_ori_n445_));
  NO2        o417(.A(ori_ori_n445_), .B(ori_ori_n443_), .Y(ori_ori_n446_));
  NA3        o418(.A(ori_ori_n446_), .B(ori_ori_n441_), .C(ori_ori_n437_), .Y(ori01));
  INV        o419(.A(ori_ori_n132_), .Y(ori_ori_n448_));
  NA2        o420(.A(ori_ori_n182_), .B(i), .Y(ori_ori_n449_));
  NA3        o421(.A(ori_ori_n449_), .B(ori_ori_n448_), .C(ori_ori_n411_), .Y(ori_ori_n450_));
  NA2        o422(.A(ori_ori_n239_), .B(ori_ori_n129_), .Y(ori_ori_n451_));
  NA2        o423(.A(ori_ori_n382_), .B(ori_ori_n451_), .Y(ori_ori_n452_));
  NA2        o424(.A(ori_ori_n452_), .B(ori_ori_n358_), .Y(ori_ori_n453_));
  NA2        o425(.A(ori_ori_n442_), .B(ori_ori_n349_), .Y(ori_ori_n454_));
  NO2        o426(.A(ori_ori_n280_), .B(ori_ori_n228_), .Y(ori_ori_n455_));
  OR2        o427(.A(ori_ori_n85_), .B(ori_ori_n83_), .Y(ori_ori_n456_));
  NA2        o428(.A(ori_ori_n456_), .B(ori_ori_n455_), .Y(ori_ori_n457_));
  NO4        o429(.A(ori_ori_n457_), .B(ori_ori_n454_), .C(ori_ori_n453_), .D(ori_ori_n450_), .Y(ori_ori_n458_));
  NA2        o430(.A(ori_ori_n131_), .B(ori_ori_n85_), .Y(ori_ori_n459_));
  NA2        o431(.A(ori_ori_n459_), .B(ori_ori_n276_), .Y(ori_ori_n460_));
  NO2        o432(.A(ori_ori_n385_), .B(ori_ori_n108_), .Y(ori_ori_n461_));
  NO2        o433(.A(ori_ori_n386_), .B(ori_ori_n241_), .Y(ori_ori_n462_));
  OAI210     o434(.A0(ori_ori_n462_), .A1(ori_ori_n461_), .B0(ori_ori_n161_), .Y(ori_ori_n463_));
  OR2        o435(.A(ori_ori_n438_), .B(c), .Y(ori_ori_n464_));
  INV        o436(.A(ori_ori_n464_), .Y(ori_ori_n465_));
  NOi21      o437(.An(ori_ori_n463_), .B(ori_ori_n465_), .Y(ori_ori_n466_));
  NO2        o438(.A(g), .B(ori_ori_n33_), .Y(ori_ori_n467_));
  AO220      o439(.A0(h), .A1(ori_ori_n261_), .B0(ori_ori_n467_), .B1(ori_ori_n295_), .Y(ori_ori_n468_));
  NA2        o440(.A(ori_ori_n468_), .B(ori_ori_n161_), .Y(ori_ori_n469_));
  NO3        o441(.A(ori_ori_n425_), .B(ori_ori_n70_), .C(ori_ori_n41_), .Y(ori_ori_n470_));
  INV        o442(.A(ori_ori_n469_), .Y(ori_ori_n471_));
  NO2        o443(.A(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n472_));
  NO4        o444(.A(ori_ori_n425_), .B(ori_ori_n472_), .C(ori_ori_n68_), .D(ori_ori_n41_), .Y(ori_ori_n473_));
  NO2        o445(.A(ori_ori_n473_), .B(ori_ori_n471_), .Y(ori_ori_n474_));
  NA4        o446(.A(ori_ori_n474_), .B(ori_ori_n466_), .C(ori_ori_n460_), .D(ori_ori_n458_), .Y(ori06));
  NO2        o447(.A(ori_ori_n100_), .B(ori_ori_n43_), .Y(ori_ori_n476_));
  OAI210     o448(.A0(ori_ori_n476_), .A1(ori_ori_n470_), .B0(ori_ori_n172_), .Y(ori_ori_n477_));
  NA2        o449(.A(ori_ori_n477_), .B(ori_ori_n463_), .Y(ori_ori_n478_));
  NO2        o450(.A(ori_ori_n478_), .B(ori_ori_n126_), .Y(ori_ori_n479_));
  AOI210     o451(.A0(i), .A1(ori_ori_n238_), .B0(ori_ori_n461_), .Y(ori_ori_n480_));
  AOI210     o452(.A0(i), .A1(ori_ori_n242_), .B0(ori_ori_n468_), .Y(ori_ori_n481_));
  AOI210     o453(.A0(ori_ori_n481_), .A1(ori_ori_n480_), .B0(ori_ori_n158_), .Y(ori_ori_n482_));
  INV        o454(.A(ori_ori_n279_), .Y(ori_ori_n483_));
  NA2        o455(.A(ori_ori_n483_), .B(ori_ori_n166_), .Y(ori_ori_n484_));
  NO2        o456(.A(ori_ori_n229_), .B(ori_ori_n66_), .Y(ori_ori_n485_));
  NO2        o457(.A(ori_ori_n210_), .B(ori_ori_n119_), .Y(ori_ori_n486_));
  NO2        o458(.A(ori_ori_n486_), .B(ori_ori_n485_), .Y(ori_ori_n487_));
  NA2        o459(.A(ori_ori_n487_), .B(ori_ori_n484_), .Y(ori_ori_n488_));
  NO2        o460(.A(ori_ori_n488_), .B(ori_ori_n482_), .Y(ori_ori_n489_));
  OAI220     o461(.A0(ori_ori_n292_), .A1(ori_ori_n119_), .B0(ori_ori_n227_), .B1(ori_ori_n229_), .Y(ori_ori_n490_));
  INV        o462(.A(ori_ori_n490_), .Y(ori_ori_n491_));
  NA2        o463(.A(ori_ori_n491_), .B(ori_ori_n444_), .Y(ori_ori_n492_));
  AN2        o464(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n493_));
  NO2        o465(.A(ori_ori_n493_), .B(ori_ori_n214_), .Y(ori_ori_n494_));
  INV        o466(.A(ori_ori_n494_), .Y(ori_ori_n495_));
  NAi21      o467(.An(j), .B(i), .Y(ori_ori_n496_));
  NO4        o468(.A(ori_ori_n472_), .B(ori_ori_n496_), .C(ori_ori_n196_), .D(ori_ori_n110_), .Y(ori_ori_n497_));
  NO3        o469(.A(ori_ori_n497_), .B(ori_ori_n495_), .C(ori_ori_n492_), .Y(ori_ori_n498_));
  NA4        o470(.A(ori_ori_n498_), .B(ori_ori_n489_), .C(ori_ori_n479_), .D(ori_ori_n474_), .Y(ori07));
  NO2        o471(.A(m), .B(h), .Y(ori_ori_n500_));
  NO2        o472(.A(ori_ori_n420_), .B(ori_ori_n138_), .Y(ori_ori_n501_));
  NO2        o473(.A(l), .B(k), .Y(ori_ori_n502_));
  NO3        o474(.A(ori_ori_n196_), .B(d), .C(c), .Y(ori_ori_n503_));
  NA2        o475(.A(ori_ori_n424_), .B(ori_ori_n213_), .Y(ori_ori_n504_));
  NO2        o476(.A(ori_ori_n504_), .B(ori_ori_n196_), .Y(ori_ori_n505_));
  INV        o477(.A(ori_ori_n505_), .Y(ori_ori_n506_));
  NA2        o478(.A(ori_ori_n500_), .B(ori_ori_n502_), .Y(ori_ori_n507_));
  INV        o479(.A(ori_ori_n507_), .Y(ori_ori_n508_));
  NA2        o480(.A(ori_ori_n426_), .B(ori_ori_n189_), .Y(ori_ori_n509_));
  NO2        o481(.A(ori_ori_n509_), .B(ori_ori_n195_), .Y(ori_ori_n510_));
  OR2        o482(.A(ori_ori_n510_), .B(ori_ori_n508_), .Y(ori_ori_n511_));
  INV        o483(.A(ori_ori_n511_), .Y(ori_ori_n512_));
  NA3        o484(.A(ori_ori_n512_), .B(ori_ori_n506_), .C(ori_ori_n35_), .Y(ori_ori_n513_));
  NO2        o485(.A(ori_ori_n179_), .B(j), .Y(ori_ori_n514_));
  NA2        o486(.A(ori_ori_n422_), .B(e), .Y(ori_ori_n515_));
  INV        o487(.A(ori_ori_n515_), .Y(ori_ori_n516_));
  NA2        o488(.A(ori_ori_n514_), .B(ori_ori_n62_), .Y(ori_ori_n517_));
  INV        o489(.A(ori_ori_n517_), .Y(ori_ori_n518_));
  NO2        o490(.A(ori_ori_n518_), .B(ori_ori_n516_), .Y(ori_ori_n519_));
  NO2        o491(.A(ori_ori_n423_), .B(h), .Y(ori_ori_n520_));
  NO2        o492(.A(ori_ori_n496_), .B(ori_ori_n68_), .Y(ori_ori_n521_));
  NA2        o493(.A(h), .B(ori_ori_n521_), .Y(ori_ori_n522_));
  INV        o494(.A(ori_ori_n522_), .Y(ori_ori_n523_));
  NO2        o495(.A(ori_ori_n523_), .B(ori_ori_n520_), .Y(ori_ori_n524_));
  NA2        o496(.A(ori_ori_n524_), .B(ori_ori_n519_), .Y(ori_ori_n525_));
  NA2        o497(.A(h), .B(ori_ori_n501_), .Y(ori_ori_n526_));
  OR2        o498(.A(h), .B(ori_ori_n233_), .Y(ori_ori_n527_));
  NO2        o499(.A(ori_ori_n527_), .B(ori_ori_n68_), .Y(ori_ori_n528_));
  NO2        o500(.A(ori_ori_n528_), .B(ori_ori_n503_), .Y(ori_ori_n529_));
  NA3        o501(.A(ori_ori_n529_), .B(ori_ori_n54_), .C(ori_ori_n526_), .Y(ori_ori_n530_));
  OR3        o502(.A(ori_ori_n530_), .B(ori_ori_n525_), .C(ori_ori_n513_), .Y(ori04));
  INV        o503(.A(h), .Y(ori_ori_n534_));
  ZERO       o504(.Y(ori02));
  ZERO       o505(.Y(ori03));
  ZERO       o506(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NO3        m0013(.A(n), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n42_));
  INV        m0014(.A(i), .Y(mai_mai_n43_));
  AN2        m0015(.A(h), .B(g), .Y(mai_mai_n44_));
  NA2        m0016(.A(mai_mai_n44_), .B(mai_mai_n43_), .Y(mai_mai_n45_));
  NAi21      m0017(.An(n), .B(m), .Y(mai_mai_n46_));
  NOi32      m0018(.An(k), .Bn(h), .C(l), .Y(mai_mai_n47_));
  NOi32      m0019(.An(k), .Bn(h), .C(g), .Y(mai_mai_n48_));
  NO2        m0020(.A(mai_mai_n48_), .B(mai_mai_n47_), .Y(mai_mai_n49_));
  NO2        m0021(.A(mai_mai_n49_), .B(mai_mai_n46_), .Y(mai_mai_n50_));
  NO2        m0022(.A(mai_mai_n46_), .B(mai_mai_n32_), .Y(mai_mai_n51_));
  INV        m0023(.A(c), .Y(mai_mai_n52_));
  NA2        m0024(.A(e), .B(b), .Y(mai_mai_n53_));
  NO2        m0025(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  INV        m0026(.A(d), .Y(mai_mai_n55_));
  NA3        m0027(.A(g), .B(mai_mai_n55_), .C(a), .Y(mai_mai_n56_));
  NAi21      m0028(.An(i), .B(h), .Y(mai_mai_n57_));
  NAi31      m0029(.An(i), .B(l), .C(j), .Y(mai_mai_n58_));
  NAi21      m0030(.An(i), .B(j), .Y(mai_mai_n59_));
  NAi32      m0031(.An(n), .Bn(k), .C(m), .Y(mai_mai_n60_));
  NAi31      m0032(.An(l), .B(m), .C(k), .Y(mai_mai_n61_));
  NAi21      m0033(.An(e), .B(h), .Y(mai_mai_n62_));
  NAi41      m0034(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n63_));
  INV        m0035(.A(m), .Y(mai_mai_n64_));
  NOi21      m0036(.An(k), .B(l), .Y(mai_mai_n65_));
  NA2        m0037(.A(mai_mai_n65_), .B(mai_mai_n64_), .Y(mai_mai_n66_));
  AN4        m0038(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n67_));
  NOi31      m0039(.An(h), .B(g), .C(f), .Y(mai_mai_n68_));
  NA2        m0040(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NAi32      m0041(.An(m), .Bn(k), .C(j), .Y(mai_mai_n70_));
  NOi32      m0042(.An(h), .Bn(g), .C(f), .Y(mai_mai_n71_));
  NA2        m0043(.A(mai_mai_n71_), .B(mai_mai_n67_), .Y(mai_mai_n72_));
  OA220      m0044(.A0(mai_mai_n72_), .A1(mai_mai_n70_), .B0(mai_mai_n69_), .B1(mai_mai_n66_), .Y(mai_mai_n73_));
  INV        m0045(.A(mai_mai_n73_), .Y(mai_mai_n74_));
  INV        m0046(.A(n), .Y(mai_mai_n75_));
  NOi32      m0047(.An(e), .Bn(b), .C(d), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  INV        m0049(.A(j), .Y(mai_mai_n78_));
  AN3        m0050(.A(m), .B(k), .C(i), .Y(mai_mai_n79_));
  NA3        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(g), .Y(mai_mai_n80_));
  NO2        m0052(.A(mai_mai_n80_), .B(f), .Y(mai_mai_n81_));
  NAi32      m0053(.An(g), .Bn(f), .C(h), .Y(mai_mai_n82_));
  NAi31      m0054(.An(j), .B(m), .C(l), .Y(mai_mai_n83_));
  NO2        m0055(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  NA2        m0056(.A(m), .B(l), .Y(mai_mai_n85_));
  NO2        m0057(.A(mai_mai_n85_), .B(f), .Y(mai_mai_n86_));
  NOi32      m0058(.An(m), .Bn(l), .C(i), .Y(mai_mai_n87_));
  NOi32      m0059(.An(m), .Bn(j), .C(k), .Y(mai_mai_n88_));
  AOI220     m0060(.A0(mai_mai_n88_), .A1(g), .B0(mai_mai_n87_), .B1(g), .Y(mai_mai_n89_));
  NO2        m0061(.A(mai_mai_n89_), .B(f), .Y(mai_mai_n90_));
  NO3        m0062(.A(mai_mai_n90_), .B(mai_mai_n84_), .C(mai_mai_n81_), .Y(mai_mai_n91_));
  NAi41      m0063(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n92_));
  AN2        m0064(.A(e), .B(b), .Y(mai_mai_n93_));
  NOi31      m0065(.An(c), .B(h), .C(f), .Y(mai_mai_n94_));
  NA2        m0066(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n95_));
  NO3        m0067(.A(mai_mai_n95_), .B(mai_mai_n92_), .C(g), .Y(mai_mai_n96_));
  NOi21      m0068(.An(i), .B(h), .Y(mai_mai_n97_));
  NA3        m0069(.A(mai_mai_n97_), .B(g), .C(mai_mai_n36_), .Y(mai_mai_n98_));
  INV        m0070(.A(a), .Y(mai_mai_n99_));
  NA2        m0071(.A(mai_mai_n93_), .B(mai_mai_n99_), .Y(mai_mai_n100_));
  INV        m0072(.A(l), .Y(mai_mai_n101_));
  NOi21      m0073(.An(m), .B(n), .Y(mai_mai_n102_));
  AN2        m0074(.A(k), .B(h), .Y(mai_mai_n103_));
  NO2        m0075(.A(mai_mai_n98_), .B(mai_mai_n77_), .Y(mai_mai_n104_));
  INV        m0076(.A(b), .Y(mai_mai_n105_));
  NA2        m0077(.A(l), .B(j), .Y(mai_mai_n106_));
  AN2        m0078(.A(k), .B(i), .Y(mai_mai_n107_));
  NA2        m0079(.A(g), .B(e), .Y(mai_mai_n108_));
  NOi32      m0080(.An(c), .Bn(a), .C(d), .Y(mai_mai_n109_));
  NA2        m0081(.A(mai_mai_n109_), .B(mai_mai_n102_), .Y(mai_mai_n110_));
  NO2        m0082(.A(mai_mai_n104_), .B(mai_mai_n96_), .Y(mai_mai_n111_));
  OAI210     m0083(.A0(mai_mai_n91_), .A1(mai_mai_n77_), .B0(mai_mai_n111_), .Y(mai_mai_n112_));
  NOi31      m0084(.An(k), .B(m), .C(j), .Y(mai_mai_n113_));
  NOi31      m0085(.An(k), .B(m), .C(i), .Y(mai_mai_n114_));
  NA3        m0086(.A(mai_mai_n114_), .B(mai_mai_n71_), .C(mai_mai_n67_), .Y(mai_mai_n115_));
  INV        m0087(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NOi32      m0088(.An(f), .Bn(b), .C(e), .Y(mai_mai_n117_));
  NAi21      m0089(.An(g), .B(h), .Y(mai_mai_n118_));
  NAi21      m0090(.An(m), .B(n), .Y(mai_mai_n119_));
  NAi21      m0091(.An(j), .B(k), .Y(mai_mai_n120_));
  NO3        m0092(.A(mai_mai_n120_), .B(mai_mai_n119_), .C(mai_mai_n118_), .Y(mai_mai_n121_));
  NAi41      m0093(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n122_));
  NAi31      m0094(.An(j), .B(k), .C(h), .Y(mai_mai_n123_));
  NO3        m0095(.A(mai_mai_n123_), .B(mai_mai_n122_), .C(mai_mai_n119_), .Y(mai_mai_n124_));
  AOI210     m0096(.A0(mai_mai_n121_), .A1(mai_mai_n117_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  NO2        m0097(.A(k), .B(j), .Y(mai_mai_n126_));
  NO2        m0098(.A(mai_mai_n126_), .B(mai_mai_n119_), .Y(mai_mai_n127_));
  AN2        m0099(.A(k), .B(j), .Y(mai_mai_n128_));
  NAi21      m0100(.An(c), .B(b), .Y(mai_mai_n129_));
  NA2        m0101(.A(f), .B(d), .Y(mai_mai_n130_));
  NO4        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(mai_mai_n128_), .D(mai_mai_n118_), .Y(mai_mai_n131_));
  NA2        m0103(.A(h), .B(c), .Y(mai_mai_n132_));
  NAi31      m0104(.An(f), .B(e), .C(b), .Y(mai_mai_n133_));
  NA2        m0105(.A(mai_mai_n131_), .B(mai_mai_n127_), .Y(mai_mai_n134_));
  NA2        m0106(.A(d), .B(b), .Y(mai_mai_n135_));
  NAi21      m0107(.An(e), .B(f), .Y(mai_mai_n136_));
  NO2        m0108(.A(mai_mai_n136_), .B(mai_mai_n135_), .Y(mai_mai_n137_));
  NA2        m0109(.A(b), .B(a), .Y(mai_mai_n138_));
  NAi21      m0110(.An(c), .B(d), .Y(mai_mai_n139_));
  NAi31      m0111(.An(l), .B(k), .C(h), .Y(mai_mai_n140_));
  NO2        m0112(.A(mai_mai_n119_), .B(mai_mai_n140_), .Y(mai_mai_n141_));
  NA2        m0113(.A(mai_mai_n141_), .B(mai_mai_n137_), .Y(mai_mai_n142_));
  NAi41      m0114(.An(mai_mai_n116_), .B(mai_mai_n142_), .C(mai_mai_n134_), .D(mai_mai_n125_), .Y(mai_mai_n143_));
  NAi31      m0115(.An(e), .B(f), .C(b), .Y(mai_mai_n144_));
  NOi21      m0116(.An(g), .B(d), .Y(mai_mai_n145_));
  NO2        m0117(.A(mai_mai_n145_), .B(mai_mai_n144_), .Y(mai_mai_n146_));
  NOi21      m0118(.An(h), .B(i), .Y(mai_mai_n147_));
  NOi21      m0119(.An(k), .B(m), .Y(mai_mai_n148_));
  NA3        m0120(.A(mai_mai_n148_), .B(mai_mai_n147_), .C(n), .Y(mai_mai_n149_));
  NOi21      m0121(.An(mai_mai_n146_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  NO2        m0122(.A(mai_mai_n130_), .B(mai_mai_n129_), .Y(mai_mai_n151_));
  NA2        m0123(.A(mai_mai_n151_), .B(h), .Y(mai_mai_n152_));
  NOi32      m0124(.An(n), .Bn(k), .C(m), .Y(mai_mai_n153_));
  NA2        m0125(.A(l), .B(i), .Y(mai_mai_n154_));
  NA2        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  NO2        m0127(.A(mai_mai_n155_), .B(mai_mai_n152_), .Y(mai_mai_n156_));
  NAi31      m0128(.An(d), .B(f), .C(c), .Y(mai_mai_n157_));
  NAi31      m0129(.An(e), .B(f), .C(c), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NA2        m0131(.A(j), .B(h), .Y(mai_mai_n160_));
  OR3        m0132(.A(n), .B(m), .C(k), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NAi32      m0134(.An(m), .Bn(k), .C(n), .Y(mai_mai_n163_));
  NO2        m0135(.A(mai_mai_n163_), .B(mai_mai_n160_), .Y(mai_mai_n164_));
  AOI220     m0136(.A0(mai_mai_n164_), .A1(mai_mai_n146_), .B0(mai_mai_n162_), .B1(mai_mai_n159_), .Y(mai_mai_n165_));
  NO2        m0137(.A(n), .B(m), .Y(mai_mai_n166_));
  NA2        m0138(.A(mai_mai_n166_), .B(mai_mai_n47_), .Y(mai_mai_n167_));
  NAi21      m0139(.An(f), .B(e), .Y(mai_mai_n168_));
  NA2        m0140(.A(d), .B(c), .Y(mai_mai_n169_));
  NAi31      m0141(.An(m), .B(n), .C(b), .Y(mai_mai_n170_));
  NAi21      m0142(.An(h), .B(f), .Y(mai_mai_n171_));
  NO2        m0143(.A(mai_mai_n170_), .B(mai_mai_n139_), .Y(mai_mai_n172_));
  NOi32      m0144(.An(f), .Bn(c), .C(d), .Y(mai_mai_n173_));
  NOi32      m0145(.An(f), .Bn(c), .C(e), .Y(mai_mai_n174_));
  NO2        m0146(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NO3        m0147(.A(n), .B(m), .C(j), .Y(mai_mai_n176_));
  NA2        m0148(.A(mai_mai_n176_), .B(mai_mai_n103_), .Y(mai_mai_n177_));
  AO210      m0149(.A0(mai_mai_n177_), .A1(mai_mai_n167_), .B0(mai_mai_n175_), .Y(mai_mai_n178_));
  NA2        m0150(.A(mai_mai_n178_), .B(mai_mai_n165_), .Y(mai_mai_n179_));
  OR4        m0151(.A(mai_mai_n179_), .B(mai_mai_n156_), .C(mai_mai_n150_), .D(mai_mai_n143_), .Y(mai_mai_n180_));
  NO4        m0152(.A(mai_mai_n180_), .B(mai_mai_n112_), .C(mai_mai_n74_), .D(mai_mai_n51_), .Y(mai_mai_n181_));
  NA3        m0153(.A(m), .B(mai_mai_n101_), .C(j), .Y(mai_mai_n182_));
  NAi31      m0154(.An(n), .B(h), .C(g), .Y(mai_mai_n183_));
  NO2        m0155(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  NOi32      m0156(.An(m), .Bn(k), .C(l), .Y(mai_mai_n185_));
  NA3        m0157(.A(mai_mai_n185_), .B(mai_mai_n78_), .C(g), .Y(mai_mai_n186_));
  NA3        m0158(.A(mai_mai_n102_), .B(i), .C(g), .Y(mai_mai_n187_));
  AN2        m0159(.A(i), .B(g), .Y(mai_mai_n188_));
  NA3        m0160(.A(mai_mai_n65_), .B(mai_mai_n188_), .C(mai_mai_n102_), .Y(mai_mai_n189_));
  NAi41      m0161(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n190_));
  INV        m0162(.A(mai_mai_n190_), .Y(mai_mai_n191_));
  INV        m0163(.A(f), .Y(mai_mai_n192_));
  INV        m0164(.A(g), .Y(mai_mai_n193_));
  NOi31      m0165(.An(i), .B(j), .C(h), .Y(mai_mai_n194_));
  NOi21      m0166(.An(l), .B(m), .Y(mai_mai_n195_));
  NA2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NO3        m0168(.A(mai_mai_n196_), .B(mai_mai_n193_), .C(mai_mai_n192_), .Y(mai_mai_n197_));
  NA2        m0169(.A(mai_mai_n197_), .B(mai_mai_n191_), .Y(mai_mai_n198_));
  INV        m0170(.A(mai_mai_n198_), .Y(mai_mai_n199_));
  NOi21      m0171(.An(n), .B(m), .Y(mai_mai_n200_));
  NOi32      m0172(.An(l), .Bn(i), .C(j), .Y(mai_mai_n201_));
  NA2        m0173(.A(mai_mai_n201_), .B(mai_mai_n200_), .Y(mai_mai_n202_));
  OA220      m0174(.A0(mai_mai_n202_), .A1(mai_mai_n95_), .B0(mai_mai_n70_), .B1(mai_mai_n69_), .Y(mai_mai_n203_));
  NAi21      m0175(.An(j), .B(h), .Y(mai_mai_n204_));
  XN2        m0176(.A(i), .B(h), .Y(mai_mai_n205_));
  NA2        m0177(.A(mai_mai_n205_), .B(mai_mai_n204_), .Y(mai_mai_n206_));
  NOi31      m0178(.An(k), .B(n), .C(m), .Y(mai_mai_n207_));
  NOi31      m0179(.An(mai_mai_n207_), .B(mai_mai_n169_), .C(mai_mai_n168_), .Y(mai_mai_n208_));
  NA2        m0180(.A(mai_mai_n208_), .B(mai_mai_n206_), .Y(mai_mai_n209_));
  NAi31      m0181(.An(f), .B(e), .C(c), .Y(mai_mai_n210_));
  NO4        m0182(.A(mai_mai_n210_), .B(mai_mai_n161_), .C(mai_mai_n160_), .D(mai_mai_n55_), .Y(mai_mai_n211_));
  NA4        m0183(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n212_));
  NAi32      m0184(.An(m), .Bn(i), .C(k), .Y(mai_mai_n213_));
  NO3        m0185(.A(mai_mai_n213_), .B(mai_mai_n82_), .C(mai_mai_n212_), .Y(mai_mai_n214_));
  INV        m0186(.A(k), .Y(mai_mai_n215_));
  NO2        m0187(.A(mai_mai_n214_), .B(mai_mai_n211_), .Y(mai_mai_n216_));
  NAi21      m0188(.An(n), .B(a), .Y(mai_mai_n217_));
  NO2        m0189(.A(mai_mai_n217_), .B(mai_mai_n135_), .Y(mai_mai_n218_));
  NAi41      m0190(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n219_));
  NO2        m0191(.A(mai_mai_n219_), .B(e), .Y(mai_mai_n220_));
  NA2        m0192(.A(mai_mai_n220_), .B(mai_mai_n218_), .Y(mai_mai_n221_));
  AN4        m0193(.A(mai_mai_n221_), .B(mai_mai_n216_), .C(mai_mai_n209_), .D(mai_mai_n203_), .Y(mai_mai_n222_));
  NAi41      m0194(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n223_));
  NO2        m0195(.A(mai_mai_n223_), .B(mai_mai_n192_), .Y(mai_mai_n224_));
  NA2        m0196(.A(mai_mai_n148_), .B(mai_mai_n97_), .Y(mai_mai_n225_));
  NAi21      m0197(.An(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  NO2        m0198(.A(n), .B(a), .Y(mai_mai_n227_));
  NAi21      m0199(.An(h), .B(i), .Y(mai_mai_n228_));
  NA2        m0200(.A(mai_mai_n166_), .B(k), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n230_), .B(mai_mai_n173_), .Y(mai_mai_n231_));
  NA2        m0203(.A(mai_mai_n231_), .B(mai_mai_n226_), .Y(mai_mai_n232_));
  NO2        m0204(.A(mai_mai_n63_), .B(mai_mai_n64_), .Y(mai_mai_n233_));
  NAi21      m0205(.An(f), .B(g), .Y(mai_mai_n234_));
  NO2        m0206(.A(mai_mai_n60_), .B(mai_mai_n106_), .Y(mai_mai_n235_));
  NO2        m0207(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n236_));
  NOi31      m0208(.An(mai_mai_n222_), .B(mai_mai_n232_), .C(mai_mai_n199_), .Y(mai_mai_n237_));
  NO3        m0209(.A(mai_mai_n184_), .B(mai_mai_n42_), .C(mai_mai_n39_), .Y(mai_mai_n238_));
  NO2        m0210(.A(mai_mai_n238_), .B(mai_mai_n100_), .Y(mai_mai_n239_));
  NAi21      m0211(.An(h), .B(g), .Y(mai_mai_n240_));
  OR4        m0212(.A(mai_mai_n240_), .B(mai_mai_n1225_), .C(mai_mai_n202_), .D(e), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n225_), .B(mai_mai_n234_), .Y(mai_mai_n242_));
  NA2        m0214(.A(mai_mai_n242_), .B(mai_mai_n67_), .Y(mai_mai_n243_));
  NAi31      m0215(.An(e), .B(d), .C(a), .Y(mai_mai_n244_));
  NA2        m0216(.A(mai_mai_n243_), .B(mai_mai_n241_), .Y(mai_mai_n245_));
  NA4        m0217(.A(mai_mai_n148_), .B(mai_mai_n71_), .C(mai_mai_n67_), .D(mai_mai_n106_), .Y(mai_mai_n246_));
  NA3        m0218(.A(mai_mai_n148_), .B(mai_mai_n147_), .C(mai_mai_n75_), .Y(mai_mai_n247_));
  NO2        m0219(.A(mai_mai_n247_), .B(mai_mai_n175_), .Y(mai_mai_n248_));
  NOi21      m0220(.An(mai_mai_n246_), .B(mai_mai_n248_), .Y(mai_mai_n249_));
  NA3        m0221(.A(e), .B(c), .C(b), .Y(mai_mai_n250_));
  NO2        m0222(.A(mai_mai_n56_), .B(mai_mai_n250_), .Y(mai_mai_n251_));
  INV        m0223(.A(mai_mai_n46_), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n251_), .B(mai_mai_n252_), .Y(mai_mai_n253_));
  NOi21      m0225(.An(l), .B(j), .Y(mai_mai_n254_));
  NA2        m0226(.A(h), .B(mai_mai_n254_), .Y(mai_mai_n255_));
  OR3        m0227(.A(mai_mai_n63_), .B(mai_mai_n64_), .C(e), .Y(mai_mai_n256_));
  AOI210     m0228(.A0(mai_mai_n1224_), .A1(mai_mai_n255_), .B0(mai_mai_n256_), .Y(mai_mai_n257_));
  INV        m0229(.A(mai_mai_n257_), .Y(mai_mai_n258_));
  NAi32      m0230(.An(j), .Bn(h), .C(i), .Y(mai_mai_n259_));
  NAi21      m0231(.An(m), .B(l), .Y(mai_mai_n260_));
  NO3        m0232(.A(mai_mai_n260_), .B(mai_mai_n259_), .C(mai_mai_n75_), .Y(mai_mai_n261_));
  NA2        m0233(.A(h), .B(g), .Y(mai_mai_n262_));
  INV        m0234(.A(mai_mai_n153_), .Y(mai_mai_n263_));
  NA2        m0235(.A(mai_mai_n261_), .B(mai_mai_n151_), .Y(mai_mai_n264_));
  NA4        m0236(.A(mai_mai_n264_), .B(mai_mai_n258_), .C(mai_mai_n253_), .D(mai_mai_n249_), .Y(mai_mai_n265_));
  NO2        m0237(.A(mai_mai_n133_), .B(d), .Y(mai_mai_n266_));
  NA2        m0238(.A(mai_mai_n266_), .B(mai_mai_n50_), .Y(mai_mai_n267_));
  NO2        m0239(.A(mai_mai_n95_), .B(mai_mai_n92_), .Y(mai_mai_n268_));
  NAi32      m0240(.An(n), .Bn(m), .C(l), .Y(mai_mai_n269_));
  NO2        m0241(.A(mai_mai_n110_), .B(mai_mai_n105_), .Y(mai_mai_n270_));
  NAi31      m0242(.An(k), .B(l), .C(j), .Y(mai_mai_n271_));
  INV        m0243(.A(mai_mai_n271_), .Y(mai_mai_n272_));
  INV        m0244(.A(mai_mai_n267_), .Y(mai_mai_n273_));
  NO4        m0245(.A(mai_mai_n273_), .B(mai_mai_n265_), .C(mai_mai_n245_), .D(mai_mai_n239_), .Y(mai_mai_n274_));
  NA2        m0246(.A(mai_mai_n230_), .B(mai_mai_n174_), .Y(mai_mai_n275_));
  NAi21      m0247(.An(m), .B(k), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n205_), .B(mai_mai_n276_), .Y(mai_mai_n277_));
  NAi41      m0249(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n278_));
  NA2        m0250(.A(e), .B(c), .Y(mai_mai_n279_));
  NO3        m0251(.A(mai_mai_n279_), .B(n), .C(d), .Y(mai_mai_n280_));
  NA2        m0252(.A(f), .B(mai_mai_n107_), .Y(mai_mai_n281_));
  NO2        m0253(.A(mai_mai_n281_), .B(mai_mai_n193_), .Y(mai_mai_n282_));
  NAi31      m0254(.An(d), .B(e), .C(b), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n119_), .B(mai_mai_n283_), .Y(mai_mai_n284_));
  NA2        m0256(.A(mai_mai_n284_), .B(mai_mai_n282_), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n285_), .B(mai_mai_n275_), .Y(mai_mai_n286_));
  NO4        m0258(.A(mai_mai_n278_), .B(mai_mai_n70_), .C(mai_mai_n62_), .D(mai_mai_n193_), .Y(mai_mai_n287_));
  NA2        m0259(.A(mai_mai_n227_), .B(mai_mai_n93_), .Y(mai_mai_n288_));
  OR2        m0260(.A(mai_mai_n288_), .B(mai_mai_n186_), .Y(mai_mai_n289_));
  NOi31      m0261(.An(l), .B(n), .C(m), .Y(mai_mai_n290_));
  NAi21      m0262(.An(mai_mai_n287_), .B(mai_mai_n289_), .Y(mai_mai_n291_));
  NAi32      m0263(.An(m), .Bn(j), .C(k), .Y(mai_mai_n292_));
  NAi41      m0264(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n293_));
  NOi31      m0265(.An(j), .B(m), .C(k), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n113_), .B(mai_mai_n294_), .Y(mai_mai_n295_));
  AN3        m0267(.A(h), .B(g), .C(f), .Y(mai_mai_n296_));
  NOi32      m0268(.An(m), .Bn(j), .C(l), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n260_), .B(mai_mai_n259_), .Y(mai_mai_n298_));
  NO2        m0270(.A(mai_mai_n196_), .B(g), .Y(mai_mai_n299_));
  NO2        m0271(.A(mai_mai_n144_), .B(mai_mai_n75_), .Y(mai_mai_n300_));
  AOI220     m0272(.A0(mai_mai_n300_), .A1(mai_mai_n299_), .B0(mai_mai_n224_), .B1(mai_mai_n298_), .Y(mai_mai_n301_));
  NA3        m0273(.A(mai_mai_n1231_), .B(mai_mai_n296_), .C(mai_mai_n191_), .Y(mai_mai_n302_));
  NA2        m0274(.A(mai_mai_n302_), .B(mai_mai_n301_), .Y(mai_mai_n303_));
  NA3        m0275(.A(h), .B(g), .C(f), .Y(mai_mai_n304_));
  NA2        m0276(.A(h), .B(e), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n305_), .B(mai_mai_n41_), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n306_), .B(mai_mai_n270_), .Y(mai_mai_n307_));
  NOi32      m0279(.An(j), .Bn(g), .C(i), .Y(mai_mai_n308_));
  NA2        m0280(.A(mai_mai_n308_), .B(mai_mai_n102_), .Y(mai_mai_n309_));
  OR2        m0281(.A(mai_mai_n100_), .B(mai_mai_n309_), .Y(mai_mai_n310_));
  NOi32      m0282(.An(e), .Bn(b), .C(a), .Y(mai_mai_n311_));
  INV        m0283(.A(mai_mai_n276_), .Y(mai_mai_n312_));
  NO3        m0284(.A(mai_mai_n278_), .B(mai_mai_n62_), .C(mai_mai_n193_), .Y(mai_mai_n313_));
  NA2        m0285(.A(mai_mai_n189_), .B(mai_mai_n35_), .Y(mai_mai_n314_));
  AOI220     m0286(.A0(mai_mai_n314_), .A1(mai_mai_n311_), .B0(mai_mai_n313_), .B1(mai_mai_n312_), .Y(mai_mai_n315_));
  NO2        m0287(.A(mai_mai_n283_), .B(n), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n188_), .B(k), .Y(mai_mai_n317_));
  NA3        m0289(.A(m), .B(mai_mai_n101_), .C(mai_mai_n192_), .Y(mai_mai_n318_));
  NA4        m0290(.A(mai_mai_n185_), .B(mai_mai_n78_), .C(g), .D(mai_mai_n192_), .Y(mai_mai_n319_));
  NAi41      m0291(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n48_), .B(mai_mai_n102_), .Y(mai_mai_n321_));
  NO2        m0293(.A(mai_mai_n321_), .B(mai_mai_n320_), .Y(mai_mai_n322_));
  AOI220     m0294(.A0(mai_mai_n322_), .A1(b), .B0(mai_mai_n185_), .B1(mai_mai_n316_), .Y(mai_mai_n323_));
  NA4        m0295(.A(mai_mai_n323_), .B(mai_mai_n315_), .C(mai_mai_n310_), .D(mai_mai_n307_), .Y(mai_mai_n324_));
  NO4        m0296(.A(mai_mai_n324_), .B(mai_mai_n303_), .C(mai_mai_n291_), .D(mai_mai_n286_), .Y(mai_mai_n325_));
  NA4        m0297(.A(mai_mai_n325_), .B(mai_mai_n274_), .C(mai_mai_n237_), .D(mai_mai_n181_), .Y(mai10));
  NA3        m0298(.A(m), .B(k), .C(i), .Y(mai_mai_n327_));
  NO3        m0299(.A(mai_mai_n327_), .B(j), .C(mai_mai_n193_), .Y(mai_mai_n328_));
  NOi21      m0300(.An(e), .B(f), .Y(mai_mai_n329_));
  NO4        m0301(.A(mai_mai_n139_), .B(mai_mai_n329_), .C(n), .D(mai_mai_n99_), .Y(mai_mai_n330_));
  NAi31      m0302(.An(b), .B(f), .C(c), .Y(mai_mai_n331_));
  INV        m0303(.A(mai_mai_n331_), .Y(mai_mai_n332_));
  NOi32      m0304(.An(k), .Bn(h), .C(j), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n333_), .B(mai_mai_n200_), .Y(mai_mai_n334_));
  NA2        m0306(.A(mai_mai_n149_), .B(mai_mai_n334_), .Y(mai_mai_n335_));
  NA2        m0307(.A(mai_mai_n335_), .B(mai_mai_n332_), .Y(mai_mai_n336_));
  AN2        m0308(.A(j), .B(h), .Y(mai_mai_n337_));
  NO3        m0309(.A(n), .B(m), .C(k), .Y(mai_mai_n338_));
  NA2        m0310(.A(mai_mai_n338_), .B(mai_mai_n337_), .Y(mai_mai_n339_));
  NO3        m0311(.A(mai_mai_n339_), .B(mai_mai_n139_), .C(mai_mai_n192_), .Y(mai_mai_n340_));
  OR2        m0312(.A(m), .B(k), .Y(mai_mai_n341_));
  NO2        m0313(.A(mai_mai_n160_), .B(mai_mai_n341_), .Y(mai_mai_n342_));
  NA4        m0314(.A(n), .B(f), .C(c), .D(mai_mai_n105_), .Y(mai_mai_n343_));
  NOi21      m0315(.An(mai_mai_n342_), .B(mai_mai_n343_), .Y(mai_mai_n344_));
  NOi32      m0316(.An(d), .Bn(a), .C(c), .Y(mai_mai_n345_));
  NA2        m0317(.A(mai_mai_n345_), .B(mai_mai_n168_), .Y(mai_mai_n346_));
  NAi31      m0318(.An(k), .B(m), .C(j), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n344_), .B(mai_mai_n340_), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n343_), .B(mai_mai_n260_), .Y(mai_mai_n349_));
  NOi32      m0321(.An(f), .Bn(d), .C(c), .Y(mai_mai_n350_));
  NA2        m0322(.A(mai_mai_n348_), .B(mai_mai_n336_), .Y(mai_mai_n351_));
  NO2        m0323(.A(mai_mai_n55_), .B(mai_mai_n105_), .Y(mai_mai_n352_));
  NA2        m0324(.A(mai_mai_n227_), .B(mai_mai_n352_), .Y(mai_mai_n353_));
  INV        m0325(.A(e), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n44_), .B(e), .Y(mai_mai_n355_));
  OAI220     m0327(.A0(mai_mai_n355_), .A1(mai_mai_n182_), .B0(mai_mai_n186_), .B1(mai_mai_n354_), .Y(mai_mai_n356_));
  INV        m0328(.A(mai_mai_n356_), .Y(mai_mai_n357_));
  NA3        m0329(.A(e), .B(mai_mai_n254_), .C(m), .Y(mai_mai_n358_));
  NOi21      m0330(.An(g), .B(h), .Y(mai_mai_n359_));
  NA3        m0331(.A(m), .B(mai_mai_n359_), .C(e), .Y(mai_mai_n360_));
  AN3        m0332(.A(h), .B(g), .C(e), .Y(mai_mai_n361_));
  AN2        m0333(.A(mai_mai_n360_), .B(mai_mai_n358_), .Y(mai_mai_n362_));
  AOI210     m0334(.A0(mai_mai_n362_), .A1(mai_mai_n357_), .B0(mai_mai_n353_), .Y(mai_mai_n363_));
  NA3        m0335(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n364_));
  NA3        m0336(.A(mai_mai_n345_), .B(mai_mai_n168_), .C(mai_mai_n75_), .Y(mai_mai_n365_));
  NAi31      m0337(.An(b), .B(c), .C(a), .Y(mai_mai_n366_));
  NO2        m0338(.A(mai_mai_n366_), .B(n), .Y(mai_mai_n367_));
  OAI210     m0339(.A0(mai_mai_n48_), .A1(mai_mai_n47_), .B0(m), .Y(mai_mai_n368_));
  NO2        m0340(.A(mai_mai_n363_), .B(mai_mai_n351_), .Y(mai_mai_n369_));
  NA2        m0341(.A(i), .B(g), .Y(mai_mai_n370_));
  NO2        m0342(.A(mai_mai_n244_), .B(c), .Y(mai_mai_n371_));
  NOi21      m0343(.An(a), .B(n), .Y(mai_mai_n372_));
  NA2        m0344(.A(d), .B(mai_mai_n372_), .Y(mai_mai_n373_));
  NA3        m0345(.A(i), .B(g), .C(f), .Y(mai_mai_n374_));
  OR2        m0346(.A(mai_mai_n374_), .B(mai_mai_n61_), .Y(mai_mai_n375_));
  NA3        m0347(.A(m), .B(mai_mai_n359_), .C(mai_mai_n168_), .Y(mai_mai_n376_));
  AOI210     m0348(.A0(mai_mai_n376_), .A1(mai_mai_n375_), .B0(mai_mai_n373_), .Y(mai_mai_n377_));
  INV        m0349(.A(mai_mai_n377_), .Y(mai_mai_n378_));
  OR2        m0350(.A(n), .B(m), .Y(mai_mai_n379_));
  NO2        m0351(.A(mai_mai_n379_), .B(mai_mai_n140_), .Y(mai_mai_n380_));
  NO2        m0352(.A(mai_mai_n169_), .B(mai_mai_n136_), .Y(mai_mai_n381_));
  OAI210     m0353(.A0(mai_mai_n380_), .A1(mai_mai_n162_), .B0(mai_mai_n381_), .Y(mai_mai_n382_));
  NO2        m0354(.A(mai_mai_n366_), .B(mai_mai_n46_), .Y(mai_mai_n383_));
  NAi21      m0355(.An(k), .B(j), .Y(mai_mai_n384_));
  NAi21      m0356(.An(e), .B(d), .Y(mai_mai_n385_));
  INV        m0357(.A(mai_mai_n385_), .Y(mai_mai_n386_));
  NO2        m0358(.A(mai_mai_n229_), .B(mai_mai_n192_), .Y(mai_mai_n387_));
  NA3        m0359(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(mai_mai_n206_), .Y(mai_mai_n388_));
  NA2        m0360(.A(mai_mai_n388_), .B(mai_mai_n382_), .Y(mai_mai_n389_));
  NOi31      m0361(.An(n), .B(m), .C(k), .Y(mai_mai_n390_));
  AOI220     m0362(.A0(mai_mai_n390_), .A1(mai_mai_n337_), .B0(mai_mai_n200_), .B1(mai_mai_n47_), .Y(mai_mai_n391_));
  NOi21      m0363(.An(mai_mai_n378_), .B(mai_mai_n389_), .Y(mai_mai_n392_));
  NOi32      m0364(.An(c), .Bn(a), .C(b), .Y(mai_mai_n393_));
  NA2        m0365(.A(mai_mai_n393_), .B(mai_mai_n102_), .Y(mai_mai_n394_));
  AN2        m0366(.A(e), .B(d), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n118_), .B(mai_mai_n41_), .Y(mai_mai_n396_));
  NO2        m0368(.A(mai_mai_n136_), .B(mai_mai_n394_), .Y(mai_mai_n397_));
  NOi21      m0369(.An(a), .B(b), .Y(mai_mai_n398_));
  NA3        m0370(.A(e), .B(d), .C(c), .Y(mai_mai_n399_));
  NAi21      m0371(.An(mai_mai_n399_), .B(mai_mai_n398_), .Y(mai_mai_n400_));
  NO2        m0372(.A(mai_mai_n365_), .B(mai_mai_n186_), .Y(mai_mai_n401_));
  NOi21      m0373(.An(mai_mai_n400_), .B(mai_mai_n401_), .Y(mai_mai_n402_));
  NO2        m0374(.A(mai_mai_n1229_), .B(mai_mai_n402_), .Y(mai_mai_n403_));
  NO4        m0375(.A(mai_mai_n171_), .B(mai_mai_n92_), .C(mai_mai_n52_), .D(b), .Y(mai_mai_n404_));
  NA2        m0376(.A(mai_mai_n332_), .B(mai_mai_n141_), .Y(mai_mai_n405_));
  OR2        m0377(.A(k), .B(j), .Y(mai_mai_n406_));
  NA2        m0378(.A(l), .B(k), .Y(mai_mai_n407_));
  NA3        m0379(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(mai_mai_n200_), .Y(mai_mai_n408_));
  AOI210     m0380(.A0(mai_mai_n213_), .A1(mai_mai_n292_), .B0(mai_mai_n75_), .Y(mai_mai_n409_));
  NOi21      m0381(.An(mai_mai_n408_), .B(mai_mai_n409_), .Y(mai_mai_n410_));
  OR3        m0382(.A(mai_mai_n410_), .B(mai_mai_n132_), .C(mai_mai_n122_), .Y(mai_mai_n411_));
  NA2        m0383(.A(mai_mai_n246_), .B(mai_mai_n115_), .Y(mai_mai_n412_));
  NO3        m0384(.A(mai_mai_n365_), .B(mai_mai_n83_), .C(mai_mai_n118_), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n413_), .B(mai_mai_n412_), .Y(mai_mai_n414_));
  NA3        m0386(.A(mai_mai_n414_), .B(mai_mai_n411_), .C(mai_mai_n405_), .Y(mai_mai_n415_));
  NO4        m0387(.A(mai_mai_n415_), .B(mai_mai_n404_), .C(mai_mai_n403_), .D(mai_mai_n397_), .Y(mai_mai_n416_));
  NOi21      m0388(.An(d), .B(e), .Y(mai_mai_n417_));
  NO2        m0389(.A(mai_mai_n171_), .B(mai_mai_n52_), .Y(mai_mai_n418_));
  NAi31      m0390(.An(j), .B(l), .C(i), .Y(mai_mai_n419_));
  OAI210     m0391(.A0(mai_mai_n419_), .A1(mai_mai_n119_), .B0(mai_mai_n92_), .Y(mai_mai_n420_));
  NA3        m0392(.A(mai_mai_n420_), .B(mai_mai_n418_), .C(mai_mai_n417_), .Y(mai_mai_n421_));
  NO2        m0393(.A(mai_mai_n346_), .B(mai_mai_n183_), .Y(mai_mai_n422_));
  NO2        m0394(.A(mai_mai_n346_), .B(mai_mai_n321_), .Y(mai_mai_n423_));
  NO3        m0395(.A(mai_mai_n423_), .B(mai_mai_n422_), .C(mai_mai_n268_), .Y(mai_mai_n424_));
  NA3        m0396(.A(mai_mai_n424_), .B(mai_mai_n421_), .C(mai_mai_n222_), .Y(mai_mai_n425_));
  NO2        m0397(.A(mai_mai_n114_), .B(mai_mai_n113_), .Y(mai_mai_n426_));
  NO2        m0398(.A(mai_mai_n426_), .B(mai_mai_n118_), .Y(mai_mai_n427_));
  XO2        m0399(.A(i), .B(h), .Y(mai_mai_n428_));
  NAi31      m0400(.An(c), .B(f), .C(d), .Y(mai_mai_n429_));
  AOI210     m0401(.A0(mai_mai_n247_), .A1(mai_mai_n177_), .B0(mai_mai_n429_), .Y(mai_mai_n430_));
  NOi21      m0402(.An(mai_mai_n73_), .B(mai_mai_n430_), .Y(mai_mai_n431_));
  NA3        m0403(.A(mai_mai_n330_), .B(mai_mai_n87_), .C(g), .Y(mai_mai_n432_));
  NA2        m0404(.A(mai_mai_n207_), .B(mai_mai_n97_), .Y(mai_mai_n433_));
  AOI210     m0405(.A0(mai_mai_n433_), .A1(mai_mai_n167_), .B0(mai_mai_n429_), .Y(mai_mai_n434_));
  NOi21      m0406(.An(mai_mai_n432_), .B(mai_mai_n434_), .Y(mai_mai_n435_));
  NA3        m0407(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n436_));
  NO2        m0408(.A(mai_mai_n436_), .B(mai_mai_n373_), .Y(mai_mai_n437_));
  INV        m0409(.A(mai_mai_n257_), .Y(mai_mai_n438_));
  NA3        m0410(.A(mai_mai_n438_), .B(mai_mai_n435_), .C(mai_mai_n431_), .Y(mai_mai_n439_));
  NO2        m0411(.A(mai_mai_n439_), .B(mai_mai_n425_), .Y(mai_mai_n440_));
  NA4        m0412(.A(mai_mai_n440_), .B(mai_mai_n416_), .C(mai_mai_n392_), .D(mai_mai_n369_), .Y(mai11));
  NO2        m0413(.A(mai_mai_n63_), .B(f), .Y(mai_mai_n442_));
  NA2        m0414(.A(j), .B(g), .Y(mai_mai_n443_));
  NAi31      m0415(.An(i), .B(m), .C(l), .Y(mai_mai_n444_));
  NA3        m0416(.A(m), .B(k), .C(j), .Y(mai_mai_n445_));
  OAI220     m0417(.A0(mai_mai_n445_), .A1(mai_mai_n118_), .B0(mai_mai_n444_), .B1(mai_mai_n443_), .Y(mai_mai_n446_));
  NA2        m0418(.A(mai_mai_n446_), .B(mai_mai_n442_), .Y(mai_mai_n447_));
  NOi32      m0419(.An(e), .Bn(b), .C(f), .Y(mai_mai_n448_));
  NA2        m0420(.A(mai_mai_n44_), .B(j), .Y(mai_mai_n449_));
  NO2        m0421(.A(mai_mai_n449_), .B(mai_mai_n263_), .Y(mai_mai_n450_));
  NAi31      m0422(.An(d), .B(e), .C(a), .Y(mai_mai_n451_));
  NO2        m0423(.A(mai_mai_n451_), .B(n), .Y(mai_mai_n452_));
  AOI220     m0424(.A0(mai_mai_n452_), .A1(mai_mai_n90_), .B0(mai_mai_n450_), .B1(mai_mai_n448_), .Y(mai_mai_n453_));
  NAi41      m0425(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n454_));
  AN2        m0426(.A(mai_mai_n454_), .B(mai_mai_n320_), .Y(mai_mai_n455_));
  AOI210     m0427(.A0(mai_mai_n455_), .A1(mai_mai_n346_), .B0(mai_mai_n240_), .Y(mai_mai_n456_));
  NAi31      m0428(.An(n), .B(m), .C(k), .Y(mai_mai_n457_));
  INV        m0429(.A(mai_mai_n457_), .Y(mai_mai_n458_));
  NO3        m0430(.A(n), .B(d), .C(mai_mai_n105_), .Y(mai_mai_n459_));
  NO2        m0431(.A(n), .B(mai_mai_n138_), .Y(mai_mai_n460_));
  NOi32      m0432(.An(g), .Bn(f), .C(i), .Y(mai_mai_n461_));
  NA2        m0433(.A(mai_mai_n446_), .B(f), .Y(mai_mai_n462_));
  NO2        m0434(.A(mai_mai_n462_), .B(n), .Y(mai_mai_n463_));
  AOI210     m0435(.A0(mai_mai_n458_), .A1(mai_mai_n456_), .B0(mai_mai_n463_), .Y(mai_mai_n464_));
  NA2        m0436(.A(mai_mai_n128_), .B(mai_mai_n34_), .Y(mai_mai_n465_));
  NOi41      m0437(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n466_));
  AN2        m0438(.A(mai_mai_n293_), .B(mai_mai_n278_), .Y(mai_mai_n467_));
  OAI220     m0439(.A0(mai_mai_n347_), .A1(i), .B0(mai_mai_n444_), .B1(mai_mai_n443_), .Y(mai_mai_n468_));
  NAi31      m0440(.An(d), .B(c), .C(a), .Y(mai_mai_n469_));
  NO2        m0441(.A(mai_mai_n469_), .B(n), .Y(mai_mai_n470_));
  NA3        m0442(.A(mai_mai_n470_), .B(mai_mai_n468_), .C(e), .Y(mai_mai_n471_));
  NO3        m0443(.A(mai_mai_n58_), .B(mai_mai_n46_), .C(mai_mai_n193_), .Y(mai_mai_n472_));
  INV        m0444(.A(mai_mai_n210_), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n472_), .B(mai_mai_n473_), .Y(mai_mai_n474_));
  NA2        m0446(.A(mai_mai_n474_), .B(mai_mai_n471_), .Y(mai_mai_n475_));
  INV        m0447(.A(mai_mai_n367_), .Y(mai_mai_n476_));
  NA2        m0448(.A(mai_mai_n468_), .B(f), .Y(mai_mai_n477_));
  NO3        m0449(.A(mai_mai_n163_), .B(mai_mai_n160_), .C(g), .Y(mai_mai_n478_));
  NA2        m0450(.A(mai_mai_n478_), .B(mai_mai_n54_), .Y(mai_mai_n479_));
  OAI210     m0451(.A0(mai_mai_n477_), .A1(mai_mai_n476_), .B0(mai_mai_n479_), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n135_), .B(c), .Y(mai_mai_n481_));
  NA3        m0453(.A(f), .B(d), .C(b), .Y(mai_mai_n482_));
  NO4        m0454(.A(mai_mai_n482_), .B(mai_mai_n163_), .C(mai_mai_n160_), .D(g), .Y(mai_mai_n483_));
  NO3        m0455(.A(mai_mai_n483_), .B(mai_mai_n480_), .C(mai_mai_n475_), .Y(mai_mai_n484_));
  AN4        m0456(.A(mai_mai_n484_), .B(mai_mai_n464_), .C(mai_mai_n453_), .D(mai_mai_n447_), .Y(mai_mai_n485_));
  INV        m0457(.A(k), .Y(mai_mai_n486_));
  NA4        m0458(.A(mai_mai_n345_), .B(mai_mai_n359_), .C(mai_mai_n168_), .D(mai_mai_n102_), .Y(mai_mai_n487_));
  NAi32      m0459(.An(h), .Bn(f), .C(g), .Y(mai_mai_n488_));
  NAi41      m0460(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n489_));
  OAI210     m0461(.A0(mai_mai_n451_), .A1(n), .B0(mai_mai_n489_), .Y(mai_mai_n490_));
  NA2        m0462(.A(mai_mai_n490_), .B(m), .Y(mai_mai_n491_));
  NAi31      m0463(.An(h), .B(g), .C(f), .Y(mai_mai_n492_));
  OR2        m0464(.A(mai_mai_n491_), .B(mai_mai_n488_), .Y(mai_mai_n493_));
  NO3        m0465(.A(mai_mai_n488_), .B(mai_mai_n63_), .C(mai_mai_n64_), .Y(mai_mai_n494_));
  NO4        m0466(.A(mai_mai_n492_), .B(n), .C(mai_mai_n138_), .D(mai_mai_n64_), .Y(mai_mai_n495_));
  OR2        m0467(.A(mai_mai_n495_), .B(mai_mai_n494_), .Y(mai_mai_n496_));
  NAi31      m0468(.An(mai_mai_n496_), .B(mai_mai_n493_), .C(mai_mai_n487_), .Y(mai_mai_n497_));
  NAi31      m0469(.An(f), .B(h), .C(g), .Y(mai_mai_n498_));
  NOi41      m0470(.An(b), .B(mai_mai_n304_), .C(mai_mai_n60_), .D(mai_mai_n106_), .Y(mai_mai_n499_));
  NOi32      m0471(.An(d), .Bn(a), .C(e), .Y(mai_mai_n500_));
  NO2        m0472(.A(n), .B(c), .Y(mai_mai_n501_));
  NA2        m0473(.A(mai_mai_n501_), .B(m), .Y(mai_mai_n502_));
  NOi32      m0474(.An(e), .Bn(a), .C(d), .Y(mai_mai_n503_));
  AOI210     m0475(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n503_), .Y(mai_mai_n504_));
  AOI210     m0476(.A0(mai_mai_n504_), .A1(mai_mai_n192_), .B0(mai_mai_n465_), .Y(mai_mai_n505_));
  AOI210     m0477(.A0(mai_mai_n505_), .A1(mai_mai_n102_), .B0(mai_mai_n499_), .Y(mai_mai_n506_));
  INV        m0478(.A(mai_mai_n506_), .Y(mai_mai_n507_));
  AOI210     m0479(.A0(mai_mai_n497_), .A1(mai_mai_n486_), .B0(mai_mai_n507_), .Y(mai_mai_n508_));
  NO3        m0480(.A(mai_mai_n276_), .B(mai_mai_n57_), .C(n), .Y(mai_mai_n509_));
  NA3        m0481(.A(mai_mai_n429_), .B(mai_mai_n158_), .C(mai_mai_n157_), .Y(mai_mai_n510_));
  INV        m0482(.A(mai_mai_n210_), .Y(mai_mai_n511_));
  OR2        m0483(.A(mai_mai_n511_), .B(mai_mai_n510_), .Y(mai_mai_n512_));
  NA2        m0484(.A(mai_mai_n65_), .B(mai_mai_n102_), .Y(mai_mai_n513_));
  NA2        m0485(.A(mai_mai_n512_), .B(mai_mai_n509_), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n514_), .B(mai_mai_n78_), .Y(mai_mai_n515_));
  NOi32      m0487(.An(e), .Bn(c), .C(f), .Y(mai_mai_n516_));
  NOi21      m0488(.An(f), .B(g), .Y(mai_mai_n517_));
  NO2        m0489(.A(mai_mai_n517_), .B(mai_mai_n190_), .Y(mai_mai_n518_));
  AOI220     m0490(.A0(mai_mai_n518_), .A1(mai_mai_n342_), .B0(mai_mai_n516_), .B1(mai_mai_n162_), .Y(mai_mai_n519_));
  NA2        m0491(.A(mai_mai_n519_), .B(mai_mai_n165_), .Y(mai_mai_n520_));
  AOI210     m0492(.A0(mai_mai_n455_), .A1(mai_mai_n346_), .B0(mai_mai_n262_), .Y(mai_mai_n521_));
  NA2        m0493(.A(mai_mai_n521_), .B(mai_mai_n235_), .Y(mai_mai_n522_));
  NOi21      m0494(.An(j), .B(l), .Y(mai_mai_n523_));
  NAi21      m0495(.An(k), .B(h), .Y(mai_mai_n524_));
  NO2        m0496(.A(mai_mai_n524_), .B(mai_mai_n234_), .Y(mai_mai_n525_));
  INV        m0497(.A(mai_mai_n525_), .Y(mai_mai_n526_));
  OR2        m0498(.A(mai_mai_n526_), .B(mai_mai_n491_), .Y(mai_mai_n527_));
  NOi31      m0499(.An(m), .B(n), .C(k), .Y(mai_mai_n528_));
  NA2        m0500(.A(mai_mai_n523_), .B(mai_mai_n528_), .Y(mai_mai_n529_));
  NO2        m0501(.A(mai_mai_n346_), .B(mai_mai_n262_), .Y(mai_mai_n530_));
  NAi21      m0502(.An(mai_mai_n529_), .B(mai_mai_n530_), .Y(mai_mai_n531_));
  INV        m0503(.A(mai_mai_n46_), .Y(mai_mai_n532_));
  NO2        m0504(.A(mai_mai_n451_), .B(mai_mai_n46_), .Y(mai_mai_n533_));
  NA3        m0505(.A(mai_mai_n531_), .B(mai_mai_n527_), .C(mai_mai_n522_), .Y(mai_mai_n534_));
  NA2        m0506(.A(mai_mai_n97_), .B(mai_mai_n36_), .Y(mai_mai_n535_));
  NO2        m0507(.A(mai_mai_n448_), .B(mai_mai_n311_), .Y(mai_mai_n536_));
  NO2        m0508(.A(mai_mai_n536_), .B(n), .Y(mai_mai_n537_));
  NAi21      m0509(.An(mai_mai_n535_), .B(mai_mai_n537_), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n449_), .B(mai_mai_n163_), .Y(mai_mai_n539_));
  NA2        m0511(.A(mai_mai_n428_), .B(mai_mai_n148_), .Y(mai_mai_n540_));
  NO3        m0512(.A(mai_mai_n343_), .B(mai_mai_n540_), .C(mai_mai_n78_), .Y(mai_mai_n541_));
  AOI210     m0513(.A0(c), .A1(mai_mai_n539_), .B0(mai_mai_n541_), .Y(mai_mai_n542_));
  NAi31      m0514(.An(m), .B(n), .C(k), .Y(mai_mai_n543_));
  NO2        m0515(.A(mai_mai_n122_), .B(mai_mai_n543_), .Y(mai_mai_n544_));
  NA2        m0516(.A(mai_mai_n544_), .B(j), .Y(mai_mai_n545_));
  NA3        m0517(.A(mai_mai_n545_), .B(mai_mai_n542_), .C(mai_mai_n538_), .Y(mai_mai_n546_));
  NO4        m0518(.A(mai_mai_n546_), .B(mai_mai_n534_), .C(mai_mai_n520_), .D(mai_mai_n515_), .Y(mai_mai_n547_));
  NAi31      m0519(.An(g), .B(h), .C(f), .Y(mai_mai_n548_));
  OR3        m0520(.A(mai_mai_n548_), .B(mai_mai_n244_), .C(n), .Y(mai_mai_n549_));
  OA210      m0521(.A0(mai_mai_n451_), .A1(n), .B0(mai_mai_n489_), .Y(mai_mai_n550_));
  NA3        m0522(.A(e), .B(mai_mai_n109_), .C(mai_mai_n75_), .Y(mai_mai_n551_));
  OAI210     m0523(.A0(mai_mai_n550_), .A1(mai_mai_n82_), .B0(mai_mai_n551_), .Y(mai_mai_n552_));
  INV        m0524(.A(mai_mai_n552_), .Y(mai_mai_n553_));
  NO2        m0525(.A(mai_mai_n553_), .B(mai_mai_n445_), .Y(mai_mai_n554_));
  OR2        m0526(.A(mai_mai_n63_), .B(mai_mai_n64_), .Y(mai_mai_n555_));
  NA2        m0527(.A(b), .B(mai_mai_n296_), .Y(mai_mai_n556_));
  OA220      m0528(.A0(mai_mai_n529_), .A1(mai_mai_n556_), .B0(mai_mai_n526_), .B1(mai_mai_n555_), .Y(mai_mai_n557_));
  AN2        m0529(.A(h), .B(f), .Y(mai_mai_n558_));
  NA2        m0530(.A(mai_mai_n558_), .B(mai_mai_n37_), .Y(mai_mai_n559_));
  NO2        m0531(.A(mai_mai_n559_), .B(mai_mai_n394_), .Y(mai_mai_n560_));
  AOI210     m0532(.A0(d), .A1(mai_mai_n366_), .B0(mai_mai_n46_), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n492_), .B(k), .Y(mai_mai_n562_));
  AOI210     m0534(.A0(mai_mai_n562_), .A1(mai_mai_n561_), .B0(mai_mai_n560_), .Y(mai_mai_n563_));
  NA2        m0535(.A(mai_mai_n563_), .B(mai_mai_n557_), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n228_), .B(f), .Y(mai_mai_n565_));
  NA2        m0537(.A(mai_mai_n284_), .B(mai_mai_n128_), .Y(mai_mai_n566_));
  AOI220     m0538(.A0(mai_mai_n1228_), .A1(mai_mai_n448_), .B0(mai_mai_n311_), .B1(mai_mai_n102_), .Y(mai_mai_n567_));
  OA220      m0539(.A0(mai_mai_n567_), .A1(mai_mai_n465_), .B0(mai_mai_n309_), .B1(mai_mai_n100_), .Y(mai_mai_n568_));
  NA2        m0540(.A(mai_mai_n566_), .B(mai_mai_n568_), .Y(mai_mai_n569_));
  NO3        m0541(.A(mai_mai_n350_), .B(mai_mai_n174_), .C(mai_mai_n173_), .Y(mai_mai_n570_));
  NA2        m0542(.A(mai_mai_n570_), .B(mai_mai_n210_), .Y(mai_mai_n571_));
  NA3        m0543(.A(mai_mai_n571_), .B(mai_mai_n230_), .C(j), .Y(mai_mai_n572_));
  NA2        m0544(.A(mai_mai_n393_), .B(mai_mai_n75_), .Y(mai_mai_n573_));
  NA3        m0545(.A(mai_mai_n572_), .B(mai_mai_n432_), .C(mai_mai_n348_), .Y(mai_mai_n574_));
  NO4        m0546(.A(mai_mai_n574_), .B(mai_mai_n569_), .C(mai_mai_n564_), .D(mai_mai_n554_), .Y(mai_mai_n575_));
  NA4        m0547(.A(mai_mai_n575_), .B(mai_mai_n547_), .C(mai_mai_n508_), .D(mai_mai_n485_), .Y(mai08));
  NO2        m0548(.A(k), .B(h), .Y(mai_mai_n577_));
  AO210      m0549(.A0(mai_mai_n228_), .A1(mai_mai_n384_), .B0(mai_mai_n577_), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n578_), .B(mai_mai_n260_), .Y(mai_mai_n579_));
  NA2        m0551(.A(mai_mai_n516_), .B(mai_mai_n75_), .Y(mai_mai_n580_));
  AOI210     m0552(.A0(mai_mai_n516_), .A1(mai_mai_n579_), .B0(mai_mai_n413_), .Y(mai_mai_n581_));
  NA2        m0553(.A(mai_mai_n75_), .B(mai_mai_n99_), .Y(mai_mai_n582_));
  NO2        m0554(.A(mai_mai_n582_), .B(mai_mai_n53_), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n327_), .B(mai_mai_n101_), .Y(mai_mai_n584_));
  NA2        m0556(.A(mai_mai_n482_), .B(mai_mai_n212_), .Y(mai_mai_n585_));
  AOI220     m0557(.A0(mai_mai_n585_), .A1(mai_mai_n299_), .B0(mai_mai_n584_), .B1(mai_mai_n583_), .Y(mai_mai_n586_));
  NA4        m0558(.A(mai_mai_n195_), .B(mai_mai_n128_), .C(mai_mai_n43_), .D(h), .Y(mai_mai_n587_));
  AN2        m0559(.A(l), .B(k), .Y(mai_mai_n588_));
  NA4        m0560(.A(mai_mai_n588_), .B(mai_mai_n97_), .C(mai_mai_n64_), .D(mai_mai_n193_), .Y(mai_mai_n589_));
  NA3        m0561(.A(mai_mai_n586_), .B(mai_mai_n581_), .C(mai_mai_n301_), .Y(mai_mai_n590_));
  NO4        m0562(.A(mai_mai_n160_), .B(mai_mai_n341_), .C(mai_mai_n101_), .D(g), .Y(mai_mai_n591_));
  AOI210     m0563(.A0(mai_mai_n591_), .A1(mai_mai_n585_), .B0(mai_mai_n437_), .Y(mai_mai_n592_));
  NO2        m0564(.A(mai_mai_n38_), .B(mai_mai_n192_), .Y(mai_mai_n593_));
  NA2        m0565(.A(mai_mai_n518_), .B(mai_mai_n298_), .Y(mai_mai_n594_));
  NA2        m0566(.A(mai_mai_n594_), .B(mai_mai_n592_), .Y(mai_mai_n595_));
  NO2        m0567(.A(e), .B(mai_mai_n45_), .Y(mai_mai_n596_));
  NO2        m0568(.A(mai_mai_n407_), .B(mai_mai_n119_), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n597_), .B(mai_mai_n596_), .Y(mai_mai_n598_));
  NO3        m0570(.A(mai_mai_n276_), .B(mai_mai_n118_), .C(mai_mai_n41_), .Y(mai_mai_n599_));
  NAi21      m0571(.An(mai_mai_n599_), .B(mai_mai_n589_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n578_), .B(mai_mai_n123_), .Y(mai_mai_n601_));
  AOI220     m0573(.A0(mai_mai_n601_), .A1(mai_mai_n349_), .B0(mai_mai_n600_), .B1(mai_mai_n67_), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n598_), .B(mai_mai_n602_), .Y(mai_mai_n603_));
  NA2        m0575(.A(mai_mai_n311_), .B(mai_mai_n42_), .Y(mai_mai_n604_));
  NA3        m0576(.A(mai_mai_n571_), .B(mai_mai_n290_), .C(mai_mai_n333_), .Y(mai_mai_n605_));
  NA2        m0577(.A(mai_mai_n588_), .B(mai_mai_n200_), .Y(mai_mai_n606_));
  NO2        m0578(.A(mai_mai_n606_), .B(mai_mai_n283_), .Y(mai_mai_n607_));
  NA2        m0579(.A(mai_mai_n607_), .B(mai_mai_n565_), .Y(mai_mai_n608_));
  NA3        m0580(.A(m), .B(l), .C(k), .Y(mai_mai_n609_));
  AOI210     m0581(.A0(mai_mai_n551_), .A1(mai_mai_n549_), .B0(mai_mai_n609_), .Y(mai_mai_n610_));
  NA4        m0582(.A(mai_mai_n102_), .B(l), .C(k), .D(mai_mai_n78_), .Y(mai_mai_n611_));
  INV        m0583(.A(mai_mai_n610_), .Y(mai_mai_n612_));
  NA4        m0584(.A(mai_mai_n612_), .B(mai_mai_n608_), .C(mai_mai_n605_), .D(mai_mai_n604_), .Y(mai_mai_n613_));
  NO4        m0585(.A(mai_mai_n613_), .B(mai_mai_n603_), .C(mai_mai_n595_), .D(mai_mai_n590_), .Y(mai_mai_n614_));
  NA2        m0586(.A(mai_mai_n533_), .B(g), .Y(mai_mai_n615_));
  BUFFER     m0587(.A(mai_mai_n615_), .Y(mai_mai_n616_));
  NO2        m0588(.A(mai_mai_n346_), .B(mai_mai_n443_), .Y(mai_mai_n617_));
  NA2        m0589(.A(mai_mai_n617_), .B(mai_mai_n102_), .Y(mai_mai_n618_));
  NA3        m0590(.A(mai_mai_n618_), .B(mai_mai_n616_), .C(mai_mai_n226_), .Y(mai_mai_n619_));
  NA2        m0591(.A(mai_mai_n588_), .B(mai_mai_n64_), .Y(mai_mai_n620_));
  NO3        m0592(.A(mai_mai_n570_), .B(mai_mai_n160_), .C(i), .Y(mai_mai_n621_));
  NOi21      m0593(.An(h), .B(j), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n622_), .B(f), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n623_), .B(mai_mai_n223_), .Y(mai_mai_n624_));
  NO2        m0596(.A(mai_mai_n624_), .B(mai_mai_n621_), .Y(mai_mai_n625_));
  NO2        m0597(.A(mai_mai_n625_), .B(mai_mai_n620_), .Y(mai_mai_n626_));
  AOI210     m0598(.A0(mai_mai_n619_), .A1(l), .B0(mai_mai_n626_), .Y(mai_mai_n627_));
  NA2        m0599(.A(mai_mai_n71_), .B(l), .Y(mai_mai_n628_));
  INV        m0600(.A(mai_mai_n33_), .Y(mai_mai_n629_));
  OR2        m0601(.A(mai_mai_n628_), .B(mai_mai_n491_), .Y(mai_mai_n630_));
  NO3        m0602(.A(mai_mai_n139_), .B(mai_mai_n46_), .C(mai_mai_n99_), .Y(mai_mai_n631_));
  NO3        m0603(.A(n), .B(mai_mai_n138_), .C(mai_mai_n64_), .Y(mai_mai_n632_));
  NO2        m0604(.A(mai_mai_n407_), .B(mai_mai_n374_), .Y(mai_mai_n633_));
  OAI210     m0605(.A0(mai_mai_n632_), .A1(mai_mai_n631_), .B0(mai_mai_n633_), .Y(mai_mai_n634_));
  INV        m0606(.A(mai_mai_n634_), .Y(mai_mai_n635_));
  NA2        m0607(.A(k), .B(j), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n260_), .B(mai_mai_n636_), .Y(mai_mai_n637_));
  AOI210     m0609(.A0(mai_mai_n448_), .A1(n), .B0(mai_mai_n466_), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n638_), .B(mai_mai_n467_), .Y(mai_mai_n639_));
  AN3        m0611(.A(mai_mai_n639_), .B(mai_mai_n637_), .C(g), .Y(mai_mai_n640_));
  NO3        m0612(.A(mai_mai_n160_), .B(mai_mai_n341_), .C(mai_mai_n101_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n641_), .B(mai_mai_n224_), .Y(mai_mai_n642_));
  NAi31      m0614(.An(mai_mai_n504_), .B(mai_mai_n84_), .C(mai_mai_n75_), .Y(mai_mai_n643_));
  NA2        m0615(.A(mai_mai_n643_), .B(mai_mai_n642_), .Y(mai_mai_n644_));
  NO2        m0616(.A(mai_mai_n609_), .B(mai_mai_n82_), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n645_), .B(mai_mai_n490_), .Y(mai_mai_n646_));
  NO2        m0618(.A(mai_mai_n492_), .B(mai_mai_n106_), .Y(mai_mai_n647_));
  OAI210     m0619(.A0(mai_mai_n647_), .A1(mai_mai_n633_), .B0(mai_mai_n561_), .Y(mai_mai_n648_));
  NA2        m0620(.A(mai_mai_n648_), .B(mai_mai_n646_), .Y(mai_mai_n649_));
  OR4        m0621(.A(mai_mai_n649_), .B(mai_mai_n644_), .C(mai_mai_n640_), .D(mai_mai_n635_), .Y(mai_mai_n650_));
  NA2        m0622(.A(mai_mai_n638_), .B(mai_mai_n467_), .Y(mai_mai_n651_));
  NA4        m0623(.A(mai_mai_n651_), .B(mai_mai_n195_), .C(mai_mai_n384_), .D(mai_mai_n34_), .Y(mai_mai_n652_));
  NO2        m0624(.A(mai_mai_n587_), .B(mai_mai_n580_), .Y(mai_mai_n653_));
  INV        m0625(.A(mai_mai_n653_), .Y(mai_mai_n654_));
  NA3        m0626(.A(mai_mai_n461_), .B(mai_mai_n254_), .C(h), .Y(mai_mai_n655_));
  NO2        m0627(.A(mai_mai_n83_), .B(mai_mai_n45_), .Y(mai_mai_n656_));
  NO2        m0628(.A(mai_mai_n628_), .B(mai_mai_n555_), .Y(mai_mai_n657_));
  AOI210     m0629(.A0(mai_mai_n656_), .A1(mai_mai_n537_), .B0(mai_mai_n657_), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n658_), .B(mai_mai_n654_), .C(mai_mai_n652_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n645_), .B(mai_mai_n218_), .Y(mai_mai_n660_));
  NO2        m0632(.A(mai_mai_n550_), .B(mai_mai_n64_), .Y(mai_mai_n661_));
  OAI210     m0633(.A0(mai_mai_n609_), .A1(mai_mai_n548_), .B0(mai_mai_n436_), .Y(mai_mai_n662_));
  NA3        m0634(.A(mai_mai_n227_), .B(mai_mai_n55_), .C(b), .Y(mai_mai_n663_));
  AOI220     m0635(.A0(mai_mai_n501_), .A1(mai_mai_n29_), .B0(mai_mai_n393_), .B1(mai_mai_n75_), .Y(mai_mai_n664_));
  NA2        m0636(.A(mai_mai_n664_), .B(mai_mai_n663_), .Y(mai_mai_n665_));
  NO2        m0637(.A(mai_mai_n655_), .B(n), .Y(mai_mai_n666_));
  AOI210     m0638(.A0(mai_mai_n665_), .A1(mai_mai_n662_), .B0(mai_mai_n666_), .Y(mai_mai_n667_));
  NA2        m0639(.A(mai_mai_n667_), .B(mai_mai_n660_), .Y(mai_mai_n668_));
  NO3        m0640(.A(mai_mai_n668_), .B(mai_mai_n659_), .C(mai_mai_n650_), .Y(mai_mai_n669_));
  OR2        m0641(.A(mai_mai_n587_), .B(mai_mai_n212_), .Y(mai_mai_n670_));
  NO3        m0642(.A(mai_mai_n295_), .B(mai_mai_n262_), .C(mai_mai_n101_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n671_), .B(mai_mai_n639_), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n44_), .B(mai_mai_n52_), .Y(mai_mai_n673_));
  NO3        m0645(.A(mai_mai_n673_), .B(mai_mai_n629_), .C(mai_mai_n244_), .Y(mai_mai_n674_));
  NO2        m0646(.A(mai_mai_n443_), .B(mai_mai_n85_), .Y(mai_mai_n675_));
  AOI210     m0647(.A0(mai_mai_n675_), .A1(mai_mai_n583_), .B0(mai_mai_n674_), .Y(mai_mai_n676_));
  NA3        m0648(.A(mai_mai_n676_), .B(mai_mai_n672_), .C(mai_mai_n670_), .Y(mai_mai_n677_));
  OR2        m0649(.A(mai_mai_n548_), .B(mai_mai_n83_), .Y(mai_mai_n678_));
  NOi31      m0650(.An(b), .B(d), .C(a), .Y(mai_mai_n679_));
  NO2        m0651(.A(mai_mai_n679_), .B(mai_mai_n500_), .Y(mai_mai_n680_));
  NO2        m0652(.A(mai_mai_n680_), .B(n), .Y(mai_mai_n681_));
  NOi21      m0653(.An(mai_mai_n664_), .B(mai_mai_n681_), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n682_), .B(mai_mai_n678_), .Y(mai_mai_n683_));
  NO2        m0655(.A(mai_mai_n283_), .B(mai_mai_n106_), .Y(mai_mai_n684_));
  NOi21      m0656(.An(mai_mai_n684_), .B(mai_mai_n149_), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n570_), .B(n), .Y(mai_mai_n686_));
  NA2        m0658(.A(mai_mai_n686_), .B(mai_mai_n579_), .Y(mai_mai_n687_));
  NO2        m0659(.A(mai_mai_n279_), .B(mai_mai_n217_), .Y(mai_mai_n688_));
  OAI210     m0660(.A0(mai_mai_n86_), .A1(mai_mai_n84_), .B0(mai_mai_n688_), .Y(mai_mai_n689_));
  NA2        m0661(.A(mai_mai_n109_), .B(mai_mai_n75_), .Y(mai_mai_n690_));
  AOI210     m0662(.A0(mai_mai_n364_), .A1(mai_mai_n358_), .B0(mai_mai_n690_), .Y(mai_mai_n691_));
  NAi21      m0663(.An(mai_mai_n691_), .B(mai_mai_n689_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n607_), .B(mai_mai_n34_), .Y(mai_mai_n693_));
  NAi21      m0665(.An(mai_mai_n611_), .B(mai_mai_n371_), .Y(mai_mai_n694_));
  NO2        m0666(.A(mai_mai_n240_), .B(i), .Y(mai_mai_n695_));
  NA2        m0667(.A(mai_mai_n591_), .B(mai_mai_n300_), .Y(mai_mai_n696_));
  OAI210     m0668(.A0(mai_mai_n495_), .A1(mai_mai_n494_), .B0(l), .Y(mai_mai_n697_));
  AN3        m0669(.A(mai_mai_n697_), .B(mai_mai_n696_), .C(mai_mai_n694_), .Y(mai_mai_n698_));
  NAi41      m0670(.An(mai_mai_n692_), .B(mai_mai_n698_), .C(mai_mai_n693_), .D(mai_mai_n687_), .Y(mai_mai_n699_));
  NO4        m0671(.A(mai_mai_n699_), .B(mai_mai_n685_), .C(mai_mai_n683_), .D(mai_mai_n677_), .Y(mai_mai_n700_));
  NA4        m0672(.A(mai_mai_n700_), .B(mai_mai_n669_), .C(mai_mai_n627_), .D(mai_mai_n614_), .Y(mai09));
  INV        m0673(.A(mai_mai_n110_), .Y(mai_mai_n702_));
  NA2        m0674(.A(f), .B(e), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n1227_), .B(g), .Y(mai_mai_n704_));
  NA4        m0676(.A(mai_mai_n271_), .B(l), .C(i), .D(j), .Y(mai_mai_n705_));
  AOI210     m0677(.A0(mai_mai_n705_), .A1(g), .B0(mai_mai_n396_), .Y(mai_mai_n706_));
  AOI210     m0678(.A0(mai_mai_n706_), .A1(mai_mai_n704_), .B0(mai_mai_n703_), .Y(mai_mai_n707_));
  NA2        m0679(.A(mai_mai_n380_), .B(e), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n707_), .B(mai_mai_n702_), .Y(mai_mai_n709_));
  NO2        m0681(.A(mai_mai_n186_), .B(mai_mai_n192_), .Y(mai_mai_n710_));
  NA3        m0682(.A(m), .B(l), .C(i), .Y(mai_mai_n711_));
  OAI220     m0683(.A0(mai_mai_n492_), .A1(mai_mai_n711_), .B0(mai_mai_n304_), .B1(mai_mai_n444_), .Y(mai_mai_n712_));
  NA4        m0684(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(g), .D(f), .Y(mai_mai_n713_));
  NAi31      m0685(.An(mai_mai_n712_), .B(mai_mai_n713_), .C(mai_mai_n375_), .Y(mai_mai_n714_));
  OR2        m0686(.A(mai_mai_n714_), .B(mai_mai_n710_), .Y(mai_mai_n715_));
  NA3        m0687(.A(mai_mai_n678_), .B(mai_mai_n477_), .C(mai_mai_n436_), .Y(mai_mai_n716_));
  OA210      m0688(.A0(mai_mai_n716_), .A1(mai_mai_n715_), .B0(mai_mai_n681_), .Y(mai_mai_n717_));
  INV        m0689(.A(mai_mai_n293_), .Y(mai_mai_n718_));
  NOi31      m0690(.An(k), .B(m), .C(l), .Y(mai_mai_n719_));
  NO2        m0691(.A(m), .B(mai_mai_n498_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n296_), .B(mai_mai_n297_), .Y(mai_mai_n721_));
  OAI210     m0693(.A0(mai_mai_n186_), .A1(mai_mai_n192_), .B0(mai_mai_n721_), .Y(mai_mai_n722_));
  AOI220     m0694(.A0(mai_mai_n722_), .A1(mai_mai_n227_), .B0(mai_mai_n720_), .B1(mai_mai_n718_), .Y(mai_mai_n723_));
  NA3        m0695(.A(mai_mai_n103_), .B(mai_mai_n172_), .C(mai_mai_n31_), .Y(mai_mai_n724_));
  NA4        m0696(.A(mai_mai_n724_), .B(mai_mai_n723_), .C(mai_mai_n519_), .D(mai_mai_n73_), .Y(mai_mai_n725_));
  NO2        m0697(.A(mai_mai_n488_), .B(mai_mai_n419_), .Y(mai_mai_n726_));
  NA2        m0698(.A(mai_mai_n726_), .B(mai_mai_n172_), .Y(mai_mai_n727_));
  NOi21      m0699(.An(f), .B(d), .Y(mai_mai_n728_));
  NA2        m0700(.A(mai_mai_n728_), .B(m), .Y(mai_mai_n729_));
  NO2        m0701(.A(mai_mai_n729_), .B(mai_mai_n49_), .Y(mai_mai_n730_));
  NOi32      m0702(.An(g), .Bn(f), .C(d), .Y(mai_mai_n731_));
  NA4        m0703(.A(mai_mai_n731_), .B(mai_mai_n501_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n732_));
  NOi21      m0704(.An(mai_mai_n272_), .B(mai_mai_n732_), .Y(mai_mai_n733_));
  AOI210     m0705(.A0(mai_mai_n730_), .A1(mai_mai_n460_), .B0(mai_mai_n733_), .Y(mai_mai_n734_));
  NA3        m0706(.A(mai_mai_n271_), .B(i), .C(j), .Y(mai_mai_n735_));
  NA3        m0707(.A(mai_mai_n398_), .B(f), .C(mai_mai_n75_), .Y(mai_mai_n736_));
  NO3        m0708(.A(mai_mai_n736_), .B(mai_mai_n64_), .C(mai_mai_n193_), .Y(mai_mai_n737_));
  NO2        m0709(.A(i), .B(mai_mai_n52_), .Y(mai_mai_n738_));
  NA2        m0710(.A(mai_mai_n735_), .B(mai_mai_n737_), .Y(mai_mai_n739_));
  NAi41      m0711(.An(mai_mai_n412_), .B(mai_mai_n739_), .C(mai_mai_n734_), .D(mai_mai_n727_), .Y(mai_mai_n740_));
  NO4        m0712(.A(mai_mai_n517_), .B(mai_mai_n119_), .C(mai_mai_n283_), .D(mai_mai_n140_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n543_), .B(mai_mai_n283_), .Y(mai_mai_n742_));
  AN2        m0714(.A(mai_mai_n742_), .B(mai_mai_n565_), .Y(mai_mai_n743_));
  NO3        m0715(.A(mai_mai_n743_), .B(mai_mai_n741_), .C(mai_mai_n214_), .Y(mai_mai_n744_));
  NA2        m0716(.A(mai_mai_n500_), .B(mai_mai_n75_), .Y(mai_mai_n745_));
  NO2        m0717(.A(mai_mai_n721_), .B(mai_mai_n745_), .Y(mai_mai_n746_));
  NO2        m0718(.A(mai_mai_n736_), .B(mai_mai_n368_), .Y(mai_mai_n747_));
  NOi41      m0719(.An(mai_mai_n203_), .B(mai_mai_n747_), .C(mai_mai_n746_), .D(mai_mai_n268_), .Y(mai_mai_n748_));
  NA2        m0720(.A(c), .B(mai_mai_n105_), .Y(mai_mai_n749_));
  OR2        m0721(.A(mai_mai_n548_), .B(mai_mai_n457_), .Y(mai_mai_n750_));
  INV        m0722(.A(mai_mai_n750_), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n1230_), .B(mai_mai_n751_), .Y(mai_mai_n752_));
  NA3        m0724(.A(mai_mai_n752_), .B(mai_mai_n748_), .C(mai_mai_n744_), .Y(mai_mai_n753_));
  NO4        m0725(.A(mai_mai_n753_), .B(mai_mai_n740_), .C(mai_mai_n725_), .D(mai_mai_n717_), .Y(mai_mai_n754_));
  OR2        m0726(.A(mai_mai_n736_), .B(mai_mai_n64_), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n1227_), .B(g), .Y(mai_mai_n756_));
  AOI210     m0728(.A0(mai_mai_n756_), .A1(mai_mai_n255_), .B0(mai_mai_n755_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n123_), .B(mai_mai_n119_), .Y(mai_mai_n758_));
  NO2        m0730(.A(mai_mai_n210_), .B(mai_mai_n204_), .Y(mai_mai_n759_));
  AOI220     m0731(.A0(mai_mai_n759_), .A1(mai_mai_n207_), .B0(mai_mai_n266_), .B1(mai_mai_n758_), .Y(mai_mai_n760_));
  NO2        m0732(.A(mai_mai_n368_), .B(mai_mai_n703_), .Y(mai_mai_n761_));
  INV        m0733(.A(mai_mai_n760_), .Y(mai_mai_n762_));
  NA2        m0734(.A(e), .B(d), .Y(mai_mai_n763_));
  OAI220     m0735(.A0(mai_mai_n763_), .A1(c), .B0(mai_mai_n279_), .B1(d), .Y(mai_mai_n764_));
  NA3        m0736(.A(mai_mai_n764_), .B(mai_mai_n387_), .C(mai_mai_n428_), .Y(mai_mai_n765_));
  AOI210     m0737(.A0(mai_mai_n433_), .A1(mai_mai_n167_), .B0(mai_mai_n210_), .Y(mai_mai_n766_));
  AOI210     m0738(.A0(mai_mai_n518_), .A1(mai_mai_n298_), .B0(mai_mai_n766_), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n737_), .B(mai_mai_n1226_), .Y(mai_mai_n768_));
  NA3        m0740(.A(mai_mai_n153_), .B(mai_mai_n76_), .C(mai_mai_n34_), .Y(mai_mai_n769_));
  NA4        m0741(.A(mai_mai_n769_), .B(mai_mai_n768_), .C(mai_mai_n767_), .D(mai_mai_n765_), .Y(mai_mai_n770_));
  NO3        m0742(.A(mai_mai_n770_), .B(mai_mai_n762_), .C(mai_mai_n757_), .Y(mai_mai_n771_));
  NA2        m0743(.A(mai_mai_n718_), .B(mai_mai_n31_), .Y(mai_mai_n772_));
  OR2        m0744(.A(mai_mai_n772_), .B(mai_mai_n196_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n517_), .B(mai_mai_n57_), .Y(mai_mai_n774_));
  AOI220     m0746(.A0(mai_mai_n774_), .A1(mai_mai_n742_), .B0(mai_mai_n509_), .B1(mai_mai_n516_), .Y(mai_mai_n775_));
  OAI210     m0747(.A0(mai_mai_n708_), .A1(mai_mai_n157_), .B0(mai_mai_n775_), .Y(mai_mai_n776_));
  OAI210     m0748(.A0(mai_mai_n1227_), .A1(mai_mai_n1226_), .B0(mai_mai_n731_), .Y(mai_mai_n777_));
  NO2        m0749(.A(mai_mai_n777_), .B(mai_mai_n502_), .Y(mai_mai_n778_));
  NO2        m0750(.A(i), .B(mai_mai_n732_), .Y(mai_mai_n779_));
  AO210      m0751(.A0(mai_mai_n227_), .A1(mai_mai_n712_), .B0(mai_mai_n779_), .Y(mai_mai_n780_));
  NOi31      m0752(.An(mai_mai_n460_), .B(mai_mai_n729_), .C(mai_mai_n255_), .Y(mai_mai_n781_));
  NO4        m0753(.A(mai_mai_n781_), .B(mai_mai_n780_), .C(mai_mai_n778_), .D(mai_mai_n776_), .Y(mai_mai_n782_));
  AO220      m0754(.A0(mai_mai_n387_), .A1(mai_mai_n622_), .B0(mai_mai_n162_), .B1(f), .Y(mai_mai_n783_));
  NA2        m0755(.A(mai_mai_n783_), .B(mai_mai_n764_), .Y(mai_mai_n784_));
  NO2        m0756(.A(mai_mai_n374_), .B(mai_mai_n61_), .Y(mai_mai_n785_));
  OAI210     m0757(.A0(mai_mai_n716_), .A1(mai_mai_n785_), .B0(mai_mai_n583_), .Y(mai_mai_n786_));
  AN4        m0758(.A(mai_mai_n786_), .B(mai_mai_n784_), .C(mai_mai_n782_), .D(mai_mai_n773_), .Y(mai_mai_n787_));
  NA4        m0759(.A(mai_mai_n787_), .B(mai_mai_n771_), .C(mai_mai_n754_), .D(mai_mai_n709_), .Y(mai12));
  NO4        m0760(.A(mai_mai_n379_), .B(mai_mai_n228_), .C(mai_mai_n486_), .D(mai_mai_n193_), .Y(mai_mai_n789_));
  NO2        m0761(.A(mai_mai_n385_), .B(mai_mai_n105_), .Y(mai_mai_n790_));
  NO2        m0762(.A(mai_mai_n548_), .B(mai_mai_n327_), .Y(mai_mai_n791_));
  NA2        m0763(.A(mai_mai_n791_), .B(mai_mai_n459_), .Y(mai_mai_n792_));
  NA2        m0764(.A(mai_mai_n792_), .B(mai_mai_n378_), .Y(mai_mai_n793_));
  AOI210     m0765(.A0(mai_mai_n213_), .A1(mai_mai_n292_), .B0(mai_mai_n183_), .Y(mai_mai_n794_));
  OR2        m0766(.A(mai_mai_n794_), .B(mai_mai_n789_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n339_), .B(mai_mai_n193_), .Y(mai_mai_n796_));
  OAI210     m0768(.A0(mai_mai_n796_), .A1(mai_mai_n795_), .B0(mai_mai_n350_), .Y(mai_mai_n797_));
  INV        m0769(.A(mai_mai_n535_), .Y(mai_mai_n798_));
  NO2        m0770(.A(mai_mai_n492_), .B(mai_mai_n711_), .Y(mai_mai_n799_));
  NA2        m0771(.A(mai_mai_n688_), .B(mai_mai_n798_), .Y(mai_mai_n800_));
  NO2        m0772(.A(mai_mai_n139_), .B(mai_mai_n217_), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n800_), .B(mai_mai_n797_), .Y(mai_mai_n802_));
  BUFFER     m0774(.A(mai_mai_n280_), .Y(mai_mai_n803_));
  NO3        m0775(.A(mai_mai_n119_), .B(mai_mai_n140_), .C(mai_mai_n193_), .Y(mai_mai_n804_));
  NA2        m0776(.A(mai_mai_n804_), .B(mai_mai_n448_), .Y(mai_mai_n805_));
  NO3        m0777(.A(mai_mai_n553_), .B(mai_mai_n83_), .C(mai_mai_n43_), .Y(mai_mai_n806_));
  NO4        m0778(.A(mai_mai_n806_), .B(mai_mai_n1223_), .C(mai_mai_n802_), .D(mai_mai_n793_), .Y(mai_mai_n807_));
  NO2        m0779(.A(mai_mai_n318_), .B(mai_mai_n317_), .Y(mai_mai_n808_));
  NA2        m0780(.A(mai_mai_n489_), .B(mai_mai_n63_), .Y(mai_mai_n809_));
  NOi21      m0781(.An(mai_mai_n34_), .B(mai_mai_n543_), .Y(mai_mai_n810_));
  AOI220     m0782(.A0(mai_mai_n810_), .A1(mai_mai_n1232_), .B0(mai_mai_n809_), .B1(mai_mai_n808_), .Y(mai_mai_n811_));
  INV        m0783(.A(mai_mai_n811_), .Y(mai_mai_n812_));
  INV        m0784(.A(mai_mai_n315_), .Y(mai_mai_n813_));
  NO2        m0785(.A(mai_mai_n813_), .B(mai_mai_n812_), .Y(mai_mai_n814_));
  NA2        m0786(.A(mai_mai_n298_), .B(g), .Y(mai_mai_n815_));
  NA2        m0787(.A(h), .B(i), .Y(mai_mai_n816_));
  NO2        m0788(.A(mai_mai_n816_), .B(mai_mai_n83_), .Y(mai_mai_n817_));
  INV        m0789(.A(mai_mai_n817_), .Y(mai_mai_n818_));
  OAI220     m0790(.A0(mai_mai_n133_), .A1(mai_mai_n815_), .B0(mai_mai_n818_), .B1(mai_mai_n288_), .Y(mai_mai_n819_));
  NO2        m0791(.A(mai_mai_n548_), .B(mai_mai_n419_), .Y(mai_mai_n820_));
  NA3        m0792(.A(mai_mai_n296_), .B(mai_mai_n523_), .C(i), .Y(mai_mai_n821_));
  OAI210     m0793(.A0(mai_mai_n374_), .A1(mai_mai_n271_), .B0(mai_mai_n821_), .Y(mai_mai_n822_));
  OAI220     m0794(.A0(mai_mai_n822_), .A1(mai_mai_n820_), .B0(mai_mai_n561_), .B1(mai_mai_n632_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n503_), .B(mai_mai_n102_), .Y(mai_mai_n824_));
  OR3        m0796(.A(mai_mai_n271_), .B(mai_mai_n370_), .C(f), .Y(mai_mai_n825_));
  NA3        m0797(.A(mai_mai_n523_), .B(mai_mai_n71_), .C(i), .Y(mai_mai_n826_));
  OA220      m0798(.A0(mai_mai_n826_), .A1(mai_mai_n824_), .B0(mai_mai_n825_), .B1(mai_mai_n491_), .Y(mai_mai_n827_));
  NA3        m0799(.A(f), .B(mai_mai_n107_), .C(g), .Y(mai_mai_n828_));
  AOI210     m0800(.A0(mai_mai_n559_), .A1(mai_mai_n828_), .B0(m), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n829_), .B(mai_mai_n280_), .Y(mai_mai_n830_));
  NA2        m0802(.A(mai_mai_n713_), .B(mai_mai_n375_), .Y(mai_mai_n831_));
  NA2        m0803(.A(mai_mai_n201_), .B(mai_mai_n68_), .Y(mai_mai_n832_));
  NA3        m0804(.A(mai_mai_n832_), .B(mai_mai_n826_), .C(mai_mai_n825_), .Y(mai_mai_n833_));
  AOI220     m0805(.A0(mai_mai_n833_), .A1(mai_mai_n233_), .B0(mai_mai_n831_), .B1(mai_mai_n75_), .Y(mai_mai_n834_));
  NA4        m0806(.A(mai_mai_n834_), .B(mai_mai_n830_), .C(mai_mai_n827_), .D(mai_mai_n823_), .Y(mai_mai_n835_));
  NO2        m0807(.A(mai_mai_n327_), .B(mai_mai_n82_), .Y(mai_mai_n836_));
  OAI210     m0808(.A0(mai_mai_n836_), .A1(mai_mai_n798_), .B0(mai_mai_n218_), .Y(mai_mai_n837_));
  NA2        m0809(.A(mai_mai_n552_), .B(mai_mai_n79_), .Y(mai_mai_n838_));
  NO2        m0810(.A(mai_mai_n391_), .B(mai_mai_n193_), .Y(mai_mai_n839_));
  AOI220     m0811(.A0(mai_mai_n839_), .A1(mai_mai_n332_), .B0(mai_mai_n803_), .B1(mai_mai_n197_), .Y(mai_mai_n840_));
  AOI220     m0812(.A0(mai_mai_n791_), .A1(mai_mai_n801_), .B0(mai_mai_n490_), .B1(mai_mai_n81_), .Y(mai_mai_n841_));
  NA4        m0813(.A(mai_mai_n841_), .B(mai_mai_n840_), .C(mai_mai_n838_), .D(mai_mai_n837_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n799_), .B(mai_mai_n459_), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n360_), .B(mai_mai_n690_), .Y(mai_mai_n844_));
  OAI210     m0816(.A0(mai_mai_n318_), .A1(mai_mai_n317_), .B0(mai_mai_n98_), .Y(mai_mai_n845_));
  AOI210     m0817(.A0(mai_mai_n845_), .A1(mai_mai_n452_), .B0(mai_mai_n844_), .Y(mai_mai_n846_));
  NA2        m0818(.A(mai_mai_n829_), .B(mai_mai_n790_), .Y(mai_mai_n847_));
  NO3        m0819(.A(mai_mai_n1221_), .B(mai_mai_n46_), .C(mai_mai_n43_), .Y(mai_mai_n848_));
  AOI220     m0820(.A0(mai_mai_n848_), .A1(mai_mai_n521_), .B0(mai_mai_n539_), .B1(mai_mai_n448_), .Y(mai_mai_n849_));
  NA4        m0821(.A(mai_mai_n849_), .B(mai_mai_n847_), .C(mai_mai_n846_), .D(mai_mai_n843_), .Y(mai_mai_n850_));
  NO4        m0822(.A(mai_mai_n850_), .B(mai_mai_n842_), .C(mai_mai_n835_), .D(mai_mai_n819_), .Y(mai_mai_n851_));
  NAi31      m0823(.An(mai_mai_n129_), .B(mai_mai_n361_), .C(n), .Y(mai_mai_n852_));
  NO2        m0824(.A(m), .B(mai_mai_n852_), .Y(mai_mai_n853_));
  NO2        m0825(.A(mai_mai_n240_), .B(mai_mai_n129_), .Y(mai_mai_n854_));
  AOI210     m0826(.A0(mai_mai_n854_), .A1(mai_mai_n420_), .B0(mai_mai_n853_), .Y(mai_mai_n855_));
  NA2        m0827(.A(mai_mai_n413_), .B(i), .Y(mai_mai_n856_));
  NA2        m0828(.A(mai_mai_n856_), .B(mai_mai_n855_), .Y(mai_mai_n857_));
  NA2        m0829(.A(mai_mai_n210_), .B(mai_mai_n158_), .Y(mai_mai_n858_));
  NO3        m0830(.A(mai_mai_n374_), .B(mai_mai_n271_), .C(mai_mai_n64_), .Y(mai_mai_n859_));
  AOI220     m0831(.A0(mai_mai_n859_), .A1(mai_mai_n372_), .B0(mai_mai_n404_), .B1(g), .Y(mai_mai_n860_));
  INV        m0832(.A(mai_mai_n860_), .Y(mai_mai_n861_));
  NA2        m0833(.A(mai_mai_n442_), .B(mai_mai_n328_), .Y(mai_mai_n862_));
  OAI220     m0834(.A0(mai_mai_n791_), .A1(mai_mai_n799_), .B0(mai_mai_n460_), .B1(mai_mai_n367_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n863_), .B(mai_mai_n862_), .Y(mai_mai_n864_));
  OAI210     m0836(.A0(mai_mai_n794_), .A1(mai_mai_n789_), .B0(mai_mai_n858_), .Y(mai_mai_n865_));
  AOI210     m0837(.A0(mai_mai_n330_), .A1(mai_mai_n328_), .B0(mai_mai_n287_), .Y(mai_mai_n866_));
  NA3        m0838(.A(mai_mai_n866_), .B(mai_mai_n865_), .C(mai_mai_n241_), .Y(mai_mai_n867_));
  OR2        m0839(.A(mai_mai_n867_), .B(mai_mai_n864_), .Y(mai_mai_n868_));
  NO3        m0840(.A(mai_mai_n868_), .B(mai_mai_n861_), .C(mai_mai_n857_), .Y(mai_mai_n869_));
  NA4        m0841(.A(mai_mai_n869_), .B(mai_mai_n851_), .C(mai_mai_n814_), .D(mai_mai_n807_), .Y(mai13));
  AN2        m0842(.A(c), .B(b), .Y(mai_mai_n871_));
  NA3        m0843(.A(mai_mai_n227_), .B(mai_mai_n871_), .C(m), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n417_), .B(f), .Y(mai_mai_n873_));
  NO3        m0845(.A(mai_mai_n873_), .B(mai_mai_n872_), .C(k), .Y(mai_mai_n874_));
  NAi32      m0846(.An(d), .Bn(c), .C(e), .Y(mai_mai_n875_));
  NA2        m0847(.A(mai_mai_n128_), .B(mai_mai_n43_), .Y(mai_mai_n876_));
  NO4        m0848(.A(mai_mai_n876_), .B(mai_mai_n875_), .C(mai_mai_n492_), .D(mai_mai_n269_), .Y(mai_mai_n877_));
  AN2        m0849(.A(d), .B(c), .Y(mai_mai_n878_));
  NA2        m0850(.A(mai_mai_n878_), .B(mai_mai_n105_), .Y(mai_mai_n879_));
  NO4        m0851(.A(mai_mai_n879_), .B(f), .C(mai_mai_n163_), .D(mai_mai_n154_), .Y(mai_mai_n880_));
  NA2        m0852(.A(mai_mai_n417_), .B(c), .Y(mai_mai_n881_));
  NO4        m0853(.A(mai_mai_n876_), .B(mai_mai_n488_), .C(mai_mai_n881_), .D(mai_mai_n269_), .Y(mai_mai_n882_));
  OR2        m0854(.A(mai_mai_n880_), .B(mai_mai_n882_), .Y(mai_mai_n883_));
  OR3        m0855(.A(mai_mai_n883_), .B(mai_mai_n877_), .C(mai_mai_n874_), .Y(mai_mai_n884_));
  NO2        m0856(.A(f), .B(mai_mai_n135_), .Y(mai_mai_n885_));
  NA2        m0857(.A(mai_mai_n885_), .B(g), .Y(mai_mai_n886_));
  OR2        m0858(.A(mai_mai_n163_), .B(mai_mai_n154_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n887_), .B(mai_mai_n886_), .Y(mai_mai_n888_));
  NO2        m0860(.A(mai_mai_n881_), .B(mai_mai_n269_), .Y(mai_mai_n889_));
  NA2        m0861(.A(mai_mai_n525_), .B(mai_mai_n1220_), .Y(mai_mai_n890_));
  NOi21      m0862(.An(mai_mai_n889_), .B(mai_mai_n890_), .Y(mai_mai_n891_));
  NO2        m0863(.A(mai_mai_n636_), .B(mai_mai_n101_), .Y(mai_mai_n892_));
  NOi41      m0864(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n893_), .B(mai_mai_n892_), .Y(mai_mai_n894_));
  NO2        m0866(.A(mai_mai_n894_), .B(mai_mai_n886_), .Y(mai_mai_n895_));
  OR3        m0867(.A(e), .B(d), .C(c), .Y(mai_mai_n896_));
  NA3        m0868(.A(k), .B(j), .C(i), .Y(mai_mai_n897_));
  NO3        m0869(.A(mai_mai_n897_), .B(mai_mai_n269_), .C(mai_mai_n82_), .Y(mai_mai_n898_));
  NOi21      m0870(.An(mai_mai_n898_), .B(mai_mai_n896_), .Y(mai_mai_n899_));
  OR4        m0871(.A(mai_mai_n899_), .B(mai_mai_n895_), .C(mai_mai_n891_), .D(mai_mai_n888_), .Y(mai_mai_n900_));
  NA3        m0872(.A(mai_mai_n395_), .B(mai_mai_n290_), .C(mai_mai_n52_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n901_), .B(mai_mai_n890_), .Y(mai_mai_n902_));
  NO3        m0874(.A(mai_mai_n901_), .B(mai_mai_n488_), .C(mai_mai_n384_), .Y(mai_mai_n903_));
  NO2        m0875(.A(f), .B(c), .Y(mai_mai_n904_));
  NOi21      m0876(.An(mai_mai_n904_), .B(mai_mai_n379_), .Y(mai_mai_n905_));
  NA2        m0877(.A(mai_mai_n905_), .B(mai_mai_n55_), .Y(mai_mai_n906_));
  NO3        m0878(.A(i), .B(h), .C(l), .Y(mai_mai_n907_));
  NOi31      m0879(.An(mai_mai_n907_), .B(mai_mai_n906_), .C(j), .Y(mai_mai_n908_));
  OR3        m0880(.A(mai_mai_n908_), .B(mai_mai_n903_), .C(mai_mai_n902_), .Y(mai_mai_n909_));
  OR3        m0881(.A(mai_mai_n909_), .B(mai_mai_n900_), .C(mai_mai_n884_), .Y(mai02));
  OR3        m0882(.A(n), .B(m), .C(i), .Y(mai_mai_n911_));
  NO4        m0883(.A(mai_mai_n911_), .B(h), .C(l), .D(mai_mai_n896_), .Y(mai_mai_n912_));
  NOi31      m0884(.An(e), .B(d), .C(c), .Y(mai_mai_n913_));
  AOI210     m0885(.A0(mai_mai_n898_), .A1(mai_mai_n913_), .B0(mai_mai_n877_), .Y(mai_mai_n914_));
  AN3        m0886(.A(g), .B(f), .C(c), .Y(mai_mai_n915_));
  INV        m0887(.A(mai_mai_n915_), .Y(mai_mai_n916_));
  OR2        m0888(.A(mai_mai_n897_), .B(mai_mai_n269_), .Y(mai_mai_n917_));
  OR2        m0889(.A(mai_mai_n917_), .B(mai_mai_n916_), .Y(mai_mai_n918_));
  NO3        m0890(.A(mai_mai_n901_), .B(mai_mai_n876_), .C(mai_mai_n488_), .Y(mai_mai_n919_));
  NO2        m0891(.A(mai_mai_n919_), .B(mai_mai_n888_), .Y(mai_mai_n920_));
  NA3        m0892(.A(l), .B(k), .C(j), .Y(mai_mai_n921_));
  NA2        m0893(.A(i), .B(h), .Y(mai_mai_n922_));
  NO3        m0894(.A(mai_mai_n922_), .B(mai_mai_n921_), .C(mai_mai_n119_), .Y(mai_mai_n923_));
  NO3        m0895(.A(mai_mai_n130_), .B(mai_mai_n250_), .C(mai_mai_n193_), .Y(mai_mai_n924_));
  AOI210     m0896(.A0(mai_mai_n924_), .A1(mai_mai_n923_), .B0(mai_mai_n891_), .Y(mai_mai_n925_));
  NA3        m0897(.A(c), .B(b), .C(a), .Y(mai_mai_n926_));
  NO3        m0898(.A(mai_mai_n926_), .B(mai_mai_n763_), .C(mai_mai_n192_), .Y(mai_mai_n927_));
  NO2        m0899(.A(mai_mai_n46_), .B(mai_mai_n101_), .Y(mai_mai_n928_));
  AOI210     m0900(.A0(mai_mai_n928_), .A1(mai_mai_n927_), .B0(mai_mai_n902_), .Y(mai_mai_n929_));
  AN4        m0901(.A(mai_mai_n929_), .B(mai_mai_n925_), .C(mai_mai_n920_), .D(mai_mai_n918_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n879_), .B(f), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n894_), .B(mai_mai_n887_), .Y(mai_mai_n932_));
  AOI210     m0904(.A0(mai_mai_n932_), .A1(mai_mai_n931_), .B0(mai_mai_n874_), .Y(mai_mai_n933_));
  NAi41      m0905(.An(mai_mai_n912_), .B(mai_mai_n933_), .C(mai_mai_n930_), .D(mai_mai_n914_), .Y(mai03));
  NA4        m0906(.A(g), .B(m), .C(mai_mai_n101_), .D(mai_mai_n192_), .Y(mai_mai_n935_));
  NOi41      m0907(.An(mai_mai_n678_), .B(mai_mai_n722_), .C(mai_mai_n714_), .D(mai_mai_n593_), .Y(mai_mai_n936_));
  OAI220     m0908(.A0(mai_mai_n936_), .A1(mai_mai_n573_), .B0(mai_mai_n935_), .B1(mai_mai_n489_), .Y(mai_mai_n937_));
  NA4        m0909(.A(i), .B(mai_mai_n913_), .C(mai_mai_n296_), .D(mai_mai_n290_), .Y(mai_mai_n938_));
  INV        m0910(.A(mai_mai_n938_), .Y(mai_mai_n939_));
  NOi31      m0911(.An(m), .B(n), .C(f), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n940_), .B(mai_mai_n48_), .Y(mai_mai_n941_));
  AN2        m0913(.A(e), .B(c), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n942_), .B(a), .Y(mai_mai_n943_));
  OAI220     m0915(.A0(mai_mai_n943_), .A1(mai_mai_n941_), .B0(mai_mai_n750_), .B1(mai_mai_n366_), .Y(mai_mai_n944_));
  NOi31      m0916(.An(mai_mai_n731_), .B(mai_mai_n872_), .C(h), .Y(mai_mai_n945_));
  NO4        m0917(.A(mai_mai_n945_), .B(mai_mai_n944_), .C(mai_mai_n939_), .D(mai_mai_n844_), .Y(mai_mai_n946_));
  INV        m0918(.A(mai_mai_n877_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n922_), .B(mai_mai_n407_), .Y(mai_mai_n948_));
  NO2        m0920(.A(mai_mai_n78_), .B(g), .Y(mai_mai_n949_));
  NO2        m0921(.A(mai_mai_n948_), .B(mai_mai_n907_), .Y(mai_mai_n950_));
  OR2        m0922(.A(mai_mai_n950_), .B(mai_mai_n906_), .Y(mai_mai_n951_));
  NA3        m0923(.A(mai_mai_n951_), .B(mai_mai_n947_), .C(mai_mai_n946_), .Y(mai_mai_n952_));
  NO4        m0924(.A(mai_mai_n952_), .B(mai_mai_n937_), .C(mai_mai_n692_), .D(mai_mai_n475_), .Y(mai_mai_n953_));
  NA2        m0925(.A(c), .B(b), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n582_), .B(mai_mai_n954_), .Y(mai_mai_n955_));
  OAI210     m0927(.A0(mai_mai_n729_), .A1(mai_mai_n706_), .B0(mai_mai_n357_), .Y(mai_mai_n956_));
  OAI210     m0928(.A0(mai_mai_n956_), .A1(mai_mai_n730_), .B0(mai_mai_n955_), .Y(mai_mai_n957_));
  NAi21      m0929(.An(mai_mai_n362_), .B(mai_mai_n955_), .Y(mai_mai_n958_));
  NA3        m0930(.A(mai_mai_n367_), .B(mai_mai_n468_), .C(f), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n959_), .B(mai_mai_n958_), .Y(mai_mai_n960_));
  NAi21      m0932(.An(f), .B(d), .Y(mai_mai_n961_));
  NO2        m0933(.A(mai_mai_n961_), .B(mai_mai_n926_), .Y(mai_mai_n962_));
  AOI210     m0934(.A0(mai_mai_n962_), .A1(mai_mai_n102_), .B0(mai_mai_n960_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n169_), .B(mai_mai_n217_), .Y(mai_mai_n964_));
  NA2        m0936(.A(mai_mai_n964_), .B(m), .Y(mai_mai_n965_));
  NO2        m0937(.A(mai_mai_n136_), .B(mai_mai_n965_), .Y(mai_mai_n966_));
  NA2        m0938(.A(mai_mai_n470_), .B(mai_mai_n356_), .Y(mai_mai_n967_));
  NO2        m0939(.A(mai_mai_n321_), .B(mai_mai_n320_), .Y(mai_mai_n968_));
  NAi21      m0940(.An(mai_mai_n968_), .B(mai_mai_n967_), .Y(mai_mai_n969_));
  NO2        m0941(.A(mai_mai_n969_), .B(mai_mai_n966_), .Y(mai_mai_n970_));
  NA4        m0942(.A(mai_mai_n970_), .B(mai_mai_n963_), .C(mai_mai_n957_), .D(mai_mai_n953_), .Y(mai00));
  NA2        m0943(.A(mai_mai_n261_), .B(mai_mai_n193_), .Y(mai_mai_n972_));
  NO2        m0944(.A(mai_mai_n972_), .B(mai_mai_n482_), .Y(mai_mai_n973_));
  AOI210     m0945(.A0(mai_mai_n761_), .A1(mai_mai_n801_), .B0(mai_mai_n939_), .Y(mai_mai_n974_));
  INV        m0946(.A(mai_mai_n919_), .Y(mai_mai_n975_));
  NA3        m0947(.A(mai_mai_n975_), .B(mai_mai_n974_), .C(mai_mai_n846_), .Y(mai_mai_n976_));
  NA3        m0948(.A(mai_mai_n719_), .B(g), .C(n), .Y(mai_mai_n977_));
  NO2        m0949(.A(mai_mai_n977_), .B(mai_mai_n879_), .Y(mai_mai_n978_));
  NO4        m0950(.A(mai_mai_n978_), .B(mai_mai_n976_), .C(mai_mai_n973_), .D(mai_mai_n900_), .Y(mai_mai_n979_));
  NA3        m0951(.A(mai_mai_n153_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n980_));
  NA2        m0952(.A(d), .B(b), .Y(mai_mai_n981_));
  NO2        m0953(.A(mai_mai_n981_), .B(mai_mai_n980_), .Y(mai_mai_n982_));
  NO3        m0954(.A(mai_mai_n982_), .B(mai_mai_n968_), .C(mai_mai_n781_), .Y(mai_mai_n983_));
  NO4        m0955(.A(mai_mai_n410_), .B(mai_mai_n305_), .C(mai_mai_n954_), .D(mai_mai_n55_), .Y(mai_mai_n984_));
  NA3        m0956(.A(mai_mai_n333_), .B(mai_mai_n200_), .C(g), .Y(mai_mai_n985_));
  OR2        m0957(.A(mai_mai_n334_), .B(mai_mai_n122_), .Y(mai_mai_n986_));
  NO2        m0958(.A(h), .B(g), .Y(mai_mai_n987_));
  NA4        m0959(.A(mai_mai_n420_), .B(mai_mai_n395_), .C(mai_mai_n987_), .D(mai_mai_n871_), .Y(mai_mai_n988_));
  NO2        m0960(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n989_));
  AOI220     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n452_), .B0(mai_mai_n804_), .B1(mai_mai_n481_), .Y(mai_mai_n990_));
  AOI220     m0962(.A0(mai_mai_n277_), .A1(mai_mai_n224_), .B0(mai_mai_n164_), .B1(mai_mai_n137_), .Y(mai_mai_n991_));
  NA4        m0963(.A(mai_mai_n991_), .B(mai_mai_n990_), .C(mai_mai_n988_), .D(mai_mai_n986_), .Y(mai_mai_n992_));
  NO2        m0964(.A(mai_mai_n992_), .B(mai_mai_n984_), .Y(mai_mai_n993_));
  AOI210     m0965(.A0(mai_mai_n224_), .A1(mai_mai_n298_), .B0(mai_mai_n483_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n994_), .B(mai_mai_n142_), .Y(mai_mai_n995_));
  NO2        m0967(.A(mai_mai_n219_), .B(mai_mai_n168_), .Y(mai_mai_n996_));
  NA2        m0968(.A(mai_mai_n996_), .B(mai_mai_n367_), .Y(mai_mai_n997_));
  NA3        m0969(.A(mai_mai_n166_), .B(mai_mai_n101_), .C(g), .Y(mai_mai_n998_));
  NA2        m0970(.A(mai_mai_n395_), .B(f), .Y(mai_mai_n999_));
  NOi31      m0971(.An(mai_mai_n738_), .B(mai_mai_n999_), .C(mai_mai_n998_), .Y(mai_mai_n1000_));
  NAi21      m0972(.An(mai_mai_n1000_), .B(mai_mai_n997_), .Y(mai_mai_n1001_));
  NO3        m0973(.A(mai_mai_n366_), .B(mai_mai_n703_), .C(n), .Y(mai_mai_n1002_));
  AOI210     m0974(.A0(mai_mai_n1002_), .A1(m), .B0(mai_mai_n912_), .Y(mai_mai_n1003_));
  NAi21      m0975(.An(mai_mai_n882_), .B(mai_mai_n1003_), .Y(mai_mai_n1004_));
  NO3        m0976(.A(mai_mai_n1004_), .B(mai_mai_n1001_), .C(mai_mai_n995_), .Y(mai_mai_n1005_));
  AN3        m0977(.A(mai_mai_n1005_), .B(mai_mai_n993_), .C(mai_mai_n983_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n452_), .B(mai_mai_n90_), .Y(mai_mai_n1007_));
  NA3        m0979(.A(mai_mai_n940_), .B(mai_mai_n503_), .C(k), .Y(mai_mai_n1008_));
  NA4        m0980(.A(mai_mai_n1008_), .B(mai_mai_n471_), .C(mai_mai_n1007_), .D(mai_mai_n221_), .Y(mai_mai_n1009_));
  OAI210     m0981(.A0(mai_mai_n394_), .A1(mai_mai_n108_), .B0(mai_mai_n732_), .Y(mai_mai_n1010_));
  AOI210     m0982(.A0(mai_mai_n470_), .A1(mai_mai_n356_), .B0(mai_mai_n1010_), .Y(mai_mai_n1011_));
  OR3        m0983(.A(mai_mai_n879_), .B(mai_mai_n240_), .C(mai_mai_n202_), .Y(mai_mai_n1012_));
  NO2        m0984(.A(mai_mai_n196_), .B(mai_mai_n193_), .Y(mai_mai_n1013_));
  INV        m0985(.A(mai_mai_n135_), .Y(mai_mai_n1014_));
  AOI220     m0986(.A0(mai_mai_n1014_), .A1(mai_mai_n242_), .B0(mai_mai_n718_), .B1(mai_mai_n1013_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n306_), .B(mai_mai_n383_), .Y(mai_mai_n1016_));
  NA4        m0988(.A(mai_mai_n1016_), .B(mai_mai_n1015_), .C(mai_mai_n1012_), .D(mai_mai_n1011_), .Y(mai_mai_n1017_));
  INV        m0989(.A(mai_mai_n691_), .Y(mai_mai_n1018_));
  NO2        m0990(.A(mai_mai_n59_), .B(h), .Y(mai_mai_n1019_));
  NO3        m0991(.A(mai_mai_n879_), .B(f), .C(mai_mai_n606_), .Y(mai_mai_n1020_));
  OAI210     m0992(.A0(mai_mai_n924_), .A1(mai_mai_n1020_), .B0(mai_mai_n1019_), .Y(mai_mai_n1021_));
  NA3        m0993(.A(mai_mai_n1021_), .B(mai_mai_n1018_), .C(mai_mai_n734_), .Y(mai_mai_n1022_));
  NO4        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1017_), .C(mai_mai_n257_), .D(mai_mai_n1009_), .Y(mai_mai_n1023_));
  NA2        m0995(.A(mai_mai_n707_), .B(mai_mai_n631_), .Y(mai_mai_n1024_));
  NA4        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1023_), .C(mai_mai_n1006_), .D(mai_mai_n979_), .Y(mai01));
  NO4        m0997(.A(mai_mai_n674_), .B(mai_mai_n666_), .C(mai_mai_n401_), .D(mai_mai_n248_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n344_), .B(i), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n1027_), .B(mai_mai_n1026_), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n775_), .B(mai_mai_n289_), .Y(mai_mai_n1029_));
  NA2        m1001(.A(mai_mai_n588_), .B(g), .Y(mai_mai_n1030_));
  NO2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1219_), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n1031_), .B(mai_mai_n532_), .Y(mai_mai_n1032_));
  INV        m1004(.A(mai_mai_n107_), .Y(mai_mai_n1033_));
  OA220      m1005(.A0(mai_mai_n1033_), .A1(mai_mai_n487_), .B0(mai_mai_n550_), .B1(mai_mai_n319_), .Y(mai_mai_n1034_));
  NAi41      m1006(.An(mai_mai_n150_), .B(mai_mai_n1034_), .C(mai_mai_n1032_), .D(mai_mai_n760_), .Y(mai_mai_n1035_));
  NO2        m1007(.A(mai_mai_n560_), .B(mai_mai_n430_), .Y(mai_mai_n1036_));
  NA4        m1008(.A(mai_mai_n588_), .B(g), .C(mai_mai_n43_), .D(mai_mai_n192_), .Y(mai_mai_n1037_));
  OA220      m1009(.A0(mai_mai_n1037_), .A1(mai_mai_n555_), .B0(mai_mai_n177_), .B1(mai_mai_n175_), .Y(mai_mai_n1038_));
  NA3        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .C(mai_mai_n125_), .Y(mai_mai_n1039_));
  NO4        m1011(.A(mai_mai_n1039_), .B(mai_mai_n1035_), .C(mai_mai_n1029_), .D(mai_mai_n1028_), .Y(mai_mai_n1040_));
  INV        m1012(.A(mai_mai_n985_), .Y(mai_mai_n1041_));
  NA2        m1013(.A(mai_mai_n1041_), .B(mai_mai_n448_), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n455_), .B(mai_mai_n346_), .Y(mai_mai_n1043_));
  NOi21      m1015(.An(mai_mai_n472_), .B(mai_mai_n486_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n1044_), .B(mai_mai_n1043_), .Y(mai_mai_n1045_));
  AOI210     m1017(.A0(mai_mai_n186_), .A1(mai_mai_n80_), .B0(mai_mai_n192_), .Y(mai_mai_n1046_));
  OAI210     m1018(.A0(mai_mai_n681_), .A1(mai_mai_n367_), .B0(mai_mai_n1046_), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n308_), .B(k), .Y(mai_mai_n1048_));
  OR2        m1020(.A(mai_mai_n1048_), .B(mai_mai_n288_), .Y(mai_mai_n1049_));
  NA4        m1021(.A(mai_mai_n1049_), .B(mai_mai_n1047_), .C(mai_mai_n1045_), .D(mai_mai_n1042_), .Y(mai_mai_n1050_));
  AOI210     m1022(.A0(mai_mai_n496_), .A1(mai_mai_n107_), .B0(mai_mai_n499_), .Y(mai_mai_n1051_));
  OAI210     m1023(.A0(mai_mai_n1033_), .A1(mai_mai_n493_), .B0(mai_mai_n1051_), .Y(mai_mai_n1052_));
  NO2        m1024(.A(mai_mai_n690_), .B(mai_mai_n186_), .Y(mai_mai_n1053_));
  INV        m1025(.A(mai_mai_n1053_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n282_), .B(mai_mai_n561_), .Y(mai_mai_n1055_));
  NA3        m1027(.A(mai_mai_n1055_), .B(mai_mai_n1054_), .C(mai_mai_n658_), .Y(mai_mai_n1056_));
  NO3        m1028(.A(mai_mai_n1056_), .B(mai_mai_n1052_), .C(mai_mai_n1050_), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n501_), .B(f), .Y(mai_mai_n1058_));
  NO2        m1030(.A(mai_mai_n1058_), .B(mai_mai_n186_), .Y(mai_mai_n1059_));
  AOI210     m1031(.A0(mai_mai_n427_), .A1(mai_mai_n54_), .B0(mai_mai_n1059_), .Y(mai_mai_n1060_));
  NO2        m1032(.A(mai_mai_n1037_), .B(mai_mai_n824_), .Y(mai_mai_n1061_));
  NO2        m1033(.A(mai_mai_n187_), .B(mai_mai_n100_), .Y(mai_mai_n1062_));
  NO3        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1061_), .C(mai_mai_n982_), .Y(mai_mai_n1063_));
  NA3        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1060_), .C(mai_mai_n630_), .Y(mai_mai_n1064_));
  NO2        m1036(.A(mai_mai_n816_), .B(mai_mai_n212_), .Y(mai_mai_n1065_));
  NO3        m1037(.A(mai_mai_n70_), .B(mai_mai_n262_), .C(mai_mai_n43_), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n1066_), .B(mai_mai_n466_), .Y(mai_mai_n1067_));
  NA2        m1039(.A(mai_mai_n1067_), .B(mai_mai_n557_), .Y(mai_mai_n1068_));
  NO2        m1040(.A(mai_mai_n319_), .B(mai_mai_n63_), .Y(mai_mai_n1069_));
  INV        m1041(.A(mai_mai_n1069_), .Y(mai_mai_n1070_));
  NA2        m1042(.A(mai_mai_n1066_), .B(n), .Y(mai_mai_n1071_));
  NA3        m1043(.A(mai_mai_n1071_), .B(mai_mai_n1070_), .C(mai_mai_n336_), .Y(mai_mai_n1072_));
  NO3        m1044(.A(mai_mai_n1072_), .B(mai_mai_n1068_), .C(mai_mai_n1064_), .Y(mai_mai_n1073_));
  NO3        m1045(.A(mai_mai_n922_), .B(mai_mai_n163_), .C(mai_mai_n78_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n511_), .B(mai_mai_n510_), .Y(mai_mai_n1075_));
  NO4        m1047(.A(mai_mai_n922_), .B(mai_mai_n1075_), .C(mai_mai_n161_), .D(mai_mai_n78_), .Y(mai_mai_n1076_));
  NO3        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1074_), .C(mai_mai_n534_), .Y(mai_mai_n1077_));
  NA4        m1049(.A(mai_mai_n1077_), .B(mai_mai_n1073_), .C(mai_mai_n1057_), .D(mai_mai_n1040_), .Y(mai06));
  NO2        m1050(.A(mai_mai_n204_), .B(mai_mai_n92_), .Y(mai_mai_n1079_));
  OAI210     m1051(.A0(mai_mai_n1079_), .A1(mai_mai_n1074_), .B0(mai_mai_n332_), .Y(mai_mai_n1080_));
  NA2        m1052(.A(mai_mai_n750_), .B(mai_mai_n1080_), .Y(mai_mai_n1081_));
  NO3        m1053(.A(mai_mai_n1081_), .B(mai_mai_n1068_), .C(mai_mai_n232_), .Y(mai_mai_n1082_));
  NO2        m1054(.A(mai_mai_n1222_), .B(mai_mai_n292_), .Y(mai_mai_n1083_));
  NO2        m1055(.A(mai_mai_n80_), .B(mai_mai_n40_), .Y(mai_mai_n1084_));
  NA2        m1056(.A(mai_mai_n1084_), .B(mai_mai_n537_), .Y(mai_mai_n1085_));
  NO2        m1057(.A(mai_mai_n433_), .B(mai_mai_n158_), .Y(mai_mai_n1086_));
  NOi21      m1058(.An(mai_mai_n124_), .B(mai_mai_n43_), .Y(mai_mai_n1087_));
  NO2        m1059(.A(mai_mai_n504_), .B(mai_mai_n941_), .Y(mai_mai_n1088_));
  NO3        m1060(.A(mai_mai_n1088_), .B(mai_mai_n1087_), .C(mai_mai_n1086_), .Y(mai_mai_n1089_));
  INV        m1061(.A(mai_mai_n499_), .Y(mai_mai_n1090_));
  NA3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1089_), .C(mai_mai_n1085_), .Y(mai_mai_n1091_));
  NO2        m1063(.A(mai_mai_n623_), .B(mai_mai_n317_), .Y(mai_mai_n1092_));
  NOi21      m1064(.An(mai_mai_n1092_), .B(mai_mai_n46_), .Y(mai_mai_n1093_));
  BUFFER     m1065(.A(mai_mai_n810_), .Y(mai_mai_n1094_));
  NO4        m1066(.A(mai_mai_n1094_), .B(mai_mai_n1093_), .C(mai_mai_n1091_), .D(mai_mai_n1083_), .Y(mai_mai_n1095_));
  NO2        m1067(.A(mai_mai_n673_), .B(mai_mai_n244_), .Y(mai_mai_n1096_));
  OAI220     m1068(.A0(mai_mai_n611_), .A1(mai_mai_n45_), .B0(mai_mai_n204_), .B1(mai_mai_n513_), .Y(mai_mai_n1097_));
  OAI210     m1069(.A0(mai_mai_n244_), .A1(c), .B0(mai_mai_n536_), .Y(mai_mai_n1098_));
  AOI220     m1070(.A0(mai_mai_n1098_), .A1(mai_mai_n1097_), .B0(mai_mai_n1096_), .B1(mai_mai_n236_), .Y(mai_mai_n1099_));
  NO3        m1071(.A(h), .B(mai_mai_n92_), .C(mai_mai_n250_), .Y(mai_mai_n1100_));
  OAI220     m1072(.A0(mai_mai_n580_), .A1(mai_mai_n225_), .B0(mai_mai_n429_), .B1(mai_mai_n433_), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n498_), .B(j), .Y(mai_mai_n1102_));
  NOi21      m1074(.An(mai_mai_n1102_), .B(mai_mai_n555_), .Y(mai_mai_n1103_));
  NO4        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1101_), .C(mai_mai_n1100_), .D(mai_mai_n944_), .Y(mai_mai_n1104_));
  NAi31      m1076(.An(mai_mai_n623_), .B(mai_mai_n75_), .C(mai_mai_n185_), .Y(mai_mai_n1105_));
  NA3        m1077(.A(mai_mai_n1105_), .B(mai_mai_n1104_), .C(mai_mai_n1099_), .Y(mai_mai_n1106_));
  OR2        m1078(.A(mai_mai_n655_), .B(mai_mai_n457_), .Y(mai_mai_n1107_));
  AOI210     m1079(.A0(g), .A1(mai_mai_n383_), .B0(mai_mai_n322_), .Y(mai_mai_n1108_));
  NA2        m1080(.A(mai_mai_n1102_), .B(mai_mai_n661_), .Y(mai_mai_n1109_));
  NA3        m1081(.A(mai_mai_n1109_), .B(mai_mai_n1108_), .C(mai_mai_n1107_), .Y(mai_mai_n1110_));
  NO3        m1082(.A(mai_mai_n743_), .B(mai_mai_n423_), .C(mai_mai_n404_), .Y(mai_mai_n1111_));
  NA2        m1083(.A(mai_mai_n1111_), .B(mai_mai_n1071_), .Y(mai_mai_n1112_));
  NAi21      m1084(.An(j), .B(i), .Y(mai_mai_n1113_));
  NO4        m1085(.A(mai_mai_n1075_), .B(mai_mai_n1113_), .C(mai_mai_n379_), .D(mai_mai_n215_), .Y(mai_mai_n1114_));
  NO4        m1086(.A(mai_mai_n1114_), .B(mai_mai_n1112_), .C(mai_mai_n1110_), .D(mai_mai_n1106_), .Y(mai_mai_n1115_));
  NA4        m1087(.A(mai_mai_n1115_), .B(mai_mai_n1095_), .C(mai_mai_n1082_), .D(mai_mai_n1077_), .Y(mai07));
  NAi21      m1088(.An(f), .B(c), .Y(mai_mai_n1117_));
  OR2        m1089(.A(e), .B(d), .Y(mai_mai_n1118_));
  OAI220     m1090(.A0(mai_mai_n1118_), .A1(mai_mai_n1117_), .B0(mai_mai_n524_), .B1(mai_mai_n279_), .Y(mai_mai_n1119_));
  NA3        m1091(.A(mai_mai_n1119_), .B(mai_mai_n1220_), .C(mai_mai_n166_), .Y(mai_mai_n1120_));
  NOi31      m1092(.An(n), .B(m), .C(b), .Y(mai_mai_n1121_));
  NO3        m1093(.A(mai_mai_n119_), .B(mai_mai_n384_), .C(h), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n78_), .B(mai_mai_n43_), .Y(mai_mai_n1123_));
  NO2        m1095(.A(mai_mai_n897_), .B(mai_mai_n269_), .Y(mai_mai_n1124_));
  NO2        m1096(.A(l), .B(k), .Y(mai_mai_n1125_));
  NOi41      m1097(.An(mai_mai_n461_), .B(mai_mai_n1125_), .C(mai_mai_n399_), .D(mai_mai_n379_), .Y(mai_mai_n1126_));
  NO2        m1098(.A(g), .B(c), .Y(mai_mai_n1127_));
  NO2        m1099(.A(mai_mai_n385_), .B(a), .Y(mai_mai_n1128_));
  NA3        m1100(.A(mai_mai_n1128_), .B(k), .C(mai_mai_n102_), .Y(mai_mai_n1129_));
  NO2        m1101(.A(i), .B(h), .Y(mai_mai_n1130_));
  NA2        m1102(.A(mai_mai_n961_), .B(h), .Y(mai_mai_n1131_));
  NA2        m1103(.A(mai_mai_n126_), .B(mai_mai_n200_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1131_), .Y(mai_mai_n1133_));
  NOi31      m1105(.An(m), .B(n), .C(b), .Y(mai_mai_n1134_));
  INV        m1106(.A(mai_mai_n1133_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n915_), .B(mai_mai_n395_), .Y(mai_mai_n1136_));
  NO4        m1108(.A(mai_mai_n1136_), .B(mai_mai_n892_), .C(mai_mai_n379_), .D(mai_mai_n43_), .Y(mai_mai_n1137_));
  OAI210     m1109(.A0(mai_mai_n169_), .A1(mai_mai_n443_), .B0(mai_mai_n893_), .Y(mai_mai_n1138_));
  INV        m1110(.A(mai_mai_n1138_), .Y(mai_mai_n1139_));
  NO2        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1137_), .Y(mai_mai_n1140_));
  AN3        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1135_), .C(mai_mai_n1129_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(mai_mai_n1121_), .B(mai_mai_n329_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n923_), .B(mai_mai_n1136_), .Y(mai_mai_n1143_));
  NO4        m1115(.A(mai_mai_n119_), .B(g), .C(f), .D(e), .Y(mai_mai_n1144_));
  OR2        m1116(.A(e), .B(a), .Y(mai_mai_n1145_));
  NA2        m1117(.A(mai_mai_n940_), .B(mai_mai_n354_), .Y(mai_mai_n1146_));
  NA4        m1118(.A(mai_mai_n1143_), .B(mai_mai_n1141_), .C(mai_mai_n1233_), .D(mai_mai_n1120_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n341_), .B(j), .Y(mai_mai_n1148_));
  NAi31      m1120(.An(mai_mai_n1130_), .B(mai_mai_n905_), .C(mai_mai_n154_), .Y(mai_mai_n1149_));
  INV        m1121(.A(mai_mai_n1149_), .Y(mai_mai_n1150_));
  NA3        m1122(.A(g), .B(mai_mai_n1148_), .C(mai_mai_n147_), .Y(mai_mai_n1151_));
  INV        m1123(.A(mai_mai_n1151_), .Y(mai_mai_n1152_));
  NO3        m1124(.A(mai_mai_n623_), .B(mai_mai_n161_), .C(e), .Y(mai_mai_n1153_));
  NO3        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1152_), .C(mai_mai_n1150_), .Y(mai_mai_n1154_));
  INV        m1126(.A(mai_mai_n46_), .Y(mai_mai_n1155_));
  AOI220     m1127(.A0(mai_mai_n1155_), .A1(mai_mai_n987_), .B0(mai_mai_n695_), .B1(mai_mai_n176_), .Y(mai_mai_n1156_));
  NO2        m1128(.A(mai_mai_n911_), .B(h), .Y(mai_mai_n1157_));
  NA2        m1129(.A(mai_mai_n166_), .B(mai_mai_n101_), .Y(mai_mai_n1158_));
  NOi21      m1130(.An(d), .B(f), .Y(mai_mai_n1159_));
  NO2        m1131(.A(mai_mai_n1118_), .B(f), .Y(mai_mai_n1160_));
  NA2        m1132(.A(mai_mai_n1156_), .B(mai_mai_n1154_), .Y(mai_mai_n1161_));
  NO3        m1133(.A(mai_mai_n915_), .B(mai_mai_n904_), .C(mai_mai_n40_), .Y(mai_mai_n1162_));
  NA2        m1134(.A(mai_mai_n1162_), .B(mai_mai_n1124_), .Y(mai_mai_n1163_));
  OAI210     m1135(.A0(mai_mai_n1144_), .A1(mai_mai_n1121_), .B0(mai_mai_n749_), .Y(mai_mai_n1164_));
  OAI220     m1136(.A0(mai_mai_n875_), .A1(mai_mai_n119_), .B0(h), .B1(mai_mai_n161_), .Y(mai_mai_n1165_));
  NA2        m1137(.A(mai_mai_n1165_), .B(mai_mai_n517_), .Y(mai_mai_n1166_));
  NA3        m1138(.A(mai_mai_n1166_), .B(mai_mai_n1164_), .C(mai_mai_n1163_), .Y(mai_mai_n1167_));
  NA2        m1139(.A(mai_mai_n1127_), .B(mai_mai_n1159_), .Y(mai_mai_n1168_));
  NO2        m1140(.A(mai_mai_n1168_), .B(m), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n139_), .B(mai_mai_n168_), .Y(mai_mai_n1170_));
  OAI210     m1142(.A0(mai_mai_n1170_), .A1(mai_mai_n99_), .B0(mai_mai_n1134_), .Y(mai_mai_n1171_));
  INV        m1143(.A(mai_mai_n1171_), .Y(mai_mai_n1172_));
  NO3        m1144(.A(mai_mai_n1172_), .B(mai_mai_n1169_), .C(mai_mai_n1167_), .Y(mai_mai_n1173_));
  NO2        m1145(.A(mai_mai_n1117_), .B(e), .Y(mai_mai_n1174_));
  OAI210     m1146(.A0(mai_mai_n1160_), .A1(mai_mai_n949_), .B0(mai_mai_n528_), .Y(mai_mai_n1175_));
  NO2        m1147(.A(mai_mai_n1175_), .B(mai_mai_n381_), .Y(mai_mai_n1176_));
  INV        m1148(.A(mai_mai_n1176_), .Y(mai_mai_n1177_));
  NO2        m1149(.A(mai_mai_n168_), .B(c), .Y(mai_mai_n1178_));
  OAI210     m1150(.A0(mai_mai_n1178_), .A1(mai_mai_n1174_), .B0(mai_mai_n166_), .Y(mai_mai_n1179_));
  AOI220     m1151(.A0(mai_mai_n1179_), .A1(mai_mai_n906_), .B0(mai_mai_n449_), .B1(mai_mai_n317_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n1145_), .B(f), .Y(mai_mai_n1181_));
  AOI210     m1153(.A0(mai_mai_n763_), .A1(mai_mai_n359_), .B0(mai_mai_n94_), .Y(mai_mai_n1182_));
  NA2        m1154(.A(mai_mai_n1181_), .B(mai_mai_n1123_), .Y(mai_mai_n1183_));
  OAI220     m1155(.A0(mai_mai_n1183_), .A1(mai_mai_n46_), .B0(mai_mai_n1182_), .B1(mai_mai_n161_), .Y(mai_mai_n1184_));
  NA2        m1156(.A(mai_mai_n1122_), .B(mai_mai_n169_), .Y(mai_mai_n1185_));
  NO2        m1157(.A(mai_mai_n46_), .B(l), .Y(mai_mai_n1186_));
  OAI210     m1158(.A0(mai_mai_n1145_), .A1(mai_mai_n728_), .B0(mai_mai_n406_), .Y(mai_mai_n1187_));
  OAI210     m1159(.A0(mai_mai_n1187_), .A1(mai_mai_n927_), .B0(mai_mai_n1186_), .Y(mai_mai_n1188_));
  NO2        m1160(.A(mai_mai_n228_), .B(g), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n905_), .B(mai_mai_n1189_), .Y(mai_mai_n1190_));
  NA3        m1162(.A(mai_mai_n1190_), .B(mai_mai_n1188_), .C(mai_mai_n1185_), .Y(mai_mai_n1191_));
  NO3        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1184_), .C(mai_mai_n1180_), .Y(mai_mai_n1192_));
  NA3        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1177_), .C(mai_mai_n1173_), .Y(mai_mai_n1193_));
  NO2        m1165(.A(mai_mai_n486_), .B(g), .Y(mai_mai_n1194_));
  NA2        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1157_), .Y(mai_mai_n1195_));
  AO210      m1167(.A0(mai_mai_n120_), .A1(l), .B0(mai_mai_n1142_), .Y(mai_mai_n1196_));
  NA2        m1168(.A(mai_mai_n1196_), .B(mai_mai_n1195_), .Y(mai_mai_n1197_));
  INV        m1169(.A(mai_mai_n1197_), .Y(mai_mai_n1198_));
  AOI210     m1170(.A0(mai_mai_n145_), .A1(mai_mai_n52_), .B0(mai_mai_n1174_), .Y(mai_mai_n1199_));
  NO2        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1158_), .Y(mai_mai_n1200_));
  NOi21      m1172(.An(mai_mai_n1122_), .B(e), .Y(mai_mai_n1201_));
  NO2        m1173(.A(mai_mai_n1201_), .B(mai_mai_n1200_), .Y(mai_mai_n1202_));
  NA2        m1174(.A(mai_mai_n55_), .B(a), .Y(mai_mai_n1203_));
  NO2        m1175(.A(mai_mai_n1146_), .B(mai_mai_n1203_), .Y(mai_mai_n1204_));
  INV        m1176(.A(mai_mai_n1204_), .Y(mai_mai_n1205_));
  NA3        m1177(.A(mai_mai_n1205_), .B(mai_mai_n1202_), .C(mai_mai_n1198_), .Y(mai_mai_n1206_));
  OR4        m1178(.A(mai_mai_n1206_), .B(mai_mai_n1193_), .C(mai_mai_n1161_), .D(mai_mai_n1147_), .Y(mai04));
  NOi21      m1179(.An(mai_mai_n1144_), .B(mai_mai_n879_), .Y(mai_mai_n1208_));
  NA2        m1180(.A(mai_mai_n1160_), .B(mai_mai_n695_), .Y(mai_mai_n1209_));
  NO2        m1181(.A(mai_mai_n1209_), .B(mai_mai_n872_), .Y(mai_mai_n1210_));
  OR3        m1182(.A(mai_mai_n1210_), .B(mai_mai_n1208_), .C(mai_mai_n895_), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n82_), .B(k), .Y(mai_mai_n1212_));
  AOI210     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n889_), .B0(mai_mai_n1000_), .Y(mai_mai_n1213_));
  NA2        m1185(.A(mai_mai_n1213_), .B(mai_mai_n1021_), .Y(mai_mai_n1214_));
  NO4        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1211_), .C(mai_mai_n903_), .D(mai_mai_n884_), .Y(mai_mai_n1215_));
  NA4        m1187(.A(mai_mai_n1215_), .B(mai_mai_n951_), .C(mai_mai_n938_), .D(mai_mai_n930_), .Y(mai05));
  INV        m1188(.A(f), .Y(mai_mai_n1219_));
  INV        m1189(.A(j), .Y(mai_mai_n1220_));
  INV        m1190(.A(j), .Y(mai_mai_n1221_));
  INV        m1191(.A(mai_mai_n1065_), .Y(mai_mai_n1222_));
  INV        m1192(.A(mai_mai_n805_), .Y(mai_mai_n1223_));
  INV        m1193(.A(g), .Y(mai_mai_n1224_));
  INV        m1194(.A(c), .Y(mai_mai_n1225_));
  INV        m1195(.A(l), .Y(mai_mai_n1226_));
  INV        m1196(.A(h), .Y(mai_mai_n1227_));
  INV        m1197(.A(m), .Y(mai_mai_n1228_));
  INV        m1198(.A(mai_mai_n102_), .Y(mai_mai_n1229_));
  INV        m1199(.A(e), .Y(mai_mai_n1230_));
  INV        m1200(.A(m), .Y(mai_mai_n1231_));
  INV        m1201(.A(f), .Y(mai_mai_n1232_));
  INV        m1202(.A(mai_mai_n1126_), .Y(mai_mai_n1233_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NAi21      u0031(.An(i), .B(h), .Y(men_men_n60_));
  NAi31      u0032(.An(i), .B(l), .C(j), .Y(men_men_n61_));
  OAI220     u0033(.A0(men_men_n61_), .A1(men_men_n49_), .B0(men_men_n60_), .B1(men_men_n44_), .Y(men_men_n62_));
  NAi31      u0034(.An(d), .B(men_men_n62_), .C(men_men_n58_), .Y(men_men_n63_));
  NAi41      u0035(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n64_));
  NA2        u0036(.A(g), .B(f), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi21      u0038(.An(i), .B(j), .Y(men_men_n67_));
  NAi32      u0039(.An(n), .Bn(k), .C(m), .Y(men_men_n68_));
  NO2        u0040(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi31      u0041(.An(l), .B(m), .C(k), .Y(men_men_n70_));
  NAi21      u0042(.An(e), .B(h), .Y(men_men_n71_));
  NAi41      u0043(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n73_));
  INV        u0045(.A(m), .Y(men_men_n74_));
  NOi21      u0046(.An(k), .B(l), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  AN4        u0048(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n77_));
  NOi31      u0049(.An(h), .B(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n77_), .Y(men_men_n79_));
  NAi32      u0051(.An(m), .Bn(k), .C(j), .Y(men_men_n80_));
  NOi32      u0052(.An(h), .Bn(g), .C(f), .Y(men_men_n81_));
  NA2        u0053(.A(men_men_n81_), .B(men_men_n77_), .Y(men_men_n82_));
  OA220      u0054(.A0(men_men_n82_), .A1(men_men_n80_), .B0(men_men_n79_), .B1(men_men_n76_), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n73_), .C(men_men_n63_), .Y(men_men_n84_));
  INV        u0056(.A(n), .Y(men_men_n85_));
  NOi32      u0057(.An(e), .Bn(b), .C(d), .Y(men_men_n86_));
  NA2        u0058(.A(men_men_n86_), .B(men_men_n85_), .Y(men_men_n87_));
  INV        u0059(.A(j), .Y(men_men_n88_));
  AN3        u0060(.A(m), .B(k), .C(i), .Y(men_men_n89_));
  NA3        u0061(.A(men_men_n89_), .B(men_men_n88_), .C(g), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(f), .Y(men_men_n91_));
  NAi32      u0063(.An(g), .Bn(f), .C(h), .Y(men_men_n92_));
  NAi31      u0064(.An(j), .B(m), .C(l), .Y(men_men_n93_));
  NO2        u0065(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NA2        u0066(.A(m), .B(l), .Y(men_men_n95_));
  NAi31      u0067(.An(k), .B(j), .C(g), .Y(men_men_n96_));
  NO3        u0068(.A(men_men_n96_), .B(men_men_n95_), .C(f), .Y(men_men_n97_));
  AN2        u0069(.A(j), .B(g), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(l), .C(i), .Y(men_men_n99_));
  NOi21      u0071(.An(g), .B(i), .Y(men_men_n100_));
  NOi32      u0072(.An(m), .Bn(j), .C(k), .Y(men_men_n101_));
  AOI220     u0073(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n99_), .B1(men_men_n98_), .Y(men_men_n102_));
  NO2        u0074(.A(men_men_n102_), .B(f), .Y(men_men_n103_));
  NO4        u0075(.A(men_men_n103_), .B(men_men_n97_), .C(men_men_n94_), .D(men_men_n91_), .Y(men_men_n104_));
  NAi41      u0076(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n105_));
  AN2        u0077(.A(e), .B(b), .Y(men_men_n106_));
  NOi31      u0078(.An(c), .B(h), .C(f), .Y(men_men_n107_));
  NA2        u0079(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NOi21      u0080(.An(g), .B(f), .Y(men_men_n109_));
  NOi21      u0081(.An(i), .B(h), .Y(men_men_n110_));
  NA3        u0082(.A(men_men_n110_), .B(men_men_n109_), .C(men_men_n36_), .Y(men_men_n111_));
  INV        u0083(.A(a), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n106_), .B(men_men_n112_), .Y(men_men_n113_));
  INV        u0085(.A(l), .Y(men_men_n114_));
  NOi21      u0086(.An(m), .B(n), .Y(men_men_n115_));
  NO2        u0087(.A(men_men_n111_), .B(men_men_n87_), .Y(men_men_n116_));
  INV        u0088(.A(b), .Y(men_men_n117_));
  NA2        u0089(.A(l), .B(j), .Y(men_men_n118_));
  AN2        u0090(.A(k), .B(i), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u0092(.A(g), .B(e), .Y(men_men_n121_));
  NOi32      u0093(.An(c), .Bn(a), .C(d), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n115_), .Y(men_men_n123_));
  NO4        u0095(.A(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n124_));
  NO2        u0096(.A(men_men_n124_), .B(men_men_n116_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n104_), .A1(men_men_n87_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n78_), .C(men_men_n77_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(i), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n81_), .C(men_men_n77_), .Y(men_men_n130_));
  NA2        u0102(.A(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NOi32      u0103(.An(f), .Bn(b), .C(e), .Y(men_men_n132_));
  NAi21      u0104(.An(g), .B(h), .Y(men_men_n133_));
  NAi21      u0105(.An(m), .B(n), .Y(men_men_n134_));
  NAi21      u0106(.An(j), .B(k), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n136_));
  NAi41      u0108(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n137_));
  NAi31      u0109(.An(j), .B(k), .C(h), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n139_));
  AOI210     u0111(.A0(men_men_n136_), .A1(men_men_n132_), .B0(men_men_n139_), .Y(men_men_n140_));
  NO2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  INV        u0113(.A(men_men_n134_), .Y(men_men_n142_));
  AN2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  NAi21      u0115(.An(c), .B(b), .Y(men_men_n144_));
  NA2        u0116(.A(f), .B(d), .Y(men_men_n145_));
  NO4        u0117(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .D(men_men_n133_), .Y(men_men_n146_));
  NA2        u0118(.A(h), .B(c), .Y(men_men_n147_));
  NAi31      u0119(.An(f), .B(e), .C(b), .Y(men_men_n148_));
  NA2        u0120(.A(men_men_n146_), .B(men_men_n142_), .Y(men_men_n149_));
  NA2        u0121(.A(d), .B(b), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(f), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NA2        u0124(.A(b), .B(a), .Y(men_men_n153_));
  NAi21      u0125(.An(c), .B(d), .Y(men_men_n154_));
  NAi31      u0126(.An(l), .B(k), .C(h), .Y(men_men_n155_));
  NO2        u0127(.A(men_men_n134_), .B(men_men_n155_), .Y(men_men_n156_));
  NA2        u0128(.A(men_men_n156_), .B(men_men_n152_), .Y(men_men_n157_));
  NAi41      u0129(.An(men_men_n131_), .B(men_men_n157_), .C(men_men_n149_), .D(men_men_n140_), .Y(men_men_n158_));
  NAi31      u0130(.An(e), .B(f), .C(b), .Y(men_men_n159_));
  NOi21      u0131(.An(g), .B(d), .Y(men_men_n160_));
  NO2        u0132(.A(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0133(.An(h), .B(i), .Y(men_men_n162_));
  NOi21      u0134(.An(k), .B(m), .Y(men_men_n163_));
  NA3        u0135(.A(men_men_n163_), .B(men_men_n162_), .C(n), .Y(men_men_n164_));
  NOi21      u0136(.An(men_men_n161_), .B(men_men_n164_), .Y(men_men_n165_));
  NOi21      u0137(.An(h), .B(g), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  NAi31      u0140(.An(l), .B(j), .C(h), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n169_), .B(men_men_n49_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n66_), .Y(men_men_n171_));
  NOi32      u0143(.An(n), .Bn(k), .C(m), .Y(men_men_n172_));
  NA2        u0144(.A(l), .B(i), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OAI210     u0146(.A0(men_men_n174_), .A1(men_men_n168_), .B0(men_men_n171_), .Y(men_men_n175_));
  NAi31      u0147(.An(e), .B(f), .C(c), .Y(men_men_n176_));
  NA2        u0148(.A(j), .B(h), .Y(men_men_n177_));
  OR3        u0149(.A(n), .B(m), .C(k), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n177_), .Y(men_men_n179_));
  NAi32      u0151(.An(m), .Bn(k), .C(n), .Y(men_men_n180_));
  NO2        u0152(.A(men_men_n180_), .B(men_men_n177_), .Y(men_men_n181_));
  AOI220     u0153(.A0(men_men_n181_), .A1(men_men_n161_), .B0(men_men_n179_), .B1(f), .Y(men_men_n182_));
  NO2        u0154(.A(n), .B(m), .Y(men_men_n183_));
  NA2        u0155(.A(men_men_n183_), .B(men_men_n50_), .Y(men_men_n184_));
  NAi21      u0156(.An(f), .B(e), .Y(men_men_n185_));
  NA2        u0157(.A(d), .B(c), .Y(men_men_n186_));
  NOi21      u0158(.An(c), .B(men_men_n184_), .Y(men_men_n187_));
  NAi21      u0159(.An(d), .B(c), .Y(men_men_n188_));
  NAi31      u0160(.An(m), .B(n), .C(b), .Y(men_men_n189_));
  NA2        u0161(.A(k), .B(i), .Y(men_men_n190_));
  NAi21      u0162(.An(h), .B(f), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NO2        u0164(.A(men_men_n189_), .B(men_men_n154_), .Y(men_men_n193_));
  NA2        u0165(.A(men_men_n193_), .B(men_men_n192_), .Y(men_men_n194_));
  NOi32      u0166(.An(f), .Bn(c), .C(e), .Y(men_men_n195_));
  NO3        u0167(.A(n), .B(m), .C(j), .Y(men_men_n196_));
  NA2        u0168(.A(men_men_n196_), .B(k), .Y(men_men_n197_));
  NAi31      u0169(.An(men_men_n187_), .B(men_men_n194_), .C(men_men_n182_), .Y(men_men_n198_));
  OR4        u0170(.A(men_men_n198_), .B(men_men_n175_), .C(men_men_n165_), .D(men_men_n158_), .Y(men_men_n199_));
  NO4        u0171(.A(men_men_n199_), .B(men_men_n126_), .C(men_men_n84_), .D(men_men_n55_), .Y(men_men_n200_));
  NA3        u0172(.A(m), .B(men_men_n114_), .C(j), .Y(men_men_n201_));
  NAi31      u0173(.An(n), .B(h), .C(g), .Y(men_men_n202_));
  NO2        u0174(.A(men_men_n202_), .B(men_men_n201_), .Y(men_men_n203_));
  NOi32      u0175(.An(m), .Bn(k), .C(l), .Y(men_men_n204_));
  NA3        u0176(.A(men_men_n204_), .B(men_men_n88_), .C(g), .Y(men_men_n205_));
  NO2        u0177(.A(men_men_n205_), .B(n), .Y(men_men_n206_));
  NOi21      u0178(.An(k), .B(j), .Y(men_men_n207_));
  NA4        u0179(.A(men_men_n207_), .B(men_men_n115_), .C(i), .D(g), .Y(men_men_n208_));
  AN2        u0180(.A(i), .B(g), .Y(men_men_n209_));
  NA3        u0181(.A(men_men_n75_), .B(men_men_n209_), .C(men_men_n115_), .Y(men_men_n210_));
  NA2        u0182(.A(men_men_n210_), .B(men_men_n208_), .Y(men_men_n211_));
  NO3        u0183(.A(men_men_n211_), .B(men_men_n206_), .C(men_men_n203_), .Y(men_men_n212_));
  NAi41      u0184(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n213_));
  INV        u0185(.A(men_men_n213_), .Y(men_men_n214_));
  INV        u0186(.A(f), .Y(men_men_n215_));
  INV        u0187(.A(g), .Y(men_men_n216_));
  NOi31      u0188(.An(i), .B(j), .C(h), .Y(men_men_n217_));
  NOi21      u0189(.An(l), .B(m), .Y(men_men_n218_));
  NA2        u0190(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n219_));
  NO3        u0191(.A(men_men_n219_), .B(men_men_n216_), .C(men_men_n215_), .Y(men_men_n220_));
  NA2        u0192(.A(men_men_n220_), .B(men_men_n214_), .Y(men_men_n221_));
  OAI210     u0193(.A0(men_men_n212_), .A1(men_men_n32_), .B0(men_men_n221_), .Y(men_men_n222_));
  NOi21      u0194(.An(n), .B(m), .Y(men_men_n223_));
  NA2        u0195(.A(i), .B(men_men_n223_), .Y(men_men_n224_));
  OA220      u0196(.A0(men_men_n224_), .A1(men_men_n108_), .B0(men_men_n80_), .B1(men_men_n79_), .Y(men_men_n225_));
  NAi21      u0197(.An(j), .B(h), .Y(men_men_n226_));
  XN2        u0198(.A(i), .B(h), .Y(men_men_n227_));
  NOi31      u0199(.An(k), .B(n), .C(m), .Y(men_men_n228_));
  NAi31      u0200(.An(f), .B(e), .C(c), .Y(men_men_n229_));
  NA4        u0201(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n230_));
  NAi32      u0202(.An(m), .Bn(i), .C(k), .Y(men_men_n231_));
  NO3        u0203(.A(men_men_n231_), .B(men_men_n92_), .C(men_men_n230_), .Y(men_men_n232_));
  INV        u0204(.A(men_men_n232_), .Y(men_men_n233_));
  NAi21      u0205(.An(n), .B(a), .Y(men_men_n234_));
  NO2        u0206(.A(men_men_n234_), .B(men_men_n150_), .Y(men_men_n235_));
  NAi41      u0207(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n236_));
  NO2        u0208(.A(men_men_n236_), .B(e), .Y(men_men_n237_));
  NO3        u0209(.A(men_men_n151_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n238_));
  OAI210     u0210(.A0(men_men_n238_), .A1(men_men_n237_), .B0(men_men_n235_), .Y(men_men_n239_));
  AN3        u0211(.A(men_men_n239_), .B(men_men_n233_), .C(men_men_n225_), .Y(men_men_n240_));
  OR2        u0212(.A(h), .B(g), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n105_), .Y(men_men_n242_));
  NA2        u0214(.A(men_men_n242_), .B(men_men_n132_), .Y(men_men_n243_));
  NAi41      u0215(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n244_));
  NO2        u0216(.A(men_men_n244_), .B(men_men_n215_), .Y(men_men_n245_));
  NA2        u0217(.A(men_men_n163_), .B(men_men_n110_), .Y(men_men_n246_));
  NAi21      u0218(.An(men_men_n246_), .B(men_men_n245_), .Y(men_men_n247_));
  NO2        u0219(.A(n), .B(a), .Y(men_men_n248_));
  NAi31      u0220(.An(men_men_n236_), .B(men_men_n248_), .C(men_men_n106_), .Y(men_men_n249_));
  AN2        u0221(.A(men_men_n249_), .B(men_men_n247_), .Y(men_men_n250_));
  NAi21      u0222(.An(h), .B(i), .Y(men_men_n251_));
  NA2        u0223(.A(men_men_n250_), .B(men_men_n243_), .Y(men_men_n252_));
  NOi21      u0224(.An(g), .B(e), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n254_));
  NA2        u0226(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NOi32      u0227(.An(l), .Bn(j), .C(i), .Y(men_men_n256_));
  AOI210     u0228(.A0(men_men_n75_), .A1(men_men_n88_), .B0(men_men_n256_), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n251_), .B(men_men_n44_), .Y(men_men_n258_));
  NAi21      u0230(.An(f), .B(g), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n64_), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n68_), .B(men_men_n118_), .Y(men_men_n261_));
  AOI220     u0233(.A0(men_men_n261_), .A1(men_men_n260_), .B0(men_men_n258_), .B1(men_men_n66_), .Y(men_men_n262_));
  OAI210     u0234(.A0(men_men_n257_), .A1(men_men_n255_), .B0(men_men_n262_), .Y(men_men_n263_));
  NO3        u0235(.A(men_men_n135_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n264_));
  NOi41      u0236(.An(men_men_n240_), .B(men_men_n263_), .C(men_men_n252_), .D(men_men_n222_), .Y(men_men_n265_));
  NO4        u0237(.A(men_men_n203_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n266_));
  NO2        u0238(.A(men_men_n266_), .B(men_men_n113_), .Y(men_men_n267_));
  NA3        u0239(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n268_));
  NAi21      u0240(.An(h), .B(g), .Y(men_men_n269_));
  OR4        u0241(.A(men_men_n269_), .B(men_men_n268_), .C(men_men_n224_), .D(e), .Y(men_men_n270_));
  NO2        u0242(.A(men_men_n246_), .B(men_men_n259_), .Y(men_men_n271_));
  NAi31      u0243(.An(g), .B(k), .C(h), .Y(men_men_n272_));
  NO3        u0244(.A(men_men_n134_), .B(men_men_n272_), .C(l), .Y(men_men_n273_));
  NAi31      u0245(.An(e), .B(d), .C(a), .Y(men_men_n274_));
  NA2        u0246(.A(men_men_n273_), .B(men_men_n132_), .Y(men_men_n275_));
  NA2        u0247(.A(men_men_n275_), .B(men_men_n270_), .Y(men_men_n276_));
  NA4        u0248(.A(men_men_n163_), .B(men_men_n81_), .C(men_men_n77_), .D(men_men_n118_), .Y(men_men_n277_));
  NA2        u0249(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n278_));
  NA3        u0250(.A(e), .B(c), .C(b), .Y(men_men_n279_));
  NO2        u0251(.A(d), .B(men_men_n279_), .Y(men_men_n280_));
  NAi32      u0252(.An(k), .Bn(i), .C(j), .Y(men_men_n281_));
  NAi31      u0253(.An(h), .B(l), .C(i), .Y(men_men_n282_));
  NA3        u0254(.A(men_men_n282_), .B(men_men_n281_), .C(men_men_n169_), .Y(men_men_n283_));
  NOi21      u0255(.An(men_men_n283_), .B(men_men_n49_), .Y(men_men_n284_));
  OAI210     u0256(.A0(men_men_n260_), .A1(men_men_n280_), .B0(men_men_n284_), .Y(men_men_n285_));
  NAi21      u0257(.An(l), .B(k), .Y(men_men_n286_));
  NO2        u0258(.A(men_men_n286_), .B(men_men_n49_), .Y(men_men_n287_));
  NOi21      u0259(.An(l), .B(j), .Y(men_men_n288_));
  NA2        u0260(.A(men_men_n166_), .B(men_men_n288_), .Y(men_men_n289_));
  NA3        u0261(.A(men_men_n119_), .B(men_men_n118_), .C(g), .Y(men_men_n290_));
  OR3        u0262(.A(men_men_n72_), .B(men_men_n74_), .C(e), .Y(men_men_n291_));
  AOI210     u0263(.A0(men_men_n290_), .A1(men_men_n289_), .B0(men_men_n291_), .Y(men_men_n292_));
  INV        u0264(.A(men_men_n292_), .Y(men_men_n293_));
  NAi32      u0265(.An(j), .Bn(h), .C(i), .Y(men_men_n294_));
  NAi21      u0266(.An(m), .B(l), .Y(men_men_n295_));
  NO2        u0267(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n296_));
  NA2        u0268(.A(h), .B(g), .Y(men_men_n297_));
  NA2        u0269(.A(men_men_n172_), .B(men_men_n45_), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n298_), .B(men_men_n297_), .Y(men_men_n299_));
  OAI210     u0271(.A0(men_men_n299_), .A1(men_men_n296_), .B0(men_men_n167_), .Y(men_men_n300_));
  NA4        u0272(.A(men_men_n300_), .B(men_men_n293_), .C(men_men_n285_), .D(men_men_n277_), .Y(men_men_n301_));
  NO2        u0273(.A(men_men_n148_), .B(d), .Y(men_men_n302_));
  NA2        u0274(.A(men_men_n302_), .B(men_men_n53_), .Y(men_men_n303_));
  NAi32      u0275(.An(n), .Bn(m), .C(l), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n304_), .B(men_men_n294_), .Y(men_men_n305_));
  INV        u0277(.A(men_men_n305_), .Y(men_men_n306_));
  NO2        u0278(.A(men_men_n123_), .B(men_men_n117_), .Y(men_men_n307_));
  NAi31      u0279(.An(k), .B(l), .C(j), .Y(men_men_n308_));
  OAI210     u0280(.A0(men_men_n286_), .A1(j), .B0(men_men_n308_), .Y(men_men_n309_));
  NOi21      u0281(.An(men_men_n309_), .B(men_men_n121_), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n310_), .B(men_men_n307_), .Y(men_men_n311_));
  NA2        u0283(.A(men_men_n311_), .B(men_men_n303_), .Y(men_men_n312_));
  NO4        u0284(.A(men_men_n312_), .B(men_men_n301_), .C(men_men_n276_), .D(men_men_n267_), .Y(men_men_n313_));
  NO2        u0285(.A(men_men_n227_), .B(m), .Y(men_men_n314_));
  NAi41      u0286(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n315_));
  NAi31      u0287(.An(i), .B(l), .C(h), .Y(men_men_n316_));
  NO4        u0288(.A(men_men_n316_), .B(e), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n317_));
  NA2        u0289(.A(e), .B(c), .Y(men_men_n318_));
  NOi21      u0290(.An(f), .B(h), .Y(men_men_n319_));
  NA2        u0291(.A(men_men_n319_), .B(men_men_n119_), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n216_), .Y(men_men_n321_));
  NAi31      u0293(.An(d), .B(e), .C(b), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n134_), .B(men_men_n322_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n321_), .Y(men_men_n324_));
  NAi21      u0296(.An(men_men_n317_), .B(men_men_n324_), .Y(men_men_n325_));
  NO4        u0297(.A(men_men_n315_), .B(men_men_n80_), .C(men_men_n71_), .D(men_men_n216_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n248_), .B(men_men_n106_), .Y(men_men_n327_));
  OR2        u0299(.A(men_men_n327_), .B(men_men_n205_), .Y(men_men_n328_));
  NOi31      u0300(.An(l), .B(n), .C(m), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n329_), .B(men_men_n217_), .Y(men_men_n330_));
  INV        u0302(.A(men_men_n330_), .Y(men_men_n331_));
  NAi32      u0303(.An(men_men_n331_), .Bn(men_men_n326_), .C(men_men_n328_), .Y(men_men_n332_));
  NAi32      u0304(.An(m), .Bn(j), .C(k), .Y(men_men_n333_));
  NAi41      u0305(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n334_));
  INV        u0306(.A(men_men_n334_), .Y(men_men_n335_));
  NOi31      u0307(.An(j), .B(m), .C(k), .Y(men_men_n336_));
  NO2        u0308(.A(men_men_n127_), .B(men_men_n336_), .Y(men_men_n337_));
  AN3        u0309(.A(h), .B(g), .C(f), .Y(men_men_n338_));
  NAi31      u0310(.An(men_men_n337_), .B(men_men_n338_), .C(men_men_n335_), .Y(men_men_n339_));
  NOi32      u0311(.An(m), .Bn(j), .C(l), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n340_), .B(men_men_n99_), .Y(men_men_n341_));
  NAi32      u0313(.An(men_men_n341_), .Bn(men_men_n202_), .C(men_men_n302_), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n219_), .B(g), .Y(men_men_n344_));
  INV        u0316(.A(men_men_n159_), .Y(men_men_n345_));
  AOI220     u0317(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n245_), .B1(men_men_n343_), .Y(men_men_n346_));
  INV        u0318(.A(men_men_n231_), .Y(men_men_n347_));
  NA3        u0319(.A(men_men_n347_), .B(men_men_n338_), .C(men_men_n214_), .Y(men_men_n348_));
  NA4        u0320(.A(men_men_n348_), .B(men_men_n346_), .C(men_men_n342_), .D(men_men_n339_), .Y(men_men_n349_));
  NA3        u0321(.A(h), .B(g), .C(f), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n350_), .B(men_men_n76_), .Y(men_men_n351_));
  NA2        u0323(.A(men_men_n334_), .B(men_men_n213_), .Y(men_men_n352_));
  NA2        u0324(.A(men_men_n166_), .B(e), .Y(men_men_n353_));
  NO2        u0325(.A(men_men_n353_), .B(men_men_n41_), .Y(men_men_n354_));
  AOI220     u0326(.A0(men_men_n354_), .A1(men_men_n307_), .B0(men_men_n352_), .B1(men_men_n351_), .Y(men_men_n355_));
  NOi32      u0327(.An(j), .Bn(g), .C(i), .Y(men_men_n356_));
  NA3        u0328(.A(men_men_n356_), .B(men_men_n286_), .C(men_men_n115_), .Y(men_men_n357_));
  AO210      u0329(.A0(men_men_n113_), .A1(men_men_n32_), .B0(men_men_n357_), .Y(men_men_n358_));
  NOi32      u0330(.An(e), .Bn(b), .C(a), .Y(men_men_n359_));
  AN2        u0331(.A(l), .B(j), .Y(men_men_n360_));
  NO2        u0332(.A(m), .B(men_men_n360_), .Y(men_men_n361_));
  NO3        u0333(.A(men_men_n315_), .B(men_men_n71_), .C(men_men_n216_), .Y(men_men_n362_));
  NA3        u0334(.A(men_men_n210_), .B(men_men_n208_), .C(men_men_n35_), .Y(men_men_n363_));
  AOI220     u0335(.A0(men_men_n363_), .A1(men_men_n359_), .B0(men_men_n362_), .B1(men_men_n361_), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n322_), .B(n), .Y(men_men_n365_));
  NA2        u0337(.A(men_men_n209_), .B(k), .Y(men_men_n366_));
  NA3        u0338(.A(m), .B(men_men_n114_), .C(men_men_n215_), .Y(men_men_n367_));
  NA4        u0339(.A(men_men_n204_), .B(men_men_n88_), .C(g), .D(men_men_n215_), .Y(men_men_n368_));
  OAI210     u0340(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n368_), .Y(men_men_n369_));
  NAi41      u0341(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n370_));
  NA2        u0342(.A(men_men_n51_), .B(men_men_n115_), .Y(men_men_n371_));
  NO2        u0343(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  AOI220     u0344(.A0(men_men_n372_), .A1(b), .B0(men_men_n369_), .B1(men_men_n365_), .Y(men_men_n373_));
  NA4        u0345(.A(men_men_n373_), .B(men_men_n364_), .C(men_men_n358_), .D(men_men_n355_), .Y(men_men_n374_));
  NO4        u0346(.A(men_men_n374_), .B(men_men_n349_), .C(men_men_n332_), .D(men_men_n325_), .Y(men_men_n375_));
  NA4        u0347(.A(men_men_n375_), .B(men_men_n313_), .C(men_men_n265_), .D(men_men_n200_), .Y(men10));
  NA3        u0348(.A(m), .B(k), .C(i), .Y(men_men_n377_));
  NO3        u0349(.A(men_men_n377_), .B(j), .C(men_men_n216_), .Y(men_men_n378_));
  NOi21      u0350(.An(e), .B(f), .Y(men_men_n379_));
  NO4        u0351(.A(men_men_n154_), .B(men_men_n379_), .C(n), .D(men_men_n112_), .Y(men_men_n380_));
  NAi31      u0352(.An(b), .B(f), .C(c), .Y(men_men_n381_));
  INV        u0353(.A(men_men_n381_), .Y(men_men_n382_));
  NOi32      u0354(.An(k), .Bn(h), .C(j), .Y(men_men_n383_));
  NA2        u0355(.A(men_men_n383_), .B(men_men_n223_), .Y(men_men_n384_));
  NA2        u0356(.A(men_men_n164_), .B(men_men_n384_), .Y(men_men_n385_));
  AOI220     u0357(.A0(men_men_n385_), .A1(men_men_n382_), .B0(men_men_n380_), .B1(men_men_n378_), .Y(men_men_n386_));
  OR2        u0358(.A(m), .B(k), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n177_), .B(men_men_n387_), .Y(men_men_n388_));
  NA3        u0360(.A(f), .B(c), .C(men_men_n117_), .Y(men_men_n389_));
  NOi32      u0361(.An(d), .Bn(a), .C(c), .Y(men_men_n390_));
  NA2        u0362(.A(men_men_n390_), .B(men_men_n185_), .Y(men_men_n391_));
  NAi21      u0363(.An(i), .B(g), .Y(men_men_n392_));
  NAi31      u0364(.An(k), .B(m), .C(j), .Y(men_men_n393_));
  NO3        u0365(.A(men_men_n393_), .B(men_men_n392_), .C(n), .Y(men_men_n394_));
  NOi21      u0366(.An(men_men_n394_), .B(men_men_n391_), .Y(men_men_n395_));
  INV        u0367(.A(men_men_n395_), .Y(men_men_n396_));
  NO2        u0368(.A(men_men_n389_), .B(men_men_n295_), .Y(men_men_n397_));
  AOI220     u0369(.A0(f), .A1(men_men_n305_), .B0(men_men_n397_), .B1(men_men_n217_), .Y(men_men_n398_));
  NA3        u0370(.A(men_men_n398_), .B(men_men_n396_), .C(men_men_n386_), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n59_), .B(men_men_n117_), .Y(men_men_n400_));
  NA2        u0372(.A(men_men_n248_), .B(men_men_n400_), .Y(men_men_n401_));
  INV        u0373(.A(e), .Y(men_men_n402_));
  NA2        u0374(.A(men_men_n46_), .B(e), .Y(men_men_n403_));
  OAI220     u0375(.A0(men_men_n403_), .A1(men_men_n201_), .B0(men_men_n205_), .B1(men_men_n402_), .Y(men_men_n404_));
  AN2        u0376(.A(g), .B(e), .Y(men_men_n405_));
  NA3        u0377(.A(men_men_n405_), .B(men_men_n204_), .C(i), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n90_), .B(men_men_n406_), .Y(men_men_n407_));
  NO2        u0379(.A(men_men_n102_), .B(men_men_n402_), .Y(men_men_n408_));
  NO3        u0380(.A(men_men_n408_), .B(men_men_n407_), .C(men_men_n404_), .Y(men_men_n409_));
  NOi32      u0381(.An(h), .Bn(e), .C(g), .Y(men_men_n410_));
  NA3        u0382(.A(men_men_n410_), .B(men_men_n288_), .C(m), .Y(men_men_n411_));
  NOi21      u0383(.An(g), .B(h), .Y(men_men_n412_));
  AN3        u0384(.A(m), .B(l), .C(i), .Y(men_men_n413_));
  NA3        u0385(.A(men_men_n413_), .B(men_men_n412_), .C(e), .Y(men_men_n414_));
  AN3        u0386(.A(h), .B(g), .C(e), .Y(men_men_n415_));
  NA2        u0387(.A(men_men_n415_), .B(men_men_n99_), .Y(men_men_n416_));
  AN3        u0388(.A(men_men_n416_), .B(men_men_n414_), .C(men_men_n411_), .Y(men_men_n417_));
  AOI210     u0389(.A0(men_men_n417_), .A1(men_men_n409_), .B0(men_men_n401_), .Y(men_men_n418_));
  NA3        u0390(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n419_), .B(men_men_n401_), .Y(men_men_n420_));
  NA3        u0392(.A(men_men_n390_), .B(men_men_n185_), .C(men_men_n85_), .Y(men_men_n421_));
  NAi31      u0393(.An(b), .B(c), .C(a), .Y(men_men_n422_));
  NO2        u0394(.A(men_men_n422_), .B(n), .Y(men_men_n423_));
  OAI210     u0395(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n424_));
  NO3        u0396(.A(men_men_n420_), .B(men_men_n418_), .C(men_men_n399_), .Y(men_men_n425_));
  NA2        u0397(.A(i), .B(g), .Y(men_men_n426_));
  NO3        u0398(.A(men_men_n274_), .B(men_men_n426_), .C(c), .Y(men_men_n427_));
  NOi21      u0399(.An(d), .B(c), .Y(men_men_n428_));
  NA2        u0400(.A(men_men_n428_), .B(a), .Y(men_men_n429_));
  NA3        u0401(.A(i), .B(g), .C(f), .Y(men_men_n430_));
  OR2        u0402(.A(men_men_n430_), .B(men_men_n70_), .Y(men_men_n431_));
  NA3        u0403(.A(men_men_n413_), .B(men_men_n412_), .C(men_men_n185_), .Y(men_men_n432_));
  AOI210     u0404(.A0(men_men_n432_), .A1(men_men_n431_), .B0(men_men_n429_), .Y(men_men_n433_));
  AOI210     u0405(.A0(men_men_n427_), .A1(men_men_n287_), .B0(men_men_n433_), .Y(men_men_n434_));
  OR2        u0406(.A(n), .B(m), .Y(men_men_n435_));
  NO2        u0407(.A(men_men_n435_), .B(men_men_n155_), .Y(men_men_n436_));
  INV        u0408(.A(men_men_n186_), .Y(men_men_n437_));
  OAI210     u0409(.A0(men_men_n436_), .A1(men_men_n179_), .B0(men_men_n437_), .Y(men_men_n438_));
  INV        u0410(.A(men_men_n371_), .Y(men_men_n439_));
  NA3        u0411(.A(men_men_n439_), .B(men_men_n359_), .C(d), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n422_), .B(men_men_n49_), .Y(men_men_n441_));
  NO3        u0413(.A(men_men_n65_), .B(men_men_n114_), .C(e), .Y(men_men_n442_));
  NAi21      u0414(.An(k), .B(j), .Y(men_men_n443_));
  NA2        u0415(.A(men_men_n251_), .B(men_men_n443_), .Y(men_men_n444_));
  NA3        u0416(.A(men_men_n444_), .B(men_men_n442_), .C(men_men_n441_), .Y(men_men_n445_));
  NAi21      u0417(.An(e), .B(d), .Y(men_men_n446_));
  NA3        u0418(.A(men_men_n445_), .B(men_men_n440_), .C(men_men_n438_), .Y(men_men_n447_));
  NOi31      u0419(.An(n), .B(m), .C(k), .Y(men_men_n448_));
  AOI220     u0420(.A0(men_men_n448_), .A1(h), .B0(men_men_n223_), .B1(men_men_n50_), .Y(men_men_n449_));
  NAi31      u0421(.An(g), .B(f), .C(c), .Y(men_men_n450_));
  OR3        u0422(.A(men_men_n450_), .B(men_men_n449_), .C(e), .Y(men_men_n451_));
  NA2        u0423(.A(men_men_n451_), .B(men_men_n306_), .Y(men_men_n452_));
  NOi41      u0424(.An(men_men_n434_), .B(men_men_n452_), .C(men_men_n447_), .D(men_men_n263_), .Y(men_men_n453_));
  NOi32      u0425(.An(c), .Bn(a), .C(b), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n115_), .Y(men_men_n455_));
  INV        u0427(.A(men_men_n272_), .Y(men_men_n456_));
  AN2        u0428(.A(e), .B(d), .Y(men_men_n457_));
  NO2        u0429(.A(men_men_n133_), .B(men_men_n41_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n65_), .B(e), .Y(men_men_n459_));
  NOi31      u0431(.An(j), .B(k), .C(i), .Y(men_men_n460_));
  NOi21      u0432(.An(men_men_n169_), .B(men_men_n460_), .Y(men_men_n461_));
  NA4        u0433(.A(men_men_n316_), .B(men_men_n461_), .C(men_men_n257_), .D(men_men_n120_), .Y(men_men_n462_));
  AOI210     u0434(.A0(men_men_n462_), .A1(men_men_n459_), .B0(men_men_n458_), .Y(men_men_n463_));
  AOI210     u0435(.A0(men_men_n463_), .A1(men_men_n272_), .B0(men_men_n455_), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n211_), .B(men_men_n206_), .Y(men_men_n465_));
  NOi21      u0437(.An(a), .B(b), .Y(men_men_n466_));
  NA3        u0438(.A(e), .B(d), .C(c), .Y(men_men_n467_));
  NAi21      u0439(.An(men_men_n467_), .B(men_men_n466_), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n421_), .B(men_men_n205_), .Y(men_men_n469_));
  NOi21      u0441(.An(men_men_n468_), .B(men_men_n469_), .Y(men_men_n470_));
  AOI210     u0442(.A0(men_men_n266_), .A1(men_men_n465_), .B0(men_men_n470_), .Y(men_men_n471_));
  OR2        u0443(.A(k), .B(j), .Y(men_men_n472_));
  NA2        u0444(.A(l), .B(k), .Y(men_men_n473_));
  NA3        u0445(.A(men_men_n473_), .B(men_men_n472_), .C(men_men_n223_), .Y(men_men_n474_));
  NA2        u0446(.A(men_men_n231_), .B(men_men_n333_), .Y(men_men_n475_));
  NOi21      u0447(.An(men_men_n474_), .B(men_men_n475_), .Y(men_men_n476_));
  OR3        u0448(.A(men_men_n476_), .B(men_men_n147_), .C(men_men_n137_), .Y(men_men_n477_));
  NA3        u0449(.A(men_men_n277_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n478_));
  NA2        u0450(.A(men_men_n390_), .B(men_men_n115_), .Y(men_men_n479_));
  NO4        u0451(.A(men_men_n479_), .B(men_men_n96_), .C(men_men_n114_), .D(e), .Y(men_men_n480_));
  NO3        u0452(.A(men_men_n421_), .B(men_men_n93_), .C(men_men_n133_), .Y(men_men_n481_));
  NO4        u0453(.A(men_men_n481_), .B(men_men_n480_), .C(men_men_n478_), .D(men_men_n317_), .Y(men_men_n482_));
  NA2        u0454(.A(men_men_n482_), .B(men_men_n477_), .Y(men_men_n483_));
  NO3        u0455(.A(men_men_n483_), .B(men_men_n471_), .C(men_men_n464_), .Y(men_men_n484_));
  NA2        u0456(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n485_));
  NO2        u0457(.A(men_men_n191_), .B(men_men_n56_), .Y(men_men_n486_));
  NAi31      u0458(.An(j), .B(l), .C(i), .Y(men_men_n487_));
  OAI210     u0459(.A0(men_men_n487_), .A1(men_men_n134_), .B0(men_men_n105_), .Y(men_men_n488_));
  NA3        u0460(.A(men_men_n488_), .B(men_men_n486_), .C(d), .Y(men_men_n489_));
  NO3        u0461(.A(men_men_n391_), .B(men_men_n341_), .C(men_men_n202_), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n391_), .B(men_men_n371_), .Y(men_men_n491_));
  NO3        u0463(.A(men_men_n491_), .B(men_men_n490_), .C(men_men_n187_), .Y(men_men_n492_));
  NA4        u0464(.A(men_men_n492_), .B(men_men_n489_), .C(men_men_n485_), .D(men_men_n240_), .Y(men_men_n493_));
  OAI210     u0465(.A0(men_men_n129_), .A1(men_men_n127_), .B0(n), .Y(men_men_n494_));
  NO2        u0466(.A(men_men_n494_), .B(men_men_n133_), .Y(men_men_n495_));
  OR2        u0467(.A(men_men_n296_), .B(men_men_n242_), .Y(men_men_n496_));
  OA210      u0468(.A0(men_men_n496_), .A1(men_men_n495_), .B0(men_men_n195_), .Y(men_men_n497_));
  XO2        u0469(.A(i), .B(h), .Y(men_men_n498_));
  NA3        u0470(.A(men_men_n498_), .B(men_men_n163_), .C(n), .Y(men_men_n499_));
  NAi41      u0471(.An(men_men_n296_), .B(men_men_n499_), .C(men_men_n449_), .D(men_men_n384_), .Y(men_men_n500_));
  NOi32      u0472(.An(men_men_n500_), .Bn(men_men_n459_), .C(men_men_n268_), .Y(men_men_n501_));
  NAi31      u0473(.An(c), .B(f), .C(d), .Y(men_men_n502_));
  BUFFER     u0474(.A(men_men_n83_), .Y(men_men_n503_));
  NA3        u0475(.A(men_men_n380_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n504_));
  NA2        u0476(.A(men_men_n228_), .B(men_men_n110_), .Y(men_men_n505_));
  AOI210     u0477(.A0(men_men_n505_), .A1(men_men_n184_), .B0(men_men_n502_), .Y(men_men_n506_));
  AOI210     u0478(.A0(men_men_n357_), .A1(men_men_n35_), .B0(men_men_n468_), .Y(men_men_n507_));
  NOi31      u0479(.An(men_men_n504_), .B(men_men_n507_), .C(men_men_n506_), .Y(men_men_n508_));
  AO220      u0480(.A0(men_men_n284_), .A1(men_men_n260_), .B0(men_men_n170_), .B1(men_men_n66_), .Y(men_men_n509_));
  NA3        u0481(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n510_));
  NO2        u0482(.A(men_men_n510_), .B(men_men_n429_), .Y(men_men_n511_));
  NO2        u0483(.A(men_men_n511_), .B(men_men_n292_), .Y(men_men_n512_));
  NAi41      u0484(.An(men_men_n509_), .B(men_men_n512_), .C(men_men_n508_), .D(men_men_n503_), .Y(men_men_n513_));
  NO4        u0485(.A(men_men_n513_), .B(men_men_n501_), .C(men_men_n497_), .D(men_men_n493_), .Y(men_men_n514_));
  NA4        u0486(.A(men_men_n514_), .B(men_men_n484_), .C(men_men_n453_), .D(men_men_n425_), .Y(men11));
  NO2        u0487(.A(men_men_n72_), .B(f), .Y(men_men_n516_));
  NA2        u0488(.A(j), .B(g), .Y(men_men_n517_));
  NAi31      u0489(.An(i), .B(m), .C(l), .Y(men_men_n518_));
  NA3        u0490(.A(m), .B(k), .C(j), .Y(men_men_n519_));
  OAI220     u0491(.A0(men_men_n519_), .A1(men_men_n133_), .B0(men_men_n518_), .B1(men_men_n517_), .Y(men_men_n520_));
  NA2        u0492(.A(men_men_n520_), .B(men_men_n516_), .Y(men_men_n521_));
  NOi32      u0493(.An(e), .Bn(b), .C(f), .Y(men_men_n522_));
  NA2        u0494(.A(men_men_n256_), .B(men_men_n115_), .Y(men_men_n523_));
  NA2        u0495(.A(men_men_n46_), .B(j), .Y(men_men_n524_));
  NO2        u0496(.A(men_men_n524_), .B(men_men_n298_), .Y(men_men_n525_));
  NAi31      u0497(.An(d), .B(e), .C(a), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n526_), .B(n), .Y(men_men_n527_));
  AOI220     u0499(.A0(men_men_n527_), .A1(men_men_n103_), .B0(men_men_n525_), .B1(men_men_n522_), .Y(men_men_n528_));
  NAi41      u0500(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n529_));
  AN2        u0501(.A(men_men_n529_), .B(men_men_n370_), .Y(men_men_n530_));
  AOI210     u0502(.A0(men_men_n530_), .A1(men_men_n391_), .B0(men_men_n269_), .Y(men_men_n531_));
  NA2        u0503(.A(j), .B(i), .Y(men_men_n532_));
  NAi31      u0504(.An(n), .B(m), .C(k), .Y(men_men_n533_));
  NO3        u0505(.A(men_men_n533_), .B(men_men_n532_), .C(men_men_n114_), .Y(men_men_n534_));
  NO4        u0506(.A(n), .B(d), .C(men_men_n117_), .D(a), .Y(men_men_n535_));
  OR2        u0507(.A(n), .B(c), .Y(men_men_n536_));
  NO2        u0508(.A(men_men_n536_), .B(men_men_n153_), .Y(men_men_n537_));
  NO2        u0509(.A(men_men_n537_), .B(men_men_n535_), .Y(men_men_n538_));
  NOi32      u0510(.An(g), .Bn(f), .C(i), .Y(men_men_n539_));
  AOI220     u0511(.A0(men_men_n539_), .A1(men_men_n101_), .B0(men_men_n520_), .B1(f), .Y(men_men_n540_));
  NO2        u0512(.A(men_men_n272_), .B(men_men_n49_), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n540_), .B(men_men_n538_), .Y(men_men_n542_));
  AOI210     u0514(.A0(men_men_n534_), .A1(men_men_n531_), .B0(men_men_n542_), .Y(men_men_n543_));
  NA2        u0515(.A(men_men_n143_), .B(men_men_n34_), .Y(men_men_n544_));
  OAI220     u0516(.A0(men_men_n544_), .A1(m), .B0(men_men_n524_), .B1(men_men_n231_), .Y(men_men_n545_));
  NOi41      u0517(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n546_));
  NAi32      u0518(.An(e), .Bn(b), .C(c), .Y(men_men_n547_));
  AN2        u0519(.A(men_men_n334_), .B(men_men_n315_), .Y(men_men_n548_));
  NA2        u0520(.A(men_men_n548_), .B(men_men_n547_), .Y(men_men_n549_));
  OA210      u0521(.A0(men_men_n549_), .A1(men_men_n546_), .B0(men_men_n545_), .Y(men_men_n550_));
  OAI220     u0522(.A0(men_men_n393_), .A1(men_men_n392_), .B0(men_men_n518_), .B1(men_men_n517_), .Y(men_men_n551_));
  NAi31      u0523(.An(d), .B(c), .C(a), .Y(men_men_n552_));
  NO2        u0524(.A(men_men_n552_), .B(n), .Y(men_men_n553_));
  NA3        u0525(.A(men_men_n553_), .B(men_men_n551_), .C(e), .Y(men_men_n554_));
  NO3        u0526(.A(men_men_n61_), .B(men_men_n49_), .C(men_men_n216_), .Y(men_men_n555_));
  NO2        u0527(.A(men_men_n229_), .B(men_men_n112_), .Y(men_men_n556_));
  OAI210     u0528(.A0(men_men_n555_), .A1(men_men_n394_), .B0(men_men_n556_), .Y(men_men_n557_));
  NA2        u0529(.A(men_men_n557_), .B(men_men_n554_), .Y(men_men_n558_));
  NO2        u0530(.A(men_men_n274_), .B(n), .Y(men_men_n559_));
  NO2        u0531(.A(men_men_n423_), .B(men_men_n559_), .Y(men_men_n560_));
  NA2        u0532(.A(men_men_n551_), .B(f), .Y(men_men_n561_));
  NAi32      u0533(.An(d), .Bn(a), .C(b), .Y(men_men_n562_));
  NO2        u0534(.A(men_men_n562_), .B(men_men_n49_), .Y(men_men_n563_));
  NA2        u0535(.A(h), .B(f), .Y(men_men_n564_));
  NO2        u0536(.A(men_men_n564_), .B(men_men_n96_), .Y(men_men_n565_));
  NO3        u0537(.A(men_men_n180_), .B(men_men_n177_), .C(g), .Y(men_men_n566_));
  AOI220     u0538(.A0(men_men_n566_), .A1(men_men_n58_), .B0(men_men_n565_), .B1(men_men_n563_), .Y(men_men_n567_));
  OAI210     u0539(.A0(men_men_n561_), .A1(men_men_n560_), .B0(men_men_n567_), .Y(men_men_n568_));
  AN3        u0540(.A(j), .B(h), .C(g), .Y(men_men_n569_));
  NO2        u0541(.A(men_men_n150_), .B(c), .Y(men_men_n570_));
  NA3        u0542(.A(men_men_n570_), .B(men_men_n569_), .C(men_men_n448_), .Y(men_men_n571_));
  NA3        u0543(.A(f), .B(d), .C(b), .Y(men_men_n572_));
  NO4        u0544(.A(men_men_n572_), .B(men_men_n180_), .C(men_men_n177_), .D(g), .Y(men_men_n573_));
  NAi21      u0545(.An(men_men_n573_), .B(men_men_n571_), .Y(men_men_n574_));
  NO4        u0546(.A(men_men_n574_), .B(men_men_n568_), .C(men_men_n558_), .D(men_men_n550_), .Y(men_men_n575_));
  AN4        u0547(.A(men_men_n575_), .B(men_men_n543_), .C(men_men_n528_), .D(men_men_n521_), .Y(men_men_n576_));
  INV        u0548(.A(k), .Y(men_men_n577_));
  NA3        u0549(.A(l), .B(men_men_n577_), .C(i), .Y(men_men_n578_));
  INV        u0550(.A(men_men_n578_), .Y(men_men_n579_));
  NA3        u0551(.A(men_men_n390_), .B(men_men_n412_), .C(men_men_n115_), .Y(men_men_n580_));
  NAi32      u0552(.An(h), .Bn(f), .C(g), .Y(men_men_n581_));
  NAi41      u0553(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n582_));
  OAI210     u0554(.A0(men_men_n526_), .A1(n), .B0(men_men_n582_), .Y(men_men_n583_));
  NA2        u0555(.A(men_men_n583_), .B(m), .Y(men_men_n584_));
  NAi31      u0556(.An(h), .B(g), .C(f), .Y(men_men_n585_));
  OR3        u0557(.A(men_men_n585_), .B(men_men_n274_), .C(men_men_n49_), .Y(men_men_n586_));
  NA4        u0558(.A(men_men_n412_), .B(men_men_n122_), .C(men_men_n115_), .D(e), .Y(men_men_n587_));
  AN2        u0559(.A(men_men_n587_), .B(men_men_n586_), .Y(men_men_n588_));
  OA210      u0560(.A0(men_men_n584_), .A1(men_men_n581_), .B0(men_men_n588_), .Y(men_men_n589_));
  NO3        u0561(.A(men_men_n581_), .B(men_men_n72_), .C(men_men_n74_), .Y(men_men_n590_));
  NO4        u0562(.A(men_men_n585_), .B(men_men_n536_), .C(men_men_n153_), .D(men_men_n74_), .Y(men_men_n591_));
  OR2        u0563(.A(men_men_n591_), .B(men_men_n590_), .Y(men_men_n592_));
  NAi31      u0564(.An(men_men_n592_), .B(men_men_n589_), .C(men_men_n580_), .Y(men_men_n593_));
  NAi31      u0565(.An(f), .B(h), .C(g), .Y(men_men_n594_));
  NO4        u0566(.A(men_men_n308_), .B(men_men_n594_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n595_));
  NOi32      u0567(.An(b), .Bn(a), .C(c), .Y(men_men_n596_));
  NOi41      u0568(.An(men_men_n596_), .B(men_men_n350_), .C(men_men_n68_), .D(men_men_n118_), .Y(men_men_n597_));
  OR2        u0569(.A(men_men_n597_), .B(men_men_n595_), .Y(men_men_n598_));
  NOi32      u0570(.An(d), .Bn(a), .C(e), .Y(men_men_n599_));
  NA2        u0571(.A(men_men_n599_), .B(men_men_n115_), .Y(men_men_n600_));
  NO2        u0572(.A(n), .B(c), .Y(men_men_n601_));
  NA3        u0573(.A(men_men_n601_), .B(men_men_n29_), .C(m), .Y(men_men_n602_));
  NAi32      u0574(.An(n), .Bn(f), .C(m), .Y(men_men_n603_));
  NA3        u0575(.A(men_men_n603_), .B(men_men_n602_), .C(men_men_n600_), .Y(men_men_n604_));
  NOi32      u0576(.An(e), .Bn(a), .C(d), .Y(men_men_n605_));
  AOI210     u0577(.A0(men_men_n29_), .A1(d), .B0(men_men_n605_), .Y(men_men_n606_));
  INV        u0578(.A(men_men_n544_), .Y(men_men_n607_));
  AOI210     u0579(.A0(men_men_n607_), .A1(men_men_n604_), .B0(men_men_n598_), .Y(men_men_n608_));
  OAI210     u0580(.A0(men_men_n247_), .A1(men_men_n88_), .B0(men_men_n608_), .Y(men_men_n609_));
  AOI210     u0581(.A0(men_men_n593_), .A1(men_men_n579_), .B0(men_men_n609_), .Y(men_men_n610_));
  NO3        u0582(.A(m), .B(men_men_n60_), .C(n), .Y(men_men_n611_));
  NA2        u0583(.A(men_men_n75_), .B(men_men_n115_), .Y(men_men_n612_));
  NO2        u0584(.A(men_men_n612_), .B(men_men_n45_), .Y(men_men_n613_));
  NA2        u0585(.A(men_men_n613_), .B(men_men_n531_), .Y(men_men_n614_));
  NO2        u0586(.A(men_men_n614_), .B(men_men_n88_), .Y(men_men_n615_));
  NA3        u0587(.A(men_men_n546_), .B(men_men_n336_), .C(men_men_n46_), .Y(men_men_n616_));
  NOi32      u0588(.An(e), .Bn(c), .C(f), .Y(men_men_n617_));
  NOi21      u0589(.An(f), .B(g), .Y(men_men_n618_));
  NO2        u0590(.A(men_men_n618_), .B(men_men_n213_), .Y(men_men_n619_));
  AOI220     u0591(.A0(men_men_n619_), .A1(men_men_n388_), .B0(men_men_n617_), .B1(men_men_n179_), .Y(men_men_n620_));
  NA3        u0592(.A(men_men_n620_), .B(men_men_n616_), .C(men_men_n182_), .Y(men_men_n621_));
  AOI210     u0593(.A0(men_men_n530_), .A1(men_men_n391_), .B0(men_men_n297_), .Y(men_men_n622_));
  NA2        u0594(.A(men_men_n622_), .B(men_men_n261_), .Y(men_men_n623_));
  NOi21      u0595(.An(j), .B(l), .Y(men_men_n624_));
  NAi21      u0596(.An(k), .B(h), .Y(men_men_n625_));
  NO2        u0597(.A(men_men_n625_), .B(men_men_n259_), .Y(men_men_n626_));
  NA2        u0598(.A(men_men_n626_), .B(men_men_n624_), .Y(men_men_n627_));
  OR2        u0599(.A(men_men_n627_), .B(men_men_n584_), .Y(men_men_n628_));
  NOi31      u0600(.An(m), .B(n), .C(k), .Y(men_men_n629_));
  NA2        u0601(.A(men_men_n624_), .B(men_men_n629_), .Y(men_men_n630_));
  AOI210     u0602(.A0(men_men_n391_), .A1(men_men_n370_), .B0(men_men_n297_), .Y(men_men_n631_));
  NAi21      u0603(.An(men_men_n630_), .B(men_men_n631_), .Y(men_men_n632_));
  NO2        u0604(.A(men_men_n274_), .B(men_men_n49_), .Y(men_men_n633_));
  NO2        u0605(.A(men_men_n308_), .B(men_men_n594_), .Y(men_men_n634_));
  NO2        u0606(.A(men_men_n526_), .B(men_men_n49_), .Y(men_men_n635_));
  AOI220     u0607(.A0(men_men_n635_), .A1(men_men_n634_), .B0(men_men_n633_), .B1(men_men_n565_), .Y(men_men_n636_));
  NA4        u0608(.A(men_men_n636_), .B(men_men_n632_), .C(men_men_n628_), .D(men_men_n623_), .Y(men_men_n637_));
  NA2        u0609(.A(men_men_n110_), .B(men_men_n36_), .Y(men_men_n638_));
  NO2        u0610(.A(k), .B(men_men_n216_), .Y(men_men_n639_));
  NO2        u0611(.A(men_men_n522_), .B(men_men_n359_), .Y(men_men_n640_));
  NO2        u0612(.A(men_men_n640_), .B(n), .Y(men_men_n641_));
  NAi31      u0613(.An(men_men_n638_), .B(men_men_n641_), .C(men_men_n639_), .Y(men_men_n642_));
  NO2        u0614(.A(men_men_n524_), .B(men_men_n180_), .Y(men_men_n643_));
  NA3        u0615(.A(men_men_n547_), .B(men_men_n268_), .C(men_men_n148_), .Y(men_men_n644_));
  NA2        u0616(.A(men_men_n498_), .B(men_men_n163_), .Y(men_men_n645_));
  NO3        u0617(.A(men_men_n389_), .B(men_men_n645_), .C(men_men_n88_), .Y(men_men_n646_));
  AOI210     u0618(.A0(men_men_n644_), .A1(men_men_n643_), .B0(men_men_n646_), .Y(men_men_n647_));
  AN3        u0619(.A(f), .B(d), .C(b), .Y(men_men_n648_));
  NO2        u0620(.A(men_men_n648_), .B(men_men_n132_), .Y(men_men_n649_));
  NA3        u0621(.A(men_men_n498_), .B(men_men_n163_), .C(men_men_n216_), .Y(men_men_n650_));
  AOI210     u0622(.A0(men_men_n649_), .A1(men_men_n230_), .B0(men_men_n650_), .Y(men_men_n651_));
  NAi31      u0623(.An(m), .B(n), .C(k), .Y(men_men_n652_));
  OR2        u0624(.A(men_men_n137_), .B(men_men_n60_), .Y(men_men_n653_));
  OAI210     u0625(.A0(men_men_n653_), .A1(men_men_n652_), .B0(men_men_n249_), .Y(men_men_n654_));
  OAI210     u0626(.A0(men_men_n654_), .A1(men_men_n651_), .B0(j), .Y(men_men_n655_));
  NA3        u0627(.A(men_men_n655_), .B(men_men_n647_), .C(men_men_n642_), .Y(men_men_n656_));
  NO4        u0628(.A(men_men_n656_), .B(men_men_n637_), .C(men_men_n621_), .D(men_men_n615_), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n380_), .B(men_men_n166_), .Y(men_men_n658_));
  NAi31      u0630(.An(g), .B(h), .C(f), .Y(men_men_n659_));
  OR3        u0631(.A(men_men_n659_), .B(men_men_n274_), .C(n), .Y(men_men_n660_));
  OA210      u0632(.A0(men_men_n526_), .A1(n), .B0(men_men_n582_), .Y(men_men_n661_));
  NA3        u0633(.A(men_men_n410_), .B(men_men_n122_), .C(men_men_n85_), .Y(men_men_n662_));
  OAI210     u0634(.A0(men_men_n661_), .A1(men_men_n92_), .B0(men_men_n662_), .Y(men_men_n663_));
  NOi21      u0635(.An(men_men_n660_), .B(men_men_n663_), .Y(men_men_n664_));
  AOI210     u0636(.A0(men_men_n664_), .A1(men_men_n658_), .B0(men_men_n519_), .Y(men_men_n665_));
  NO3        u0637(.A(g), .B(men_men_n215_), .C(men_men_n56_), .Y(men_men_n666_));
  NAi21      u0638(.An(h), .B(j), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n388_), .B(men_men_n666_), .Y(men_men_n668_));
  NA2        u0640(.A(men_men_n596_), .B(men_men_n338_), .Y(men_men_n669_));
  OA220      u0641(.A0(men_men_n630_), .A1(men_men_n669_), .B0(men_men_n627_), .B1(men_men_n72_), .Y(men_men_n670_));
  NA3        u0642(.A(men_men_n516_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n671_));
  NA2        u0643(.A(h), .B(men_men_n37_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n101_), .B(men_men_n46_), .Y(men_men_n673_));
  OAI220     u0645(.A0(men_men_n673_), .A1(men_men_n327_), .B0(men_men_n672_), .B1(men_men_n455_), .Y(men_men_n674_));
  AOI210     u0646(.A0(men_men_n562_), .A1(men_men_n422_), .B0(men_men_n49_), .Y(men_men_n675_));
  OAI220     u0647(.A0(men_men_n585_), .A1(men_men_n578_), .B0(men_men_n320_), .B1(men_men_n517_), .Y(men_men_n676_));
  AOI210     u0648(.A0(men_men_n676_), .A1(men_men_n675_), .B0(men_men_n674_), .Y(men_men_n677_));
  NA4        u0649(.A(men_men_n677_), .B(men_men_n671_), .C(men_men_n670_), .D(men_men_n668_), .Y(men_men_n678_));
  NO2        u0650(.A(men_men_n251_), .B(f), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n618_), .B(men_men_n60_), .Y(men_men_n680_));
  NO3        u0652(.A(men_men_n680_), .B(men_men_n679_), .C(men_men_n34_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n323_), .B(men_men_n143_), .Y(men_men_n682_));
  NA2        u0654(.A(men_men_n134_), .B(men_men_n49_), .Y(men_men_n683_));
  AOI220     u0655(.A0(men_men_n683_), .A1(men_men_n522_), .B0(men_men_n359_), .B1(men_men_n115_), .Y(men_men_n684_));
  OA220      u0656(.A0(men_men_n684_), .A1(men_men_n544_), .B0(men_men_n357_), .B1(men_men_n113_), .Y(men_men_n685_));
  OAI210     u0657(.A0(men_men_n682_), .A1(men_men_n681_), .B0(men_men_n685_), .Y(men_men_n686_));
  NO3        u0658(.A(men_men_n450_), .B(men_men_n177_), .C(i), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n454_), .B(men_men_n85_), .Y(men_men_n688_));
  NO4        u0660(.A(men_men_n519_), .B(men_men_n688_), .C(men_men_n133_), .D(men_men_n215_), .Y(men_men_n689_));
  INV        u0661(.A(men_men_n689_), .Y(men_men_n690_));
  NA3        u0662(.A(men_men_n690_), .B(men_men_n504_), .C(men_men_n396_), .Y(men_men_n691_));
  NO4        u0663(.A(men_men_n691_), .B(men_men_n686_), .C(men_men_n678_), .D(men_men_n665_), .Y(men_men_n692_));
  NA4        u0664(.A(men_men_n692_), .B(men_men_n657_), .C(men_men_n610_), .D(men_men_n576_), .Y(men08));
  NO2        u0665(.A(k), .B(h), .Y(men_men_n694_));
  AO210      u0666(.A0(men_men_n251_), .A1(men_men_n443_), .B0(men_men_n694_), .Y(men_men_n695_));
  NO2        u0667(.A(men_men_n695_), .B(men_men_n295_), .Y(men_men_n696_));
  INV        u0668(.A(men_men_n617_), .Y(men_men_n697_));
  AOI210     u0669(.A0(men_men_n1517_), .A1(men_men_n696_), .B0(men_men_n481_), .Y(men_men_n698_));
  NA2        u0670(.A(men_men_n85_), .B(men_men_n112_), .Y(men_men_n699_));
  NO2        u0671(.A(men_men_n699_), .B(men_men_n57_), .Y(men_men_n700_));
  NO4        u0672(.A(men_men_n377_), .B(men_men_n114_), .C(j), .D(men_men_n216_), .Y(men_men_n701_));
  AOI220     u0673(.A0(b), .A1(men_men_n344_), .B0(men_men_n701_), .B1(men_men_n700_), .Y(men_men_n702_));
  AOI210     u0674(.A0(men_men_n572_), .A1(men_men_n159_), .B0(men_men_n85_), .Y(men_men_n703_));
  NA4        u0675(.A(men_men_n218_), .B(men_men_n143_), .C(men_men_n45_), .D(h), .Y(men_men_n704_));
  AN2        u0676(.A(l), .B(k), .Y(men_men_n705_));
  NA4        u0677(.A(men_men_n705_), .B(men_men_n110_), .C(men_men_n74_), .D(men_men_n216_), .Y(men_men_n706_));
  OAI210     u0678(.A0(men_men_n704_), .A1(g), .B0(men_men_n706_), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n707_), .B(men_men_n703_), .Y(men_men_n708_));
  NA4        u0680(.A(men_men_n708_), .B(men_men_n702_), .C(men_men_n698_), .D(men_men_n346_), .Y(men_men_n709_));
  AN2        u0681(.A(men_men_n527_), .B(men_men_n97_), .Y(men_men_n710_));
  NO4        u0682(.A(men_men_n177_), .B(men_men_n387_), .C(men_men_n114_), .D(g), .Y(men_men_n711_));
  AOI210     u0683(.A0(men_men_n711_), .A1(b), .B0(men_men_n511_), .Y(men_men_n712_));
  NO2        u0684(.A(men_men_n38_), .B(men_men_n215_), .Y(men_men_n713_));
  AOI220     u0685(.A0(men_men_n619_), .A1(men_men_n343_), .B0(men_men_n713_), .B1(men_men_n559_), .Y(men_men_n714_));
  NAi31      u0686(.An(men_men_n710_), .B(men_men_n714_), .C(men_men_n712_), .Y(men_men_n715_));
  NO2        u0687(.A(men_men_n530_), .B(men_men_n35_), .Y(men_men_n716_));
  OAI210     u0688(.A0(men_men_n547_), .A1(men_men_n47_), .B0(men_men_n653_), .Y(men_men_n717_));
  NO2        u0689(.A(men_men_n473_), .B(men_men_n134_), .Y(men_men_n718_));
  AOI210     u0690(.A0(men_men_n718_), .A1(men_men_n717_), .B0(men_men_n716_), .Y(men_men_n719_));
  NO3        u0691(.A(m), .B(men_men_n133_), .C(men_men_n41_), .Y(men_men_n720_));
  NAi21      u0692(.An(men_men_n720_), .B(men_men_n706_), .Y(men_men_n721_));
  NA2        u0693(.A(men_men_n721_), .B(men_men_n77_), .Y(men_men_n722_));
  OAI210     u0694(.A0(men_men_n719_), .A1(men_men_n88_), .B0(men_men_n722_), .Y(men_men_n723_));
  NA2        u0695(.A(men_men_n359_), .B(men_men_n43_), .Y(men_men_n724_));
  NA2        u0696(.A(men_men_n705_), .B(men_men_n223_), .Y(men_men_n725_));
  NO2        u0697(.A(men_men_n725_), .B(men_men_n322_), .Y(men_men_n726_));
  AOI210     u0698(.A0(men_men_n726_), .A1(men_men_n679_), .B0(men_men_n480_), .Y(men_men_n727_));
  NA3        u0699(.A(m), .B(l), .C(k), .Y(men_men_n728_));
  AOI210     u0700(.A0(men_men_n662_), .A1(men_men_n660_), .B0(men_men_n728_), .Y(men_men_n729_));
  NO2        u0701(.A(men_men_n529_), .B(men_men_n269_), .Y(men_men_n730_));
  NOi21      u0702(.An(men_men_n730_), .B(men_men_n523_), .Y(men_men_n731_));
  NA4        u0703(.A(men_men_n115_), .B(l), .C(k), .D(men_men_n88_), .Y(men_men_n732_));
  NA3        u0704(.A(men_men_n122_), .B(men_men_n405_), .C(i), .Y(men_men_n733_));
  NO2        u0705(.A(men_men_n733_), .B(men_men_n732_), .Y(men_men_n734_));
  NO3        u0706(.A(men_men_n734_), .B(men_men_n731_), .C(men_men_n729_), .Y(men_men_n735_));
  NA3        u0707(.A(men_men_n735_), .B(men_men_n727_), .C(men_men_n724_), .Y(men_men_n736_));
  NO4        u0708(.A(men_men_n736_), .B(men_men_n723_), .C(men_men_n715_), .D(men_men_n709_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n619_), .B(men_men_n388_), .Y(men_men_n738_));
  NOi31      u0710(.An(g), .B(h), .C(f), .Y(men_men_n739_));
  NA2        u0711(.A(men_men_n635_), .B(men_men_n739_), .Y(men_men_n740_));
  AO210      u0712(.A0(men_men_n740_), .A1(men_men_n586_), .B0(men_men_n532_), .Y(men_men_n741_));
  NO3        u0713(.A(men_men_n391_), .B(men_men_n517_), .C(h), .Y(men_men_n742_));
  AOI210     u0714(.A0(men_men_n742_), .A1(men_men_n115_), .B0(men_men_n491_), .Y(men_men_n743_));
  NA4        u0715(.A(men_men_n743_), .B(men_men_n741_), .C(men_men_n738_), .D(men_men_n250_), .Y(men_men_n744_));
  NA2        u0716(.A(men_men_n705_), .B(men_men_n74_), .Y(men_men_n745_));
  NOi21      u0717(.An(h), .B(j), .Y(men_men_n746_));
  NA2        u0718(.A(men_men_n746_), .B(f), .Y(men_men_n747_));
  NO2        u0719(.A(men_men_n747_), .B(men_men_n244_), .Y(men_men_n748_));
  NO2        u0720(.A(men_men_n748_), .B(men_men_n687_), .Y(men_men_n749_));
  OAI220     u0721(.A0(men_men_n749_), .A1(men_men_n745_), .B0(men_men_n588_), .B1(men_men_n61_), .Y(men_men_n750_));
  AOI210     u0722(.A0(men_men_n744_), .A1(l), .B0(men_men_n750_), .Y(men_men_n751_));
  NO2        u0723(.A(j), .B(i), .Y(men_men_n752_));
  NA3        u0724(.A(men_men_n752_), .B(men_men_n81_), .C(l), .Y(men_men_n753_));
  NA2        u0725(.A(men_men_n752_), .B(men_men_n33_), .Y(men_men_n754_));
  NA2        u0726(.A(men_men_n415_), .B(men_men_n122_), .Y(men_men_n755_));
  OA220      u0727(.A0(men_men_n755_), .A1(men_men_n754_), .B0(men_men_n753_), .B1(men_men_n584_), .Y(men_men_n756_));
  NO3        u0728(.A(men_men_n154_), .B(men_men_n49_), .C(men_men_n112_), .Y(men_men_n757_));
  NO3        u0729(.A(men_men_n536_), .B(men_men_n153_), .C(men_men_n74_), .Y(men_men_n758_));
  NO3        u0730(.A(men_men_n473_), .B(men_men_n430_), .C(j), .Y(men_men_n759_));
  OAI210     u0731(.A0(men_men_n758_), .A1(men_men_n757_), .B0(men_men_n759_), .Y(men_men_n760_));
  OAI210     u0732(.A0(men_men_n740_), .A1(men_men_n61_), .B0(men_men_n760_), .Y(men_men_n761_));
  NA2        u0733(.A(k), .B(j), .Y(men_men_n762_));
  NO3        u0734(.A(men_men_n295_), .B(men_men_n762_), .C(men_men_n40_), .Y(men_men_n763_));
  AOI210     u0735(.A0(men_men_n522_), .A1(n), .B0(men_men_n546_), .Y(men_men_n764_));
  NA2        u0736(.A(men_men_n764_), .B(men_men_n548_), .Y(men_men_n765_));
  AN3        u0737(.A(men_men_n765_), .B(men_men_n763_), .C(men_men_n100_), .Y(men_men_n766_));
  NO3        u0738(.A(men_men_n177_), .B(men_men_n387_), .C(men_men_n114_), .Y(men_men_n767_));
  AOI220     u0739(.A0(men_men_n767_), .A1(men_men_n245_), .B0(c), .B1(men_men_n305_), .Y(men_men_n768_));
  NAi21      u0740(.An(men_men_n606_), .B(men_men_n94_), .Y(men_men_n769_));
  NA2        u0741(.A(men_men_n769_), .B(men_men_n768_), .Y(men_men_n770_));
  NO2        u0742(.A(men_men_n295_), .B(men_men_n138_), .Y(men_men_n771_));
  AOI220     u0743(.A0(men_men_n771_), .A1(men_men_n619_), .B0(men_men_n720_), .B1(men_men_n703_), .Y(men_men_n772_));
  NO2        u0744(.A(men_men_n728_), .B(men_men_n92_), .Y(men_men_n773_));
  NA2        u0745(.A(men_men_n773_), .B(men_men_n583_), .Y(men_men_n774_));
  NO2        u0746(.A(men_men_n585_), .B(men_men_n118_), .Y(men_men_n775_));
  OAI210     u0747(.A0(men_men_n775_), .A1(men_men_n759_), .B0(men_men_n675_), .Y(men_men_n776_));
  NA3        u0748(.A(men_men_n776_), .B(men_men_n774_), .C(men_men_n772_), .Y(men_men_n777_));
  OR4        u0749(.A(men_men_n777_), .B(men_men_n770_), .C(men_men_n766_), .D(men_men_n761_), .Y(men_men_n778_));
  NA3        u0750(.A(men_men_n764_), .B(men_men_n548_), .C(men_men_n547_), .Y(men_men_n779_));
  NA3        u0751(.A(men_men_n779_), .B(men_men_n218_), .C(men_men_n34_), .Y(men_men_n780_));
  NO4        u0752(.A(men_men_n473_), .B(men_men_n426_), .C(j), .D(f), .Y(men_men_n781_));
  OAI220     u0753(.A0(men_men_n704_), .A1(men_men_n697_), .B0(men_men_n327_), .B1(men_men_n38_), .Y(men_men_n782_));
  AOI210     u0754(.A0(men_men_n781_), .A1(men_men_n254_), .B0(men_men_n782_), .Y(men_men_n783_));
  NA3        u0755(.A(men_men_n539_), .B(men_men_n288_), .C(h), .Y(men_men_n784_));
  NOi21      u0756(.An(men_men_n675_), .B(men_men_n784_), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n93_), .B(men_men_n47_), .Y(men_men_n786_));
  OAI220     u0758(.A0(men_men_n784_), .A1(men_men_n602_), .B0(men_men_n753_), .B1(men_men_n72_), .Y(men_men_n787_));
  AOI210     u0759(.A0(men_men_n786_), .A1(men_men_n641_), .B0(men_men_n787_), .Y(men_men_n788_));
  NAi41      u0760(.An(men_men_n785_), .B(men_men_n788_), .C(men_men_n783_), .D(men_men_n780_), .Y(men_men_n789_));
  OR2        u0761(.A(men_men_n773_), .B(men_men_n97_), .Y(men_men_n790_));
  AOI220     u0762(.A0(men_men_n790_), .A1(men_men_n235_), .B0(men_men_n759_), .B1(men_men_n633_), .Y(men_men_n791_));
  NO2        u0763(.A(men_men_n661_), .B(men_men_n74_), .Y(men_men_n792_));
  AOI210     u0764(.A0(men_men_n781_), .A1(men_men_n792_), .B0(men_men_n331_), .Y(men_men_n793_));
  OAI210     u0765(.A0(men_men_n728_), .A1(men_men_n659_), .B0(men_men_n510_), .Y(men_men_n794_));
  NA3        u0766(.A(men_men_n248_), .B(men_men_n59_), .C(b), .Y(men_men_n795_));
  AOI220     u0767(.A0(men_men_n601_), .A1(men_men_n29_), .B0(men_men_n454_), .B1(men_men_n85_), .Y(men_men_n796_));
  NA2        u0768(.A(men_men_n796_), .B(men_men_n795_), .Y(men_men_n797_));
  NO2        u0769(.A(men_men_n784_), .B(men_men_n479_), .Y(men_men_n798_));
  AOI210     u0770(.A0(men_men_n797_), .A1(men_men_n794_), .B0(men_men_n798_), .Y(men_men_n799_));
  NA3        u0771(.A(men_men_n799_), .B(men_men_n793_), .C(men_men_n791_), .Y(men_men_n800_));
  NOi41      u0772(.An(men_men_n756_), .B(men_men_n800_), .C(men_men_n789_), .D(men_men_n778_), .Y(men_men_n801_));
  NO3        u0773(.A(men_men_n337_), .B(men_men_n297_), .C(men_men_n114_), .Y(men_men_n802_));
  NA2        u0774(.A(men_men_n802_), .B(men_men_n765_), .Y(men_men_n803_));
  NA2        u0775(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n804_));
  NO3        u0776(.A(men_men_n804_), .B(men_men_n754_), .C(men_men_n274_), .Y(men_men_n805_));
  NO3        u0777(.A(men_men_n517_), .B(men_men_n95_), .C(h), .Y(men_men_n806_));
  AOI210     u0778(.A0(men_men_n806_), .A1(men_men_n700_), .B0(men_men_n805_), .Y(men_men_n807_));
  NA3        u0779(.A(men_men_n807_), .B(men_men_n803_), .C(men_men_n398_), .Y(men_men_n808_));
  OR2        u0780(.A(men_men_n659_), .B(men_men_n93_), .Y(men_men_n809_));
  NOi31      u0781(.An(b), .B(d), .C(a), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n810_), .B(men_men_n599_), .Y(men_men_n811_));
  NO2        u0783(.A(men_men_n811_), .B(n), .Y(men_men_n812_));
  NOi21      u0784(.An(men_men_n796_), .B(men_men_n812_), .Y(men_men_n813_));
  OAI220     u0785(.A0(men_men_n813_), .A1(men_men_n809_), .B0(men_men_n784_), .B1(men_men_n600_), .Y(men_men_n814_));
  INV        u0786(.A(men_men_n547_), .Y(men_men_n815_));
  NO3        u0787(.A(men_men_n618_), .B(men_men_n322_), .C(men_men_n118_), .Y(men_men_n816_));
  NOi21      u0788(.An(men_men_n816_), .B(men_men_n164_), .Y(men_men_n817_));
  AOI210     u0789(.A0(men_men_n802_), .A1(men_men_n815_), .B0(men_men_n817_), .Y(men_men_n818_));
  OAI210     u0790(.A0(men_men_n704_), .A1(men_men_n389_), .B0(men_men_n818_), .Y(men_men_n819_));
  NA2        u0791(.A(men_men_n771_), .B(men_men_n666_), .Y(men_men_n820_));
  NO2        u0792(.A(men_men_n318_), .B(men_men_n234_), .Y(men_men_n821_));
  OAI210     u0793(.A0(men_men_n97_), .A1(men_men_n94_), .B0(men_men_n821_), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n122_), .B(men_men_n85_), .Y(men_men_n823_));
  AOI210     u0795(.A0(men_men_n419_), .A1(men_men_n411_), .B0(men_men_n823_), .Y(men_men_n824_));
  NAi21      u0796(.An(men_men_n824_), .B(men_men_n822_), .Y(men_men_n825_));
  NA2        u0797(.A(men_men_n726_), .B(men_men_n34_), .Y(men_men_n826_));
  NAi21      u0798(.An(men_men_n732_), .B(men_men_n427_), .Y(men_men_n827_));
  OAI210     u0799(.A0(men_men_n591_), .A1(men_men_n590_), .B0(men_men_n360_), .Y(men_men_n828_));
  AN2        u0800(.A(men_men_n828_), .B(men_men_n827_), .Y(men_men_n829_));
  NAi41      u0801(.An(men_men_n825_), .B(men_men_n829_), .C(men_men_n826_), .D(men_men_n820_), .Y(men_men_n830_));
  NO4        u0802(.A(men_men_n830_), .B(men_men_n819_), .C(men_men_n814_), .D(men_men_n808_), .Y(men_men_n831_));
  NA4        u0803(.A(men_men_n831_), .B(men_men_n801_), .C(men_men_n751_), .D(men_men_n737_), .Y(men09));
  INV        u0804(.A(men_men_n123_), .Y(men_men_n833_));
  NA2        u0805(.A(f), .B(e), .Y(men_men_n834_));
  NO2        u0806(.A(men_men_n227_), .B(men_men_n114_), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n835_), .B(g), .Y(men_men_n836_));
  NA4        u0808(.A(men_men_n308_), .B(men_men_n461_), .C(men_men_n257_), .D(men_men_n120_), .Y(men_men_n837_));
  AOI210     u0809(.A0(men_men_n837_), .A1(g), .B0(men_men_n458_), .Y(men_men_n838_));
  AOI210     u0810(.A0(men_men_n838_), .A1(men_men_n836_), .B0(men_men_n834_), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n436_), .B(e), .Y(men_men_n840_));
  INV        u0812(.A(men_men_n840_), .Y(men_men_n841_));
  AOI210     u0813(.A0(men_men_n839_), .A1(men_men_n833_), .B0(men_men_n841_), .Y(men_men_n842_));
  NO2        u0814(.A(men_men_n205_), .B(men_men_n215_), .Y(men_men_n843_));
  NA3        u0815(.A(m), .B(l), .C(i), .Y(men_men_n844_));
  OAI220     u0816(.A0(men_men_n585_), .A1(men_men_n844_), .B0(men_men_n350_), .B1(men_men_n518_), .Y(men_men_n845_));
  NA4        u0817(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(f), .Y(men_men_n846_));
  NAi31      u0818(.An(men_men_n845_), .B(men_men_n846_), .C(men_men_n431_), .Y(men_men_n847_));
  OA210      u0819(.A0(men_men_n847_), .A1(men_men_n843_), .B0(men_men_n559_), .Y(men_men_n848_));
  NA3        u0820(.A(men_men_n809_), .B(men_men_n561_), .C(men_men_n510_), .Y(men_men_n849_));
  OA210      u0821(.A0(men_men_n849_), .A1(men_men_n848_), .B0(men_men_n812_), .Y(men_men_n850_));
  INV        u0822(.A(men_men_n334_), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n852_));
  NOi31      u0824(.An(k), .B(m), .C(l), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n336_), .B(men_men_n853_), .Y(men_men_n854_));
  AOI210     u0826(.A0(men_men_n854_), .A1(men_men_n852_), .B0(men_men_n594_), .Y(men_men_n855_));
  NA2        u0827(.A(men_men_n795_), .B(men_men_n327_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n338_), .B(men_men_n340_), .Y(men_men_n857_));
  OAI210     u0829(.A0(men_men_n205_), .A1(men_men_n215_), .B0(men_men_n857_), .Y(men_men_n858_));
  AOI220     u0830(.A0(men_men_n858_), .A1(men_men_n856_), .B0(men_men_n855_), .B1(men_men_n851_), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n173_), .B(k), .Y(men_men_n860_));
  NA2        u0832(.A(men_men_n860_), .B(men_men_n695_), .Y(men_men_n861_));
  NA3        u0833(.A(men_men_n861_), .B(men_men_n193_), .C(men_men_n31_), .Y(men_men_n862_));
  NA4        u0834(.A(men_men_n862_), .B(men_men_n859_), .C(men_men_n620_), .D(men_men_n83_), .Y(men_men_n863_));
  NO2        u0835(.A(men_men_n581_), .B(men_men_n487_), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n864_), .B(men_men_n193_), .Y(men_men_n865_));
  NO2        u0837(.A(d), .B(men_men_n52_), .Y(men_men_n866_));
  NOi32      u0838(.An(g), .Bn(f), .C(d), .Y(men_men_n867_));
  NA4        u0839(.A(men_men_n867_), .B(men_men_n601_), .C(men_men_n29_), .D(m), .Y(men_men_n868_));
  NOi21      u0840(.An(men_men_n309_), .B(men_men_n868_), .Y(men_men_n869_));
  AOI210     u0841(.A0(men_men_n866_), .A1(men_men_n537_), .B0(men_men_n869_), .Y(men_men_n870_));
  NA3        u0842(.A(men_men_n308_), .B(men_men_n257_), .C(men_men_n120_), .Y(men_men_n871_));
  AN2        u0843(.A(f), .B(d), .Y(men_men_n872_));
  NA3        u0844(.A(men_men_n466_), .B(men_men_n872_), .C(men_men_n85_), .Y(men_men_n873_));
  NO3        u0845(.A(men_men_n873_), .B(men_men_n74_), .C(men_men_n216_), .Y(men_men_n874_));
  INV        u0846(.A(men_men_n281_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n871_), .B(men_men_n874_), .Y(men_men_n876_));
  NAi41      u0848(.An(men_men_n478_), .B(men_men_n876_), .C(men_men_n870_), .D(men_men_n865_), .Y(men_men_n877_));
  NO4        u0849(.A(men_men_n618_), .B(men_men_n134_), .C(men_men_n322_), .D(men_men_n155_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n652_), .B(men_men_n322_), .Y(men_men_n879_));
  AN2        u0851(.A(men_men_n879_), .B(men_men_n679_), .Y(men_men_n880_));
  NO3        u0852(.A(men_men_n880_), .B(men_men_n878_), .C(men_men_n232_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n599_), .B(men_men_n85_), .Y(men_men_n882_));
  OAI220     u0854(.A0(men_men_n857_), .A1(men_men_n882_), .B0(men_men_n795_), .B1(men_men_n431_), .Y(men_men_n883_));
  NA3        u0855(.A(men_men_n163_), .B(men_men_n110_), .C(men_men_n109_), .Y(men_men_n884_));
  OAI220     u0856(.A0(men_men_n873_), .A1(men_men_n424_), .B0(men_men_n334_), .B1(men_men_n884_), .Y(men_men_n885_));
  NOi31      u0857(.An(men_men_n225_), .B(men_men_n885_), .C(men_men_n883_), .Y(men_men_n886_));
  NA2        u0858(.A(c), .B(men_men_n117_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n887_), .B(men_men_n402_), .Y(men_men_n888_));
  NA3        u0860(.A(men_men_n888_), .B(men_men_n500_), .C(f), .Y(men_men_n889_));
  OR2        u0861(.A(men_men_n659_), .B(men_men_n533_), .Y(men_men_n890_));
  INV        u0862(.A(men_men_n890_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n811_), .B(men_men_n113_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n892_), .B(men_men_n891_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n889_), .C(men_men_n886_), .D(men_men_n881_), .Y(men_men_n894_));
  NO4        u0866(.A(men_men_n894_), .B(men_men_n877_), .C(men_men_n863_), .D(men_men_n850_), .Y(men_men_n895_));
  BUFFER     u0867(.A(men_men_n873_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n835_), .B(g), .Y(men_men_n897_));
  AOI210     u0869(.A0(men_men_n897_), .A1(men_men_n289_), .B0(men_men_n896_), .Y(men_men_n898_));
  AOI210     u0870(.A0(men_men_n795_), .A1(men_men_n327_), .B0(men_men_n846_), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n900_));
  NA2        u0872(.A(men_men_n302_), .B(men_men_n900_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n424_), .B(men_men_n834_), .Y(men_men_n902_));
  NA2        u0874(.A(men_men_n902_), .B(men_men_n553_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n903_), .B(men_men_n901_), .Y(men_men_n904_));
  NA2        u0876(.A(e), .B(d), .Y(men_men_n905_));
  NA2        u0877(.A(men_men_n619_), .B(men_men_n343_), .Y(men_men_n906_));
  NA2        u0878(.A(men_men_n281_), .B(men_men_n169_), .Y(men_men_n907_));
  NA2        u0879(.A(men_men_n874_), .B(men_men_n907_), .Y(men_men_n908_));
  NA3        u0880(.A(men_men_n172_), .B(men_men_n86_), .C(men_men_n34_), .Y(men_men_n909_));
  NA3        u0881(.A(men_men_n909_), .B(men_men_n908_), .C(men_men_n906_), .Y(men_men_n910_));
  NO4        u0882(.A(men_men_n910_), .B(men_men_n904_), .C(men_men_n899_), .D(men_men_n898_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n851_), .B(men_men_n31_), .Y(men_men_n912_));
  OR2        u0884(.A(men_men_n912_), .B(men_men_n219_), .Y(men_men_n913_));
  NO2        u0885(.A(men_men_n297_), .B(j), .Y(men_men_n914_));
  AOI220     u0886(.A0(men_men_n914_), .A1(men_men_n879_), .B0(men_men_n611_), .B1(men_men_n617_), .Y(men_men_n915_));
  OAI210     u0887(.A0(men_men_n840_), .A1(d), .B0(men_men_n915_), .Y(men_men_n916_));
  OAI210     u0888(.A0(men_men_n835_), .A1(men_men_n907_), .B0(men_men_n867_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n917_), .B(men_men_n602_), .Y(men_men_n918_));
  AOI210     u0890(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n256_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n919_), .B(men_men_n868_), .Y(men_men_n920_));
  AO210      u0892(.A0(men_men_n856_), .A1(men_men_n845_), .B0(men_men_n920_), .Y(men_men_n921_));
  NOi31      u0893(.An(men_men_n537_), .B(d), .C(men_men_n289_), .Y(men_men_n922_));
  NO4        u0894(.A(men_men_n922_), .B(men_men_n921_), .C(men_men_n918_), .D(men_men_n916_), .Y(men_men_n923_));
  NO2        u0895(.A(men_men_n430_), .B(men_men_n70_), .Y(men_men_n924_));
  OAI210     u0896(.A0(men_men_n849_), .A1(men_men_n924_), .B0(men_men_n700_), .Y(men_men_n925_));
  AN4        u0897(.A(men_men_n925_), .B(men_men_n330_), .C(men_men_n923_), .D(men_men_n913_), .Y(men_men_n926_));
  NA4        u0898(.A(men_men_n926_), .B(men_men_n911_), .C(men_men_n895_), .D(men_men_n842_), .Y(men12));
  NO2        u0899(.A(men_men_n446_), .B(c), .Y(men_men_n928_));
  NO4        u0900(.A(men_men_n435_), .B(men_men_n251_), .C(men_men_n577_), .D(men_men_n216_), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n929_), .B(men_men_n928_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n537_), .B(men_men_n924_), .Y(men_men_n931_));
  NO2        u0903(.A(men_men_n446_), .B(men_men_n117_), .Y(men_men_n932_));
  NO2        u0904(.A(men_men_n852_), .B(men_men_n350_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n659_), .B(men_men_n377_), .Y(men_men_n934_));
  AOI220     u0906(.A0(men_men_n934_), .A1(men_men_n535_), .B0(men_men_n933_), .B1(men_men_n932_), .Y(men_men_n935_));
  NA4        u0907(.A(men_men_n935_), .B(men_men_n931_), .C(men_men_n930_), .D(men_men_n434_), .Y(men_men_n936_));
  AOI210     u0908(.A0(men_men_n231_), .A1(men_men_n333_), .B0(men_men_n202_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n330_), .B(men_men_n216_), .Y(men_men_n938_));
  NA2        u0910(.A(men_men_n938_), .B(f), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n638_), .B(men_men_n259_), .Y(men_men_n940_));
  NO2        u0912(.A(men_men_n585_), .B(men_men_n844_), .Y(men_men_n941_));
  AOI220     u0913(.A0(men_men_n941_), .A1(men_men_n559_), .B0(men_men_n821_), .B1(men_men_n940_), .Y(men_men_n942_));
  NO2        u0914(.A(men_men_n154_), .B(men_men_n234_), .Y(men_men_n943_));
  NA3        u0915(.A(men_men_n943_), .B(men_men_n237_), .C(i), .Y(men_men_n944_));
  NA3        u0916(.A(men_men_n944_), .B(men_men_n942_), .C(men_men_n939_), .Y(men_men_n945_));
  OR2        u0917(.A(men_men_n1519_), .B(men_men_n932_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n946_), .B(men_men_n351_), .Y(men_men_n947_));
  NO3        u0919(.A(men_men_n134_), .B(men_men_n155_), .C(men_men_n216_), .Y(men_men_n948_));
  NA2        u0920(.A(men_men_n948_), .B(men_men_n522_), .Y(men_men_n949_));
  NA3        u0921(.A(men_men_n436_), .B(men_men_n428_), .C(g), .Y(men_men_n950_));
  NA3        u0922(.A(men_men_n950_), .B(men_men_n949_), .C(men_men_n947_), .Y(men_men_n951_));
  NO3        u0923(.A(men_men_n664_), .B(men_men_n93_), .C(men_men_n45_), .Y(men_men_n952_));
  NO4        u0924(.A(men_men_n952_), .B(men_men_n951_), .C(men_men_n945_), .D(men_men_n936_), .Y(men_men_n953_));
  NO2        u0925(.A(men_men_n367_), .B(men_men_n366_), .Y(men_men_n954_));
  NA2        u0926(.A(men_men_n582_), .B(men_men_n72_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n547_), .B(men_men_n148_), .Y(men_men_n956_));
  NOi21      u0928(.An(men_men_n34_), .B(men_men_n652_), .Y(men_men_n957_));
  AOI220     u0929(.A0(men_men_n957_), .A1(men_men_n956_), .B0(men_men_n955_), .B1(men_men_n954_), .Y(men_men_n958_));
  OAI210     u0930(.A0(men_men_n249_), .A1(men_men_n45_), .B0(men_men_n958_), .Y(men_men_n959_));
  NA2        u0931(.A(men_men_n427_), .B(men_men_n261_), .Y(men_men_n960_));
  NO3        u0932(.A(men_men_n823_), .B(men_men_n90_), .C(men_men_n402_), .Y(men_men_n961_));
  NAi21      u0933(.An(men_men_n961_), .B(men_men_n960_), .Y(men_men_n962_));
  NO2        u0934(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n963_));
  NO2        u0935(.A(men_men_n494_), .B(men_men_n297_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n964_), .B(men_men_n363_), .Y(men_men_n965_));
  NO2        u0937(.A(men_men_n965_), .B(men_men_n148_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n629_), .B(men_men_n360_), .Y(men_men_n967_));
  OAI210     u0939(.A0(men_men_n733_), .A1(men_men_n967_), .B0(men_men_n364_), .Y(men_men_n968_));
  NO4        u0940(.A(men_men_n968_), .B(men_men_n966_), .C(men_men_n962_), .D(men_men_n959_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n343_), .B(g), .Y(men_men_n970_));
  NA2        u0942(.A(men_men_n166_), .B(i), .Y(men_men_n971_));
  OAI220     u0943(.A0(men_men_n1520_), .A1(men_men_n201_), .B0(men_men_n971_), .B1(men_men_n93_), .Y(men_men_n972_));
  AOI210     u0944(.A0(men_men_n413_), .A1(men_men_n37_), .B0(men_men_n972_), .Y(men_men_n973_));
  NO2        u0945(.A(men_men_n148_), .B(men_men_n85_), .Y(men_men_n974_));
  OR2        u0946(.A(men_men_n974_), .B(men_men_n546_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n547_), .B(men_men_n381_), .Y(men_men_n976_));
  NO2        u0948(.A(men_men_n976_), .B(men_men_n975_), .Y(men_men_n977_));
  OAI220     u0949(.A0(men_men_n977_), .A1(men_men_n970_), .B0(men_men_n973_), .B1(men_men_n327_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n659_), .B(men_men_n487_), .Y(men_men_n979_));
  NA3        u0951(.A(men_men_n338_), .B(men_men_n624_), .C(i), .Y(men_men_n980_));
  OAI210     u0952(.A0(men_men_n430_), .A1(men_men_n308_), .B0(men_men_n980_), .Y(men_men_n981_));
  OAI220     u0953(.A0(men_men_n981_), .A1(men_men_n979_), .B0(men_men_n675_), .B1(men_men_n758_), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n605_), .B(men_men_n115_), .Y(men_men_n983_));
  OR3        u0955(.A(men_men_n308_), .B(men_men_n426_), .C(f), .Y(men_men_n984_));
  NA3        u0956(.A(men_men_n624_), .B(men_men_n81_), .C(i), .Y(men_men_n985_));
  OA220      u0957(.A0(men_men_n985_), .A1(men_men_n983_), .B0(men_men_n984_), .B1(men_men_n584_), .Y(men_men_n986_));
  NA2        u0958(.A(men_men_n933_), .B(men_men_n1519_), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n688_), .B(men_men_n882_), .Y(men_men_n988_));
  NA2        u0960(.A(men_men_n846_), .B(men_men_n431_), .Y(men_men_n989_));
  NA2        u0961(.A(i), .B(men_men_n78_), .Y(men_men_n990_));
  NA3        u0962(.A(men_men_n990_), .B(men_men_n985_), .C(men_men_n984_), .Y(men_men_n991_));
  AOI220     u0963(.A0(men_men_n991_), .A1(men_men_n254_), .B0(men_men_n989_), .B1(men_men_n988_), .Y(men_men_n992_));
  NA4        u0964(.A(men_men_n992_), .B(men_men_n987_), .C(men_men_n986_), .D(men_men_n982_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n940_), .B(men_men_n235_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n663_), .B(men_men_n89_), .Y(men_men_n995_));
  NO2        u0967(.A(men_men_n449_), .B(men_men_n216_), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n946_), .B(men_men_n220_), .Y(men_men_n997_));
  AOI220     u0969(.A0(men_men_n934_), .A1(men_men_n943_), .B0(men_men_n583_), .B1(men_men_n91_), .Y(men_men_n998_));
  NA4        u0970(.A(men_men_n998_), .B(men_men_n997_), .C(men_men_n995_), .D(men_men_n994_), .Y(men_men_n999_));
  OAI210     u0971(.A0(men_men_n989_), .A1(men_men_n941_), .B0(men_men_n535_), .Y(men_men_n1000_));
  AOI210     u0972(.A0(men_men_n414_), .A1(men_men_n406_), .B0(men_men_n823_), .Y(men_men_n1001_));
  OAI210     u0973(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n111_), .Y(men_men_n1002_));
  AOI210     u0974(.A0(men_men_n1002_), .A1(men_men_n527_), .B0(men_men_n1001_), .Y(men_men_n1003_));
  NO3        u0975(.A(l), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1004_));
  AOI220     u0976(.A0(men_men_n1004_), .A1(men_men_n622_), .B0(men_men_n643_), .B1(men_men_n522_), .Y(men_men_n1005_));
  NA3        u0977(.A(men_men_n1005_), .B(men_men_n1003_), .C(men_men_n1000_), .Y(men_men_n1006_));
  NO4        u0978(.A(men_men_n1006_), .B(men_men_n999_), .C(men_men_n993_), .D(men_men_n978_), .Y(men_men_n1007_));
  NAi31      u0979(.An(men_men_n144_), .B(men_men_n415_), .C(n), .Y(men_men_n1008_));
  NO3        u0980(.A(men_men_n127_), .B(men_men_n336_), .C(men_men_n853_), .Y(men_men_n1009_));
  NO2        u0981(.A(men_men_n1009_), .B(men_men_n1008_), .Y(men_men_n1010_));
  NO3        u0982(.A(men_men_n269_), .B(men_men_n144_), .C(men_men_n402_), .Y(men_men_n1011_));
  AOI210     u0983(.A0(men_men_n1011_), .A1(men_men_n488_), .B0(men_men_n1010_), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n481_), .B(i), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n1013_), .B(men_men_n1012_), .Y(men_men_n1014_));
  NA2        u0986(.A(men_men_n229_), .B(men_men_n176_), .Y(men_men_n1015_));
  NO3        u0987(.A(men_men_n305_), .B(men_men_n436_), .C(men_men_n179_), .Y(men_men_n1016_));
  NOi31      u0988(.An(men_men_n1015_), .B(men_men_n1016_), .C(men_men_n216_), .Y(men_men_n1017_));
  NAi21      u0989(.An(men_men_n547_), .B(men_men_n996_), .Y(men_men_n1018_));
  NA2        u0990(.A(men_men_n429_), .B(men_men_n882_), .Y(men_men_n1019_));
  NO3        u0991(.A(men_men_n430_), .B(men_men_n308_), .C(men_men_n74_), .Y(men_men_n1020_));
  NA2        u0992(.A(men_men_n1020_), .B(men_men_n1019_), .Y(men_men_n1021_));
  NA2        u0993(.A(men_men_n1021_), .B(men_men_n1018_), .Y(men_men_n1022_));
  OAI220     u0994(.A0(men_men_n1008_), .A1(men_men_n231_), .B0(men_men_n980_), .B1(men_men_n600_), .Y(men_men_n1023_));
  NO2        u0995(.A(men_men_n660_), .B(men_men_n377_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n937_), .B(men_men_n928_), .Y(men_men_n1025_));
  NO3        u0997(.A(men_men_n536_), .B(men_men_n153_), .C(men_men_n215_), .Y(men_men_n1026_));
  OAI210     u0998(.A0(men_men_n1026_), .A1(men_men_n516_), .B0(men_men_n378_), .Y(men_men_n1027_));
  OAI220     u0999(.A0(men_men_n934_), .A1(men_men_n941_), .B0(men_men_n537_), .B1(men_men_n423_), .Y(men_men_n1028_));
  NA4        u1000(.A(men_men_n1028_), .B(men_men_n1027_), .C(men_men_n1025_), .D(men_men_n616_), .Y(men_men_n1029_));
  NA3        u1001(.A(men_men_n976_), .B(men_men_n475_), .C(men_men_n46_), .Y(men_men_n1030_));
  AOI210     u1002(.A0(men_men_n380_), .A1(men_men_n378_), .B0(men_men_n326_), .Y(men_men_n1031_));
  NA3        u1003(.A(men_men_n1031_), .B(men_men_n1030_), .C(men_men_n270_), .Y(men_men_n1032_));
  OR4        u1004(.A(men_men_n1032_), .B(men_men_n1029_), .C(men_men_n1024_), .D(men_men_n1023_), .Y(men_men_n1033_));
  NO4        u1005(.A(men_men_n1033_), .B(men_men_n1022_), .C(men_men_n1017_), .D(men_men_n1014_), .Y(men_men_n1034_));
  NA4        u1006(.A(men_men_n1034_), .B(men_men_n1007_), .C(men_men_n969_), .D(men_men_n953_), .Y(men13));
  NA2        u1007(.A(men_men_n46_), .B(men_men_n88_), .Y(men_men_n1036_));
  NA3        u1008(.A(men_men_n248_), .B(c), .C(m), .Y(men_men_n1037_));
  NO4        u1009(.A(e), .B(men_men_n1037_), .C(men_men_n1036_), .D(men_men_n578_), .Y(men_men_n1038_));
  NA2        u1010(.A(men_men_n261_), .B(c), .Y(men_men_n1039_));
  NO4        u1011(.A(men_men_n1039_), .B(e), .C(men_men_n971_), .D(a), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n143_), .B(men_men_n45_), .Y(men_men_n1041_));
  NO4        u1013(.A(men_men_n1041_), .B(d), .C(men_men_n585_), .D(men_men_n304_), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n667_), .B(men_men_n226_), .Y(men_men_n1043_));
  NA2        u1015(.A(men_men_n405_), .B(men_men_n215_), .Y(men_men_n1044_));
  AN2        u1016(.A(d), .B(c), .Y(men_men_n1045_));
  NA2        u1017(.A(men_men_n1045_), .B(men_men_n117_), .Y(men_men_n1046_));
  NO3        u1018(.A(men_men_n1046_), .B(men_men_n1044_), .C(men_men_n180_), .Y(men_men_n1047_));
  NO3        u1019(.A(men_men_n1041_), .B(men_men_n581_), .C(men_men_n304_), .Y(men_men_n1048_));
  AO210      u1020(.A0(men_men_n1047_), .A1(men_men_n1043_), .B0(men_men_n1048_), .Y(men_men_n1049_));
  OR4        u1021(.A(men_men_n1049_), .B(men_men_n1042_), .C(men_men_n1040_), .D(men_men_n1038_), .Y(men_men_n1050_));
  NAi32      u1022(.An(f), .Bn(e), .C(c), .Y(men_men_n1051_));
  NO2        u1023(.A(men_men_n1051_), .B(men_men_n150_), .Y(men_men_n1052_));
  NA2        u1024(.A(men_men_n1052_), .B(g), .Y(men_men_n1053_));
  OR2        u1025(.A(men_men_n226_), .B(men_men_n180_), .Y(men_men_n1054_));
  NO2        u1026(.A(men_men_n1054_), .B(men_men_n1053_), .Y(men_men_n1055_));
  INV        u1027(.A(men_men_n304_), .Y(men_men_n1056_));
  NO2        u1028(.A(j), .B(men_men_n45_), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n626_), .B(men_men_n1057_), .Y(men_men_n1058_));
  NOi21      u1030(.An(men_men_n1056_), .B(men_men_n1058_), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n762_), .B(men_men_n114_), .Y(men_men_n1060_));
  NOi41      u1032(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1061_));
  NO2        u1033(.A(men_men_n1518_), .B(men_men_n1053_), .Y(men_men_n1062_));
  NA3        u1034(.A(k), .B(j), .C(i), .Y(men_men_n1063_));
  NO3        u1035(.A(men_men_n1063_), .B(men_men_n304_), .C(men_men_n92_), .Y(men_men_n1064_));
  OR4        u1036(.A(men_men_n1064_), .B(men_men_n1062_), .C(men_men_n1059_), .D(men_men_n1055_), .Y(men_men_n1065_));
  NA3        u1037(.A(men_men_n457_), .B(men_men_n329_), .C(men_men_n56_), .Y(men_men_n1066_));
  NO3        u1038(.A(men_men_n1066_), .B(men_men_n581_), .C(men_men_n45_), .Y(men_men_n1067_));
  INV        u1039(.A(men_men_n435_), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n1068_), .B(men_men_n59_), .Y(men_men_n1069_));
  NO3        u1041(.A(k), .B(men_men_n241_), .C(l), .Y(men_men_n1070_));
  NOi21      u1042(.An(men_men_n1070_), .B(men_men_n1069_), .Y(men_men_n1071_));
  OR2        u1043(.A(men_men_n1071_), .B(men_men_n1067_), .Y(men_men_n1072_));
  OR3        u1044(.A(men_men_n1072_), .B(men_men_n1065_), .C(men_men_n1050_), .Y(men02));
  OR2        u1045(.A(l), .B(k), .Y(men_men_n1074_));
  OR3        u1046(.A(h), .B(g), .C(f), .Y(men_men_n1075_));
  OR3        u1047(.A(n), .B(m), .C(i), .Y(men_men_n1076_));
  NO4        u1048(.A(men_men_n1076_), .B(men_men_n1075_), .C(men_men_n1074_), .D(e), .Y(men_men_n1077_));
  NO2        u1049(.A(men_men_n1064_), .B(men_men_n1042_), .Y(men_men_n1078_));
  NA3        u1050(.A(c), .B(men_men_n457_), .C(h), .Y(men_men_n1079_));
  OR2        u1051(.A(men_men_n304_), .B(men_men_n1079_), .Y(men_men_n1080_));
  NO3        u1052(.A(men_men_n1066_), .B(men_men_n1041_), .C(men_men_n581_), .Y(men_men_n1081_));
  NO2        u1053(.A(men_men_n1081_), .B(men_men_n1055_), .Y(men_men_n1082_));
  NA3        u1054(.A(l), .B(k), .C(j), .Y(men_men_n1083_));
  NA2        u1055(.A(i), .B(h), .Y(men_men_n1084_));
  NO2        u1056(.A(men_men_n1084_), .B(men_men_n1083_), .Y(men_men_n1085_));
  NO3        u1057(.A(men_men_n145_), .B(men_men_n279_), .C(men_men_n216_), .Y(men_men_n1086_));
  AOI210     u1058(.A0(men_men_n1086_), .A1(men_men_n1085_), .B0(men_men_n1059_), .Y(men_men_n1087_));
  NA3        u1059(.A(c), .B(b), .C(a), .Y(men_men_n1088_));
  NO3        u1060(.A(men_men_n1088_), .B(men_men_n905_), .C(men_men_n215_), .Y(men_men_n1089_));
  AN3        u1061(.A(men_men_n1087_), .B(men_men_n1082_), .C(men_men_n1080_), .Y(men_men_n1090_));
  NO2        u1062(.A(men_men_n1046_), .B(men_men_n1044_), .Y(men_men_n1091_));
  NA2        u1063(.A(men_men_n1518_), .B(men_men_n1054_), .Y(men_men_n1092_));
  AOI210     u1064(.A0(men_men_n1092_), .A1(men_men_n1091_), .B0(men_men_n1038_), .Y(men_men_n1093_));
  NAi41      u1065(.An(men_men_n1077_), .B(men_men_n1093_), .C(men_men_n1090_), .D(men_men_n1078_), .Y(men03));
  NO2        u1066(.A(men_men_n518_), .B(men_men_n594_), .Y(men_men_n1095_));
  NA4        u1067(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(men_men_n215_), .Y(men_men_n1096_));
  NA4        u1068(.A(men_men_n569_), .B(m), .C(men_men_n114_), .D(men_men_n215_), .Y(men_men_n1097_));
  NA3        u1069(.A(men_men_n1097_), .B(men_men_n368_), .C(men_men_n1096_), .Y(men_men_n1098_));
  NO3        u1070(.A(men_men_n1098_), .B(men_men_n1095_), .C(men_men_n1002_), .Y(men_men_n1099_));
  NOi41      u1071(.An(men_men_n809_), .B(men_men_n858_), .C(men_men_n847_), .D(men_men_n713_), .Y(men_men_n1100_));
  OAI220     u1072(.A0(men_men_n1100_), .A1(men_men_n688_), .B0(men_men_n1099_), .B1(men_men_n582_), .Y(men_men_n1101_));
  NOi31      u1073(.An(i), .B(k), .C(j), .Y(men_men_n1102_));
  NA4        u1074(.A(men_men_n1102_), .B(e), .C(men_men_n338_), .D(men_men_n329_), .Y(men_men_n1103_));
  OAI210     u1075(.A0(men_men_n823_), .A1(men_men_n416_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  NOi31      u1076(.An(m), .B(n), .C(f), .Y(men_men_n1105_));
  NA2        u1077(.A(men_men_n1105_), .B(men_men_n51_), .Y(men_men_n1106_));
  AN2        u1078(.A(e), .B(c), .Y(men_men_n1107_));
  NA2        u1079(.A(men_men_n1107_), .B(a), .Y(men_men_n1108_));
  OAI220     u1080(.A0(men_men_n1108_), .A1(men_men_n1106_), .B0(men_men_n890_), .B1(men_men_n422_), .Y(men_men_n1109_));
  NA2        u1081(.A(men_men_n498_), .B(l), .Y(men_men_n1110_));
  NOi31      u1082(.An(men_men_n867_), .B(men_men_n1037_), .C(men_men_n1110_), .Y(men_men_n1111_));
  NO4        u1083(.A(men_men_n1111_), .B(men_men_n1109_), .C(men_men_n1104_), .D(men_men_n1001_), .Y(men_men_n1112_));
  NO2        u1084(.A(men_men_n279_), .B(a), .Y(men_men_n1113_));
  INV        u1085(.A(men_men_n1042_), .Y(men_men_n1114_));
  NO2        u1086(.A(men_men_n88_), .B(g), .Y(men_men_n1115_));
  AOI210     u1087(.A0(men_men_n1115_), .A1(i), .B0(men_men_n1070_), .Y(men_men_n1116_));
  OR2        u1088(.A(men_men_n1116_), .B(men_men_n1069_), .Y(men_men_n1117_));
  NA3        u1089(.A(men_men_n1117_), .B(men_men_n1114_), .C(men_men_n1112_), .Y(men_men_n1118_));
  NO4        u1090(.A(men_men_n1118_), .B(men_men_n1101_), .C(men_men_n825_), .D(men_men_n558_), .Y(men_men_n1119_));
  NA2        u1091(.A(c), .B(b), .Y(men_men_n1120_));
  NO2        u1092(.A(men_men_n699_), .B(men_men_n1120_), .Y(men_men_n1121_));
  OAI210     u1093(.A0(d), .A1(men_men_n838_), .B0(men_men_n409_), .Y(men_men_n1122_));
  OAI210     u1094(.A0(men_men_n1122_), .A1(men_men_n866_), .B0(men_men_n1121_), .Y(men_men_n1123_));
  NAi21      u1095(.An(men_men_n417_), .B(men_men_n1121_), .Y(men_men_n1124_));
  NA2        u1096(.A(men_men_n423_), .B(men_men_n551_), .Y(men_men_n1125_));
  OAI210     u1097(.A0(men_men_n541_), .A1(men_men_n39_), .B0(men_men_n1113_), .Y(men_men_n1126_));
  NA3        u1098(.A(men_men_n1126_), .B(men_men_n1125_), .C(men_men_n1124_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n257_), .B(men_men_n120_), .Y(men_men_n1128_));
  OAI210     u1100(.A0(men_men_n1128_), .A1(men_men_n283_), .B0(g), .Y(men_men_n1129_));
  NAi21      u1101(.An(f), .B(d), .Y(men_men_n1130_));
  NO2        u1102(.A(men_men_n1130_), .B(men_men_n1088_), .Y(men_men_n1131_));
  INV        u1103(.A(men_men_n1131_), .Y(men_men_n1132_));
  AOI210     u1104(.A0(men_men_n1129_), .A1(men_men_n289_), .B0(men_men_n1132_), .Y(men_men_n1133_));
  AOI210     u1105(.A0(men_men_n1133_), .A1(men_men_n115_), .B0(men_men_n1127_), .Y(men_men_n1134_));
  INV        u1106(.A(men_men_n458_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n186_), .B(men_men_n234_), .Y(men_men_n1136_));
  NA2        u1108(.A(men_men_n1136_), .B(m), .Y(men_men_n1137_));
  NA3        u1109(.A(men_men_n919_), .B(men_men_n1110_), .C(men_men_n461_), .Y(men_men_n1138_));
  OAI210     u1110(.A0(men_men_n1138_), .A1(men_men_n309_), .B0(men_men_n459_), .Y(men_men_n1139_));
  AOI210     u1111(.A0(men_men_n1139_), .A1(men_men_n1135_), .B0(men_men_n1137_), .Y(men_men_n1140_));
  NA2        u1112(.A(men_men_n553_), .B(men_men_n404_), .Y(men_men_n1141_));
  NA2        u1113(.A(men_men_n162_), .B(men_men_n33_), .Y(men_men_n1142_));
  AOI210     u1114(.A0(men_men_n967_), .A1(men_men_n1142_), .B0(men_men_n216_), .Y(men_men_n1143_));
  NA2        u1115(.A(men_men_n1143_), .B(men_men_n1131_), .Y(men_men_n1144_));
  NO2        u1116(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n1145_));
  AOI210     u1117(.A0(men_men_n1136_), .A1(men_men_n51_), .B0(men_men_n961_), .Y(men_men_n1146_));
  NAi41      u1118(.An(men_men_n1145_), .B(men_men_n1146_), .C(men_men_n1144_), .D(men_men_n1141_), .Y(men_men_n1147_));
  NO2        u1119(.A(men_men_n1147_), .B(men_men_n1140_), .Y(men_men_n1148_));
  NA4        u1120(.A(men_men_n1148_), .B(men_men_n1134_), .C(men_men_n1123_), .D(men_men_n1119_), .Y(men00));
  NO2        u1121(.A(men_men_n296_), .B(men_men_n273_), .Y(men_men_n1150_));
  NO2        u1122(.A(men_men_n1150_), .B(men_men_n572_), .Y(men_men_n1151_));
  AOI210     u1123(.A0(men_men_n902_), .A1(men_men_n943_), .B0(men_men_n1104_), .Y(men_men_n1152_));
  NO2        u1124(.A(men_men_n961_), .B(men_men_n710_), .Y(men_men_n1153_));
  NA3        u1125(.A(men_men_n1153_), .B(men_men_n1152_), .C(men_men_n1003_), .Y(men_men_n1154_));
  NA2        u1126(.A(men_men_n500_), .B(f), .Y(men_men_n1155_));
  OAI210     u1127(.A0(men_men_n1009_), .A1(men_men_n40_), .B0(men_men_n645_), .Y(men_men_n1156_));
  NA2        u1128(.A(men_men_n1156_), .B(men_men_n253_), .Y(men_men_n1157_));
  AOI210     u1129(.A0(men_men_n1157_), .A1(men_men_n1155_), .B0(men_men_n1046_), .Y(men_men_n1158_));
  NO4        u1130(.A(men_men_n1158_), .B(men_men_n1154_), .C(men_men_n1151_), .D(men_men_n1065_), .Y(men_men_n1159_));
  NA3        u1131(.A(men_men_n172_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1160_));
  NA3        u1132(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1161_));
  NOi31      u1133(.An(n), .B(m), .C(i), .Y(men_men_n1162_));
  NA3        u1134(.A(men_men_n1162_), .B(men_men_n648_), .C(men_men_n51_), .Y(men_men_n1163_));
  OAI210     u1135(.A0(men_men_n1161_), .A1(men_men_n1160_), .B0(men_men_n1163_), .Y(men_men_n1164_));
  INV        u1136(.A(men_men_n571_), .Y(men_men_n1165_));
  NO4        u1137(.A(men_men_n1165_), .B(men_men_n1164_), .C(men_men_n1145_), .D(men_men_n922_), .Y(men_men_n1166_));
  NO3        u1138(.A(men_men_n476_), .B(men_men_n353_), .C(men_men_n1120_), .Y(men_men_n1167_));
  NA3        u1139(.A(men_men_n383_), .B(men_men_n223_), .C(g), .Y(men_men_n1168_));
  OA220      u1140(.A0(men_men_n1168_), .A1(men_men_n1161_), .B0(men_men_n384_), .B1(men_men_n137_), .Y(men_men_n1169_));
  NO2        u1141(.A(h), .B(g), .Y(men_men_n1170_));
  NA4        u1142(.A(men_men_n488_), .B(men_men_n457_), .C(men_men_n1170_), .D(c), .Y(men_men_n1171_));
  OAI220     u1143(.A0(men_men_n518_), .A1(men_men_n594_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n1172_));
  AOI220     u1144(.A0(men_men_n1172_), .A1(men_men_n527_), .B0(men_men_n948_), .B1(men_men_n570_), .Y(men_men_n1173_));
  AOI220     u1145(.A0(men_men_n314_), .A1(men_men_n245_), .B0(men_men_n181_), .B1(men_men_n152_), .Y(men_men_n1174_));
  NA4        u1146(.A(men_men_n1174_), .B(men_men_n1173_), .C(men_men_n1171_), .D(men_men_n1169_), .Y(men_men_n1175_));
  NO3        u1147(.A(men_men_n1175_), .B(men_men_n1167_), .C(men_men_n263_), .Y(men_men_n1176_));
  INV        u1148(.A(men_men_n317_), .Y(men_men_n1177_));
  NA2        u1149(.A(men_men_n1177_), .B(men_men_n157_), .Y(men_men_n1178_));
  NO2        u1150(.A(men_men_n236_), .B(men_men_n185_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n1179_), .B(men_men_n423_), .Y(men_men_n1180_));
  NA3        u1152(.A(men_men_n183_), .B(men_men_n114_), .C(g), .Y(men_men_n1181_));
  NA3        u1153(.A(men_men_n457_), .B(men_men_n40_), .C(f), .Y(men_men_n1182_));
  NOi31      u1154(.An(men_men_n875_), .B(men_men_n1182_), .C(men_men_n1181_), .Y(men_men_n1183_));
  NAi31      u1155(.An(men_men_n189_), .B(men_men_n864_), .C(men_men_n457_), .Y(men_men_n1184_));
  NAi31      u1156(.An(men_men_n1183_), .B(men_men_n1184_), .C(men_men_n1180_), .Y(men_men_n1185_));
  NO2        u1157(.A(men_men_n272_), .B(men_men_n74_), .Y(men_men_n1186_));
  NO3        u1158(.A(men_men_n422_), .B(men_men_n834_), .C(n), .Y(men_men_n1187_));
  AOI210     u1159(.A0(men_men_n1187_), .A1(men_men_n1186_), .B0(men_men_n1077_), .Y(men_men_n1188_));
  NAi31      u1160(.An(men_men_n1048_), .B(men_men_n1188_), .C(men_men_n73_), .Y(men_men_n1189_));
  NO4        u1161(.A(men_men_n1189_), .B(men_men_n1185_), .C(men_men_n1178_), .D(men_men_n509_), .Y(men_men_n1190_));
  AN3        u1162(.A(men_men_n1190_), .B(men_men_n1176_), .C(men_men_n1166_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n527_), .B(men_men_n103_), .Y(men_men_n1192_));
  NA3        u1164(.A(men_men_n1105_), .B(men_men_n605_), .C(men_men_n456_), .Y(men_men_n1193_));
  NA4        u1165(.A(men_men_n1193_), .B(men_men_n554_), .C(men_men_n1192_), .D(men_men_n239_), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n1098_), .B(men_men_n527_), .Y(men_men_n1195_));
  NA4        u1167(.A(men_men_n648_), .B(men_men_n207_), .C(men_men_n223_), .D(men_men_n166_), .Y(men_men_n1196_));
  NA3        u1168(.A(men_men_n1196_), .B(men_men_n1195_), .C(men_men_n293_), .Y(men_men_n1197_));
  OAI210     u1169(.A0(men_men_n455_), .A1(men_men_n121_), .B0(men_men_n868_), .Y(men_men_n1198_));
  AOI220     u1170(.A0(men_men_n1198_), .A1(men_men_n1138_), .B0(men_men_n553_), .B1(men_men_n404_), .Y(men_men_n1199_));
  OR4        u1171(.A(men_men_n1046_), .B(men_men_n269_), .C(men_men_n224_), .D(e), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n219_), .B(men_men_n216_), .Y(men_men_n1201_));
  NA2        u1173(.A(n), .B(e), .Y(men_men_n1202_));
  NO2        u1174(.A(men_men_n1202_), .B(men_men_n150_), .Y(men_men_n1203_));
  AOI220     u1175(.A0(men_men_n1203_), .A1(men_men_n271_), .B0(men_men_n851_), .B1(men_men_n1201_), .Y(men_men_n1204_));
  OAI210     u1176(.A0(men_men_n354_), .A1(men_men_n310_), .B0(men_men_n441_), .Y(men_men_n1205_));
  NA4        u1177(.A(men_men_n1205_), .B(men_men_n1204_), .C(men_men_n1200_), .D(men_men_n1199_), .Y(men_men_n1206_));
  AOI210     u1178(.A0(men_men_n1203_), .A1(men_men_n855_), .B0(men_men_n824_), .Y(men_men_n1207_));
  AOI220     u1179(.A0(men_men_n957_), .A1(men_men_n570_), .B0(men_men_n648_), .B1(men_men_n242_), .Y(men_men_n1208_));
  NO2        u1180(.A(men_men_n67_), .B(h), .Y(men_men_n1209_));
  NO3        u1181(.A(men_men_n1046_), .B(men_men_n1044_), .C(men_men_n725_), .Y(men_men_n1210_));
  NO2        u1182(.A(men_men_n1074_), .B(men_men_n134_), .Y(men_men_n1211_));
  AN2        u1183(.A(men_men_n1211_), .B(men_men_n1086_), .Y(men_men_n1212_));
  OAI210     u1184(.A0(men_men_n1212_), .A1(men_men_n1210_), .B0(men_men_n1209_), .Y(men_men_n1213_));
  NA4        u1185(.A(men_men_n1213_), .B(men_men_n1208_), .C(men_men_n1207_), .D(men_men_n870_), .Y(men_men_n1214_));
  NO4        u1186(.A(men_men_n1214_), .B(men_men_n1206_), .C(men_men_n1197_), .D(men_men_n1194_), .Y(men_men_n1215_));
  NA2        u1187(.A(men_men_n839_), .B(men_men_n757_), .Y(men_men_n1216_));
  NA4        u1188(.A(men_men_n1216_), .B(men_men_n1215_), .C(men_men_n1191_), .D(men_men_n1159_), .Y(men01));
  AN2        u1189(.A(men_men_n1027_), .B(men_men_n1025_), .Y(men_men_n1218_));
  NO3        u1190(.A(men_men_n805_), .B(men_men_n798_), .C(men_men_n469_), .Y(men_men_n1219_));
  NO2        u1191(.A(men_men_n587_), .B(men_men_n286_), .Y(men_men_n1220_));
  INV        u1192(.A(men_men_n1220_), .Y(men_men_n1221_));
  NA3        u1193(.A(men_men_n1221_), .B(men_men_n1219_), .C(men_men_n1218_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n583_), .B(men_men_n91_), .Y(men_men_n1223_));
  NA2        u1195(.A(men_men_n547_), .B(men_men_n268_), .Y(men_men_n1224_));
  NA2        u1196(.A(men_men_n964_), .B(men_men_n1224_), .Y(men_men_n1225_));
  NA4        u1197(.A(men_men_n1225_), .B(men_men_n1223_), .C(men_men_n915_), .D(men_men_n328_), .Y(men_men_n1226_));
  NA2        u1198(.A(men_men_n705_), .B(men_men_n98_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n1227_), .B(i), .Y(men_men_n1228_));
  OAI210     u1200(.A0(men_men_n784_), .A1(men_men_n600_), .B0(men_men_n1196_), .Y(men_men_n1229_));
  AOI210     u1201(.A0(men_men_n1228_), .A1(men_men_n633_), .B0(men_men_n1229_), .Y(men_men_n1230_));
  NA2        u1202(.A(men_men_n119_), .B(l), .Y(men_men_n1231_));
  OA220      u1203(.A0(men_men_n1231_), .A1(men_men_n580_), .B0(men_men_n661_), .B1(men_men_n368_), .Y(men_men_n1232_));
  NAi41      u1204(.An(men_men_n165_), .B(men_men_n1232_), .C(men_men_n1230_), .D(men_men_n901_), .Y(men_men_n1233_));
  NO2        u1205(.A(men_men_n785_), .B(men_men_n674_), .Y(men_men_n1234_));
  NA4        u1206(.A(men_men_n705_), .B(men_men_n98_), .C(men_men_n45_), .D(men_men_n215_), .Y(men_men_n1235_));
  NA2        u1207(.A(men_men_n1234_), .B(men_men_n140_), .Y(men_men_n1236_));
  NO4        u1208(.A(men_men_n1236_), .B(men_men_n1233_), .C(men_men_n1226_), .D(men_men_n1222_), .Y(men_men_n1237_));
  NA2        u1209(.A(men_men_n1168_), .B(men_men_n208_), .Y(men_men_n1238_));
  OAI210     u1210(.A0(men_men_n1238_), .A1(men_men_n299_), .B0(men_men_n522_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n530_), .B(men_men_n391_), .Y(men_men_n1240_));
  AOI210     u1212(.A0(men_men_n586_), .A1(men_men_n580_), .B0(l), .Y(men_men_n1241_));
  AOI210     u1213(.A0(men_men_n555_), .A1(men_men_n1240_), .B0(men_men_n1241_), .Y(men_men_n1242_));
  AOI210     u1214(.A0(men_men_n205_), .A1(men_men_n90_), .B0(men_men_n215_), .Y(men_men_n1243_));
  OAI210     u1215(.A0(men_men_n812_), .A1(men_men_n423_), .B0(men_men_n1243_), .Y(men_men_n1244_));
  AN3        u1216(.A(m), .B(l), .C(k), .Y(men_men_n1245_));
  OAI210     u1217(.A0(men_men_n356_), .A1(men_men_n34_), .B0(men_men_n1245_), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n204_), .B(men_men_n34_), .Y(men_men_n1247_));
  AO210      u1219(.A0(men_men_n1247_), .A1(men_men_n1246_), .B0(men_men_n327_), .Y(men_men_n1248_));
  NA4        u1220(.A(men_men_n1248_), .B(men_men_n1244_), .C(men_men_n1242_), .D(men_men_n1239_), .Y(men_men_n1249_));
  AOI210     u1221(.A0(men_men_n592_), .A1(men_men_n119_), .B0(men_men_n598_), .Y(men_men_n1250_));
  OAI210     u1222(.A0(men_men_n1231_), .A1(men_men_n589_), .B0(men_men_n1250_), .Y(men_men_n1251_));
  NA2        u1223(.A(men_men_n278_), .B(men_men_n197_), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n1252_), .B(men_men_n666_), .Y(men_men_n1253_));
  NO3        u1225(.A(men_men_n823_), .B(men_men_n205_), .C(men_men_n402_), .Y(men_men_n1254_));
  NO2        u1226(.A(men_men_n1254_), .B(men_men_n961_), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n1228_), .A1(men_men_n321_), .B0(men_men_n675_), .Y(men_men_n1256_));
  NA4        u1228(.A(men_men_n1256_), .B(men_men_n1255_), .C(men_men_n1253_), .D(men_men_n788_), .Y(men_men_n1257_));
  NO3        u1229(.A(men_men_n1257_), .B(men_men_n1251_), .C(men_men_n1249_), .Y(men_men_n1258_));
  NA3        u1230(.A(men_men_n601_), .B(men_men_n29_), .C(f), .Y(men_men_n1259_));
  NO2        u1231(.A(men_men_n1259_), .B(men_men_n205_), .Y(men_men_n1260_));
  AOI210     u1232(.A0(men_men_n495_), .A1(men_men_n58_), .B0(men_men_n1260_), .Y(men_men_n1261_));
  OR3        u1233(.A(men_men_n1227_), .B(men_men_n602_), .C(i), .Y(men_men_n1262_));
  NA3        u1234(.A(men_men_n739_), .B(men_men_n75_), .C(i), .Y(men_men_n1263_));
  AOI210     u1235(.A0(men_men_n1263_), .A1(men_men_n1235_), .B0(men_men_n983_), .Y(men_men_n1264_));
  NO2        u1236(.A(men_men_n208_), .B(men_men_n113_), .Y(men_men_n1265_));
  NO3        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .C(men_men_n1164_), .Y(men_men_n1266_));
  NA4        u1238(.A(men_men_n1266_), .B(men_men_n1262_), .C(men_men_n1261_), .D(men_men_n756_), .Y(men_men_n1267_));
  NA2        u1239(.A(men_men_n565_), .B(men_men_n563_), .Y(men_men_n1268_));
  NO3        u1240(.A(men_men_n80_), .B(men_men_n297_), .C(men_men_n45_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n546_), .Y(men_men_n1270_));
  NA3        u1242(.A(men_men_n1270_), .B(men_men_n1268_), .C(men_men_n670_), .Y(men_men_n1271_));
  OR2        u1243(.A(men_men_n1168_), .B(men_men_n1161_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n368_), .B(men_men_n72_), .Y(men_men_n1273_));
  AOI210     u1245(.A0(men_men_n730_), .A1(men_men_n613_), .B0(men_men_n1273_), .Y(men_men_n1274_));
  NA2        u1246(.A(men_men_n1269_), .B(men_men_n815_), .Y(men_men_n1275_));
  NA4        u1247(.A(men_men_n1275_), .B(men_men_n1274_), .C(men_men_n1272_), .D(men_men_n386_), .Y(men_men_n1276_));
  NO3        u1248(.A(men_men_n1276_), .B(men_men_n1271_), .C(men_men_n1267_), .Y(men_men_n1277_));
  AO220      u1249(.A0(i), .A1(men_men_n619_), .B0(men_men_n1521_), .B1(men_men_n703_), .Y(men_men_n1278_));
  NA2        u1250(.A(men_men_n450_), .B(men_men_n137_), .Y(men_men_n1279_));
  NO3        u1251(.A(men_men_n1084_), .B(men_men_n180_), .C(men_men_n88_), .Y(men_men_n1280_));
  AOI220     u1252(.A0(men_men_n1280_), .A1(men_men_n1279_), .B0(men_men_n1269_), .B1(men_men_n974_), .Y(men_men_n1281_));
  INV        u1253(.A(men_men_n1281_), .Y(men_men_n1282_));
  NO3        u1254(.A(men_men_n450_), .B(men_men_n178_), .C(men_men_n88_), .Y(men_men_n1283_));
  NO3        u1255(.A(men_men_n1283_), .B(men_men_n1282_), .C(men_men_n637_), .Y(men_men_n1284_));
  NA4        u1256(.A(men_men_n1284_), .B(men_men_n1277_), .C(men_men_n1258_), .D(men_men_n1237_), .Y(men06));
  NO2        u1257(.A(men_men_n403_), .B(men_men_n552_), .Y(men_men_n1286_));
  NO2        u1258(.A(men_men_n732_), .B(i), .Y(men_men_n1287_));
  OAI210     u1259(.A0(men_men_n1287_), .A1(men_men_n264_), .B0(men_men_n1286_), .Y(men_men_n1288_));
  NO3        u1260(.A(men_men_n596_), .B(men_men_n810_), .C(men_men_n599_), .Y(men_men_n1289_));
  OR2        u1261(.A(men_men_n1289_), .B(men_men_n890_), .Y(men_men_n1290_));
  NA2        u1262(.A(men_men_n1290_), .B(men_men_n1288_), .Y(men_men_n1291_));
  NO3        u1263(.A(men_men_n1291_), .B(men_men_n1271_), .C(men_men_n252_), .Y(men_men_n1292_));
  NO2        u1264(.A(men_men_n297_), .B(men_men_n45_), .Y(men_men_n1293_));
  NA2        u1265(.A(men_men_n1293_), .B(men_men_n975_), .Y(men_men_n1294_));
  AOI210     u1266(.A0(men_men_n1293_), .A1(men_men_n549_), .B0(men_men_n1278_), .Y(men_men_n1295_));
  AOI210     u1267(.A0(men_men_n1295_), .A1(men_men_n1294_), .B0(men_men_n333_), .Y(men_men_n1296_));
  OAI210     u1268(.A0(men_men_n90_), .A1(men_men_n40_), .B0(men_men_n673_), .Y(men_men_n1297_));
  NA2        u1269(.A(men_men_n1297_), .B(men_men_n641_), .Y(men_men_n1298_));
  NO2        u1270(.A(men_men_n606_), .B(men_men_n1106_), .Y(men_men_n1299_));
  OAI210     u1271(.A0(men_men_n450_), .A1(men_men_n246_), .B0(men_men_n909_), .Y(men_men_n1300_));
  NO3        u1272(.A(men_men_n1300_), .B(men_men_n1299_), .C(men_men_n139_), .Y(men_men_n1301_));
  OR2        u1273(.A(men_men_n597_), .B(men_men_n595_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n367_), .B(men_men_n138_), .Y(men_men_n1303_));
  AOI210     u1275(.A0(men_men_n1303_), .A1(men_men_n583_), .B0(men_men_n1302_), .Y(men_men_n1304_));
  NA3        u1276(.A(men_men_n1304_), .B(men_men_n1301_), .C(men_men_n1298_), .Y(men_men_n1305_));
  NO2        u1277(.A(men_men_n747_), .B(men_men_n366_), .Y(men_men_n1306_));
  NO3        u1278(.A(men_men_n675_), .B(men_men_n758_), .C(men_men_n633_), .Y(men_men_n1307_));
  NOi21      u1279(.An(men_men_n1306_), .B(men_men_n1307_), .Y(men_men_n1308_));
  AN2        u1280(.A(men_men_n957_), .B(men_men_n644_), .Y(men_men_n1309_));
  NO4        u1281(.A(men_men_n1309_), .B(men_men_n1308_), .C(men_men_n1305_), .D(men_men_n1296_), .Y(men_men_n1310_));
  NO2        u1282(.A(men_men_n804_), .B(men_men_n274_), .Y(men_men_n1311_));
  OAI220     u1283(.A0(men_men_n732_), .A1(men_men_n47_), .B0(men_men_n226_), .B1(men_men_n612_), .Y(men_men_n1312_));
  OAI210     u1284(.A0(men_men_n274_), .A1(c), .B0(men_men_n640_), .Y(men_men_n1313_));
  AOI220     u1285(.A0(men_men_n1313_), .A1(men_men_n1312_), .B0(men_men_n1311_), .B1(men_men_n264_), .Y(men_men_n1314_));
  NO3        u1286(.A(men_men_n241_), .B(men_men_n105_), .C(men_men_n279_), .Y(men_men_n1315_));
  OAI210     u1287(.A0(l), .A1(i), .B0(k), .Y(men_men_n1316_));
  NO3        u1288(.A(men_men_n1316_), .B(men_men_n594_), .C(j), .Y(men_men_n1317_));
  NOi21      u1289(.An(men_men_n1317_), .B(men_men_n72_), .Y(men_men_n1318_));
  NO3        u1290(.A(men_men_n1318_), .B(men_men_n1315_), .C(men_men_n1109_), .Y(men_men_n1319_));
  NA4        u1291(.A(men_men_n796_), .B(men_men_n795_), .C(men_men_n429_), .D(men_men_n882_), .Y(men_men_n1320_));
  NAi31      u1292(.An(men_men_n747_), .B(men_men_n1320_), .C(men_men_n204_), .Y(men_men_n1321_));
  NA4        u1293(.A(men_men_n1321_), .B(men_men_n1319_), .C(men_men_n1314_), .D(men_men_n1208_), .Y(men_men_n1322_));
  NOi31      u1294(.An(men_men_n1289_), .B(men_men_n454_), .C(men_men_n390_), .Y(men_men_n1323_));
  OR3        u1295(.A(men_men_n1323_), .B(men_men_n784_), .C(men_men_n533_), .Y(men_men_n1324_));
  OR3        u1296(.A(men_men_n370_), .B(men_men_n226_), .C(men_men_n612_), .Y(men_men_n1325_));
  AOI210     u1297(.A0(men_men_n565_), .A1(men_men_n441_), .B0(men_men_n372_), .Y(men_men_n1326_));
  NA2        u1298(.A(men_men_n1317_), .B(men_men_n792_), .Y(men_men_n1327_));
  NA4        u1299(.A(men_men_n1327_), .B(men_men_n1326_), .C(men_men_n1325_), .D(men_men_n1324_), .Y(men_men_n1328_));
  AOI220     u1300(.A0(men_men_n1306_), .A1(men_men_n757_), .B0(men_men_n1303_), .B1(men_men_n235_), .Y(men_men_n1329_));
  NO3        u1301(.A(men_men_n929_), .B(men_men_n880_), .C(men_men_n491_), .Y(men_men_n1330_));
  NA3        u1302(.A(men_men_n1330_), .B(men_men_n1329_), .C(men_men_n1275_), .Y(men_men_n1331_));
  NO3        u1303(.A(men_men_n450_), .B(j), .C(men_men_n435_), .Y(men_men_n1332_));
  NO4        u1304(.A(men_men_n1332_), .B(men_men_n1331_), .C(men_men_n1328_), .D(men_men_n1322_), .Y(men_men_n1333_));
  NA4        u1305(.A(men_men_n1333_), .B(men_men_n1310_), .C(men_men_n1292_), .D(men_men_n1284_), .Y(men07));
  NOi21      u1306(.An(j), .B(k), .Y(men_men_n1335_));
  NAi32      u1307(.An(m), .Bn(b), .C(n), .Y(men_men_n1336_));
  NO3        u1308(.A(men_men_n1336_), .B(g), .C(f), .Y(men_men_n1337_));
  OAI210     u1309(.A0(men_men_n316_), .A1(men_men_n472_), .B0(men_men_n1337_), .Y(men_men_n1338_));
  NAi21      u1310(.An(f), .B(c), .Y(men_men_n1339_));
  OR2        u1311(.A(e), .B(d), .Y(men_men_n1340_));
  NOi31      u1312(.An(n), .B(m), .C(b), .Y(men_men_n1341_));
  INV        u1313(.A(men_men_n1338_), .Y(men_men_n1342_));
  NOi41      u1314(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1343_));
  NA3        u1315(.A(men_men_n1343_), .B(men_men_n872_), .C(men_men_n405_), .Y(men_men_n1344_));
  INV        u1316(.A(men_men_n1344_), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n1086_), .B(men_men_n223_), .Y(men_men_n1346_));
  NO2        u1318(.A(men_men_n1346_), .B(men_men_n60_), .Y(men_men_n1347_));
  NO2        u1319(.A(k), .B(i), .Y(men_men_n1348_));
  NA2        u1320(.A(men_men_n88_), .B(men_men_n45_), .Y(men_men_n1349_));
  NO2        u1321(.A(men_men_n1051_), .B(men_men_n435_), .Y(men_men_n1350_));
  NA3        u1322(.A(men_men_n1350_), .B(men_men_n1349_), .C(men_men_n216_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n1063_), .B(men_men_n304_), .Y(men_men_n1352_));
  NA2        u1324(.A(men_men_n534_), .B(men_men_n81_), .Y(men_men_n1353_));
  NA2        u1325(.A(men_men_n1209_), .B(men_men_n287_), .Y(men_men_n1354_));
  NA3        u1326(.A(men_men_n1354_), .B(men_men_n1353_), .C(men_men_n1351_), .Y(men_men_n1355_));
  NO4        u1327(.A(men_men_n1355_), .B(men_men_n1347_), .C(men_men_n1345_), .D(men_men_n1342_), .Y(men_men_n1356_));
  NO3        u1328(.A(e), .B(d), .C(c), .Y(men_men_n1357_));
  OAI210     u1329(.A0(men_men_n134_), .A1(men_men_n216_), .B0(men_men_n603_), .Y(men_men_n1358_));
  NA2        u1330(.A(men_men_n1358_), .B(men_men_n1357_), .Y(men_men_n1359_));
  INV        u1331(.A(men_men_n1359_), .Y(men_men_n1360_));
  OR2        u1332(.A(h), .B(f), .Y(men_men_n1361_));
  NO3        u1333(.A(n), .B(m), .C(i), .Y(men_men_n1362_));
  OAI210     u1334(.A0(men_men_n1107_), .A1(men_men_n160_), .B0(men_men_n1362_), .Y(men_men_n1363_));
  NO2        u1335(.A(i), .B(g), .Y(men_men_n1364_));
  OR3        u1336(.A(men_men_n1364_), .B(men_men_n1336_), .C(men_men_n71_), .Y(men_men_n1365_));
  OAI220     u1337(.A0(men_men_n1365_), .A1(men_men_n472_), .B0(men_men_n1363_), .B1(men_men_n1361_), .Y(men_men_n1366_));
  NA3        u1338(.A(men_men_n694_), .B(men_men_n683_), .C(men_men_n114_), .Y(men_men_n1367_));
  NA3        u1339(.A(men_men_n1341_), .B(men_men_n1060_), .C(h), .Y(men_men_n1368_));
  AOI210     u1340(.A0(men_men_n1368_), .A1(men_men_n1367_), .B0(men_men_n45_), .Y(men_men_n1369_));
  NA2        u1341(.A(men_men_n1362_), .B(men_men_n639_), .Y(men_men_n1370_));
  NO3        u1342(.A(men_men_n435_), .B(d), .C(c), .Y(men_men_n1371_));
  NO3        u1343(.A(men_men_n1369_), .B(men_men_n1366_), .C(men_men_n1360_), .Y(men_men_n1372_));
  NO2        u1344(.A(men_men_n151_), .B(h), .Y(men_men_n1373_));
  NO2        u1345(.A(g), .B(c), .Y(men_men_n1374_));
  NA3        u1346(.A(men_men_n1374_), .B(men_men_n145_), .C(men_men_n190_), .Y(men_men_n1375_));
  NO2        u1347(.A(men_men_n1375_), .B(men_men_n1515_), .Y(men_men_n1376_));
  NA2        u1348(.A(men_men_n1376_), .B(men_men_n183_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n446_), .B(a), .Y(men_men_n1378_));
  NA3        u1350(.A(men_men_n1378_), .B(men_men_n1516_), .C(men_men_n115_), .Y(men_men_n1379_));
  NO2        u1351(.A(i), .B(h), .Y(men_men_n1380_));
  NA2        u1352(.A(men_men_n1380_), .B(men_men_n223_), .Y(men_men_n1381_));
  AOI210     u1353(.A0(men_men_n253_), .A1(men_men_n117_), .B0(men_men_n522_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n1382_), .B(men_men_n1381_), .Y(men_men_n1383_));
  NO2        u1355(.A(men_men_n754_), .B(men_men_n191_), .Y(men_men_n1384_));
  NOi31      u1356(.An(m), .B(n), .C(b), .Y(men_men_n1385_));
  NOi31      u1357(.An(f), .B(d), .C(c), .Y(men_men_n1386_));
  NA2        u1358(.A(men_men_n1386_), .B(men_men_n1385_), .Y(men_men_n1387_));
  INV        u1359(.A(men_men_n1387_), .Y(men_men_n1388_));
  NO3        u1360(.A(men_men_n1388_), .B(men_men_n1384_), .C(men_men_n1383_), .Y(men_men_n1389_));
  NO3        u1361(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1390_));
  AN3        u1362(.A(men_men_n1389_), .B(men_men_n1379_), .C(men_men_n1377_), .Y(men_men_n1391_));
  NA2        u1363(.A(men_men_n1341_), .B(men_men_n379_), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n1392_), .B(men_men_n1043_), .Y(men_men_n1393_));
  NO2        u1365(.A(men_men_n191_), .B(b), .Y(men_men_n1394_));
  NA2        u1366(.A(men_men_n1162_), .B(men_men_n1394_), .Y(men_men_n1395_));
  NO2        u1367(.A(i), .B(men_men_n215_), .Y(men_men_n1396_));
  NA4        u1368(.A(men_men_n1136_), .B(men_men_n1396_), .C(men_men_n106_), .D(m), .Y(men_men_n1397_));
  NAi31      u1369(.An(men_men_n1393_), .B(men_men_n1397_), .C(men_men_n1395_), .Y(men_men_n1398_));
  NO4        u1370(.A(men_men_n134_), .B(g), .C(f), .D(e), .Y(men_men_n1399_));
  NA3        u1371(.A(men_men_n1348_), .B(men_men_n288_), .C(h), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n196_), .B(men_men_n100_), .Y(men_men_n1401_));
  NA2        u1373(.A(men_men_n30_), .B(h), .Y(men_men_n1402_));
  NO2        u1374(.A(men_men_n1402_), .B(men_men_n1076_), .Y(men_men_n1403_));
  NOi41      u1375(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1404_));
  NA2        u1376(.A(men_men_n1404_), .B(men_men_n115_), .Y(men_men_n1405_));
  INV        u1377(.A(men_men_n1405_), .Y(men_men_n1406_));
  OR3        u1378(.A(men_men_n533_), .B(men_men_n532_), .C(men_men_n114_), .Y(men_men_n1407_));
  NA2        u1379(.A(men_men_n1105_), .B(men_men_n402_), .Y(men_men_n1408_));
  OAI220     u1380(.A0(men_men_n1408_), .A1(men_men_n428_), .B0(men_men_n1407_), .B1(men_men_n297_), .Y(men_men_n1409_));
  AO210      u1381(.A0(men_men_n1409_), .A1(men_men_n117_), .B0(men_men_n1406_), .Y(men_men_n1410_));
  NO3        u1382(.A(men_men_n1410_), .B(men_men_n1403_), .C(men_men_n1398_), .Y(men_men_n1411_));
  NA4        u1383(.A(men_men_n1411_), .B(men_men_n1391_), .C(men_men_n1372_), .D(men_men_n1356_), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1120_), .B(men_men_n112_), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n379_), .B(men_men_n56_), .Y(men_men_n1414_));
  NO2        u1386(.A(men_men_n1414_), .B(men_men_n1370_), .Y(men_men_n1415_));
  NA2        u1387(.A(men_men_n217_), .B(men_men_n183_), .Y(men_men_n1416_));
  AOI210     u1388(.A0(men_men_n1416_), .A1(men_men_n1181_), .B0(men_men_n1414_), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n1079_), .B(men_men_n1076_), .Y(men_men_n1418_));
  NO3        u1390(.A(men_men_n1418_), .B(men_men_n1417_), .C(men_men_n1415_), .Y(men_men_n1419_));
  NA3        u1391(.A(men_men_n1390_), .B(men_men_n1340_), .C(men_men_n1105_), .Y(men_men_n1420_));
  NO3        u1392(.A(men_men_n1076_), .B(men_men_n577_), .C(g), .Y(men_men_n1421_));
  INV        u1393(.A(men_men_n1421_), .Y(men_men_n1422_));
  AOI210     u1394(.A0(men_men_n1422_), .A1(men_men_n1401_), .B0(men_men_n1051_), .Y(men_men_n1423_));
  INV        u1395(.A(men_men_n49_), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n1424_), .B(men_men_n1170_), .Y(men_men_n1425_));
  INV        u1397(.A(men_men_n1425_), .Y(men_men_n1426_));
  OAI220     u1398(.A0(men_men_n667_), .A1(g), .B0(men_men_n226_), .B1(c), .Y(men_men_n1427_));
  AOI210     u1399(.A0(men_men_n1394_), .A1(men_men_n41_), .B0(men_men_n1427_), .Y(men_men_n1428_));
  NO2        u1400(.A(men_men_n134_), .B(l), .Y(men_men_n1429_));
  NO2        u1401(.A(men_men_n226_), .B(k), .Y(men_men_n1430_));
  OAI210     u1402(.A0(men_men_n1430_), .A1(men_men_n1380_), .B0(men_men_n1429_), .Y(men_men_n1431_));
  OAI220     u1403(.A0(men_men_n1431_), .A1(men_men_n31_), .B0(men_men_n1428_), .B1(men_men_n180_), .Y(men_men_n1432_));
  NO3        u1404(.A(men_men_n1407_), .B(men_men_n457_), .C(men_men_n350_), .Y(men_men_n1433_));
  NO4        u1405(.A(men_men_n1433_), .B(men_men_n1432_), .C(men_men_n1426_), .D(men_men_n1423_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n49_), .B(men_men_n577_), .Y(men_men_n1435_));
  NO3        u1407(.A(men_men_n1088_), .B(men_men_n1340_), .C(men_men_n49_), .Y(men_men_n1436_));
  NA2        u1408(.A(men_men_n1089_), .B(men_men_n1435_), .Y(men_men_n1437_));
  NO2        u1409(.A(men_men_n1076_), .B(h), .Y(men_men_n1438_));
  NA3        u1410(.A(men_men_n1438_), .B(d), .C(men_men_n1044_), .Y(men_men_n1439_));
  OAI220     u1411(.A0(men_men_n1439_), .A1(c), .B0(men_men_n1437_), .B1(j), .Y(men_men_n1440_));
  NA3        u1412(.A(men_men_n1413_), .B(men_men_n457_), .C(f), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n1335_), .B(men_men_n42_), .Y(men_men_n1442_));
  AOI210     u1414(.A0(men_men_n115_), .A1(men_men_n40_), .B0(men_men_n1442_), .Y(men_men_n1443_));
  NO2        u1415(.A(men_men_n1443_), .B(men_men_n1441_), .Y(men_men_n1444_));
  AOI210     u1416(.A0(men_men_n517_), .A1(h), .B0(men_men_n68_), .Y(men_men_n1445_));
  NA2        u1417(.A(men_men_n1445_), .B(men_men_n1378_), .Y(men_men_n1446_));
  NO2        u1418(.A(j), .B(men_men_n178_), .Y(men_men_n1447_));
  NOi21      u1419(.An(d), .B(f), .Y(men_men_n1448_));
  NO3        u1420(.A(men_men_n1386_), .B(men_men_n1448_), .C(men_men_n40_), .Y(men_men_n1449_));
  NA2        u1421(.A(men_men_n1449_), .B(men_men_n1447_), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1378_), .B(men_men_n1442_), .Y(men_men_n1451_));
  NO2        u1423(.A(men_men_n297_), .B(c), .Y(men_men_n1452_));
  NA2        u1424(.A(men_men_n1452_), .B(men_men_n534_), .Y(men_men_n1453_));
  NA4        u1425(.A(men_men_n1453_), .B(men_men_n1451_), .C(men_men_n1450_), .D(men_men_n1446_), .Y(men_men_n1454_));
  NO3        u1426(.A(men_men_n1454_), .B(men_men_n1444_), .C(men_men_n1440_), .Y(men_men_n1455_));
  NA4        u1427(.A(men_men_n1455_), .B(men_men_n1434_), .C(men_men_n1420_), .D(men_men_n1419_), .Y(men_men_n1456_));
  OAI220     u1428(.A0(men_men_n457_), .A1(men_men_n297_), .B0(men_men_n133_), .B1(men_men_n59_), .Y(men_men_n1457_));
  NA2        u1429(.A(men_men_n1457_), .B(men_men_n1352_), .Y(men_men_n1458_));
  OAI210     u1430(.A0(men_men_n1399_), .A1(men_men_n1341_), .B0(men_men_n887_), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n1459_), .B(men_men_n1458_), .Y(men_men_n1460_));
  NA2        u1432(.A(men_men_n1374_), .B(men_men_n1448_), .Y(men_men_n1461_));
  NO2        u1433(.A(men_men_n1461_), .B(m), .Y(men_men_n1462_));
  NA3        u1434(.A(men_men_n1086_), .B(men_men_n110_), .C(men_men_n223_), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n112_), .B(men_men_n1385_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n1464_), .B(men_men_n1463_), .Y(men_men_n1465_));
  NO3        u1437(.A(men_men_n1465_), .B(men_men_n1462_), .C(men_men_n1460_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n1339_), .B(e), .Y(men_men_n1467_));
  NA2        u1439(.A(men_men_n1467_), .B(men_men_n400_), .Y(men_men_n1468_));
  OR3        u1440(.A(men_men_n1430_), .B(men_men_n1209_), .C(men_men_n134_), .Y(men_men_n1469_));
  NO2        u1441(.A(men_men_n1469_), .B(men_men_n1468_), .Y(men_men_n1470_));
  NO3        u1442(.A(men_men_n1407_), .B(men_men_n350_), .C(a), .Y(men_men_n1471_));
  NO2        u1443(.A(men_men_n1471_), .B(men_men_n1470_), .Y(men_men_n1472_));
  NA2        u1444(.A(men_men_n532_), .B(g), .Y(men_men_n1473_));
  AOI210     u1445(.A0(men_men_n1473_), .A1(men_men_n1371_), .B0(men_men_n1436_), .Y(men_men_n1474_));
  NA2        u1446(.A(men_men_n1115_), .B(a), .Y(men_men_n1475_));
  OAI220     u1447(.A0(men_men_n1475_), .A1(men_men_n68_), .B0(men_men_n1474_), .B1(men_men_n215_), .Y(men_men_n1476_));
  NA4        u1448(.A(men_men_n1086_), .B(men_men_n1083_), .C(men_men_n223_), .D(men_men_n67_), .Y(men_men_n1477_));
  NO2        u1449(.A(m), .B(i), .Y(men_men_n1478_));
  NA2        u1450(.A(men_men_n1478_), .B(men_men_n1373_), .Y(men_men_n1479_));
  NA2        u1451(.A(men_men_n1479_), .B(men_men_n1477_), .Y(men_men_n1480_));
  NO2        u1452(.A(men_men_n1480_), .B(men_men_n1476_), .Y(men_men_n1481_));
  NA3        u1453(.A(men_men_n1481_), .B(men_men_n1472_), .C(men_men_n1466_), .Y(men_men_n1482_));
  NA3        u1454(.A(men_men_n963_), .B(men_men_n141_), .C(men_men_n46_), .Y(men_men_n1483_));
  AOI210     u1455(.A0(men_men_n152_), .A1(c), .B0(men_men_n1483_), .Y(men_men_n1484_));
  OAI210     u1456(.A0(men_men_n577_), .A1(g), .B0(men_men_n188_), .Y(men_men_n1485_));
  NA2        u1457(.A(men_men_n1485_), .B(men_men_n1438_), .Y(men_men_n1486_));
  NO2        u1458(.A(men_men_n71_), .B(c), .Y(men_men_n1487_));
  NO4        u1459(.A(men_men_n1361_), .B(men_men_n189_), .C(men_men_n443_), .D(men_men_n45_), .Y(men_men_n1488_));
  AOI210     u1460(.A0(men_men_n1447_), .A1(men_men_n1487_), .B0(men_men_n1488_), .Y(men_men_n1489_));
  NA2        u1461(.A(men_men_n1489_), .B(men_men_n1486_), .Y(men_men_n1490_));
  NO2        u1462(.A(men_men_n1490_), .B(men_men_n1484_), .Y(men_men_n1491_));
  NO4        u1463(.A(men_men_n226_), .B(men_men_n189_), .C(men_men_n253_), .D(k), .Y(men_men_n1492_));
  NO2        u1464(.A(men_men_n1483_), .B(men_men_n112_), .Y(men_men_n1493_));
  NO2        u1465(.A(men_men_n1493_), .B(men_men_n1492_), .Y(men_men_n1494_));
  AN2        u1466(.A(men_men_n1086_), .B(men_men_n1074_), .Y(men_men_n1495_));
  NA2        u1467(.A(men_men_n1057_), .B(men_men_n163_), .Y(men_men_n1496_));
  NOi31      u1468(.An(men_men_n30_), .B(men_men_n1496_), .C(n), .Y(men_men_n1497_));
  AOI210     u1469(.A0(men_men_n1495_), .A1(men_men_n1162_), .B0(men_men_n1497_), .Y(men_men_n1498_));
  NO2        u1470(.A(men_men_n1441_), .B(men_men_n68_), .Y(men_men_n1499_));
  NO2        u1471(.A(men_men_n1348_), .B(men_men_n119_), .Y(men_men_n1500_));
  NO2        u1472(.A(men_men_n1500_), .B(men_men_n1392_), .Y(men_men_n1501_));
  NO2        u1473(.A(men_men_n1501_), .B(men_men_n1499_), .Y(men_men_n1502_));
  NA4        u1474(.A(men_men_n1502_), .B(men_men_n1498_), .C(men_men_n1494_), .D(men_men_n1491_), .Y(men_men_n1503_));
  OR4        u1475(.A(men_men_n1503_), .B(men_men_n1482_), .C(men_men_n1456_), .D(men_men_n1412_), .Y(men04));
  NOi31      u1476(.An(men_men_n1399_), .B(men_men_n1400_), .C(men_men_n1046_), .Y(men_men_n1505_));
  NO4        u1477(.A(men_men_n269_), .B(men_men_n1037_), .C(men_men_n473_), .D(j), .Y(men_men_n1506_));
  OR3        u1478(.A(men_men_n1506_), .B(men_men_n1505_), .C(men_men_n1062_), .Y(men_men_n1507_));
  NO3        u1479(.A(men_men_n1349_), .B(men_men_n92_), .C(k), .Y(men_men_n1508_));
  AOI210     u1480(.A0(men_men_n1508_), .A1(men_men_n1056_), .B0(men_men_n1183_), .Y(men_men_n1509_));
  NA2        u1481(.A(men_men_n1509_), .B(men_men_n1213_), .Y(men_men_n1510_));
  NO4        u1482(.A(men_men_n1510_), .B(men_men_n1507_), .C(men_men_n1067_), .D(men_men_n1050_), .Y(men_men_n1511_));
  NA4        u1483(.A(men_men_n1511_), .B(men_men_n1117_), .C(men_men_n1103_), .D(men_men_n1090_), .Y(men05));
  INV        u1484(.A(l), .Y(men_men_n1515_));
  INV        u1485(.A(i), .Y(men_men_n1516_));
  INV        u1486(.A(men_men_n450_), .Y(men_men_n1517_));
  INV        u1487(.A(men_men_n1061_), .Y(men_men_n1518_));
  INV        u1488(.A(n), .Y(men_men_n1519_));
  INV        u1489(.A(i), .Y(men_men_n1520_));
  INV        u1490(.A(g), .Y(men_men_n1521_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule