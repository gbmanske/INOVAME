//  Package: package
//
package pkg;
    //  Group: Typedefs
    

    //  Group: Parameters
    `include "my_txn.sv"

    
endpackage: pkg
