//Benchmark atmr_intb_466_0.0625

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n328_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n350_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n417_, mai_mai_n418_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n355_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO2        o027(.A(ori_ori_n49_), .B(x11), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  AOI210     o039(.A0(x11), .A1(ori_ori_n48_), .B0(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o040(.A(ori_ori_n59_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n64_), .B(ori_ori_n24_), .Y(ori_ori_n65_));
  OAI220     o043(.A0(ori_ori_n65_), .A1(ori_ori_n63_), .B0(ori_ori_n62_), .B1(ori_ori_n60_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n30_), .B(x11), .Y(ori_ori_n67_));
  AOI220     o045(.A0(ori_ori_n67_), .A1(ori_ori_n59_), .B0(ori_ori_n66_), .B1(ori_ori_n31_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n69_));
  NA2        o047(.A(x09), .B(x05), .Y(ori_ori_n70_));
  NA2        o048(.A(x10), .B(x06), .Y(ori_ori_n71_));
  NA2        o049(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n72_), .A1(x07), .B0(x03), .Y(ori_ori_n74_));
  NOi31      o052(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n75_));
  INV        o053(.A(x07), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n24_), .Y(ori_ori_n77_));
  NO2        o055(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n36_), .Y(ori_ori_n79_));
  OAI210     o057(.A0(ori_ori_n78_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n80_));
  AOI210     o058(.A0(ori_ori_n79_), .A1(ori_ori_n48_), .B0(ori_ori_n80_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n82_));
  NO2        o060(.A(x08), .B(x01), .Y(ori_ori_n83_));
  OAI210     o061(.A0(ori_ori_n83_), .A1(ori_ori_n82_), .B0(ori_ori_n35_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n81_), .C(ori_ori_n77_), .Y(ori_ori_n85_));
  AN2        o063(.A(ori_ori_n85_), .B(ori_ori_n74_), .Y(ori_ori_n86_));
  INV        o064(.A(ori_ori_n84_), .Y(ori_ori_n87_));
  NA2        o065(.A(x11), .B(x00), .Y(ori_ori_n88_));
  NO2        o066(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n89_));
  NOi21      o067(.An(ori_ori_n88_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  NOi21      o068(.An(x01), .B(x10), .Y(ori_ori_n91_));
  NO2        o069(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n92_));
  NO3        o070(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(x06), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n93_), .B(ori_ori_n27_), .Y(ori_ori_n94_));
  OAI210     o072(.A0(ori_ori_n377_), .A1(x07), .B0(ori_ori_n94_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n86_), .C(ori_ori_n69_), .Y(ori01));
  INV        o074(.A(x12), .Y(ori_ori_n97_));
  INV        o075(.A(x13), .Y(ori_ori_n98_));
  NA2        o076(.A(x08), .B(x04), .Y(ori_ori_n99_));
  NO2        o077(.A(x10), .B(x01), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NA2        o080(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n104_));
  INV        o082(.A(x13), .Y(ori_ori_n105_));
  NA2        o083(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n106_));
  NA2        o084(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n107_), .B(x05), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n110_));
  NA2        o088(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n111_), .B(ori_ori_n110_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n114_));
  NA3        o092(.A(ori_ori_n114_), .B(ori_ori_n113_), .C(x13), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n116_));
  NOi31      o094(.An(ori_ori_n115_), .B(ori_ori_n116_), .C(ori_ori_n112_), .Y(ori_ori_n117_));
  NO3        o095(.A(ori_ori_n117_), .B(x06), .C(x03), .Y(ori_ori_n118_));
  INV        o096(.A(ori_ori_n118_), .Y(ori_ori_n119_));
  NA2        o097(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n120_));
  OAI210     o098(.A0(ori_ori_n83_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n123_));
  NO2        o101(.A(x09), .B(x05), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(ori_ori_n47_), .Y(ori_ori_n125_));
  AOI210     o103(.A0(ori_ori_n125_), .A1(ori_ori_n102_), .B0(ori_ori_n49_), .Y(ori_ori_n126_));
  NA2        o104(.A(x09), .B(x00), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n104_), .B(ori_ori_n127_), .Y(ori_ori_n128_));
  INV        o106(.A(ori_ori_n126_), .Y(ori_ori_n129_));
  NO2        o107(.A(x03), .B(x02), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n84_), .B(ori_ori_n98_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n131_), .B(ori_ori_n130_), .Y(ori_ori_n132_));
  OA210      o110(.A0(ori_ori_n129_), .A1(x11), .B0(ori_ori_n132_), .Y(ori_ori_n133_));
  OAI210     o111(.A0(ori_ori_n119_), .A1(ori_ori_n23_), .B0(ori_ori_n133_), .Y(ori_ori_n134_));
  NAi21      o112(.An(x06), .B(x10), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n98_), .B(x01), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n137_), .B(x08), .Y(ori_ori_n138_));
  OAI210     o116(.A0(x05), .A1(ori_ori_n138_), .B0(ori_ori_n51_), .Y(ori_ori_n139_));
  AOI210     o117(.A0(ori_ori_n139_), .A1(ori_ori_n136_), .B0(ori_ori_n48_), .Y(ori_ori_n140_));
  AOI210     o118(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n140_), .B(ori_ori_n141_), .Y(ori_ori_n142_));
  NA2        o120(.A(x04), .B(x02), .Y(ori_ori_n143_));
  INV        o121(.A(x05), .Y(ori_ori_n144_));
  NO2        o122(.A(x09), .B(x01), .Y(ori_ori_n145_));
  NO3        o123(.A(ori_ori_n145_), .B(ori_ori_n100_), .C(ori_ori_n31_), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n146_), .B(x00), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n104_), .B(x08), .Y(ori_ori_n148_));
  NAi21      o126(.An(ori_ori_n143_), .B(ori_ori_n376_), .Y(ori_ori_n149_));
  INV        o127(.A(ori_ori_n25_), .Y(ori_ori_n150_));
  NAi21      o128(.An(x13), .B(x00), .Y(ori_ori_n151_));
  AOI220     o129(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(ori_ori_n152_));
  AN2        o130(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n153_));
  NO2        o131(.A(ori_ori_n92_), .B(x06), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n151_), .B(ori_ori_n36_), .Y(ori_ori_n155_));
  INV        o133(.A(ori_ori_n155_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n154_), .B(ori_ori_n153_), .Y(ori_ori_n157_));
  NA2        o135(.A(ori_ori_n157_), .B(ori_ori_n150_), .Y(ori_ori_n158_));
  NOi21      o136(.An(x09), .B(x00), .Y(ori_ori_n159_));
  NO3        o137(.A(ori_ori_n82_), .B(ori_ori_n159_), .C(ori_ori_n47_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n111_), .Y(ori_ori_n161_));
  NA2        o139(.A(x06), .B(x05), .Y(ori_ori_n162_));
  OAI210     o140(.A0(ori_ori_n162_), .A1(ori_ori_n35_), .B0(ori_ori_n97_), .Y(ori_ori_n163_));
  AOI210     o141(.A0(x08), .A1(ori_ori_n58_), .B0(ori_ori_n163_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n164_), .B(ori_ori_n161_), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n98_), .B(x12), .Y(ori_ori_n166_));
  AOI210     o144(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n91_), .B(ori_ori_n51_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n169_));
  NA2        o147(.A(ori_ori_n169_), .B(x02), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n167_), .B(ori_ori_n165_), .Y(ori_ori_n171_));
  NA4        o149(.A(ori_ori_n171_), .B(ori_ori_n158_), .C(ori_ori_n149_), .D(ori_ori_n142_), .Y(ori_ori_n172_));
  AOI210     o150(.A0(ori_ori_n134_), .A1(ori_ori_n97_), .B0(ori_ori_n172_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n174_), .B(ori_ori_n121_), .Y(ori_ori_n175_));
  AOI210     o153(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n110_), .B(x06), .Y(ori_ori_n177_));
  AOI210     o155(.A0(ori_ori_n176_), .A1(ori_ori_n175_), .B0(ori_ori_n177_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n178_), .B(x12), .Y(ori_ori_n179_));
  INV        o157(.A(ori_ori_n75_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n91_), .B(x06), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n182_));
  NO3        o160(.A(ori_ori_n182_), .B(ori_ori_n181_), .C(ori_ori_n41_), .Y(ori_ori_n183_));
  INV        o161(.A(ori_ori_n123_), .Y(ori_ori_n184_));
  OAI210     o162(.A0(ori_ori_n184_), .A1(ori_ori_n183_), .B0(x02), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n185_), .A1(ori_ori_n57_), .B0(ori_ori_n23_), .Y(ori_ori_n186_));
  OAI210     o164(.A0(ori_ori_n179_), .A1(ori_ori_n57_), .B0(ori_ori_n186_), .Y(ori_ori_n187_));
  INV        o165(.A(ori_ori_n123_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n189_));
  OAI210     o167(.A0(ori_ori_n78_), .A1(ori_ori_n36_), .B0(ori_ori_n106_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n98_), .B(x03), .Y(ori_ori_n191_));
  AOI220     o169(.A0(ori_ori_n191_), .A1(ori_ori_n190_), .B0(ori_ori_n75_), .B1(ori_ori_n189_), .Y(ori_ori_n192_));
  NA2        o170(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n193_));
  INV        o171(.A(ori_ori_n135_), .Y(ori_ori_n194_));
  NOi21      o172(.An(x13), .B(x04), .Y(ori_ori_n195_));
  NO3        o173(.A(ori_ori_n195_), .B(ori_ori_n75_), .C(ori_ori_n159_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n196_), .B(x05), .Y(ori_ori_n197_));
  AOI220     o175(.A0(ori_ori_n197_), .A1(ori_ori_n193_), .B0(ori_ori_n194_), .B1(ori_ori_n57_), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n192_), .B(ori_ori_n198_), .Y(ori_ori_n199_));
  INV        o177(.A(ori_ori_n89_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n200_), .B(x12), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n202_));
  AOI210     o180(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n203_));
  NO2        o181(.A(x06), .B(x00), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n204_), .B(ori_ori_n203_), .C(ori_ori_n41_), .Y(ori_ori_n205_));
  OAI210     o183(.A0(ori_ori_n99_), .A1(ori_ori_n127_), .B0(ori_ori_n71_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(ori_ori_n205_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n208_));
  NA2        o186(.A(ori_ori_n208_), .B(x03), .Y(ori_ori_n209_));
  OR2        o187(.A(ori_ori_n209_), .B(ori_ori_n207_), .Y(ori_ori_n210_));
  NA2        o188(.A(x13), .B(ori_ori_n97_), .Y(ori_ori_n211_));
  NA3        o189(.A(ori_ori_n211_), .B(ori_ori_n163_), .C(ori_ori_n90_), .Y(ori_ori_n212_));
  OAI210     o190(.A0(ori_ori_n210_), .A1(ori_ori_n202_), .B0(ori_ori_n212_), .Y(ori_ori_n213_));
  AOI210     o191(.A0(ori_ori_n201_), .A1(ori_ori_n199_), .B0(ori_ori_n213_), .Y(ori_ori_n214_));
  AOI210     o192(.A0(ori_ori_n214_), .A1(ori_ori_n187_), .B0(x07), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n70_), .B(ori_ori_n29_), .Y(ori_ori_n216_));
  NOi31      o194(.An(ori_ori_n120_), .B(ori_ori_n195_), .C(ori_ori_n159_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n217_), .B(ori_ori_n216_), .Y(ori_ori_n218_));
  NO2        o196(.A(x08), .B(x05), .Y(ori_ori_n219_));
  NO2        o197(.A(x12), .B(x02), .Y(ori_ori_n220_));
  INV        o198(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n221_), .B(ori_ori_n200_), .Y(ori_ori_n222_));
  OA210      o200(.A0(ori_ori_n75_), .A1(ori_ori_n218_), .B0(ori_ori_n222_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n224_), .B(x01), .Y(ori_ori_n225_));
  NOi21      o203(.An(ori_ori_n83_), .B(ori_ori_n106_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(ori_ori_n225_), .Y(ori_ori_n227_));
  AOI210     o205(.A0(ori_ori_n227_), .A1(ori_ori_n115_), .B0(ori_ori_n29_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n98_), .B(x04), .Y(ori_ori_n229_));
  NO2        o207(.A(x02), .B(ori_ori_n105_), .Y(ori_ori_n230_));
  NO3        o208(.A(ori_ori_n88_), .B(x12), .C(x03), .Y(ori_ori_n231_));
  OAI210     o209(.A0(ori_ori_n230_), .A1(ori_ori_n228_), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  AOI210     o210(.A0(ori_ori_n168_), .A1(ori_ori_n162_), .B0(ori_ori_n99_), .Y(ori_ori_n233_));
  NOi21      o211(.An(ori_ori_n216_), .B(ori_ori_n181_), .Y(ori_ori_n234_));
  NO2        o212(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n235_));
  OAI210     o213(.A0(ori_ori_n234_), .A1(ori_ori_n233_), .B0(ori_ori_n235_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n237_));
  NO3        o215(.A(ori_ori_n237_), .B(ori_ori_n182_), .C(ori_ori_n154_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n202_), .B(ori_ori_n28_), .Y(ori_ori_n239_));
  OAI210     o217(.A0(ori_ori_n238_), .A1(ori_ori_n188_), .B0(ori_ori_n239_), .Y(ori_ori_n240_));
  NA3        o218(.A(ori_ori_n240_), .B(ori_ori_n236_), .C(ori_ori_n232_), .Y(ori_ori_n241_));
  NO3        o219(.A(ori_ori_n241_), .B(ori_ori_n223_), .C(ori_ori_n215_), .Y(ori_ori_n242_));
  OAI210     o220(.A0(ori_ori_n173_), .A1(ori_ori_n61_), .B0(ori_ori_n242_), .Y(ori02));
  NOi21      o221(.An(ori_ori_n196_), .B(ori_ori_n145_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n98_), .B(ori_ori_n35_), .Y(ori_ori_n245_));
  NA3        o223(.A(ori_ori_n245_), .B(x08), .C(ori_ori_n56_), .Y(ori_ori_n246_));
  OAI210     o224(.A0(ori_ori_n244_), .A1(ori_ori_n32_), .B0(ori_ori_n246_), .Y(ori_ori_n247_));
  NA2        o225(.A(ori_ori_n247_), .B(ori_ori_n144_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n131_), .B(ori_ori_n130_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n249_), .A1(ori_ori_n248_), .B0(ori_ori_n48_), .Y(ori_ori_n250_));
  NO2        o228(.A(x05), .B(x02), .Y(ori_ori_n251_));
  OAI210     o229(.A0(ori_ori_n175_), .A1(ori_ori_n159_), .B0(ori_ori_n251_), .Y(ori_ori_n252_));
  AOI220     o230(.A0(ori_ori_n219_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n253_));
  NOi21      o231(.An(ori_ori_n245_), .B(ori_ori_n253_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n195_), .A1(ori_ori_n78_), .B0(ori_ori_n254_), .Y(ori_ori_n255_));
  AOI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n252_), .B0(ori_ori_n123_), .Y(ori_ori_n256_));
  NAi21      o234(.An(ori_ori_n197_), .B(ori_ori_n192_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n208_), .B(ori_ori_n47_), .Y(ori_ori_n258_));
  NA2        o236(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  AN2        o237(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n260_));
  OAI210     o238(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n261_));
  NA2        o239(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n262_));
  BUFFER     o240(.A(ori_ori_n125_), .Y(ori_ori_n263_));
  AOI210     o241(.A0(ori_ori_n263_), .A1(ori_ori_n121_), .B0(ori_ori_n261_), .Y(ori_ori_n264_));
  OAI210     o242(.A0(ori_ori_n264_), .A1(ori_ori_n260_), .B0(ori_ori_n92_), .Y(ori_ori_n265_));
  NA3        o243(.A(ori_ori_n92_), .B(ori_ori_n83_), .C(ori_ori_n189_), .Y(ori_ori_n266_));
  NA3        o244(.A(ori_ori_n91_), .B(ori_ori_n82_), .C(ori_ori_n42_), .Y(ori_ori_n267_));
  AOI210     o245(.A0(ori_ori_n267_), .A1(ori_ori_n266_), .B0(x04), .Y(ori_ori_n268_));
  INV        o246(.A(ori_ori_n130_), .Y(ori_ori_n269_));
  NO2        o247(.A(ori_ori_n269_), .B(ori_ori_n112_), .Y(ori_ori_n270_));
  AOI210     o248(.A0(ori_ori_n270_), .A1(x13), .B0(ori_ori_n268_), .Y(ori_ori_n271_));
  NA3        o249(.A(ori_ori_n271_), .B(ori_ori_n265_), .C(ori_ori_n259_), .Y(ori_ori_n272_));
  NO3        o250(.A(ori_ori_n272_), .B(ori_ori_n256_), .C(ori_ori_n250_), .Y(ori_ori_n273_));
  NA2        o251(.A(ori_ori_n122_), .B(x03), .Y(ori_ori_n274_));
  INV        o252(.A(ori_ori_n151_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n35_), .B(ori_ori_n36_), .Y(ori_ori_n276_));
  AOI220     o254(.A0(ori_ori_n276_), .A1(ori_ori_n275_), .B0(ori_ori_n169_), .B1(x08), .Y(ori_ori_n277_));
  OAI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n237_), .B0(ori_ori_n274_), .Y(ori_ori_n278_));
  NA2        o256(.A(ori_ori_n278_), .B(ori_ori_n100_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n143_), .B(ori_ori_n137_), .Y(ori_ori_n280_));
  AN2        o258(.A(ori_ori_n280_), .B(ori_ori_n148_), .Y(ori_ori_n281_));
  INV        o259(.A(ori_ori_n56_), .Y(ori_ori_n282_));
  OAI220     o260(.A0(ori_ori_n229_), .A1(ori_ori_n282_), .B0(ori_ori_n113_), .B1(ori_ori_n28_), .Y(ori_ori_n283_));
  OAI210     o261(.A0(ori_ori_n283_), .A1(ori_ori_n281_), .B0(ori_ori_n101_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n229_), .B(ori_ori_n97_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n97_), .B(ori_ori_n41_), .Y(ori_ori_n286_));
  NA3        o264(.A(ori_ori_n286_), .B(ori_ori_n285_), .C(ori_ori_n112_), .Y(ori_ori_n287_));
  NA4        o265(.A(ori_ori_n287_), .B(ori_ori_n284_), .C(ori_ori_n279_), .D(ori_ori_n48_), .Y(ori_ori_n288_));
  INV        o266(.A(ori_ori_n169_), .Y(ori_ori_n289_));
  NO2        o267(.A(ori_ori_n378_), .B(ori_ori_n31_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n290_), .B(x02), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n166_), .B(x04), .Y(ori_ori_n292_));
  NO2        o270(.A(ori_ori_n152_), .B(ori_ori_n31_), .Y(ori_ori_n293_));
  NA2        o271(.A(ori_ori_n293_), .B(ori_ori_n92_), .Y(ori_ori_n294_));
  NO3        o272(.A(ori_ori_n166_), .B(ori_ori_n136_), .C(ori_ori_n52_), .Y(ori_ori_n295_));
  OAI210     o273(.A0(x12), .A1(ori_ori_n160_), .B0(ori_ori_n295_), .Y(ori_ori_n296_));
  NA4        o274(.A(ori_ori_n296_), .B(ori_ori_n294_), .C(ori_ori_n291_), .D(x06), .Y(ori_ori_n297_));
  NA2        o275(.A(x09), .B(x03), .Y(ori_ori_n298_));
  OAI220     o276(.A0(ori_ori_n298_), .A1(ori_ori_n111_), .B0(ori_ori_n174_), .B1(ori_ori_n64_), .Y(ori_ori_n299_));
  NO3        o277(.A(ori_ori_n237_), .B(ori_ori_n110_), .C(x08), .Y(ori_ori_n300_));
  AOI210     o278(.A0(x01), .A1(ori_ori_n188_), .B0(ori_ori_n300_), .Y(ori_ori_n301_));
  NO2        o279(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n302_));
  NO3        o280(.A(ori_ori_n104_), .B(ori_ori_n111_), .C(ori_ori_n38_), .Y(ori_ori_n303_));
  AOI210     o281(.A0(ori_ori_n295_), .A1(ori_ori_n302_), .B0(ori_ori_n303_), .Y(ori_ori_n304_));
  OAI210     o282(.A0(ori_ori_n301_), .A1(ori_ori_n28_), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  AO220      o283(.A0(ori_ori_n305_), .A1(x04), .B0(ori_ori_n299_), .B1(x05), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n297_), .A1(ori_ori_n288_), .B0(ori_ori_n306_), .Y(ori_ori_n307_));
  OAI210     o285(.A0(ori_ori_n273_), .A1(x12), .B0(ori_ori_n307_), .Y(ori03));
  OR2        o286(.A(ori_ori_n42_), .B(ori_ori_n189_), .Y(ori_ori_n309_));
  AOI210     o287(.A0(ori_ori_n131_), .A1(ori_ori_n97_), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n166_), .B(ori_ori_n130_), .Y(ori_ori_n311_));
  NA2        o289(.A(ori_ori_n311_), .B(ori_ori_n170_), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n310_), .B0(x05), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n309_), .B(x05), .Y(ori_ori_n314_));
  AOI210     o292(.A0(ori_ori_n121_), .A1(ori_ori_n180_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  AOI210     o293(.A0(ori_ori_n191_), .A1(ori_ori_n79_), .B0(ori_ori_n108_), .Y(ori_ori_n316_));
  OAI220     o294(.A0(ori_ori_n316_), .A1(ori_ori_n59_), .B0(ori_ori_n262_), .B1(ori_ori_n253_), .Y(ori_ori_n317_));
  OAI210     o295(.A0(ori_ori_n317_), .A1(ori_ori_n315_), .B0(ori_ori_n97_), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n125_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n145_), .B(ori_ori_n116_), .Y(ori_ori_n320_));
  OAI220     o298(.A0(ori_ori_n320_), .A1(ori_ori_n37_), .B0(ori_ori_n128_), .B1(x13), .Y(ori_ori_n321_));
  OAI210     o299(.A0(ori_ori_n321_), .A1(ori_ori_n319_), .B0(x04), .Y(ori_ori_n322_));
  NO3        o300(.A(ori_ori_n286_), .B(ori_ori_n84_), .C(ori_ori_n59_), .Y(ori_ori_n323_));
  AOI210     o301(.A0(ori_ori_n156_), .A1(ori_ori_n97_), .B0(ori_ori_n125_), .Y(ori_ori_n324_));
  OA210      o302(.A0(ori_ori_n138_), .A1(x12), .B0(ori_ori_n116_), .Y(ori_ori_n325_));
  NO3        o303(.A(ori_ori_n325_), .B(ori_ori_n324_), .C(ori_ori_n323_), .Y(ori_ori_n326_));
  NA4        o304(.A(ori_ori_n326_), .B(ori_ori_n322_), .C(ori_ori_n318_), .D(ori_ori_n313_), .Y(ori04));
  NO2        o305(.A(ori_ori_n87_), .B(ori_ori_n39_), .Y(ori_ori_n328_));
  XO2        o306(.A(ori_ori_n328_), .B(ori_ori_n211_), .Y(ori05));
  AOI210     o307(.A0(ori_ori_n70_), .A1(ori_ori_n52_), .B0(ori_ori_n177_), .Y(ori_ori_n330_));
  AOI210     o308(.A0(ori_ori_n330_), .A1(ori_ori_n261_), .B0(ori_ori_n25_), .Y(ori_ori_n331_));
  NA3        o309(.A(ori_ori_n123_), .B(ori_ori_n113_), .C(ori_ori_n31_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n194_), .B(ori_ori_n57_), .Y(ori_ori_n333_));
  AOI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n332_), .B0(ori_ori_n24_), .Y(ori_ori_n334_));
  OAI210     o312(.A0(ori_ori_n334_), .A1(ori_ori_n331_), .B0(ori_ori_n97_), .Y(ori_ori_n335_));
  OAI210     o313(.A0(ori_ori_n26_), .A1(ori_ori_n97_), .B0(x07), .Y(ori_ori_n336_));
  INV        o314(.A(ori_ori_n336_), .Y(ori_ori_n337_));
  NO3        o315(.A(x02), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n338_));
  OR2        o316(.A(x03), .B(ori_ori_n202_), .Y(ori_ori_n339_));
  NA2        o317(.A(ori_ori_n204_), .B(ori_ori_n200_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n340_), .B(ori_ori_n339_), .Y(ori_ori_n341_));
  OAI210     o319(.A0(ori_ori_n341_), .A1(ori_ori_n338_), .B0(ori_ori_n97_), .Y(ori_ori_n342_));
  NA2        o320(.A(ori_ori_n33_), .B(ori_ori_n97_), .Y(ori_ori_n343_));
  AOI210     o321(.A0(ori_ori_n343_), .A1(ori_ori_n89_), .B0(x07), .Y(ori_ori_n344_));
  AOI220     o322(.A0(ori_ori_n344_), .A1(ori_ori_n342_), .B0(ori_ori_n337_), .B1(ori_ori_n335_), .Y(ori_ori_n345_));
  AOI210     o323(.A0(ori_ori_n292_), .A1(ori_ori_n103_), .B0(ori_ori_n220_), .Y(ori_ori_n346_));
  NOi21      o324(.An(ori_ori_n274_), .B(ori_ori_n116_), .Y(ori_ori_n347_));
  NO2        o325(.A(ori_ori_n347_), .B(ori_ori_n221_), .Y(ori_ori_n348_));
  OAI210     o326(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n349_));
  AOI210     o327(.A0(ori_ori_n211_), .A1(ori_ori_n47_), .B0(ori_ori_n349_), .Y(ori_ori_n350_));
  NO4        o328(.A(ori_ori_n350_), .B(ori_ori_n348_), .C(ori_ori_n346_), .D(x08), .Y(ori_ori_n351_));
  NO2        o329(.A(ori_ori_n113_), .B(ori_ori_n28_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n225_), .Y(ori_ori_n353_));
  OR3        o331(.A(ori_ori_n353_), .B(x12), .C(x03), .Y(ori_ori_n354_));
  NA3        o332(.A(ori_ori_n289_), .B(ori_ori_n109_), .C(x12), .Y(ori_ori_n355_));
  AO210      o333(.A0(ori_ori_n289_), .A1(ori_ori_n109_), .B0(ori_ori_n211_), .Y(ori_ori_n356_));
  NA4        o334(.A(ori_ori_n356_), .B(ori_ori_n355_), .C(ori_ori_n354_), .D(x08), .Y(ori_ori_n357_));
  INV        o335(.A(ori_ori_n357_), .Y(ori_ori_n358_));
  NO2        o336(.A(ori_ori_n351_), .B(ori_ori_n358_), .Y(ori_ori_n359_));
  NO2        o337(.A(ori_ori_n124_), .B(ori_ori_n43_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n360_), .B(ori_ori_n155_), .Y(ori_ori_n361_));
  NA3        o339(.A(ori_ori_n353_), .B(ori_ori_n347_), .C(ori_ori_n285_), .Y(ori_ori_n362_));
  INV        o340(.A(x14), .Y(ori_ori_n363_));
  NO3        o341(.A(ori_ori_n137_), .B(ori_ori_n73_), .C(ori_ori_n57_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NA3        o343(.A(ori_ori_n365_), .B(ori_ori_n362_), .C(ori_ori_n361_), .Y(ori_ori_n366_));
  NA2        o344(.A(ori_ori_n343_), .B(ori_ori_n61_), .Y(ori_ori_n367_));
  NOi21      o345(.An(ori_ori_n229_), .B(ori_ori_n128_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n235_), .B(ori_ori_n194_), .Y(ori_ori_n369_));
  OAI210     o347(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n369_), .Y(ori_ori_n370_));
  OAI210     o348(.A0(ori_ori_n370_), .A1(ori_ori_n368_), .B0(ori_ori_n97_), .Y(ori_ori_n371_));
  OAI210     o349(.A0(ori_ori_n367_), .A1(ori_ori_n88_), .B0(ori_ori_n371_), .Y(ori_ori_n372_));
  NO4        o350(.A(ori_ori_n372_), .B(ori_ori_n366_), .C(ori_ori_n359_), .D(ori_ori_n345_), .Y(ori06));
  INV        o351(.A(ori_ori_n147_), .Y(ori_ori_n376_));
  INV        o352(.A(ori_ori_n90_), .Y(ori_ori_n377_));
  INV        o353(.A(x05), .Y(ori_ori_n378_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n59_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n63_), .B(mai_mai_n24_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n66_));
  OAI210     m044(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  AOI220     m045(.A0(mai_mai_n67_), .A1(mai_mai_n59_), .B0(mai_mai_n65_), .B1(mai_mai_n31_), .Y(mai_mai_n68_));
  AOI210     m046(.A0(mai_mai_n68_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x09), .B(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x10), .B(x06), .Y(mai_mai_n71_));
  NA3        m049(.A(mai_mai_n71_), .B(mai_mai_n70_), .C(mai_mai_n28_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n61_), .B(mai_mai_n41_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n72_), .A1(x11), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  NO2        m053(.A(x10), .B(x09), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n417_), .B(mai_mai_n24_), .Y(mai_mai_n77_));
  NO2        m055(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n78_), .B(mai_mai_n36_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n78_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n80_));
  NO2        m058(.A(mai_mai_n48_), .B(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m059(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n82_));
  NO2        m060(.A(x08), .B(x01), .Y(mai_mai_n83_));
  OAI210     m061(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n35_), .Y(mai_mai_n84_));
  NA2        m062(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n84_), .B(mai_mai_n81_), .C(mai_mai_n77_), .Y(mai_mai_n86_));
  AN2        m064(.A(mai_mai_n86_), .B(mai_mai_n74_), .Y(mai_mai_n87_));
  INV        m065(.A(mai_mai_n84_), .Y(mai_mai_n88_));
  NO2        m066(.A(x06), .B(x05), .Y(mai_mai_n89_));
  NA2        m067(.A(x11), .B(x00), .Y(mai_mai_n90_));
  NO2        m068(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n91_));
  NOi21      m069(.An(mai_mai_n90_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  AOI210     m070(.A0(mai_mai_n89_), .A1(mai_mai_n88_), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  NOi21      m071(.An(x01), .B(x10), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n95_));
  NO3        m073(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(x06), .Y(mai_mai_n96_));
  NA2        m074(.A(mai_mai_n96_), .B(mai_mai_n27_), .Y(mai_mai_n97_));
  OAI210     m075(.A0(mai_mai_n93_), .A1(x07), .B0(mai_mai_n97_), .Y(mai_mai_n98_));
  NO3        m076(.A(mai_mai_n98_), .B(mai_mai_n87_), .C(mai_mai_n69_), .Y(mai01));
  INV        m077(.A(x12), .Y(mai_mai_n100_));
  INV        m078(.A(x13), .Y(mai_mai_n101_));
  NA2        m079(.A(x04), .B(mai_mai_n89_), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n94_), .B(mai_mai_n28_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n70_), .Y(mai_mai_n104_));
  NO2        m082(.A(x10), .B(x01), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(mai_mai_n105_), .Y(mai_mai_n107_));
  NA2        m085(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n108_));
  NO3        m086(.A(mai_mai_n108_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n109_));
  AOI210     m087(.A0(mai_mai_n109_), .A1(mai_mai_n107_), .B0(mai_mai_n104_), .Y(mai_mai_n110_));
  AOI210     m088(.A0(mai_mai_n110_), .A1(mai_mai_n102_), .B0(mai_mai_n101_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n112_));
  NOi21      m090(.An(mai_mai_n112_), .B(mai_mai_n58_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n114_));
  NA3        m092(.A(x08), .B(mai_mai_n114_), .C(x06), .Y(mai_mai_n115_));
  INV        m093(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n83_), .B(x13), .Y(mai_mai_n117_));
  NA2        m095(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n118_), .B(x05), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n120_));
  NO2        m098(.A(x00), .B(mai_mai_n71_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n122_));
  NA2        m100(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(mai_mai_n122_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(x13), .Y(mai_mai_n126_));
  NO2        m104(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n127_));
  NOi41      m105(.An(mai_mai_n126_), .B(mai_mai_n127_), .C(mai_mai_n57_), .D(mai_mai_n124_), .Y(mai_mai_n128_));
  NO3        m106(.A(mai_mai_n128_), .B(x06), .C(x03), .Y(mai_mai_n129_));
  NO4        m107(.A(mai_mai_n129_), .B(mai_mai_n121_), .C(mai_mai_n116_), .D(mai_mai_n111_), .Y(mai_mai_n130_));
  NA2        m108(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n131_));
  OAI210     m109(.A0(mai_mai_n83_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n35_), .B(mai_mai_n47_), .Y(mai_mai_n134_));
  OA210      m112(.A0(x00), .A1(mai_mai_n76_), .B0(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n137_));
  AOI210     m115(.A0(mai_mai_n137_), .A1(mai_mai_n49_), .B0(mai_mai_n136_), .Y(mai_mai_n138_));
  OA210      m116(.A0(mai_mai_n138_), .A1(mai_mai_n135_), .B0(mai_mai_n133_), .Y(mai_mai_n139_));
  NO2        m117(.A(x09), .B(x05), .Y(mai_mai_n140_));
  NA2        m118(.A(mai_mai_n140_), .B(mai_mai_n47_), .Y(mai_mai_n141_));
  AOI210     m119(.A0(mai_mai_n141_), .A1(mai_mai_n107_), .B0(mai_mai_n49_), .Y(mai_mai_n142_));
  NA2        m120(.A(x09), .B(x00), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n112_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n75_), .B(mai_mai_n51_), .Y(mai_mai_n145_));
  AOI210     m123(.A0(mai_mai_n145_), .A1(mai_mai_n144_), .B0(mai_mai_n137_), .Y(mai_mai_n146_));
  NO3        m124(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n139_), .Y(mai_mai_n147_));
  NO2        m125(.A(x03), .B(x02), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n84_), .B(mai_mai_n101_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n149_), .A1(mai_mai_n113_), .B0(mai_mai_n148_), .Y(mai_mai_n150_));
  OA210      m128(.A0(mai_mai_n147_), .A1(x11), .B0(mai_mai_n150_), .Y(mai_mai_n151_));
  OAI210     m129(.A0(mai_mai_n130_), .A1(mai_mai_n23_), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  NA2        m130(.A(mai_mai_n107_), .B(mai_mai_n40_), .Y(mai_mai_n153_));
  NAi21      m131(.An(x06), .B(x10), .Y(mai_mai_n154_));
  NOi21      m132(.An(x01), .B(x13), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n154_), .Y(mai_mai_n156_));
  BUFFER     m134(.A(mai_mai_n156_), .Y(mai_mai_n157_));
  AOI210     m135(.A0(mai_mai_n157_), .A1(mai_mai_n153_), .B0(mai_mai_n41_), .Y(mai_mai_n158_));
  NO2        m136(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n101_), .B(x01), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(x08), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n159_), .B(mai_mai_n48_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n163_));
  OAI210     m141(.A0(mai_mai_n162_), .A1(mai_mai_n158_), .B0(mai_mai_n163_), .Y(mai_mai_n164_));
  NA2        m142(.A(x04), .B(x02), .Y(mai_mai_n165_));
  NA2        m143(.A(x10), .B(x05), .Y(mai_mai_n166_));
  NO2        m144(.A(x09), .B(x01), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n105_), .B(mai_mai_n31_), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n168_), .B(x00), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n112_), .B(x08), .Y(mai_mai_n170_));
  NA3        m148(.A(mai_mai_n155_), .B(mai_mai_n154_), .C(mai_mai_n51_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n94_), .B(x05), .Y(mai_mai_n172_));
  OAI210     m150(.A0(mai_mai_n172_), .A1(x08), .B0(mai_mai_n171_), .Y(mai_mai_n173_));
  AOI210     m151(.A0(mai_mai_n170_), .A1(x06), .B0(mai_mai_n173_), .Y(mai_mai_n174_));
  OAI210     m152(.A0(mai_mai_n174_), .A1(x11), .B0(mai_mai_n169_), .Y(mai_mai_n175_));
  NAi21      m153(.An(mai_mai_n165_), .B(mai_mai_n175_), .Y(mai_mai_n176_));
  INV        m154(.A(mai_mai_n25_), .Y(mai_mai_n177_));
  NAi21      m155(.An(x13), .B(x00), .Y(mai_mai_n178_));
  AOI210     m156(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n178_), .Y(mai_mai_n179_));
  BUFFER     m157(.A(mai_mai_n179_), .Y(mai_mai_n180_));
  BUFFER     m158(.A(mai_mai_n70_), .Y(mai_mai_n181_));
  NO2        m159(.A(mai_mai_n95_), .B(x06), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n178_), .B(mai_mai_n36_), .Y(mai_mai_n183_));
  INV        m161(.A(mai_mai_n183_), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n185_));
  OAI210     m163(.A0(mai_mai_n185_), .A1(mai_mai_n180_), .B0(mai_mai_n177_), .Y(mai_mai_n186_));
  NOi21      m164(.An(x09), .B(x00), .Y(mai_mai_n187_));
  NO3        m165(.A(mai_mai_n82_), .B(mai_mai_n187_), .C(mai_mai_n47_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(mai_mai_n123_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n100_), .B(mai_mai_n189_), .Y(mai_mai_n190_));
  NO2        m168(.A(mai_mai_n101_), .B(x12), .Y(mai_mai_n191_));
  AOI210     m169(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n191_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n94_), .B(mai_mai_n51_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(x02), .Y(mai_mai_n195_));
  NO2        m173(.A(mai_mai_n195_), .B(mai_mai_n193_), .Y(mai_mai_n196_));
  AOI210     m174(.A0(mai_mai_n192_), .A1(mai_mai_n190_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  NA4        m175(.A(mai_mai_n197_), .B(mai_mai_n186_), .C(mai_mai_n176_), .D(mai_mai_n164_), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n152_), .A1(mai_mai_n100_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n72_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n200_), .B(mai_mai_n133_), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n202_));
  NA2        m180(.A(mai_mai_n202_), .B(mai_mai_n132_), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n122_), .B(x06), .Y(mai_mai_n205_));
  AOI210     m183(.A0(mai_mai_n204_), .A1(mai_mai_n203_), .B0(mai_mai_n205_), .Y(mai_mai_n206_));
  AOI210     m184(.A0(mai_mai_n206_), .A1(mai_mai_n201_), .B0(x12), .Y(mai_mai_n207_));
  INV        m185(.A(mai_mai_n75_), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n156_), .B(mai_mai_n57_), .Y(mai_mai_n209_));
  NA2        m187(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n94_), .B(x06), .Y(mai_mai_n211_));
  AOI210     m189(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n212_));
  NO3        m190(.A(mai_mai_n212_), .B(mai_mai_n211_), .C(mai_mai_n41_), .Y(mai_mai_n213_));
  NA4        m191(.A(mai_mai_n154_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n214_), .B(mai_mai_n137_), .Y(mai_mai_n215_));
  OAI210     m193(.A0(mai_mai_n215_), .A1(mai_mai_n213_), .B0(x02), .Y(mai_mai_n216_));
  AOI210     m194(.A0(mai_mai_n216_), .A1(mai_mai_n210_), .B0(mai_mai_n23_), .Y(mai_mai_n217_));
  OAI210     m195(.A0(mai_mai_n207_), .A1(mai_mai_n57_), .B0(mai_mai_n217_), .Y(mai_mai_n218_));
  INV        m196(.A(mai_mai_n137_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n220_));
  OAI210     m198(.A0(mai_mai_n78_), .A1(mai_mai_n36_), .B0(x04), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n101_), .B(x03), .Y(mai_mai_n222_));
  AOI220     m200(.A0(mai_mai_n222_), .A1(mai_mai_n221_), .B0(mai_mai_n75_), .B1(mai_mai_n220_), .Y(mai_mai_n223_));
  INV        m201(.A(mai_mai_n154_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(mai_mai_n57_), .Y(mai_mai_n225_));
  OAI210     m203(.A0(mai_mai_n223_), .A1(mai_mai_n219_), .B0(mai_mai_n225_), .Y(mai_mai_n226_));
  INV        m204(.A(mai_mai_n91_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n227_), .B(x12), .Y(mai_mai_n228_));
  NA2        m206(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n230_));
  INV        m208(.A(mai_mai_n179_), .Y(mai_mai_n231_));
  AOI210     m209(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n232_));
  NO2        m210(.A(x06), .B(x00), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n234_));
  INV        m212(.A(x03), .Y(mai_mai_n235_));
  OA210      m213(.A0(mai_mai_n235_), .A1(mai_mai_n71_), .B0(mai_mai_n231_), .Y(mai_mai_n236_));
  NA2        m214(.A(x13), .B(mai_mai_n100_), .Y(mai_mai_n237_));
  NA3        m215(.A(mai_mai_n237_), .B(x12), .C(mai_mai_n92_), .Y(mai_mai_n238_));
  OAI210     m216(.A0(mai_mai_n236_), .A1(mai_mai_n229_), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  AOI210     m217(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n239_), .Y(mai_mai_n240_));
  AOI210     m218(.A0(mai_mai_n240_), .A1(mai_mai_n218_), .B0(x07), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n70_), .B(mai_mai_n29_), .Y(mai_mai_n242_));
  AOI210     m220(.A0(mai_mai_n131_), .A1(mai_mai_n145_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  NO2        m221(.A(mai_mai_n101_), .B(x06), .Y(mai_mai_n244_));
  INV        m222(.A(mai_mai_n244_), .Y(mai_mai_n245_));
  NO2        m223(.A(x08), .B(x05), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n246_), .B(mai_mai_n232_), .Y(mai_mai_n247_));
  OAI210     m225(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n248_));
  OAI210     m226(.A0(mai_mai_n247_), .A1(mai_mai_n245_), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  NO2        m227(.A(x12), .B(x02), .Y(mai_mai_n250_));
  INV        m228(.A(mai_mai_n250_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n251_), .B(mai_mai_n227_), .Y(mai_mai_n252_));
  OA210      m230(.A0(mai_mai_n249_), .A1(mai_mai_n243_), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n254_), .B(x01), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n126_), .B(mai_mai_n29_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n244_), .B(mai_mai_n221_), .Y(mai_mai_n257_));
  NA2        m235(.A(mai_mai_n101_), .B(x04), .Y(mai_mai_n258_));
  OAI210     m236(.A0(x02), .A1(mai_mai_n117_), .B0(mai_mai_n257_), .Y(mai_mai_n259_));
  NO3        m237(.A(mai_mai_n90_), .B(x12), .C(x03), .Y(mai_mai_n260_));
  OAI210     m238(.A0(mai_mai_n259_), .A1(mai_mai_n256_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  NOi21      m239(.An(mai_mai_n242_), .B(mai_mai_n211_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n262_), .B(mai_mai_n263_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n265_));
  NO3        m243(.A(mai_mai_n265_), .B(mai_mai_n212_), .C(mai_mai_n182_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n229_), .B(mai_mai_n28_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n266_), .A1(mai_mai_n219_), .B0(mai_mai_n267_), .Y(mai_mai_n268_));
  NA3        m246(.A(mai_mai_n268_), .B(mai_mai_n264_), .C(mai_mai_n261_), .Y(mai_mai_n269_));
  NO3        m247(.A(mai_mai_n269_), .B(mai_mai_n253_), .C(mai_mai_n241_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n199_), .A1(mai_mai_n61_), .B0(mai_mai_n270_), .Y(mai02));
  AOI210     m249(.A0(mai_mai_n131_), .A1(mai_mai_n84_), .B0(mai_mai_n125_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n101_), .B(mai_mai_n35_), .Y(mai_mai_n273_));
  NO2        m251(.A(x00), .B(mai_mai_n32_), .Y(mai_mai_n274_));
  OAI210     m252(.A0(mai_mai_n274_), .A1(mai_mai_n272_), .B0(mai_mai_n166_), .Y(mai_mai_n275_));
  INV        m253(.A(mai_mai_n166_), .Y(mai_mai_n276_));
  AOI210     m254(.A0(mai_mai_n114_), .A1(mai_mai_n85_), .B0(mai_mai_n212_), .Y(mai_mai_n277_));
  OAI220     m255(.A0(mai_mai_n277_), .A1(mai_mai_n101_), .B0(mai_mai_n84_), .B1(mai_mai_n51_), .Y(mai_mai_n278_));
  AOI220     m256(.A0(mai_mai_n278_), .A1(mai_mai_n276_), .B0(mai_mai_n149_), .B1(mai_mai_n148_), .Y(mai_mai_n279_));
  AOI210     m257(.A0(mai_mai_n279_), .A1(mai_mai_n275_), .B0(mai_mai_n48_), .Y(mai_mai_n280_));
  NO2        m258(.A(x05), .B(x02), .Y(mai_mai_n281_));
  OAI210     m259(.A0(mai_mai_n203_), .A1(mai_mai_n187_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  AOI220     m260(.A0(mai_mai_n246_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n283_));
  NOi21      m261(.An(mai_mai_n273_), .B(mai_mai_n283_), .Y(mai_mai_n284_));
  AOI210     m262(.A0(x13), .A1(mai_mai_n78_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  AOI210     m263(.A0(mai_mai_n285_), .A1(mai_mai_n282_), .B0(mai_mai_n137_), .Y(mai_mai_n286_));
  INV        m264(.A(mai_mai_n223_), .Y(mai_mai_n287_));
  NO2        m265(.A(mai_mai_n234_), .B(mai_mai_n47_), .Y(mai_mai_n288_));
  NA2        m266(.A(mai_mai_n288_), .B(mai_mai_n287_), .Y(mai_mai_n289_));
  AN2        m267(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n290_));
  OAI210     m268(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n291_));
  NA2        m269(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n292_));
  AOI210     m270(.A0(mai_mai_n292_), .A1(mai_mai_n132_), .B0(mai_mai_n291_), .Y(mai_mai_n293_));
  OAI210     m271(.A0(mai_mai_n293_), .A1(mai_mai_n290_), .B0(mai_mai_n95_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n247_), .B(mai_mai_n103_), .Y(mai_mai_n295_));
  NA2        m273(.A(mai_mai_n295_), .B(x13), .Y(mai_mai_n296_));
  NA3        m274(.A(mai_mai_n296_), .B(mai_mai_n294_), .C(mai_mai_n289_), .Y(mai_mai_n297_));
  NO3        m275(.A(mai_mai_n297_), .B(mai_mai_n286_), .C(mai_mai_n280_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n136_), .B(x03), .Y(mai_mai_n299_));
  OAI210     m277(.A0(mai_mai_n178_), .A1(mai_mai_n265_), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n300_), .B(mai_mai_n105_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n165_), .B(mai_mai_n160_), .Y(mai_mai_n302_));
  AN2        m280(.A(mai_mai_n302_), .B(mai_mai_n170_), .Y(mai_mai_n303_));
  INV        m281(.A(mai_mai_n56_), .Y(mai_mai_n304_));
  OAI220     m282(.A0(mai_mai_n258_), .A1(mai_mai_n304_), .B0(mai_mai_n125_), .B1(mai_mai_n28_), .Y(mai_mai_n305_));
  OAI210     m283(.A0(mai_mai_n305_), .A1(mai_mai_n303_), .B0(mai_mai_n106_), .Y(mai_mai_n306_));
  NA2        m284(.A(mai_mai_n258_), .B(mai_mai_n100_), .Y(mai_mai_n307_));
  NA2        m285(.A(mai_mai_n100_), .B(mai_mai_n41_), .Y(mai_mai_n308_));
  NA3        m286(.A(mai_mai_n308_), .B(mai_mai_n307_), .C(mai_mai_n124_), .Y(mai_mai_n309_));
  NA4        m287(.A(mai_mai_n309_), .B(mai_mai_n306_), .C(mai_mai_n301_), .D(mai_mai_n48_), .Y(mai_mai_n310_));
  INV        m288(.A(mai_mai_n194_), .Y(mai_mai_n311_));
  NO2        m289(.A(mai_mai_n161_), .B(mai_mai_n40_), .Y(mai_mai_n312_));
  NA2        m290(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n313_));
  OAI220     m291(.A0(mai_mai_n313_), .A1(mai_mai_n312_), .B0(mai_mai_n311_), .B1(mai_mai_n59_), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n314_), .B(x02), .Y(mai_mai_n315_));
  INV        m293(.A(mai_mai_n230_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n191_), .B(x04), .Y(mai_mai_n317_));
  NO3        m295(.A(mai_mai_n191_), .B(mai_mai_n159_), .C(mai_mai_n52_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n143_), .A1(mai_mai_n36_), .B0(mai_mai_n100_), .Y(mai_mai_n319_));
  OAI210     m297(.A0(mai_mai_n319_), .A1(mai_mai_n188_), .B0(mai_mai_n318_), .Y(mai_mai_n320_));
  NA3        m298(.A(mai_mai_n320_), .B(mai_mai_n315_), .C(x06), .Y(mai_mai_n321_));
  NA2        m299(.A(x09), .B(x03), .Y(mai_mai_n322_));
  OAI220     m300(.A0(mai_mai_n322_), .A1(mai_mai_n123_), .B0(mai_mai_n202_), .B1(mai_mai_n63_), .Y(mai_mai_n323_));
  NO2        m301(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n318_), .B(mai_mai_n324_), .Y(mai_mai_n325_));
  INV        m303(.A(mai_mai_n325_), .Y(mai_mai_n326_));
  AO220      m304(.A0(mai_mai_n326_), .A1(x04), .B0(mai_mai_n323_), .B1(x05), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n310_), .B0(mai_mai_n327_), .Y(mai_mai_n328_));
  OAI210     m306(.A0(mai_mai_n298_), .A1(x12), .B0(mai_mai_n328_), .Y(mai03));
  OR2        m307(.A(mai_mai_n42_), .B(mai_mai_n220_), .Y(mai_mai_n330_));
  AOI210     m308(.A0(mai_mai_n149_), .A1(mai_mai_n100_), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  AO210      m309(.A0(mai_mai_n316_), .A1(mai_mai_n85_), .B0(mai_mai_n317_), .Y(mai_mai_n332_));
  NA2        m310(.A(mai_mai_n191_), .B(mai_mai_n148_), .Y(mai_mai_n333_));
  NA3        m311(.A(mai_mai_n333_), .B(mai_mai_n332_), .C(mai_mai_n195_), .Y(mai_mai_n334_));
  OAI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n331_), .B0(x05), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n330_), .B(x05), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n132_), .A1(mai_mai_n208_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  AOI210     m315(.A0(mai_mai_n222_), .A1(mai_mai_n79_), .B0(mai_mai_n119_), .Y(mai_mai_n338_));
  OAI220     m316(.A0(mai_mai_n338_), .A1(mai_mai_n59_), .B0(mai_mai_n292_), .B1(mai_mai_n283_), .Y(mai_mai_n339_));
  OAI210     m317(.A0(mai_mai_n339_), .A1(mai_mai_n337_), .B0(mai_mai_n100_), .Y(mai_mai_n340_));
  AOI210     m318(.A0(mai_mai_n141_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n341_));
  NO2        m319(.A(mai_mai_n167_), .B(mai_mai_n127_), .Y(mai_mai_n342_));
  OAI220     m320(.A0(mai_mai_n342_), .A1(mai_mai_n37_), .B0(mai_mai_n144_), .B1(x13), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(x04), .Y(mai_mai_n344_));
  NO3        m322(.A(mai_mai_n308_), .B(mai_mai_n84_), .C(mai_mai_n59_), .Y(mai_mai_n345_));
  AOI210     m323(.A0(mai_mai_n184_), .A1(mai_mai_n100_), .B0(mai_mai_n141_), .Y(mai_mai_n346_));
  OA210      m324(.A0(mai_mai_n161_), .A1(x12), .B0(mai_mai_n127_), .Y(mai_mai_n347_));
  NO3        m325(.A(mai_mai_n347_), .B(mai_mai_n346_), .C(mai_mai_n345_), .Y(mai_mai_n348_));
  NA4        m326(.A(mai_mai_n348_), .B(mai_mai_n344_), .C(mai_mai_n340_), .D(mai_mai_n335_), .Y(mai04));
  NO2        m327(.A(mai_mai_n88_), .B(mai_mai_n39_), .Y(mai_mai_n350_));
  XO2        m328(.A(mai_mai_n350_), .B(mai_mai_n237_), .Y(mai05));
  AOI210     m329(.A0(mai_mai_n70_), .A1(mai_mai_n52_), .B0(mai_mai_n205_), .Y(mai_mai_n352_));
  AOI210     m330(.A0(mai_mai_n352_), .A1(mai_mai_n291_), .B0(mai_mai_n25_), .Y(mai_mai_n353_));
  NO2        m331(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n354_));
  OAI210     m332(.A0(mai_mai_n354_), .A1(mai_mai_n353_), .B0(mai_mai_n100_), .Y(mai_mai_n355_));
  NA2        m333(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n356_));
  NA2        m334(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n357_));
  NA2        m335(.A(mai_mai_n242_), .B(x03), .Y(mai_mai_n358_));
  OAI220     m336(.A0(mai_mai_n358_), .A1(mai_mai_n357_), .B0(mai_mai_n356_), .B1(mai_mai_n80_), .Y(mai_mai_n359_));
  OAI210     m337(.A0(mai_mai_n26_), .A1(mai_mai_n100_), .B0(x07), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n359_), .A1(x06), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  AOI220     m339(.A0(mai_mai_n80_), .A1(mai_mai_n31_), .B0(mai_mai_n52_), .B1(mai_mai_n51_), .Y(mai_mai_n362_));
  NO3        m340(.A(mai_mai_n362_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n363_));
  AOI210     m341(.A0(mai_mai_n418_), .A1(mai_mai_n358_), .B0(mai_mai_n244_), .Y(mai_mai_n364_));
  OR2        m342(.A(mai_mai_n364_), .B(mai_mai_n229_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n155_), .B(x05), .Y(mai_mai_n366_));
  NA3        m344(.A(mai_mai_n366_), .B(mai_mai_n233_), .C(mai_mai_n227_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n368_));
  OAI210     m346(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n369_));
  OR3        m347(.A(mai_mai_n369_), .B(mai_mai_n368_), .C(mai_mai_n44_), .Y(mai_mai_n370_));
  NA3        m348(.A(mai_mai_n370_), .B(mai_mai_n367_), .C(mai_mai_n365_), .Y(mai_mai_n371_));
  OAI210     m349(.A0(mai_mai_n371_), .A1(mai_mai_n363_), .B0(mai_mai_n100_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n33_), .B(mai_mai_n100_), .Y(mai_mai_n373_));
  AOI210     m351(.A0(mai_mai_n373_), .A1(mai_mai_n91_), .B0(x07), .Y(mai_mai_n374_));
  AOI220     m352(.A0(mai_mai_n374_), .A1(mai_mai_n372_), .B0(mai_mai_n361_), .B1(mai_mai_n355_), .Y(mai_mai_n375_));
  NA3        m353(.A(mai_mai_n23_), .B(mai_mai_n61_), .C(mai_mai_n48_), .Y(mai_mai_n376_));
  AO210      m354(.A0(mai_mai_n376_), .A1(mai_mai_n254_), .B0(mai_mai_n251_), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n73_), .B(mai_mai_n136_), .Y(mai_mai_n378_));
  OR2        m356(.A(mai_mai_n378_), .B(x03), .Y(mai_mai_n379_));
  NA2        m357(.A(mai_mai_n324_), .B(mai_mai_n61_), .Y(mai_mai_n380_));
  NO3        m358(.A(mai_mai_n324_), .B(mai_mai_n140_), .C(mai_mai_n28_), .Y(mai_mai_n381_));
  AOI220     m359(.A0(mai_mai_n381_), .A1(mai_mai_n379_), .B0(mai_mai_n377_), .B1(mai_mai_n47_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n382_), .B(mai_mai_n101_), .Y(mai_mai_n383_));
  AOI210     m361(.A0(mai_mai_n317_), .A1(mai_mai_n108_), .B0(mai_mai_n250_), .Y(mai_mai_n384_));
  NOi21      m362(.An(mai_mai_n299_), .B(mai_mai_n127_), .Y(mai_mai_n385_));
  OAI210     m363(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n386_));
  AOI210     m364(.A0(mai_mai_n237_), .A1(mai_mai_n47_), .B0(mai_mai_n386_), .Y(mai_mai_n387_));
  NO3        m365(.A(mai_mai_n387_), .B(mai_mai_n384_), .C(x08), .Y(mai_mai_n388_));
  NA2        m366(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n389_), .B(x03), .Y(mai_mai_n390_));
  NO2        m368(.A(x13), .B(x12), .Y(mai_mai_n391_));
  NO2        m369(.A(mai_mai_n125_), .B(mai_mai_n28_), .Y(mai_mai_n392_));
  NO2        m370(.A(mai_mai_n392_), .B(mai_mai_n255_), .Y(mai_mai_n393_));
  NA3        m371(.A(mai_mai_n311_), .B(mai_mai_n120_), .C(x12), .Y(mai_mai_n394_));
  AO210      m372(.A0(mai_mai_n311_), .A1(mai_mai_n120_), .B0(mai_mai_n237_), .Y(mai_mai_n395_));
  NA3        m373(.A(mai_mai_n395_), .B(mai_mai_n394_), .C(x08), .Y(mai_mai_n396_));
  AOI210     m374(.A0(mai_mai_n391_), .A1(mai_mai_n390_), .B0(mai_mai_n396_), .Y(mai_mai_n397_));
  AOI210     m375(.A0(mai_mai_n388_), .A1(mai_mai_n383_), .B0(mai_mai_n397_), .Y(mai_mai_n398_));
  OAI210     m376(.A0(mai_mai_n380_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n166_), .B(mai_mai_n357_), .Y(mai_mai_n400_));
  OAI210     m378(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n183_), .Y(mai_mai_n401_));
  NA3        m379(.A(mai_mai_n393_), .B(mai_mai_n385_), .C(mai_mai_n307_), .Y(mai_mai_n402_));
  INV        m380(.A(x14), .Y(mai_mai_n403_));
  NO3        m381(.A(mai_mai_n299_), .B(mai_mai_n103_), .C(x11), .Y(mai_mai_n404_));
  NO3        m382(.A(mai_mai_n160_), .B(mai_mai_n73_), .C(mai_mai_n57_), .Y(mai_mai_n405_));
  NO3        m383(.A(mai_mai_n376_), .B(mai_mai_n308_), .C(mai_mai_n178_), .Y(mai_mai_n406_));
  NO4        m384(.A(mai_mai_n406_), .B(mai_mai_n405_), .C(mai_mai_n404_), .D(mai_mai_n403_), .Y(mai_mai_n407_));
  NA3        m385(.A(mai_mai_n407_), .B(mai_mai_n402_), .C(mai_mai_n401_), .Y(mai_mai_n408_));
  AOI220     m386(.A0(mai_mai_n373_), .A1(mai_mai_n61_), .B0(mai_mai_n392_), .B1(mai_mai_n159_), .Y(mai_mai_n409_));
  NOi21      m387(.An(mai_mai_n258_), .B(mai_mai_n144_), .Y(mai_mai_n410_));
  NO2        m388(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n411_));
  OAI210     m389(.A0(mai_mai_n411_), .A1(mai_mai_n410_), .B0(mai_mai_n100_), .Y(mai_mai_n412_));
  OAI210     m390(.A0(mai_mai_n409_), .A1(mai_mai_n90_), .B0(mai_mai_n412_), .Y(mai_mai_n413_));
  NO4        m391(.A(mai_mai_n413_), .B(mai_mai_n408_), .C(mai_mai_n398_), .D(mai_mai_n375_), .Y(mai06));
  INV        m392(.A(x07), .Y(mai_mai_n417_));
  INV        m393(.A(x02), .Y(mai_mai_n418_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  INV        u027(.A(x09), .Y(men_men_n50_));
  NO2        u028(.A(x10), .B(x02), .Y(men_men_n51_));
  NOi21      u029(.An(x01), .B(x09), .Y(men_men_n52_));
  INV        u030(.A(x00), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n54_), .B(men_men_n52_), .Y(men_men_n55_));
  NA2        u033(.A(x09), .B(men_men_n53_), .Y(men_men_n56_));
  INV        u034(.A(x07), .Y(men_men_n57_));
  AOI220     u035(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n57_), .Y(men_men_n58_));
  INV        u036(.A(men_men_n55_), .Y(men_men_n59_));
  NA2        u037(.A(men_men_n29_), .B(x02), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n60_), .B(men_men_n24_), .Y(men_men_n61_));
  OAI220     u039(.A0(men_men_n61_), .A1(men_men_n59_), .B0(men_men_n58_), .B1(men_men_n56_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n57_), .B(men_men_n48_), .Y(men_men_n63_));
  OAI210     u041(.A0(men_men_n30_), .A1(x11), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u042(.A0(men_men_n64_), .A1(men_men_n55_), .B0(men_men_n62_), .B1(men_men_n31_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n65_), .B(x05), .Y(men_men_n66_));
  NA2        u044(.A(x10), .B(x09), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n57_), .B(men_men_n23_), .Y(men_men_n68_));
  NA2        u046(.A(x09), .B(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x06), .Y(men_men_n70_));
  NA3        u048(.A(men_men_n70_), .B(men_men_n69_), .C(men_men_n28_), .Y(men_men_n71_));
  OAI210     u049(.A0(men_men_n71_), .A1(men_men_n68_), .B0(x03), .Y(men_men_n72_));
  NOi31      u050(.An(x08), .B(x04), .C(x00), .Y(men_men_n73_));
  INV        u051(.A(men_men_n24_), .Y(men_men_n74_));
  NO2        u052(.A(x09), .B(men_men_n41_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n75_), .B(men_men_n36_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n77_));
  INV        u055(.A(men_men_n77_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n36_), .B(x00), .Y(men_men_n79_));
  NO2        u057(.A(x08), .B(x01), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n80_), .A1(men_men_n79_), .B0(men_men_n35_), .Y(men_men_n81_));
  NA2        u059(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n82_));
  NO3        u060(.A(men_men_n81_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n83_));
  AN2        u061(.A(men_men_n83_), .B(men_men_n72_), .Y(men_men_n84_));
  INV        u062(.A(men_men_n81_), .Y(men_men_n85_));
  NO2        u063(.A(x06), .B(x05), .Y(men_men_n86_));
  NA2        u064(.A(x11), .B(x00), .Y(men_men_n87_));
  NO2        u065(.A(x11), .B(men_men_n47_), .Y(men_men_n88_));
  NOi21      u066(.An(men_men_n87_), .B(men_men_n88_), .Y(men_men_n89_));
  NOi21      u067(.An(x01), .B(x10), .Y(men_men_n90_));
  NO2        u068(.A(men_men_n29_), .B(men_men_n53_), .Y(men_men_n91_));
  NO3        u069(.A(men_men_n91_), .B(men_men_n90_), .C(x06), .Y(men_men_n92_));
  NA2        u070(.A(men_men_n92_), .B(men_men_n27_), .Y(men_men_n93_));
  OAI210     u071(.A0(men_men_n423_), .A1(x07), .B0(men_men_n93_), .Y(men_men_n94_));
  NO3        u072(.A(men_men_n94_), .B(men_men_n84_), .C(men_men_n66_), .Y(men01));
  INV        u073(.A(x12), .Y(men_men_n96_));
  INV        u074(.A(x13), .Y(men_men_n97_));
  NA2        u075(.A(men_men_n86_), .B(x01), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n98_), .B(men_men_n67_), .Y(men_men_n99_));
  NA2        u077(.A(x08), .B(x04), .Y(men_men_n100_));
  NO2        u078(.A(men_men_n100_), .B(men_men_n53_), .Y(men_men_n101_));
  NA2        u079(.A(men_men_n101_), .B(men_men_n99_), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n90_), .B(men_men_n28_), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n103_), .B(men_men_n69_), .Y(men_men_n104_));
  NO2        u082(.A(x10), .B(x01), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n29_), .B(x00), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NA2        u085(.A(x04), .B(men_men_n28_), .Y(men_men_n108_));
  NO3        u086(.A(men_men_n108_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n109_));
  AOI210     u087(.A0(men_men_n109_), .A1(men_men_n107_), .B0(men_men_n104_), .Y(men_men_n110_));
  AOI210     u088(.A0(men_men_n110_), .A1(men_men_n102_), .B0(men_men_n97_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n52_), .B(x05), .Y(men_men_n112_));
  NOi21      u090(.An(men_men_n112_), .B(men_men_n54_), .Y(men_men_n113_));
  NA3        u091(.A(x13), .B(men_men_n425_), .C(x06), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n114_), .B(men_men_n113_), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n80_), .B(x13), .Y(men_men_n116_));
  NA2        u094(.A(x09), .B(men_men_n35_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u096(.A(x13), .B(men_men_n35_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(x05), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(men_men_n118_), .Y(men_men_n121_));
  NA2        u099(.A(men_men_n35_), .B(men_men_n53_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n122_), .B(men_men_n97_), .Y(men_men_n123_));
  AOI210     u101(.A0(men_men_n123_), .A1(men_men_n76_), .B0(men_men_n113_), .Y(men_men_n124_));
  AOI210     u102(.A0(men_men_n124_), .A1(men_men_n121_), .B0(men_men_n70_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n126_));
  NA2        u104(.A(x10), .B(men_men_n53_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n50_), .B(x05), .Y(men_men_n129_));
  NO3        u107(.A(men_men_n122_), .B(men_men_n75_), .C(men_men_n36_), .Y(men_men_n130_));
  NO2        u108(.A(men_men_n56_), .B(x05), .Y(men_men_n131_));
  NO3        u109(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n132_), .B(x06), .C(x03), .Y(men_men_n133_));
  NO4        u111(.A(men_men_n133_), .B(men_men_n125_), .C(men_men_n115_), .D(men_men_n111_), .Y(men_men_n134_));
  NA2        u112(.A(x13), .B(men_men_n36_), .Y(men_men_n135_));
  OAI210     u113(.A0(men_men_n80_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n136_), .B(men_men_n135_), .Y(men_men_n137_));
  NO2        u115(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n29_), .B(x06), .Y(men_men_n139_));
  AOI210     u117(.A0(men_men_n139_), .A1(men_men_n49_), .B0(men_men_n138_), .Y(men_men_n140_));
  NO2        u118(.A(x09), .B(x05), .Y(men_men_n141_));
  NA2        u119(.A(men_men_n141_), .B(men_men_n47_), .Y(men_men_n142_));
  NA2        u120(.A(x09), .B(x00), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n112_), .B(men_men_n143_), .Y(men_men_n144_));
  INV        u122(.A(men_men_n73_), .Y(men_men_n145_));
  NO2        u123(.A(x03), .B(x02), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n81_), .B(men_men_n97_), .Y(men_men_n147_));
  OAI210     u125(.A0(men_men_n147_), .A1(men_men_n113_), .B0(men_men_n146_), .Y(men_men_n148_));
  OA210      u126(.A0(men_men_n427_), .A1(x11), .B0(men_men_n148_), .Y(men_men_n149_));
  OAI210     u127(.A0(men_men_n134_), .A1(men_men_n23_), .B0(men_men_n149_), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n107_), .B(men_men_n40_), .Y(men_men_n151_));
  NAi21      u129(.An(x06), .B(x10), .Y(men_men_n152_));
  NA2        u130(.A(x01), .B(men_men_n152_), .Y(men_men_n153_));
  OR2        u131(.A(men_men_n153_), .B(x08), .Y(men_men_n154_));
  AOI210     u132(.A0(men_men_n154_), .A1(men_men_n151_), .B0(men_men_n41_), .Y(men_men_n155_));
  NO2        u133(.A(men_men_n29_), .B(x03), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n97_), .B(x01), .Y(men_men_n157_));
  NO2        u135(.A(men_men_n157_), .B(x08), .Y(men_men_n158_));
  AOI210     u136(.A0(x09), .A1(men_men_n156_), .B0(men_men_n48_), .Y(men_men_n159_));
  AOI210     u137(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n160_));
  OAI210     u138(.A0(men_men_n159_), .A1(men_men_n155_), .B0(men_men_n160_), .Y(men_men_n161_));
  NA2        u139(.A(x04), .B(x02), .Y(men_men_n162_));
  NA2        u140(.A(x10), .B(x05), .Y(men_men_n163_));
  NA2        u141(.A(x09), .B(x06), .Y(men_men_n164_));
  NO2        u142(.A(x09), .B(x01), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n424_), .B(x11), .Y(men_men_n166_));
  NAi21      u144(.An(men_men_n162_), .B(men_men_n166_), .Y(men_men_n167_));
  INV        u145(.A(men_men_n25_), .Y(men_men_n168_));
  NAi21      u146(.An(x13), .B(x00), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n169_), .Y(men_men_n170_));
  AOI220     u148(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n163_), .A1(men_men_n35_), .B0(men_men_n171_), .Y(men_men_n172_));
  AN2        u150(.A(men_men_n172_), .B(men_men_n170_), .Y(men_men_n173_));
  BUFFER     u151(.A(men_men_n70_), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n169_), .B(men_men_n36_), .Y(men_men_n175_));
  INV        u153(.A(men_men_n175_), .Y(men_men_n176_));
  OAI210     u154(.A0(men_men_n176_), .A1(men_men_n164_), .B0(men_men_n174_), .Y(men_men_n177_));
  OAI210     u155(.A0(men_men_n177_), .A1(men_men_n173_), .B0(men_men_n168_), .Y(men_men_n178_));
  NOi21      u156(.An(x09), .B(x00), .Y(men_men_n179_));
  NO3        u157(.A(men_men_n79_), .B(men_men_n179_), .C(men_men_n47_), .Y(men_men_n180_));
  INV        u158(.A(men_men_n180_), .Y(men_men_n181_));
  NA2        u159(.A(x10), .B(x08), .Y(men_men_n182_));
  INV        u160(.A(men_men_n182_), .Y(men_men_n183_));
  NA2        u161(.A(x06), .B(x05), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(men_men_n35_), .B0(men_men_n96_), .Y(men_men_n185_));
  AOI210     u163(.A0(men_men_n183_), .A1(men_men_n54_), .B0(men_men_n185_), .Y(men_men_n186_));
  NA2        u164(.A(men_men_n186_), .B(men_men_n181_), .Y(men_men_n187_));
  NO2        u165(.A(men_men_n97_), .B(x12), .Y(men_men_n188_));
  AOI210     u166(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n188_), .Y(men_men_n189_));
  NA2        u167(.A(men_men_n90_), .B(men_men_n50_), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n191_), .B(x02), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n192_), .B(men_men_n190_), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n189_), .A1(men_men_n187_), .B0(men_men_n193_), .Y(men_men_n194_));
  NA4        u172(.A(men_men_n194_), .B(men_men_n178_), .C(men_men_n167_), .D(men_men_n161_), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n150_), .A1(men_men_n96_), .B0(men_men_n195_), .Y(men_men_n196_));
  INV        u174(.A(men_men_n71_), .Y(men_men_n197_));
  NA2        u175(.A(men_men_n197_), .B(men_men_n137_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n199_));
  NO2        u177(.A(men_men_n126_), .B(x06), .Y(men_men_n200_));
  INV        u178(.A(men_men_n200_), .Y(men_men_n201_));
  AOI210     u179(.A0(men_men_n201_), .A1(men_men_n198_), .B0(x12), .Y(men_men_n202_));
  INV        u180(.A(men_men_n73_), .Y(men_men_n203_));
  NO2        u181(.A(x05), .B(men_men_n50_), .Y(men_men_n204_));
  OAI210     u182(.A0(men_men_n204_), .A1(men_men_n153_), .B0(men_men_n53_), .Y(men_men_n205_));
  NA2        u183(.A(men_men_n205_), .B(men_men_n203_), .Y(men_men_n206_));
  INV        u184(.A(men_men_n139_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(x02), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n208_), .A1(men_men_n206_), .B0(men_men_n23_), .Y(men_men_n209_));
  OAI210     u187(.A0(men_men_n202_), .A1(men_men_n53_), .B0(men_men_n209_), .Y(men_men_n210_));
  INV        u188(.A(men_men_n139_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n50_), .B(x03), .Y(men_men_n212_));
  OAI210     u190(.A0(men_men_n75_), .A1(men_men_n36_), .B0(men_men_n117_), .Y(men_men_n213_));
  NO2        u191(.A(men_men_n97_), .B(x03), .Y(men_men_n214_));
  NA2        u192(.A(men_men_n32_), .B(x06), .Y(men_men_n215_));
  INV        u193(.A(men_men_n152_), .Y(men_men_n216_));
  NOi21      u194(.An(x13), .B(x04), .Y(men_men_n217_));
  NO3        u195(.A(men_men_n217_), .B(men_men_n73_), .C(men_men_n179_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n218_), .B(x05), .Y(men_men_n219_));
  AOI220     u197(.A0(men_men_n219_), .A1(men_men_n215_), .B0(men_men_n216_), .B1(men_men_n53_), .Y(men_men_n220_));
  INV        u198(.A(men_men_n220_), .Y(men_men_n221_));
  INV        u199(.A(men_men_n88_), .Y(men_men_n222_));
  NO2        u200(.A(men_men_n222_), .B(x12), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n225_), .A1(men_men_n172_), .B0(men_men_n170_), .Y(men_men_n226_));
  AOI210     u204(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n227_), .B(men_men_n41_), .Y(men_men_n228_));
  OAI210     u206(.A0(men_men_n100_), .A1(men_men_n143_), .B0(men_men_n70_), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  NA2        u208(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n231_), .B(x03), .Y(men_men_n232_));
  OA210      u210(.A0(men_men_n232_), .A1(men_men_n230_), .B0(men_men_n226_), .Y(men_men_n233_));
  NA2        u211(.A(x13), .B(men_men_n96_), .Y(men_men_n234_));
  NA3        u212(.A(men_men_n234_), .B(men_men_n185_), .C(men_men_n89_), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n233_), .A1(men_men_n224_), .B0(men_men_n235_), .Y(men_men_n236_));
  AOI210     u214(.A0(men_men_n223_), .A1(men_men_n221_), .B0(men_men_n236_), .Y(men_men_n237_));
  AOI210     u215(.A0(men_men_n237_), .A1(men_men_n210_), .B0(x07), .Y(men_men_n238_));
  NA2        u216(.A(men_men_n69_), .B(men_men_n29_), .Y(men_men_n239_));
  NO2        u217(.A(men_men_n217_), .B(men_men_n179_), .Y(men_men_n240_));
  AOI210     u218(.A0(men_men_n240_), .A1(men_men_n145_), .B0(men_men_n239_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n97_), .B(x06), .Y(men_men_n242_));
  INV        u220(.A(men_men_n242_), .Y(men_men_n243_));
  NO2        u221(.A(x08), .B(x05), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n244_), .B(men_men_n227_), .Y(men_men_n245_));
  NA2        u223(.A(x13), .B(men_men_n31_), .Y(men_men_n246_));
  OAI210     u224(.A0(men_men_n245_), .A1(men_men_n243_), .B0(men_men_n246_), .Y(men_men_n247_));
  NO2        u225(.A(x12), .B(x02), .Y(men_men_n248_));
  INV        u226(.A(men_men_n248_), .Y(men_men_n249_));
  NO2        u227(.A(men_men_n249_), .B(men_men_n222_), .Y(men_men_n250_));
  OA210      u228(.A0(men_men_n247_), .A1(men_men_n241_), .B0(men_men_n250_), .Y(men_men_n251_));
  NA2        u229(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(x01), .Y(men_men_n253_));
  NOi21      u231(.An(men_men_n80_), .B(men_men_n117_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NO2        u233(.A(men_men_n255_), .B(men_men_n29_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n242_), .B(men_men_n213_), .Y(men_men_n257_));
  NA2        u235(.A(men_men_n97_), .B(x04), .Y(men_men_n258_));
  NA2        u236(.A(men_men_n258_), .B(men_men_n28_), .Y(men_men_n259_));
  OAI210     u237(.A0(men_men_n259_), .A1(men_men_n116_), .B0(men_men_n257_), .Y(men_men_n260_));
  NO3        u238(.A(men_men_n87_), .B(x12), .C(x03), .Y(men_men_n261_));
  OAI210     u239(.A0(men_men_n260_), .A1(men_men_n256_), .B0(men_men_n261_), .Y(men_men_n262_));
  AOI210     u240(.A0(men_men_n190_), .A1(men_men_n184_), .B0(men_men_n100_), .Y(men_men_n263_));
  NOi21      u241(.An(men_men_n239_), .B(men_men_n426_), .Y(men_men_n264_));
  NO2        u242(.A(men_men_n25_), .B(x00), .Y(men_men_n265_));
  OAI210     u243(.A0(men_men_n264_), .A1(men_men_n263_), .B0(men_men_n265_), .Y(men_men_n266_));
  NO2        u244(.A(men_men_n54_), .B(x05), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n224_), .B(men_men_n28_), .Y(men_men_n268_));
  NA2        u246(.A(men_men_n211_), .B(men_men_n268_), .Y(men_men_n269_));
  NA3        u247(.A(men_men_n269_), .B(men_men_n266_), .C(men_men_n262_), .Y(men_men_n270_));
  NO3        u248(.A(men_men_n270_), .B(men_men_n251_), .C(men_men_n238_), .Y(men_men_n271_));
  OAI210     u249(.A0(men_men_n196_), .A1(men_men_n57_), .B0(men_men_n271_), .Y(men02));
  AOI210     u250(.A0(men_men_n135_), .A1(men_men_n81_), .B0(men_men_n129_), .Y(men_men_n273_));
  NOi21      u251(.An(men_men_n218_), .B(men_men_n165_), .Y(men_men_n274_));
  NA3        u252(.A(x13), .B(men_men_n183_), .C(men_men_n52_), .Y(men_men_n275_));
  OAI210     u253(.A0(men_men_n274_), .A1(men_men_n32_), .B0(men_men_n275_), .Y(men_men_n276_));
  OAI210     u254(.A0(men_men_n276_), .A1(men_men_n273_), .B0(men_men_n163_), .Y(men_men_n277_));
  INV        u255(.A(men_men_n163_), .Y(men_men_n278_));
  OAI220     u256(.A0(men_men_n50_), .A1(men_men_n97_), .B0(men_men_n81_), .B1(men_men_n50_), .Y(men_men_n279_));
  AOI220     u257(.A0(men_men_n279_), .A1(men_men_n278_), .B0(men_men_n147_), .B1(men_men_n146_), .Y(men_men_n280_));
  AOI210     u258(.A0(men_men_n280_), .A1(men_men_n277_), .B0(men_men_n48_), .Y(men_men_n281_));
  NO2        u259(.A(x05), .B(x02), .Y(men_men_n282_));
  OAI210     u260(.A0(men_men_n47_), .A1(men_men_n179_), .B0(men_men_n282_), .Y(men_men_n283_));
  AOI220     u261(.A0(men_men_n244_), .A1(men_men_n54_), .B0(men_men_n52_), .B1(men_men_n36_), .Y(men_men_n284_));
  NO2        u262(.A(men_men_n283_), .B(men_men_n139_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n231_), .B(men_men_n47_), .Y(men_men_n286_));
  NA2        u264(.A(men_men_n286_), .B(men_men_n219_), .Y(men_men_n287_));
  OAI210     u265(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n288_));
  NA2        u266(.A(x13), .B(men_men_n28_), .Y(men_men_n289_));
  OA210      u267(.A0(men_men_n289_), .A1(x08), .B0(men_men_n142_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n290_), .A1(men_men_n136_), .B0(men_men_n288_), .Y(men_men_n291_));
  NA2        u269(.A(men_men_n291_), .B(men_men_n91_), .Y(men_men_n292_));
  NA3        u270(.A(men_men_n91_), .B(men_men_n80_), .C(men_men_n212_), .Y(men_men_n293_));
  NA3        u271(.A(men_men_n90_), .B(men_men_n79_), .C(men_men_n42_), .Y(men_men_n294_));
  AOI210     u272(.A0(men_men_n294_), .A1(men_men_n293_), .B0(x04), .Y(men_men_n295_));
  INV        u273(.A(men_men_n146_), .Y(men_men_n296_));
  OAI220     u274(.A0(men_men_n245_), .A1(men_men_n103_), .B0(men_men_n296_), .B1(men_men_n128_), .Y(men_men_n297_));
  AOI210     u275(.A0(men_men_n297_), .A1(x13), .B0(men_men_n295_), .Y(men_men_n298_));
  NA3        u276(.A(men_men_n298_), .B(men_men_n292_), .C(men_men_n287_), .Y(men_men_n299_));
  NO3        u277(.A(men_men_n299_), .B(men_men_n285_), .C(men_men_n281_), .Y(men_men_n300_));
  NA2        u278(.A(men_men_n138_), .B(x03), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n35_), .A1(men_men_n267_), .B0(men_men_n301_), .Y(men_men_n302_));
  NA2        u280(.A(men_men_n302_), .B(men_men_n105_), .Y(men_men_n303_));
  NO2        u281(.A(men_men_n129_), .B(men_men_n28_), .Y(men_men_n304_));
  NA2        u282(.A(men_men_n304_), .B(men_men_n106_), .Y(men_men_n305_));
  NA2        u283(.A(men_men_n258_), .B(men_men_n96_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n96_), .B(men_men_n41_), .Y(men_men_n307_));
  NA3        u285(.A(men_men_n307_), .B(men_men_n306_), .C(men_men_n128_), .Y(men_men_n308_));
  NA4        u286(.A(men_men_n308_), .B(men_men_n305_), .C(men_men_n303_), .D(men_men_n48_), .Y(men_men_n309_));
  INV        u287(.A(men_men_n191_), .Y(men_men_n310_));
  NO2        u288(.A(men_men_n158_), .B(men_men_n40_), .Y(men_men_n311_));
  NA2        u289(.A(men_men_n32_), .B(x05), .Y(men_men_n312_));
  OAI220     u290(.A0(men_men_n312_), .A1(men_men_n311_), .B0(men_men_n310_), .B1(men_men_n55_), .Y(men_men_n313_));
  NA2        u291(.A(men_men_n313_), .B(x02), .Y(men_men_n314_));
  INV        u292(.A(men_men_n225_), .Y(men_men_n315_));
  NA2        u293(.A(men_men_n188_), .B(x04), .Y(men_men_n316_));
  NO2        u294(.A(men_men_n316_), .B(men_men_n315_), .Y(men_men_n317_));
  NO3        u295(.A(men_men_n171_), .B(x13), .C(men_men_n31_), .Y(men_men_n318_));
  OAI210     u296(.A0(men_men_n318_), .A1(men_men_n317_), .B0(men_men_n91_), .Y(men_men_n319_));
  NO3        u297(.A(men_men_n188_), .B(men_men_n156_), .C(men_men_n51_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n143_), .A1(men_men_n36_), .B0(men_men_n96_), .Y(men_men_n321_));
  OAI210     u299(.A0(men_men_n321_), .A1(men_men_n180_), .B0(men_men_n320_), .Y(men_men_n322_));
  NA4        u300(.A(men_men_n322_), .B(men_men_n319_), .C(men_men_n314_), .D(x06), .Y(men_men_n323_));
  NA2        u301(.A(x09), .B(x03), .Y(men_men_n324_));
  OAI220     u302(.A0(men_men_n324_), .A1(men_men_n127_), .B0(men_men_n199_), .B1(men_men_n60_), .Y(men_men_n325_));
  OAI220     u303(.A0(men_men_n157_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n326_));
  NO3        u304(.A(men_men_n267_), .B(men_men_n126_), .C(x08), .Y(men_men_n327_));
  AOI210     u305(.A0(men_men_n326_), .A1(men_men_n211_), .B0(men_men_n327_), .Y(men_men_n328_));
  NO3        u306(.A(men_men_n112_), .B(men_men_n127_), .C(men_men_n38_), .Y(men_men_n329_));
  INV        u307(.A(men_men_n329_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n328_), .A1(men_men_n28_), .B0(men_men_n330_), .Y(men_men_n331_));
  AO220      u309(.A0(men_men_n331_), .A1(x04), .B0(men_men_n325_), .B1(x05), .Y(men_men_n332_));
  AOI210     u310(.A0(men_men_n323_), .A1(men_men_n309_), .B0(men_men_n332_), .Y(men_men_n333_));
  OAI210     u311(.A0(men_men_n300_), .A1(x12), .B0(men_men_n333_), .Y(men03));
  OR2        u312(.A(men_men_n42_), .B(men_men_n212_), .Y(men_men_n335_));
  AOI210     u313(.A0(men_men_n147_), .A1(men_men_n96_), .B0(men_men_n335_), .Y(men_men_n336_));
  AO210      u314(.A0(men_men_n315_), .A1(men_men_n82_), .B0(men_men_n316_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n188_), .B(men_men_n146_), .Y(men_men_n338_));
  NA3        u316(.A(men_men_n338_), .B(men_men_n337_), .C(men_men_n192_), .Y(men_men_n339_));
  OAI210     u317(.A0(men_men_n339_), .A1(men_men_n336_), .B0(x05), .Y(men_men_n340_));
  NA2        u318(.A(men_men_n335_), .B(x05), .Y(men_men_n341_));
  AOI210     u319(.A0(men_men_n136_), .A1(men_men_n203_), .B0(men_men_n341_), .Y(men_men_n342_));
  AOI210     u320(.A0(men_men_n214_), .A1(men_men_n76_), .B0(men_men_n120_), .Y(men_men_n343_));
  OAI220     u321(.A0(men_men_n343_), .A1(men_men_n55_), .B0(men_men_n289_), .B1(men_men_n284_), .Y(men_men_n344_));
  OAI210     u322(.A0(men_men_n344_), .A1(men_men_n342_), .B0(men_men_n96_), .Y(men_men_n345_));
  AOI210     u323(.A0(men_men_n142_), .A1(men_men_n56_), .B0(men_men_n38_), .Y(men_men_n346_));
  NO2        u324(.A(men_men_n165_), .B(men_men_n131_), .Y(men_men_n347_));
  OAI220     u325(.A0(men_men_n347_), .A1(men_men_n37_), .B0(men_men_n144_), .B1(x13), .Y(men_men_n348_));
  OAI210     u326(.A0(men_men_n348_), .A1(men_men_n346_), .B0(x04), .Y(men_men_n349_));
  NO3        u327(.A(men_men_n307_), .B(men_men_n81_), .C(men_men_n55_), .Y(men_men_n350_));
  AOI210     u328(.A0(men_men_n176_), .A1(men_men_n96_), .B0(men_men_n142_), .Y(men_men_n351_));
  OA210      u329(.A0(men_men_n158_), .A1(x12), .B0(men_men_n131_), .Y(men_men_n352_));
  NO3        u330(.A(men_men_n352_), .B(men_men_n351_), .C(men_men_n350_), .Y(men_men_n353_));
  NA4        u331(.A(men_men_n353_), .B(men_men_n349_), .C(men_men_n345_), .D(men_men_n340_), .Y(men04));
  NO2        u332(.A(men_men_n85_), .B(men_men_n39_), .Y(men_men_n355_));
  XO2        u333(.A(men_men_n355_), .B(men_men_n234_), .Y(men05));
  NA2        u334(.A(men_men_n129_), .B(men_men_n31_), .Y(men_men_n357_));
  AOI210     u335(.A0(x05), .A1(men_men_n357_), .B0(men_men_n24_), .Y(men_men_n358_));
  NA2        u336(.A(men_men_n358_), .B(men_men_n96_), .Y(men_men_n359_));
  NA2        u337(.A(x11), .B(men_men_n31_), .Y(men_men_n360_));
  NA2        u338(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n361_));
  NA2        u339(.A(men_men_n239_), .B(x03), .Y(men_men_n362_));
  OAI220     u340(.A0(men_men_n362_), .A1(men_men_n361_), .B0(men_men_n360_), .B1(men_men_n77_), .Y(men_men_n363_));
  OAI210     u341(.A0(men_men_n26_), .A1(men_men_n96_), .B0(x07), .Y(men_men_n364_));
  AOI210     u342(.A0(men_men_n363_), .A1(x06), .B0(men_men_n364_), .Y(men_men_n365_));
  NA2        u343(.A(men_men_n77_), .B(men_men_n31_), .Y(men_men_n366_));
  NO3        u344(.A(men_men_n366_), .B(men_men_n23_), .C(x00), .Y(men_men_n367_));
  NA2        u345(.A(men_men_n67_), .B(x02), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n368_), .A1(men_men_n362_), .B0(men_men_n242_), .Y(men_men_n369_));
  OR2        u347(.A(men_men_n369_), .B(men_men_n224_), .Y(men_men_n370_));
  NO2        u348(.A(men_men_n23_), .B(x10), .Y(men_men_n371_));
  OAI210     u349(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n372_));
  OR3        u350(.A(men_men_n372_), .B(men_men_n371_), .C(men_men_n44_), .Y(men_men_n373_));
  NA2        u351(.A(men_men_n373_), .B(men_men_n370_), .Y(men_men_n374_));
  OAI210     u352(.A0(men_men_n374_), .A1(men_men_n367_), .B0(men_men_n96_), .Y(men_men_n375_));
  NA2        u353(.A(men_men_n33_), .B(men_men_n96_), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n376_), .A1(men_men_n88_), .B0(x07), .Y(men_men_n377_));
  AOI220     u355(.A0(men_men_n377_), .A1(men_men_n375_), .B0(men_men_n365_), .B1(men_men_n359_), .Y(men_men_n378_));
  AO210      u356(.A0(x06), .A1(men_men_n252_), .B0(men_men_n249_), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n371_), .A1(x07), .B0(men_men_n138_), .Y(men_men_n380_));
  OR2        u358(.A(men_men_n380_), .B(x03), .Y(men_men_n381_));
  NO2        u359(.A(x07), .B(x11), .Y(men_men_n382_));
  NO3        u360(.A(men_men_n382_), .B(men_men_n141_), .C(men_men_n28_), .Y(men_men_n383_));
  AOI220     u361(.A0(men_men_n383_), .A1(men_men_n381_), .B0(men_men_n379_), .B1(men_men_n47_), .Y(men_men_n384_));
  NO3        u362(.A(men_men_n307_), .B(men_men_n32_), .C(x11), .Y(men_men_n385_));
  OAI210     u363(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n97_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n316_), .A1(men_men_n108_), .B0(men_men_n248_), .Y(men_men_n387_));
  NOi21      u365(.An(men_men_n301_), .B(men_men_n131_), .Y(men_men_n388_));
  NO2        u366(.A(men_men_n388_), .B(men_men_n249_), .Y(men_men_n389_));
  OAI210     u367(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n234_), .A1(men_men_n47_), .B0(men_men_n390_), .Y(men_men_n391_));
  NO4        u369(.A(men_men_n391_), .B(men_men_n389_), .C(men_men_n387_), .D(x08), .Y(men_men_n392_));
  AOI210     u370(.A0(men_men_n371_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n393_));
  OAI210     u371(.A0(x05), .A1(men_men_n393_), .B0(men_men_n360_), .Y(men_men_n394_));
  NO2        u372(.A(x13), .B(x12), .Y(men_men_n395_));
  NO2        u373(.A(men_men_n129_), .B(men_men_n28_), .Y(men_men_n396_));
  NO2        u374(.A(men_men_n396_), .B(men_men_n253_), .Y(men_men_n397_));
  OR3        u375(.A(men_men_n397_), .B(x12), .C(x03), .Y(men_men_n398_));
  NA3        u376(.A(men_men_n310_), .B(men_men_n122_), .C(x12), .Y(men_men_n399_));
  AO210      u377(.A0(men_men_n310_), .A1(men_men_n122_), .B0(men_men_n234_), .Y(men_men_n400_));
  NA4        u378(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n398_), .D(x08), .Y(men_men_n401_));
  AOI210     u379(.A0(men_men_n395_), .A1(men_men_n394_), .B0(men_men_n401_), .Y(men_men_n402_));
  AOI210     u380(.A0(men_men_n392_), .A1(men_men_n386_), .B0(men_men_n402_), .Y(men_men_n403_));
  INV        u381(.A(x07), .Y(men_men_n404_));
  OAI220     u382(.A0(men_men_n404_), .A1(men_men_n361_), .B0(men_men_n141_), .B1(men_men_n43_), .Y(men_men_n405_));
  OAI210     u383(.A0(men_men_n405_), .A1(x11), .B0(men_men_n175_), .Y(men_men_n406_));
  NA3        u384(.A(men_men_n397_), .B(men_men_n388_), .C(men_men_n306_), .Y(men_men_n407_));
  INV        u385(.A(x14), .Y(men_men_n408_));
  NO3        u386(.A(men_men_n301_), .B(men_men_n103_), .C(x11), .Y(men_men_n409_));
  NO3        u387(.A(x06), .B(men_men_n307_), .C(men_men_n169_), .Y(men_men_n410_));
  NO3        u388(.A(men_men_n410_), .B(men_men_n409_), .C(men_men_n408_), .Y(men_men_n411_));
  NA3        u389(.A(men_men_n411_), .B(men_men_n407_), .C(men_men_n406_), .Y(men_men_n412_));
  AOI220     u390(.A0(men_men_n376_), .A1(men_men_n57_), .B0(men_men_n396_), .B1(men_men_n156_), .Y(men_men_n413_));
  NOi21      u391(.An(men_men_n258_), .B(men_men_n144_), .Y(men_men_n414_));
  NO3        u392(.A(men_men_n126_), .B(men_men_n24_), .C(x06), .Y(men_men_n415_));
  AOI210     u393(.A0(men_men_n265_), .A1(men_men_n216_), .B0(men_men_n415_), .Y(men_men_n416_));
  OAI210     u394(.A0(men_men_n44_), .A1(x04), .B0(men_men_n416_), .Y(men_men_n417_));
  OAI210     u395(.A0(men_men_n417_), .A1(men_men_n414_), .B0(men_men_n96_), .Y(men_men_n418_));
  OAI210     u396(.A0(men_men_n413_), .A1(men_men_n87_), .B0(men_men_n418_), .Y(men_men_n419_));
  NO4        u397(.A(men_men_n419_), .B(men_men_n412_), .C(men_men_n403_), .D(men_men_n378_), .Y(men06));
  INV        u398(.A(men_men_n89_), .Y(men_men_n423_));
  INV        u399(.A(x01), .Y(men_men_n424_));
  INV        u400(.A(x02), .Y(men_men_n425_));
  INV        u401(.A(x06), .Y(men_men_n426_));
  INV        u402(.A(men_men_n140_), .Y(men_men_n427_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule