library verilog;
use verilog.vl_types.all;
entity testeflecha_vlg_vec_tst is
end testeflecha_vlg_vec_tst;
