//Benchmark atmr_misex3_1774_0.25

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n33_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  INV        o00(.A(n), .Y(ori_ori_n29_));
  OR2        o01(.A(ori_ori_n33_), .B(ori_ori_n29_), .Y(ori04));
  INV        o02(.A(m), .Y(ori_ori_n33_));
  ZERO       o03(.Y(ori10));
  ZERO       o04(.Y(ori11));
  ZERO       o05(.Y(ori08));
  ZERO       o06(.Y(ori09));
  ZERO       o07(.Y(ori12));
  ZERO       o08(.Y(ori13));
  ZERO       o09(.Y(ori02));
  ZERO       o10(.Y(ori03));
  ZERO       o11(.Y(ori00));
  ZERO       o12(.Y(ori01));
  ZERO       o13(.Y(ori06));
  ZERO       o14(.Y(ori07));
  ZERO       o15(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(m), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(m), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(m), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(m), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(m), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(m), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  NA2        m0034(.A(m), .B(f), .Y(mai_mai_n63_));
  NAi21      m0035(.An(i), .B(j), .Y(mai_mai_n64_));
  NAi32      m0036(.An(n), .Bn(k), .C(m), .Y(mai_mai_n65_));
  NAi31      m0037(.An(l), .B(m), .C(k), .Y(mai_mai_n66_));
  NAi21      m0038(.An(e), .B(h), .Y(mai_mai_n67_));
  NAi41      m0039(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n68_));
  INV        m0040(.A(m), .Y(mai_mai_n69_));
  NOi21      m0041(.An(k), .B(l), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n70_), .B(mai_mai_n69_), .Y(mai_mai_n71_));
  AN4        m0043(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n72_));
  NOi31      m0044(.An(h), .B(m), .C(f), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NAi32      m0046(.An(m), .Bn(k), .C(j), .Y(mai_mai_n75_));
  NOi32      m0047(.An(h), .Bn(m), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n72_), .Y(mai_mai_n77_));
  OA220      m0049(.A0(mai_mai_n77_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .B1(mai_mai_n71_), .Y(mai_mai_n78_));
  INV        m0050(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  INV        m0051(.A(n), .Y(mai_mai_n80_));
  NOi32      m0052(.An(e), .Bn(b), .C(d), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  INV        m0054(.A(j), .Y(mai_mai_n83_));
  AN3        m0055(.A(m), .B(k), .C(i), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(m), .Y(mai_mai_n85_));
  NO2        m0057(.A(mai_mai_n85_), .B(f), .Y(mai_mai_n86_));
  NAi32      m0058(.An(m), .Bn(f), .C(h), .Y(mai_mai_n87_));
  NAi31      m0059(.An(j), .B(m), .C(l), .Y(mai_mai_n88_));
  NO2        m0060(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n89_));
  NA2        m0061(.A(m), .B(l), .Y(mai_mai_n90_));
  NAi31      m0062(.An(k), .B(j), .C(m), .Y(mai_mai_n91_));
  NO3        m0063(.A(mai_mai_n91_), .B(mai_mai_n90_), .C(f), .Y(mai_mai_n92_));
  AN2        m0064(.A(j), .B(m), .Y(mai_mai_n93_));
  NOi32      m0065(.An(m), .Bn(l), .C(i), .Y(mai_mai_n94_));
  NOi21      m0066(.An(m), .B(i), .Y(mai_mai_n95_));
  NOi32      m0067(.An(m), .Bn(j), .C(k), .Y(mai_mai_n96_));
  AOI220     m0068(.A0(mai_mai_n96_), .A1(mai_mai_n95_), .B0(mai_mai_n94_), .B1(mai_mai_n93_), .Y(mai_mai_n97_));
  NO2        m0069(.A(mai_mai_n97_), .B(f), .Y(mai_mai_n98_));
  NO4        m0070(.A(mai_mai_n98_), .B(mai_mai_n92_), .C(mai_mai_n89_), .D(mai_mai_n86_), .Y(mai_mai_n99_));
  NAi41      m0071(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n100_));
  AN2        m0072(.A(e), .B(b), .Y(mai_mai_n101_));
  NOi31      m0073(.An(c), .B(h), .C(f), .Y(mai_mai_n102_));
  NA2        m0074(.A(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  NO3        m0075(.A(mai_mai_n103_), .B(mai_mai_n100_), .C(m), .Y(mai_mai_n104_));
  NOi21      m0076(.An(m), .B(f), .Y(mai_mai_n105_));
  NOi21      m0077(.An(i), .B(h), .Y(mai_mai_n106_));
  NA3        m0078(.A(mai_mai_n106_), .B(mai_mai_n105_), .C(mai_mai_n36_), .Y(mai_mai_n107_));
  INV        m0079(.A(a), .Y(mai_mai_n108_));
  NA2        m0080(.A(mai_mai_n101_), .B(mai_mai_n108_), .Y(mai_mai_n109_));
  INV        m0081(.A(l), .Y(mai_mai_n110_));
  NOi21      m0082(.An(m), .B(n), .Y(mai_mai_n111_));
  AN2        m0083(.A(k), .B(h), .Y(mai_mai_n112_));
  NO2        m0084(.A(mai_mai_n107_), .B(mai_mai_n82_), .Y(mai_mai_n113_));
  INV        m0085(.A(b), .Y(mai_mai_n114_));
  NA2        m0086(.A(l), .B(j), .Y(mai_mai_n115_));
  AN2        m0087(.A(k), .B(i), .Y(mai_mai_n116_));
  NA2        m0088(.A(m), .B(e), .Y(mai_mai_n117_));
  NOi32      m0089(.An(c), .Bn(a), .C(d), .Y(mai_mai_n118_));
  NA2        m0090(.A(mai_mai_n118_), .B(mai_mai_n111_), .Y(mai_mai_n119_));
  NO2        m0091(.A(mai_mai_n113_), .B(mai_mai_n104_), .Y(mai_mai_n120_));
  OAI210     m0092(.A0(mai_mai_n99_), .A1(mai_mai_n82_), .B0(mai_mai_n120_), .Y(mai_mai_n121_));
  NOi31      m0093(.An(k), .B(m), .C(j), .Y(mai_mai_n122_));
  NA3        m0094(.A(mai_mai_n122_), .B(mai_mai_n73_), .C(mai_mai_n72_), .Y(mai_mai_n123_));
  NOi31      m0095(.An(k), .B(m), .C(i), .Y(mai_mai_n124_));
  NA3        m0096(.A(mai_mai_n124_), .B(mai_mai_n76_), .C(mai_mai_n72_), .Y(mai_mai_n125_));
  NA2        m0097(.A(mai_mai_n125_), .B(mai_mai_n123_), .Y(mai_mai_n126_));
  NOi32      m0098(.An(f), .Bn(b), .C(e), .Y(mai_mai_n127_));
  NAi21      m0099(.An(m), .B(h), .Y(mai_mai_n128_));
  NAi21      m0100(.An(m), .B(n), .Y(mai_mai_n129_));
  NAi21      m0101(.An(j), .B(k), .Y(mai_mai_n130_));
  NO3        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(mai_mai_n128_), .Y(mai_mai_n131_));
  NAi41      m0103(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n132_));
  NAi31      m0104(.An(j), .B(k), .C(h), .Y(mai_mai_n133_));
  NO3        m0105(.A(mai_mai_n133_), .B(mai_mai_n132_), .C(mai_mai_n129_), .Y(mai_mai_n134_));
  AOI210     m0106(.A0(mai_mai_n131_), .A1(mai_mai_n127_), .B0(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m0107(.A(k), .B(j), .Y(mai_mai_n136_));
  NO2        m0108(.A(mai_mai_n136_), .B(mai_mai_n129_), .Y(mai_mai_n137_));
  AN2        m0109(.A(k), .B(j), .Y(mai_mai_n138_));
  NAi21      m0110(.An(c), .B(b), .Y(mai_mai_n139_));
  NA2        m0111(.A(f), .B(d), .Y(mai_mai_n140_));
  NO4        m0112(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n138_), .D(mai_mai_n128_), .Y(mai_mai_n141_));
  NA2        m0113(.A(h), .B(c), .Y(mai_mai_n142_));
  NAi31      m0114(.An(f), .B(e), .C(b), .Y(mai_mai_n143_));
  NA2        m0115(.A(mai_mai_n141_), .B(mai_mai_n137_), .Y(mai_mai_n144_));
  NA2        m0116(.A(d), .B(b), .Y(mai_mai_n145_));
  NAi21      m0117(.An(e), .B(f), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NA2        m0119(.A(b), .B(a), .Y(mai_mai_n148_));
  NAi21      m0120(.An(e), .B(m), .Y(mai_mai_n149_));
  NAi21      m0121(.An(c), .B(d), .Y(mai_mai_n150_));
  NAi31      m0122(.An(l), .B(k), .C(h), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n129_), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  NA2        m0124(.A(mai_mai_n152_), .B(mai_mai_n147_), .Y(mai_mai_n153_));
  NAi41      m0125(.An(mai_mai_n126_), .B(mai_mai_n153_), .C(mai_mai_n144_), .D(mai_mai_n135_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(b), .Y(mai_mai_n155_));
  NOi21      m0127(.An(m), .B(d), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  NOi21      m0129(.An(h), .B(i), .Y(mai_mai_n158_));
  NOi21      m0130(.An(k), .B(m), .Y(mai_mai_n159_));
  NA3        m0131(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n160_));
  NOi21      m0132(.An(mai_mai_n157_), .B(mai_mai_n160_), .Y(mai_mai_n161_));
  NOi21      m0133(.An(h), .B(m), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  INV        m0136(.A(mai_mai_n49_), .Y(mai_mai_n165_));
  NOi32      m0137(.An(n), .Bn(k), .C(m), .Y(mai_mai_n166_));
  NA2        m0138(.A(l), .B(i), .Y(mai_mai_n167_));
  NA2        m0139(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  NO2        m0140(.A(mai_mai_n168_), .B(mai_mai_n164_), .Y(mai_mai_n169_));
  NAi31      m0141(.An(d), .B(f), .C(c), .Y(mai_mai_n170_));
  NAi31      m0142(.An(e), .B(f), .C(c), .Y(mai_mai_n171_));
  NA2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NA2        m0144(.A(j), .B(h), .Y(mai_mai_n173_));
  OR3        m0145(.A(n), .B(m), .C(k), .Y(mai_mai_n174_));
  NO2        m0146(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NAi32      m0147(.An(m), .Bn(k), .C(n), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  AOI220     m0149(.A0(mai_mai_n177_), .A1(mai_mai_n157_), .B0(mai_mai_n175_), .B1(mai_mai_n172_), .Y(mai_mai_n178_));
  NO2        m0150(.A(n), .B(m), .Y(mai_mai_n179_));
  NA2        m0151(.A(mai_mai_n179_), .B(mai_mai_n50_), .Y(mai_mai_n180_));
  NAi21      m0152(.An(f), .B(e), .Y(mai_mai_n181_));
  NA2        m0153(.A(d), .B(c), .Y(mai_mai_n182_));
  NO2        m0154(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  NOi21      m0155(.An(mai_mai_n183_), .B(mai_mai_n180_), .Y(mai_mai_n184_));
  NAi31      m0156(.An(m), .B(n), .C(b), .Y(mai_mai_n185_));
  NA2        m0157(.A(k), .B(i), .Y(mai_mai_n186_));
  NAi21      m0158(.An(h), .B(f), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n187_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  NO2        m0160(.A(mai_mai_n185_), .B(mai_mai_n150_), .Y(mai_mai_n189_));
  NA2        m0161(.A(mai_mai_n189_), .B(mai_mai_n188_), .Y(mai_mai_n190_));
  NOi32      m0162(.An(f), .Bn(c), .C(d), .Y(mai_mai_n191_));
  NOi32      m0163(.An(f), .Bn(c), .C(e), .Y(mai_mai_n192_));
  NO2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NO3        m0165(.A(n), .B(m), .C(j), .Y(mai_mai_n194_));
  NA2        m0166(.A(mai_mai_n194_), .B(mai_mai_n112_), .Y(mai_mai_n195_));
  AO210      m0167(.A0(mai_mai_n195_), .A1(mai_mai_n180_), .B0(mai_mai_n193_), .Y(mai_mai_n196_));
  NAi41      m0168(.An(mai_mai_n184_), .B(mai_mai_n196_), .C(mai_mai_n190_), .D(mai_mai_n178_), .Y(mai_mai_n197_));
  OR4        m0169(.A(mai_mai_n197_), .B(mai_mai_n169_), .C(mai_mai_n161_), .D(mai_mai_n154_), .Y(mai_mai_n198_));
  NO4        m0170(.A(mai_mai_n198_), .B(mai_mai_n121_), .C(mai_mai_n79_), .D(mai_mai_n55_), .Y(mai_mai_n199_));
  NA3        m0171(.A(m), .B(mai_mai_n110_), .C(j), .Y(mai_mai_n200_));
  NAi31      m0172(.An(n), .B(h), .C(m), .Y(mai_mai_n201_));
  NO2        m0173(.A(mai_mai_n201_), .B(mai_mai_n200_), .Y(mai_mai_n202_));
  NOi32      m0174(.An(m), .Bn(k), .C(l), .Y(mai_mai_n203_));
  NA3        m0175(.A(mai_mai_n203_), .B(mai_mai_n83_), .C(m), .Y(mai_mai_n204_));
  NO2        m0176(.A(mai_mai_n204_), .B(n), .Y(mai_mai_n205_));
  NOi21      m0177(.An(k), .B(j), .Y(mai_mai_n206_));
  NA4        m0178(.A(mai_mai_n206_), .B(mai_mai_n111_), .C(i), .D(m), .Y(mai_mai_n207_));
  AN2        m0179(.A(i), .B(m), .Y(mai_mai_n208_));
  NA3        m0180(.A(mai_mai_n70_), .B(mai_mai_n208_), .C(mai_mai_n111_), .Y(mai_mai_n209_));
  NA2        m0181(.A(mai_mai_n209_), .B(mai_mai_n207_), .Y(mai_mai_n210_));
  NO3        m0182(.A(mai_mai_n210_), .B(mai_mai_n205_), .C(mai_mai_n202_), .Y(mai_mai_n211_));
  NAi41      m0183(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n212_));
  INV        m0184(.A(mai_mai_n212_), .Y(mai_mai_n213_));
  INV        m0185(.A(f), .Y(mai_mai_n214_));
  INV        m0186(.A(m), .Y(mai_mai_n215_));
  NOi31      m0187(.An(i), .B(j), .C(h), .Y(mai_mai_n216_));
  NOi21      m0188(.An(l), .B(m), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  NO3        m0190(.A(mai_mai_n218_), .B(mai_mai_n215_), .C(mai_mai_n214_), .Y(mai_mai_n219_));
  NA2        m0191(.A(mai_mai_n219_), .B(mai_mai_n213_), .Y(mai_mai_n220_));
  OAI210     m0192(.A0(mai_mai_n211_), .A1(mai_mai_n32_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  NOi21      m0193(.An(n), .B(m), .Y(mai_mai_n222_));
  NOi32      m0194(.An(l), .Bn(i), .C(j), .Y(mai_mai_n223_));
  NA2        m0195(.A(mai_mai_n223_), .B(mai_mai_n222_), .Y(mai_mai_n224_));
  OA220      m0196(.A0(mai_mai_n224_), .A1(mai_mai_n103_), .B0(mai_mai_n75_), .B1(mai_mai_n74_), .Y(mai_mai_n225_));
  NAi21      m0197(.An(j), .B(h), .Y(mai_mai_n226_));
  XN2        m0198(.A(i), .B(h), .Y(mai_mai_n227_));
  NA2        m0199(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  NOi31      m0200(.An(k), .B(n), .C(m), .Y(mai_mai_n229_));
  NOi31      m0201(.An(mai_mai_n229_), .B(mai_mai_n182_), .C(mai_mai_n181_), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n230_), .B(mai_mai_n228_), .Y(mai_mai_n231_));
  NAi31      m0203(.An(f), .B(e), .C(c), .Y(mai_mai_n232_));
  NO4        m0204(.A(mai_mai_n232_), .B(mai_mai_n174_), .C(mai_mai_n173_), .D(mai_mai_n59_), .Y(mai_mai_n233_));
  NA4        m0205(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n234_));
  NAi32      m0206(.An(m), .Bn(i), .C(k), .Y(mai_mai_n235_));
  NO3        m0207(.A(mai_mai_n235_), .B(mai_mai_n87_), .C(mai_mai_n234_), .Y(mai_mai_n236_));
  NA2        m0208(.A(k), .B(h), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n236_), .B(mai_mai_n233_), .Y(mai_mai_n238_));
  NAi21      m0210(.An(n), .B(a), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(mai_mai_n145_), .Y(mai_mai_n240_));
  NAi41      m0212(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n241_), .B(e), .Y(mai_mai_n242_));
  NO3        m0214(.A(mai_mai_n146_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n243_));
  OAI210     m0215(.A0(mai_mai_n243_), .A1(mai_mai_n242_), .B0(mai_mai_n240_), .Y(mai_mai_n244_));
  AN4        m0216(.A(mai_mai_n244_), .B(mai_mai_n238_), .C(mai_mai_n231_), .D(mai_mai_n225_), .Y(mai_mai_n245_));
  OR2        m0217(.A(h), .B(m), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n246_), .B(mai_mai_n100_), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n247_), .B(mai_mai_n127_), .Y(mai_mai_n248_));
  NAi41      m0220(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n249_), .B(mai_mai_n214_), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n159_), .B(mai_mai_n106_), .Y(mai_mai_n251_));
  NAi21      m0223(.An(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  NO2        m0224(.A(n), .B(a), .Y(mai_mai_n253_));
  NAi31      m0225(.An(mai_mai_n241_), .B(mai_mai_n253_), .C(mai_mai_n101_), .Y(mai_mai_n254_));
  AN2        m0226(.A(mai_mai_n254_), .B(mai_mai_n252_), .Y(mai_mai_n255_));
  NAi21      m0227(.An(h), .B(i), .Y(mai_mai_n256_));
  NA2        m0228(.A(mai_mai_n179_), .B(k), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n256_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n258_), .B(mai_mai_n191_), .Y(mai_mai_n259_));
  NA3        m0231(.A(mai_mai_n259_), .B(mai_mai_n255_), .C(mai_mai_n248_), .Y(mai_mai_n260_));
  NOi21      m0232(.An(m), .B(e), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n68_), .B(mai_mai_n69_), .Y(mai_mai_n262_));
  NOi32      m0234(.An(l), .Bn(j), .C(i), .Y(mai_mai_n263_));
  INV        m0235(.A(mai_mai_n44_), .Y(mai_mai_n264_));
  NAi21      m0236(.An(f), .B(m), .Y(mai_mai_n265_));
  NO2        m0237(.A(mai_mai_n65_), .B(mai_mai_n115_), .Y(mai_mai_n266_));
  NA2        m0238(.A(mai_mai_n266_), .B(mai_mai_n264_), .Y(mai_mai_n267_));
  INV        m0239(.A(mai_mai_n267_), .Y(mai_mai_n268_));
  NO3        m0240(.A(mai_mai_n130_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n269_));
  NOi41      m0241(.An(mai_mai_n245_), .B(mai_mai_n268_), .C(mai_mai_n260_), .D(mai_mai_n221_), .Y(mai_mai_n270_));
  NO4        m0242(.A(mai_mai_n202_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n271_));
  NO2        m0243(.A(mai_mai_n271_), .B(mai_mai_n109_), .Y(mai_mai_n272_));
  NA3        m0244(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n273_));
  NAi21      m0245(.An(h), .B(m), .Y(mai_mai_n274_));
  OR4        m0246(.A(mai_mai_n274_), .B(mai_mai_n273_), .C(mai_mai_n224_), .D(e), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n251_), .B(mai_mai_n265_), .Y(mai_mai_n276_));
  NA2        m0248(.A(mai_mai_n276_), .B(mai_mai_n72_), .Y(mai_mai_n277_));
  NAi31      m0249(.An(m), .B(k), .C(h), .Y(mai_mai_n278_));
  NO3        m0250(.A(mai_mai_n129_), .B(mai_mai_n278_), .C(l), .Y(mai_mai_n279_));
  NAi31      m0251(.An(e), .B(d), .C(a), .Y(mai_mai_n280_));
  NA2        m0252(.A(mai_mai_n279_), .B(mai_mai_n127_), .Y(mai_mai_n281_));
  NA3        m0253(.A(mai_mai_n281_), .B(mai_mai_n277_), .C(mai_mai_n275_), .Y(mai_mai_n282_));
  NA4        m0254(.A(mai_mai_n159_), .B(mai_mai_n76_), .C(mai_mai_n72_), .D(mai_mai_n115_), .Y(mai_mai_n283_));
  NA3        m0255(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(mai_mai_n80_), .Y(mai_mai_n284_));
  NO2        m0256(.A(mai_mai_n284_), .B(mai_mai_n193_), .Y(mai_mai_n285_));
  NOi21      m0257(.An(mai_mai_n283_), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  NA3        m0258(.A(e), .B(c), .C(b), .Y(mai_mai_n287_));
  NO2        m0259(.A(mai_mai_n60_), .B(mai_mai_n287_), .Y(mai_mai_n288_));
  NAi32      m0260(.An(k), .Bn(i), .C(j), .Y(mai_mai_n289_));
  INV        m0261(.A(mai_mai_n49_), .Y(mai_mai_n290_));
  NA2        m0262(.A(mai_mai_n288_), .B(mai_mai_n290_), .Y(mai_mai_n291_));
  NAi21      m0263(.An(l), .B(k), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n292_), .B(mai_mai_n49_), .Y(mai_mai_n293_));
  NOi21      m0265(.An(l), .B(j), .Y(mai_mai_n294_));
  NA2        m0266(.A(mai_mai_n162_), .B(mai_mai_n294_), .Y(mai_mai_n295_));
  OR3        m0267(.A(mai_mai_n68_), .B(mai_mai_n69_), .C(e), .Y(mai_mai_n296_));
  AOI210     m0268(.A0(mai_mai_n1549_), .A1(mai_mai_n295_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  INV        m0269(.A(mai_mai_n297_), .Y(mai_mai_n298_));
  NAi32      m0270(.An(j), .Bn(h), .C(i), .Y(mai_mai_n299_));
  NAi21      m0271(.An(m), .B(l), .Y(mai_mai_n300_));
  NO3        m0272(.A(mai_mai_n300_), .B(mai_mai_n299_), .C(mai_mai_n80_), .Y(mai_mai_n301_));
  NA2        m0273(.A(h), .B(m), .Y(mai_mai_n302_));
  NA2        m0274(.A(mai_mai_n166_), .B(mai_mai_n45_), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n303_), .B(mai_mai_n302_), .Y(mai_mai_n304_));
  OAI210     m0276(.A0(mai_mai_n304_), .A1(mai_mai_n301_), .B0(mai_mai_n163_), .Y(mai_mai_n305_));
  NA4        m0277(.A(mai_mai_n305_), .B(mai_mai_n298_), .C(mai_mai_n291_), .D(mai_mai_n286_), .Y(mai_mai_n306_));
  NO2        m0278(.A(mai_mai_n143_), .B(d), .Y(mai_mai_n307_));
  NA2        m0279(.A(mai_mai_n307_), .B(mai_mai_n53_), .Y(mai_mai_n308_));
  NO2        m0280(.A(mai_mai_n103_), .B(mai_mai_n100_), .Y(mai_mai_n309_));
  NAi32      m0281(.An(n), .Bn(m), .C(l), .Y(mai_mai_n310_));
  NO2        m0282(.A(mai_mai_n310_), .B(mai_mai_n299_), .Y(mai_mai_n311_));
  NA2        m0283(.A(mai_mai_n311_), .B(mai_mai_n183_), .Y(mai_mai_n312_));
  NO2        m0284(.A(mai_mai_n119_), .B(mai_mai_n114_), .Y(mai_mai_n313_));
  INV        m0285(.A(mai_mai_n117_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n312_), .B(mai_mai_n308_), .Y(mai_mai_n315_));
  NO4        m0287(.A(mai_mai_n315_), .B(mai_mai_n306_), .C(mai_mai_n282_), .D(mai_mai_n272_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n258_), .B(mai_mai_n192_), .Y(mai_mai_n317_));
  NAi21      m0289(.An(m), .B(k), .Y(mai_mai_n318_));
  NO2        m0290(.A(mai_mai_n227_), .B(mai_mai_n318_), .Y(mai_mai_n319_));
  NAi41      m0291(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n320_));
  NO2        m0292(.A(mai_mai_n320_), .B(mai_mai_n149_), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n321_), .B(mai_mai_n319_), .Y(mai_mai_n322_));
  NO4        m0294(.A(i), .B(mai_mai_n149_), .C(mai_mai_n68_), .D(mai_mai_n69_), .Y(mai_mai_n323_));
  NA2        m0295(.A(e), .B(c), .Y(mai_mai_n324_));
  NO3        m0296(.A(mai_mai_n324_), .B(n), .C(d), .Y(mai_mai_n325_));
  NOi21      m0297(.An(f), .B(h), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n326_), .B(mai_mai_n116_), .Y(mai_mai_n327_));
  NO2        m0299(.A(mai_mai_n327_), .B(mai_mai_n215_), .Y(mai_mai_n328_));
  NAi31      m0300(.An(d), .B(e), .C(b), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n129_), .B(mai_mai_n329_), .Y(mai_mai_n330_));
  NA2        m0302(.A(mai_mai_n330_), .B(mai_mai_n328_), .Y(mai_mai_n331_));
  NAi41      m0303(.An(mai_mai_n323_), .B(mai_mai_n331_), .C(mai_mai_n322_), .D(mai_mai_n317_), .Y(mai_mai_n332_));
  NO4        m0304(.A(mai_mai_n320_), .B(mai_mai_n75_), .C(mai_mai_n67_), .D(mai_mai_n215_), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n253_), .B(mai_mai_n101_), .Y(mai_mai_n334_));
  OR2        m0306(.A(mai_mai_n334_), .B(mai_mai_n204_), .Y(mai_mai_n335_));
  NOi31      m0307(.An(l), .B(n), .C(m), .Y(mai_mai_n336_));
  NA2        m0308(.A(mai_mai_n336_), .B(mai_mai_n216_), .Y(mai_mai_n337_));
  NO2        m0309(.A(mai_mai_n337_), .B(mai_mai_n193_), .Y(mai_mai_n338_));
  NAi32      m0310(.An(mai_mai_n338_), .Bn(mai_mai_n333_), .C(mai_mai_n335_), .Y(mai_mai_n339_));
  NAi32      m0311(.An(m), .Bn(j), .C(k), .Y(mai_mai_n340_));
  NAi41      m0312(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n341_));
  NA2        m0313(.A(mai_mai_n212_), .B(mai_mai_n341_), .Y(mai_mai_n342_));
  NOi31      m0314(.An(j), .B(m), .C(k), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n122_), .B(mai_mai_n343_), .Y(mai_mai_n344_));
  AN3        m0316(.A(h), .B(m), .C(f), .Y(mai_mai_n345_));
  NAi31      m0317(.An(mai_mai_n344_), .B(mai_mai_n345_), .C(mai_mai_n342_), .Y(mai_mai_n346_));
  NOi32      m0318(.An(m), .Bn(j), .C(l), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n347_), .B(mai_mai_n94_), .Y(mai_mai_n348_));
  NAi32      m0320(.An(mai_mai_n348_), .Bn(mai_mai_n201_), .C(mai_mai_n307_), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n350_));
  NO2        m0322(.A(mai_mai_n218_), .B(m), .Y(mai_mai_n351_));
  NO2        m0323(.A(mai_mai_n155_), .B(mai_mai_n80_), .Y(mai_mai_n352_));
  AOI220     m0324(.A0(mai_mai_n352_), .A1(mai_mai_n351_), .B0(mai_mai_n250_), .B1(mai_mai_n350_), .Y(mai_mai_n353_));
  INV        m0325(.A(mai_mai_n235_), .Y(mai_mai_n354_));
  NA3        m0326(.A(mai_mai_n354_), .B(mai_mai_n345_), .C(mai_mai_n213_), .Y(mai_mai_n355_));
  NA4        m0327(.A(mai_mai_n355_), .B(mai_mai_n353_), .C(mai_mai_n349_), .D(mai_mai_n346_), .Y(mai_mai_n356_));
  NA3        m0328(.A(h), .B(m), .C(f), .Y(mai_mai_n357_));
  NO2        m0329(.A(mai_mai_n357_), .B(mai_mai_n71_), .Y(mai_mai_n358_));
  NA2        m0330(.A(mai_mai_n341_), .B(mai_mai_n212_), .Y(mai_mai_n359_));
  NA2        m0331(.A(mai_mai_n162_), .B(e), .Y(mai_mai_n360_));
  NO2        m0332(.A(mai_mai_n360_), .B(mai_mai_n41_), .Y(mai_mai_n361_));
  AOI220     m0333(.A0(mai_mai_n361_), .A1(mai_mai_n313_), .B0(mai_mai_n359_), .B1(mai_mai_n358_), .Y(mai_mai_n362_));
  NOi32      m0334(.An(j), .Bn(m), .C(i), .Y(mai_mai_n363_));
  NA3        m0335(.A(mai_mai_n363_), .B(mai_mai_n292_), .C(mai_mai_n111_), .Y(mai_mai_n364_));
  AO210      m0336(.A0(mai_mai_n109_), .A1(mai_mai_n32_), .B0(mai_mai_n364_), .Y(mai_mai_n365_));
  NOi32      m0337(.An(e), .Bn(b), .C(a), .Y(mai_mai_n366_));
  AN2        m0338(.A(l), .B(j), .Y(mai_mai_n367_));
  NO2        m0339(.A(mai_mai_n318_), .B(mai_mai_n367_), .Y(mai_mai_n368_));
  NO3        m0340(.A(mai_mai_n320_), .B(mai_mai_n67_), .C(mai_mai_n215_), .Y(mai_mai_n369_));
  NA3        m0341(.A(mai_mai_n209_), .B(mai_mai_n207_), .C(mai_mai_n35_), .Y(mai_mai_n370_));
  AOI220     m0342(.A0(mai_mai_n370_), .A1(mai_mai_n366_), .B0(mai_mai_n369_), .B1(mai_mai_n368_), .Y(mai_mai_n371_));
  NO2        m0343(.A(mai_mai_n329_), .B(n), .Y(mai_mai_n372_));
  NA2        m0344(.A(mai_mai_n208_), .B(k), .Y(mai_mai_n373_));
  NA3        m0345(.A(m), .B(mai_mai_n110_), .C(mai_mai_n214_), .Y(mai_mai_n374_));
  NA4        m0346(.A(mai_mai_n203_), .B(mai_mai_n83_), .C(m), .D(mai_mai_n214_), .Y(mai_mai_n375_));
  OAI210     m0347(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n375_), .Y(mai_mai_n376_));
  NAi41      m0348(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n377_));
  NA2        m0349(.A(mai_mai_n51_), .B(mai_mai_n111_), .Y(mai_mai_n378_));
  NO2        m0350(.A(mai_mai_n378_), .B(mai_mai_n377_), .Y(mai_mai_n379_));
  AOI220     m0351(.A0(mai_mai_n379_), .A1(b), .B0(mai_mai_n376_), .B1(mai_mai_n372_), .Y(mai_mai_n380_));
  NA4        m0352(.A(mai_mai_n380_), .B(mai_mai_n371_), .C(mai_mai_n365_), .D(mai_mai_n362_), .Y(mai_mai_n381_));
  NO4        m0353(.A(mai_mai_n381_), .B(mai_mai_n356_), .C(mai_mai_n339_), .D(mai_mai_n332_), .Y(mai_mai_n382_));
  NA4        m0354(.A(mai_mai_n382_), .B(mai_mai_n316_), .C(mai_mai_n270_), .D(mai_mai_n199_), .Y(mai10));
  NA3        m0355(.A(m), .B(k), .C(i), .Y(mai_mai_n384_));
  NO3        m0356(.A(mai_mai_n384_), .B(j), .C(mai_mai_n215_), .Y(mai_mai_n385_));
  NOi21      m0357(.An(e), .B(f), .Y(mai_mai_n386_));
  NO4        m0358(.A(mai_mai_n150_), .B(mai_mai_n386_), .C(n), .D(mai_mai_n108_), .Y(mai_mai_n387_));
  NAi31      m0359(.An(b), .B(f), .C(c), .Y(mai_mai_n388_));
  INV        m0360(.A(mai_mai_n388_), .Y(mai_mai_n389_));
  NOi32      m0361(.An(k), .Bn(h), .C(j), .Y(mai_mai_n390_));
  NA2        m0362(.A(mai_mai_n390_), .B(mai_mai_n222_), .Y(mai_mai_n391_));
  NA2        m0363(.A(mai_mai_n160_), .B(mai_mai_n391_), .Y(mai_mai_n392_));
  AOI220     m0364(.A0(mai_mai_n392_), .A1(mai_mai_n389_), .B0(mai_mai_n387_), .B1(mai_mai_n385_), .Y(mai_mai_n393_));
  AN2        m0365(.A(j), .B(h), .Y(mai_mai_n394_));
  NO3        m0366(.A(n), .B(m), .C(k), .Y(mai_mai_n395_));
  NA2        m0367(.A(mai_mai_n395_), .B(mai_mai_n394_), .Y(mai_mai_n396_));
  NO3        m0368(.A(mai_mai_n396_), .B(mai_mai_n150_), .C(mai_mai_n214_), .Y(mai_mai_n397_));
  OR2        m0369(.A(m), .B(k), .Y(mai_mai_n398_));
  NO2        m0370(.A(mai_mai_n173_), .B(mai_mai_n398_), .Y(mai_mai_n399_));
  NA4        m0371(.A(n), .B(f), .C(c), .D(mai_mai_n114_), .Y(mai_mai_n400_));
  NOi21      m0372(.An(mai_mai_n399_), .B(mai_mai_n400_), .Y(mai_mai_n401_));
  NOi32      m0373(.An(d), .Bn(a), .C(c), .Y(mai_mai_n402_));
  NA2        m0374(.A(mai_mai_n402_), .B(mai_mai_n181_), .Y(mai_mai_n403_));
  NAi21      m0375(.An(i), .B(m), .Y(mai_mai_n404_));
  NAi31      m0376(.An(k), .B(m), .C(j), .Y(mai_mai_n405_));
  NO3        m0377(.A(mai_mai_n405_), .B(mai_mai_n404_), .C(n), .Y(mai_mai_n406_));
  NOi21      m0378(.An(mai_mai_n406_), .B(mai_mai_n403_), .Y(mai_mai_n407_));
  NO3        m0379(.A(mai_mai_n407_), .B(mai_mai_n401_), .C(mai_mai_n397_), .Y(mai_mai_n408_));
  NO2        m0380(.A(mai_mai_n400_), .B(mai_mai_n300_), .Y(mai_mai_n409_));
  NOi32      m0381(.An(f), .Bn(d), .C(c), .Y(mai_mai_n410_));
  AOI220     m0382(.A0(mai_mai_n410_), .A1(mai_mai_n311_), .B0(mai_mai_n409_), .B1(mai_mai_n216_), .Y(mai_mai_n411_));
  NA3        m0383(.A(mai_mai_n411_), .B(mai_mai_n408_), .C(mai_mai_n393_), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n59_), .B(mai_mai_n114_), .Y(mai_mai_n413_));
  NA2        m0385(.A(mai_mai_n253_), .B(mai_mai_n413_), .Y(mai_mai_n414_));
  INV        m0386(.A(e), .Y(mai_mai_n415_));
  NA2        m0387(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n416_));
  OAI220     m0388(.A0(mai_mai_n416_), .A1(mai_mai_n200_), .B0(mai_mai_n204_), .B1(mai_mai_n415_), .Y(mai_mai_n417_));
  AN2        m0389(.A(m), .B(e), .Y(mai_mai_n418_));
  NA3        m0390(.A(mai_mai_n418_), .B(mai_mai_n203_), .C(i), .Y(mai_mai_n419_));
  OAI210     m0391(.A0(mai_mai_n85_), .A1(mai_mai_n415_), .B0(mai_mai_n419_), .Y(mai_mai_n420_));
  NO2        m0392(.A(mai_mai_n97_), .B(mai_mai_n415_), .Y(mai_mai_n421_));
  NO3        m0393(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(mai_mai_n417_), .Y(mai_mai_n422_));
  NOi32      m0394(.An(h), .Bn(e), .C(m), .Y(mai_mai_n423_));
  NA3        m0395(.A(mai_mai_n423_), .B(mai_mai_n294_), .C(m), .Y(mai_mai_n424_));
  NOi21      m0396(.An(m), .B(h), .Y(mai_mai_n425_));
  AN3        m0397(.A(m), .B(l), .C(i), .Y(mai_mai_n426_));
  NA3        m0398(.A(mai_mai_n426_), .B(mai_mai_n425_), .C(e), .Y(mai_mai_n427_));
  AN3        m0399(.A(h), .B(m), .C(e), .Y(mai_mai_n428_));
  NA2        m0400(.A(mai_mai_n428_), .B(mai_mai_n94_), .Y(mai_mai_n429_));
  AN3        m0401(.A(mai_mai_n429_), .B(mai_mai_n427_), .C(mai_mai_n424_), .Y(mai_mai_n430_));
  AOI210     m0402(.A0(mai_mai_n430_), .A1(mai_mai_n422_), .B0(mai_mai_n414_), .Y(mai_mai_n431_));
  NA3        m0403(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n432_));
  NO2        m0404(.A(mai_mai_n432_), .B(mai_mai_n414_), .Y(mai_mai_n433_));
  NA3        m0405(.A(mai_mai_n402_), .B(mai_mai_n181_), .C(mai_mai_n80_), .Y(mai_mai_n434_));
  NAi31      m0406(.An(b), .B(c), .C(a), .Y(mai_mai_n435_));
  NO2        m0407(.A(mai_mai_n435_), .B(n), .Y(mai_mai_n436_));
  OAI210     m0408(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n437_));
  NO2        m0409(.A(mai_mai_n437_), .B(mai_mai_n146_), .Y(mai_mai_n438_));
  NA2        m0410(.A(mai_mai_n438_), .B(mai_mai_n436_), .Y(mai_mai_n439_));
  INV        m0411(.A(mai_mai_n439_), .Y(mai_mai_n440_));
  NO4        m0412(.A(mai_mai_n440_), .B(mai_mai_n433_), .C(mai_mai_n431_), .D(mai_mai_n412_), .Y(mai_mai_n441_));
  NA2        m0413(.A(i), .B(m), .Y(mai_mai_n442_));
  NO3        m0414(.A(mai_mai_n280_), .B(mai_mai_n442_), .C(c), .Y(mai_mai_n443_));
  NOi21      m0415(.An(a), .B(n), .Y(mai_mai_n444_));
  NOi21      m0416(.An(d), .B(c), .Y(mai_mai_n445_));
  NA2        m0417(.A(mai_mai_n445_), .B(mai_mai_n444_), .Y(mai_mai_n446_));
  NA3        m0418(.A(i), .B(m), .C(f), .Y(mai_mai_n447_));
  OR2        m0419(.A(mai_mai_n447_), .B(mai_mai_n66_), .Y(mai_mai_n448_));
  NA3        m0420(.A(mai_mai_n426_), .B(mai_mai_n425_), .C(mai_mai_n181_), .Y(mai_mai_n449_));
  AOI210     m0421(.A0(mai_mai_n449_), .A1(mai_mai_n448_), .B0(mai_mai_n446_), .Y(mai_mai_n450_));
  AOI210     m0422(.A0(mai_mai_n443_), .A1(mai_mai_n293_), .B0(mai_mai_n450_), .Y(mai_mai_n451_));
  OR2        m0423(.A(n), .B(m), .Y(mai_mai_n452_));
  NO2        m0424(.A(mai_mai_n452_), .B(mai_mai_n151_), .Y(mai_mai_n453_));
  NO2        m0425(.A(mai_mai_n182_), .B(mai_mai_n146_), .Y(mai_mai_n454_));
  OAI210     m0426(.A0(mai_mai_n453_), .A1(mai_mai_n175_), .B0(mai_mai_n454_), .Y(mai_mai_n455_));
  INV        m0427(.A(mai_mai_n378_), .Y(mai_mai_n456_));
  NA3        m0428(.A(mai_mai_n456_), .B(mai_mai_n366_), .C(d), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n435_), .B(mai_mai_n49_), .Y(mai_mai_n458_));
  NAi21      m0430(.An(k), .B(j), .Y(mai_mai_n459_));
  NAi21      m0431(.An(e), .B(d), .Y(mai_mai_n460_));
  INV        m0432(.A(mai_mai_n460_), .Y(mai_mai_n461_));
  NO2        m0433(.A(mai_mai_n257_), .B(mai_mai_n214_), .Y(mai_mai_n462_));
  NA3        m0434(.A(mai_mai_n462_), .B(mai_mai_n461_), .C(mai_mai_n228_), .Y(mai_mai_n463_));
  NA3        m0435(.A(mai_mai_n463_), .B(mai_mai_n457_), .C(mai_mai_n455_), .Y(mai_mai_n464_));
  NO2        m0436(.A(mai_mai_n337_), .B(mai_mai_n214_), .Y(mai_mai_n465_));
  NA2        m0437(.A(mai_mai_n465_), .B(mai_mai_n461_), .Y(mai_mai_n466_));
  NOi31      m0438(.An(n), .B(m), .C(k), .Y(mai_mai_n467_));
  AOI220     m0439(.A0(mai_mai_n467_), .A1(mai_mai_n394_), .B0(mai_mai_n222_), .B1(mai_mai_n50_), .Y(mai_mai_n468_));
  NAi31      m0440(.An(m), .B(f), .C(c), .Y(mai_mai_n469_));
  OR3        m0441(.A(mai_mai_n469_), .B(mai_mai_n468_), .C(e), .Y(mai_mai_n470_));
  NA3        m0442(.A(mai_mai_n470_), .B(mai_mai_n466_), .C(mai_mai_n312_), .Y(mai_mai_n471_));
  NOi41      m0443(.An(mai_mai_n451_), .B(mai_mai_n471_), .C(mai_mai_n464_), .D(mai_mai_n268_), .Y(mai_mai_n472_));
  NOi32      m0444(.An(c), .Bn(a), .C(b), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n473_), .B(mai_mai_n111_), .Y(mai_mai_n474_));
  INV        m0446(.A(mai_mai_n278_), .Y(mai_mai_n475_));
  AN2        m0447(.A(e), .B(d), .Y(mai_mai_n476_));
  NA2        m0448(.A(mai_mai_n476_), .B(mai_mai_n475_), .Y(mai_mai_n477_));
  INV        m0449(.A(mai_mai_n146_), .Y(mai_mai_n478_));
  NO2        m0450(.A(mai_mai_n128_), .B(mai_mai_n41_), .Y(mai_mai_n479_));
  NO2        m0451(.A(mai_mai_n63_), .B(e), .Y(mai_mai_n480_));
  AOI210     m0452(.A0(mai_mai_n479_), .A1(mai_mai_n478_), .B0(mai_mai_n480_), .Y(mai_mai_n481_));
  AOI210     m0453(.A0(mai_mai_n481_), .A1(mai_mai_n477_), .B0(mai_mai_n474_), .Y(mai_mai_n482_));
  NO2        m0454(.A(mai_mai_n210_), .B(mai_mai_n205_), .Y(mai_mai_n483_));
  NOi21      m0455(.An(a), .B(b), .Y(mai_mai_n484_));
  NA3        m0456(.A(e), .B(d), .C(c), .Y(mai_mai_n485_));
  NAi21      m0457(.An(mai_mai_n485_), .B(mai_mai_n484_), .Y(mai_mai_n486_));
  NO2        m0458(.A(mai_mai_n434_), .B(mai_mai_n204_), .Y(mai_mai_n487_));
  NOi21      m0459(.An(mai_mai_n486_), .B(mai_mai_n487_), .Y(mai_mai_n488_));
  AOI210     m0460(.A0(mai_mai_n271_), .A1(mai_mai_n483_), .B0(mai_mai_n488_), .Y(mai_mai_n489_));
  NO4        m0461(.A(mai_mai_n187_), .B(mai_mai_n100_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n490_));
  NA2        m0462(.A(mai_mai_n389_), .B(mai_mai_n152_), .Y(mai_mai_n491_));
  OR2        m0463(.A(k), .B(j), .Y(mai_mai_n492_));
  NA2        m0464(.A(l), .B(k), .Y(mai_mai_n493_));
  NA3        m0465(.A(mai_mai_n493_), .B(mai_mai_n492_), .C(mai_mai_n222_), .Y(mai_mai_n494_));
  AOI210     m0466(.A0(mai_mai_n235_), .A1(mai_mai_n340_), .B0(mai_mai_n80_), .Y(mai_mai_n495_));
  NOi21      m0467(.An(mai_mai_n494_), .B(mai_mai_n495_), .Y(mai_mai_n496_));
  OR3        m0468(.A(mai_mai_n496_), .B(mai_mai_n142_), .C(mai_mai_n132_), .Y(mai_mai_n497_));
  NA3        m0469(.A(mai_mai_n283_), .B(mai_mai_n125_), .C(mai_mai_n123_), .Y(mai_mai_n498_));
  NA2        m0470(.A(mai_mai_n402_), .B(mai_mai_n111_), .Y(mai_mai_n499_));
  NO4        m0471(.A(mai_mai_n499_), .B(mai_mai_n91_), .C(mai_mai_n110_), .D(e), .Y(mai_mai_n500_));
  NO3        m0472(.A(mai_mai_n434_), .B(mai_mai_n88_), .C(mai_mai_n128_), .Y(mai_mai_n501_));
  NO4        m0473(.A(mai_mai_n501_), .B(mai_mai_n500_), .C(mai_mai_n498_), .D(mai_mai_n323_), .Y(mai_mai_n502_));
  NA3        m0474(.A(mai_mai_n502_), .B(mai_mai_n497_), .C(mai_mai_n491_), .Y(mai_mai_n503_));
  NO4        m0475(.A(mai_mai_n503_), .B(mai_mai_n490_), .C(mai_mai_n489_), .D(mai_mai_n482_), .Y(mai_mai_n504_));
  NOi21      m0476(.An(d), .B(e), .Y(mai_mai_n505_));
  NO2        m0477(.A(mai_mai_n187_), .B(mai_mai_n56_), .Y(mai_mai_n506_));
  NAi31      m0478(.An(j), .B(l), .C(i), .Y(mai_mai_n507_));
  OAI210     m0479(.A0(mai_mai_n507_), .A1(mai_mai_n129_), .B0(mai_mai_n100_), .Y(mai_mai_n508_));
  NA4        m0480(.A(mai_mai_n508_), .B(mai_mai_n506_), .C(mai_mai_n505_), .D(b), .Y(mai_mai_n509_));
  NO3        m0481(.A(mai_mai_n403_), .B(mai_mai_n348_), .C(mai_mai_n201_), .Y(mai_mai_n510_));
  NO2        m0482(.A(mai_mai_n403_), .B(mai_mai_n378_), .Y(mai_mai_n511_));
  NO4        m0483(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n184_), .D(mai_mai_n309_), .Y(mai_mai_n512_));
  NA3        m0484(.A(mai_mai_n512_), .B(mai_mai_n509_), .C(mai_mai_n245_), .Y(mai_mai_n513_));
  OAI210     m0485(.A0(mai_mai_n124_), .A1(mai_mai_n122_), .B0(n), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n514_), .B(mai_mai_n128_), .Y(mai_mai_n515_));
  AO210      m0487(.A0(mai_mai_n301_), .A1(mai_mai_n215_), .B0(mai_mai_n247_), .Y(mai_mai_n516_));
  OA210      m0488(.A0(mai_mai_n516_), .A1(mai_mai_n515_), .B0(mai_mai_n192_), .Y(mai_mai_n517_));
  XO2        m0489(.A(i), .B(h), .Y(mai_mai_n518_));
  NA3        m0490(.A(mai_mai_n518_), .B(mai_mai_n159_), .C(n), .Y(mai_mai_n519_));
  NAi41      m0491(.An(mai_mai_n301_), .B(mai_mai_n519_), .C(mai_mai_n468_), .D(mai_mai_n391_), .Y(mai_mai_n520_));
  NOi32      m0492(.An(mai_mai_n520_), .Bn(mai_mai_n480_), .C(mai_mai_n273_), .Y(mai_mai_n521_));
  NAi31      m0493(.An(c), .B(f), .C(d), .Y(mai_mai_n522_));
  AOI210     m0494(.A0(mai_mai_n284_), .A1(mai_mai_n195_), .B0(mai_mai_n522_), .Y(mai_mai_n523_));
  NOi21      m0495(.An(mai_mai_n78_), .B(mai_mai_n523_), .Y(mai_mai_n524_));
  NA3        m0496(.A(mai_mai_n387_), .B(mai_mai_n94_), .C(mai_mai_n93_), .Y(mai_mai_n525_));
  NA2        m0497(.A(mai_mai_n229_), .B(mai_mai_n106_), .Y(mai_mai_n526_));
  AOI210     m0498(.A0(mai_mai_n526_), .A1(mai_mai_n180_), .B0(mai_mai_n522_), .Y(mai_mai_n527_));
  AOI210     m0499(.A0(mai_mai_n364_), .A1(mai_mai_n35_), .B0(mai_mai_n486_), .Y(mai_mai_n528_));
  NOi31      m0500(.An(mai_mai_n525_), .B(mai_mai_n528_), .C(mai_mai_n527_), .Y(mai_mai_n529_));
  AN2        m0501(.A(mai_mai_n290_), .B(mai_mai_n165_), .Y(mai_mai_n530_));
  NA3        m0502(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n531_));
  NO2        m0503(.A(mai_mai_n531_), .B(mai_mai_n446_), .Y(mai_mai_n532_));
  NO2        m0504(.A(mai_mai_n532_), .B(mai_mai_n297_), .Y(mai_mai_n533_));
  NAi41      m0505(.An(mai_mai_n530_), .B(mai_mai_n533_), .C(mai_mai_n529_), .D(mai_mai_n524_), .Y(mai_mai_n534_));
  NO4        m0506(.A(mai_mai_n534_), .B(mai_mai_n521_), .C(mai_mai_n517_), .D(mai_mai_n513_), .Y(mai_mai_n535_));
  NA4        m0507(.A(mai_mai_n535_), .B(mai_mai_n504_), .C(mai_mai_n472_), .D(mai_mai_n441_), .Y(mai11));
  NO2        m0508(.A(mai_mai_n68_), .B(f), .Y(mai_mai_n537_));
  NA2        m0509(.A(j), .B(m), .Y(mai_mai_n538_));
  NAi31      m0510(.An(i), .B(m), .C(l), .Y(mai_mai_n539_));
  NA3        m0511(.A(m), .B(k), .C(j), .Y(mai_mai_n540_));
  OAI220     m0512(.A0(mai_mai_n540_), .A1(mai_mai_n128_), .B0(mai_mai_n539_), .B1(mai_mai_n538_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n541_), .B(mai_mai_n537_), .Y(mai_mai_n542_));
  NOi32      m0514(.An(e), .Bn(b), .C(f), .Y(mai_mai_n543_));
  NA2        m0515(.A(mai_mai_n263_), .B(mai_mai_n111_), .Y(mai_mai_n544_));
  NA2        m0516(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n545_));
  NO2        m0517(.A(mai_mai_n545_), .B(mai_mai_n303_), .Y(mai_mai_n546_));
  NAi31      m0518(.An(d), .B(e), .C(a), .Y(mai_mai_n547_));
  NO2        m0519(.A(mai_mai_n547_), .B(n), .Y(mai_mai_n548_));
  AOI220     m0520(.A0(mai_mai_n548_), .A1(mai_mai_n98_), .B0(mai_mai_n546_), .B1(mai_mai_n543_), .Y(mai_mai_n549_));
  NAi41      m0521(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n550_));
  AN2        m0522(.A(mai_mai_n550_), .B(mai_mai_n377_), .Y(mai_mai_n551_));
  AOI210     m0523(.A0(mai_mai_n551_), .A1(mai_mai_n403_), .B0(mai_mai_n274_), .Y(mai_mai_n552_));
  NA2        m0524(.A(j), .B(i), .Y(mai_mai_n553_));
  NAi31      m0525(.An(n), .B(m), .C(k), .Y(mai_mai_n554_));
  NO2        m0526(.A(mai_mai_n554_), .B(mai_mai_n553_), .Y(mai_mai_n555_));
  NO4        m0527(.A(n), .B(d), .C(mai_mai_n114_), .D(a), .Y(mai_mai_n556_));
  OR2        m0528(.A(n), .B(c), .Y(mai_mai_n557_));
  NO2        m0529(.A(mai_mai_n557_), .B(mai_mai_n148_), .Y(mai_mai_n558_));
  NO2        m0530(.A(mai_mai_n558_), .B(mai_mai_n556_), .Y(mai_mai_n559_));
  NOi32      m0531(.An(m), .Bn(f), .C(i), .Y(mai_mai_n560_));
  AOI220     m0532(.A0(mai_mai_n560_), .A1(mai_mai_n96_), .B0(mai_mai_n541_), .B1(f), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n278_), .B(mai_mai_n49_), .Y(mai_mai_n562_));
  NO2        m0534(.A(mai_mai_n561_), .B(mai_mai_n559_), .Y(mai_mai_n563_));
  AOI210     m0535(.A0(mai_mai_n555_), .A1(mai_mai_n552_), .B0(mai_mai_n563_), .Y(mai_mai_n564_));
  NA2        m0536(.A(mai_mai_n138_), .B(mai_mai_n34_), .Y(mai_mai_n565_));
  OAI220     m0537(.A0(mai_mai_n565_), .A1(m), .B0(mai_mai_n545_), .B1(mai_mai_n235_), .Y(mai_mai_n566_));
  NOi41      m0538(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n567_));
  NAi32      m0539(.An(e), .Bn(b), .C(c), .Y(mai_mai_n568_));
  OR2        m0540(.A(mai_mai_n568_), .B(mai_mai_n80_), .Y(mai_mai_n569_));
  AN2        m0541(.A(mai_mai_n341_), .B(mai_mai_n320_), .Y(mai_mai_n570_));
  NA2        m0542(.A(mai_mai_n570_), .B(mai_mai_n569_), .Y(mai_mai_n571_));
  OA210      m0543(.A0(mai_mai_n571_), .A1(mai_mai_n567_), .B0(mai_mai_n566_), .Y(mai_mai_n572_));
  OAI220     m0544(.A0(mai_mai_n405_), .A1(mai_mai_n404_), .B0(mai_mai_n539_), .B1(mai_mai_n538_), .Y(mai_mai_n573_));
  NAi31      m0545(.An(d), .B(c), .C(a), .Y(mai_mai_n574_));
  NO2        m0546(.A(mai_mai_n574_), .B(n), .Y(mai_mai_n575_));
  NA3        m0547(.A(mai_mai_n575_), .B(mai_mai_n573_), .C(e), .Y(mai_mai_n576_));
  NO3        m0548(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n215_), .Y(mai_mai_n577_));
  NO2        m0549(.A(mai_mai_n232_), .B(mai_mai_n108_), .Y(mai_mai_n578_));
  OAI210     m0550(.A0(mai_mai_n577_), .A1(mai_mai_n406_), .B0(mai_mai_n578_), .Y(mai_mai_n579_));
  NA2        m0551(.A(mai_mai_n579_), .B(mai_mai_n576_), .Y(mai_mai_n580_));
  NO2        m0552(.A(mai_mai_n280_), .B(n), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n436_), .B(mai_mai_n581_), .Y(mai_mai_n582_));
  NA2        m0554(.A(mai_mai_n573_), .B(f), .Y(mai_mai_n583_));
  NAi32      m0555(.An(d), .Bn(a), .C(b), .Y(mai_mai_n584_));
  NO2        m0556(.A(mai_mai_n584_), .B(mai_mai_n49_), .Y(mai_mai_n585_));
  NA2        m0557(.A(h), .B(f), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n586_), .B(mai_mai_n91_), .Y(mai_mai_n587_));
  NO3        m0559(.A(mai_mai_n176_), .B(mai_mai_n173_), .C(m), .Y(mai_mai_n588_));
  AOI220     m0560(.A0(mai_mai_n588_), .A1(mai_mai_n58_), .B0(mai_mai_n587_), .B1(mai_mai_n585_), .Y(mai_mai_n589_));
  OAI210     m0561(.A0(mai_mai_n583_), .A1(mai_mai_n582_), .B0(mai_mai_n589_), .Y(mai_mai_n590_));
  AN3        m0562(.A(j), .B(h), .C(m), .Y(mai_mai_n591_));
  NO2        m0563(.A(mai_mai_n145_), .B(c), .Y(mai_mai_n592_));
  NA3        m0564(.A(mai_mai_n592_), .B(mai_mai_n591_), .C(mai_mai_n467_), .Y(mai_mai_n593_));
  NA3        m0565(.A(f), .B(d), .C(b), .Y(mai_mai_n594_));
  NO4        m0566(.A(mai_mai_n594_), .B(mai_mai_n176_), .C(mai_mai_n173_), .D(m), .Y(mai_mai_n595_));
  NAi21      m0567(.An(mai_mai_n595_), .B(mai_mai_n593_), .Y(mai_mai_n596_));
  NO4        m0568(.A(mai_mai_n596_), .B(mai_mai_n590_), .C(mai_mai_n580_), .D(mai_mai_n572_), .Y(mai_mai_n597_));
  AN4        m0569(.A(mai_mai_n597_), .B(mai_mai_n564_), .C(mai_mai_n549_), .D(mai_mai_n542_), .Y(mai_mai_n598_));
  INV        m0570(.A(k), .Y(mai_mai_n599_));
  NA3        m0571(.A(l), .B(mai_mai_n599_), .C(i), .Y(mai_mai_n600_));
  INV        m0572(.A(mai_mai_n600_), .Y(mai_mai_n601_));
  NA4        m0573(.A(mai_mai_n402_), .B(mai_mai_n425_), .C(mai_mai_n181_), .D(mai_mai_n111_), .Y(mai_mai_n602_));
  NAi32      m0574(.An(h), .Bn(f), .C(m), .Y(mai_mai_n603_));
  NAi41      m0575(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n604_));
  OAI210     m0576(.A0(mai_mai_n547_), .A1(n), .B0(mai_mai_n604_), .Y(mai_mai_n605_));
  NA2        m0577(.A(mai_mai_n605_), .B(m), .Y(mai_mai_n606_));
  NAi31      m0578(.An(h), .B(m), .C(f), .Y(mai_mai_n607_));
  OR3        m0579(.A(mai_mai_n607_), .B(mai_mai_n280_), .C(mai_mai_n49_), .Y(mai_mai_n608_));
  NA4        m0580(.A(mai_mai_n425_), .B(mai_mai_n118_), .C(mai_mai_n111_), .D(e), .Y(mai_mai_n609_));
  AN2        m0581(.A(mai_mai_n609_), .B(mai_mai_n608_), .Y(mai_mai_n610_));
  OA210      m0582(.A0(mai_mai_n606_), .A1(mai_mai_n603_), .B0(mai_mai_n610_), .Y(mai_mai_n611_));
  NO3        m0583(.A(mai_mai_n603_), .B(mai_mai_n68_), .C(mai_mai_n69_), .Y(mai_mai_n612_));
  NO4        m0584(.A(mai_mai_n607_), .B(mai_mai_n557_), .C(mai_mai_n148_), .D(mai_mai_n69_), .Y(mai_mai_n613_));
  OR2        m0585(.A(mai_mai_n613_), .B(mai_mai_n612_), .Y(mai_mai_n614_));
  NAi31      m0586(.An(mai_mai_n614_), .B(mai_mai_n611_), .C(mai_mai_n602_), .Y(mai_mai_n615_));
  NAi31      m0587(.An(f), .B(h), .C(m), .Y(mai_mai_n616_));
  NOi32      m0588(.An(b), .Bn(a), .C(c), .Y(mai_mai_n617_));
  NOi32      m0589(.An(d), .Bn(a), .C(e), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n618_), .B(mai_mai_n111_), .Y(mai_mai_n619_));
  NO2        m0591(.A(n), .B(c), .Y(mai_mai_n620_));
  NA3        m0592(.A(mai_mai_n620_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n621_));
  NAi32      m0593(.An(n), .Bn(f), .C(m), .Y(mai_mai_n622_));
  NA3        m0594(.A(mai_mai_n622_), .B(mai_mai_n621_), .C(mai_mai_n619_), .Y(mai_mai_n623_));
  NOi32      m0595(.An(e), .Bn(a), .C(d), .Y(mai_mai_n624_));
  AOI210     m0596(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n624_), .Y(mai_mai_n625_));
  AOI210     m0597(.A0(mai_mai_n625_), .A1(mai_mai_n214_), .B0(mai_mai_n565_), .Y(mai_mai_n626_));
  NA2        m0598(.A(mai_mai_n626_), .B(mai_mai_n623_), .Y(mai_mai_n627_));
  OAI210     m0599(.A0(mai_mai_n252_), .A1(mai_mai_n83_), .B0(mai_mai_n627_), .Y(mai_mai_n628_));
  AOI210     m0600(.A0(mai_mai_n615_), .A1(mai_mai_n601_), .B0(mai_mai_n628_), .Y(mai_mai_n629_));
  NO3        m0601(.A(mai_mai_n318_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n630_));
  NA3        m0602(.A(mai_mai_n522_), .B(mai_mai_n171_), .C(mai_mai_n170_), .Y(mai_mai_n631_));
  NA2        m0603(.A(mai_mai_n469_), .B(mai_mai_n232_), .Y(mai_mai_n632_));
  OR2        m0604(.A(mai_mai_n632_), .B(mai_mai_n631_), .Y(mai_mai_n633_));
  NA2        m0605(.A(mai_mai_n70_), .B(mai_mai_n111_), .Y(mai_mai_n634_));
  NO2        m0606(.A(mai_mai_n634_), .B(mai_mai_n45_), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n633_), .B(mai_mai_n630_), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n636_), .B(mai_mai_n83_), .Y(mai_mai_n637_));
  NA3        m0609(.A(mai_mai_n567_), .B(mai_mai_n343_), .C(mai_mai_n46_), .Y(mai_mai_n638_));
  NOi32      m0610(.An(e), .Bn(c), .C(f), .Y(mai_mai_n639_));
  NOi21      m0611(.An(f), .B(m), .Y(mai_mai_n640_));
  NO2        m0612(.A(mai_mai_n640_), .B(mai_mai_n212_), .Y(mai_mai_n641_));
  AOI220     m0613(.A0(mai_mai_n641_), .A1(mai_mai_n399_), .B0(mai_mai_n639_), .B1(mai_mai_n175_), .Y(mai_mai_n642_));
  NA3        m0614(.A(mai_mai_n642_), .B(mai_mai_n638_), .C(mai_mai_n178_), .Y(mai_mai_n643_));
  AOI210     m0615(.A0(mai_mai_n551_), .A1(mai_mai_n403_), .B0(mai_mai_n302_), .Y(mai_mai_n644_));
  NAi21      m0616(.An(k), .B(h), .Y(mai_mai_n645_));
  NO2        m0617(.A(mai_mai_n645_), .B(mai_mai_n265_), .Y(mai_mai_n646_));
  NA2        m0618(.A(mai_mai_n646_), .B(j), .Y(mai_mai_n647_));
  OR2        m0619(.A(mai_mai_n647_), .B(mai_mai_n606_), .Y(mai_mai_n648_));
  NOi31      m0620(.An(m), .B(n), .C(k), .Y(mai_mai_n649_));
  NA2        m0621(.A(j), .B(mai_mai_n649_), .Y(mai_mai_n650_));
  AOI210     m0622(.A0(mai_mai_n403_), .A1(mai_mai_n377_), .B0(mai_mai_n302_), .Y(mai_mai_n651_));
  NAi21      m0623(.An(mai_mai_n650_), .B(mai_mai_n651_), .Y(mai_mai_n652_));
  NO2        m0624(.A(mai_mai_n280_), .B(mai_mai_n49_), .Y(mai_mai_n653_));
  NO2        m0625(.A(mai_mai_n547_), .B(mai_mai_n49_), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n653_), .B(mai_mai_n587_), .Y(mai_mai_n655_));
  NA3        m0627(.A(mai_mai_n655_), .B(mai_mai_n652_), .C(mai_mai_n648_), .Y(mai_mai_n656_));
  NA2        m0628(.A(mai_mai_n106_), .B(mai_mai_n36_), .Y(mai_mai_n657_));
  NO2        m0629(.A(k), .B(mai_mai_n215_), .Y(mai_mai_n658_));
  NO2        m0630(.A(mai_mai_n543_), .B(mai_mai_n366_), .Y(mai_mai_n659_));
  NO2        m0631(.A(mai_mai_n659_), .B(n), .Y(mai_mai_n660_));
  NAi31      m0632(.An(mai_mai_n657_), .B(mai_mai_n660_), .C(mai_mai_n658_), .Y(mai_mai_n661_));
  NO2        m0633(.A(mai_mai_n545_), .B(mai_mai_n176_), .Y(mai_mai_n662_));
  NA3        m0634(.A(mai_mai_n568_), .B(mai_mai_n273_), .C(mai_mai_n143_), .Y(mai_mai_n663_));
  NA2        m0635(.A(mai_mai_n518_), .B(mai_mai_n159_), .Y(mai_mai_n664_));
  NO3        m0636(.A(mai_mai_n400_), .B(mai_mai_n664_), .C(mai_mai_n83_), .Y(mai_mai_n665_));
  AOI210     m0637(.A0(mai_mai_n663_), .A1(mai_mai_n662_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  AN3        m0638(.A(f), .B(d), .C(b), .Y(mai_mai_n667_));
  OAI210     m0639(.A0(mai_mai_n667_), .A1(mai_mai_n127_), .B0(n), .Y(mai_mai_n668_));
  NA3        m0640(.A(mai_mai_n518_), .B(mai_mai_n159_), .C(mai_mai_n215_), .Y(mai_mai_n669_));
  AOI210     m0641(.A0(mai_mai_n668_), .A1(mai_mai_n234_), .B0(mai_mai_n669_), .Y(mai_mai_n670_));
  NAi31      m0642(.An(m), .B(n), .C(k), .Y(mai_mai_n671_));
  OR2        m0643(.A(mai_mai_n132_), .B(mai_mai_n61_), .Y(mai_mai_n672_));
  OAI210     m0644(.A0(mai_mai_n672_), .A1(mai_mai_n671_), .B0(mai_mai_n254_), .Y(mai_mai_n673_));
  OAI210     m0645(.A0(mai_mai_n673_), .A1(mai_mai_n670_), .B0(j), .Y(mai_mai_n674_));
  NA3        m0646(.A(mai_mai_n674_), .B(mai_mai_n666_), .C(mai_mai_n661_), .Y(mai_mai_n675_));
  NO4        m0647(.A(mai_mai_n675_), .B(mai_mai_n656_), .C(mai_mai_n643_), .D(mai_mai_n637_), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n387_), .B(mai_mai_n162_), .Y(mai_mai_n677_));
  NAi31      m0649(.An(m), .B(h), .C(f), .Y(mai_mai_n678_));
  OR3        m0650(.A(mai_mai_n678_), .B(mai_mai_n280_), .C(n), .Y(mai_mai_n679_));
  OA210      m0651(.A0(mai_mai_n547_), .A1(n), .B0(mai_mai_n604_), .Y(mai_mai_n680_));
  NA3        m0652(.A(mai_mai_n423_), .B(mai_mai_n118_), .C(mai_mai_n80_), .Y(mai_mai_n681_));
  OAI210     m0653(.A0(mai_mai_n680_), .A1(mai_mai_n87_), .B0(mai_mai_n681_), .Y(mai_mai_n682_));
  NOi21      m0654(.An(mai_mai_n679_), .B(mai_mai_n682_), .Y(mai_mai_n683_));
  AOI210     m0655(.A0(mai_mai_n683_), .A1(mai_mai_n677_), .B0(mai_mai_n540_), .Y(mai_mai_n684_));
  NO3        m0656(.A(m), .B(mai_mai_n214_), .C(mai_mai_n56_), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n526_), .B(mai_mai_n83_), .Y(mai_mai_n686_));
  OAI210     m0658(.A0(mai_mai_n686_), .A1(mai_mai_n399_), .B0(mai_mai_n685_), .Y(mai_mai_n687_));
  OR2        m0659(.A(mai_mai_n68_), .B(mai_mai_n69_), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n617_), .B(mai_mai_n345_), .Y(mai_mai_n689_));
  OA220      m0661(.A0(mai_mai_n650_), .A1(mai_mai_n689_), .B0(mai_mai_n647_), .B1(mai_mai_n688_), .Y(mai_mai_n690_));
  NA3        m0662(.A(mai_mai_n537_), .B(mai_mai_n96_), .C(mai_mai_n95_), .Y(mai_mai_n691_));
  AN2        m0663(.A(h), .B(f), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n692_), .B(mai_mai_n37_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n96_), .B(mai_mai_n46_), .Y(mai_mai_n694_));
  OAI220     m0666(.A0(mai_mai_n694_), .A1(mai_mai_n334_), .B0(mai_mai_n693_), .B1(mai_mai_n474_), .Y(mai_mai_n695_));
  AOI210     m0667(.A0(mai_mai_n584_), .A1(mai_mai_n435_), .B0(mai_mai_n49_), .Y(mai_mai_n696_));
  OAI220     m0668(.A0(mai_mai_n607_), .A1(mai_mai_n600_), .B0(mai_mai_n327_), .B1(mai_mai_n538_), .Y(mai_mai_n697_));
  AOI210     m0669(.A0(mai_mai_n697_), .A1(mai_mai_n696_), .B0(mai_mai_n695_), .Y(mai_mai_n698_));
  NA4        m0670(.A(mai_mai_n698_), .B(mai_mai_n691_), .C(mai_mai_n690_), .D(mai_mai_n687_), .Y(mai_mai_n699_));
  NO2        m0671(.A(mai_mai_n256_), .B(f), .Y(mai_mai_n700_));
  NO2        m0672(.A(mai_mai_n640_), .B(mai_mai_n61_), .Y(mai_mai_n701_));
  NO3        m0673(.A(mai_mai_n701_), .B(mai_mai_n700_), .C(mai_mai_n34_), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n330_), .B(mai_mai_n138_), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n129_), .B(mai_mai_n49_), .Y(mai_mai_n704_));
  AOI220     m0676(.A0(mai_mai_n704_), .A1(mai_mai_n543_), .B0(mai_mai_n366_), .B1(mai_mai_n111_), .Y(mai_mai_n705_));
  OA220      m0677(.A0(mai_mai_n705_), .A1(mai_mai_n565_), .B0(mai_mai_n364_), .B1(mai_mai_n109_), .Y(mai_mai_n706_));
  OAI210     m0678(.A0(mai_mai_n703_), .A1(mai_mai_n702_), .B0(mai_mai_n706_), .Y(mai_mai_n707_));
  NO3        m0679(.A(mai_mai_n410_), .B(mai_mai_n192_), .C(mai_mai_n191_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n708_), .B(mai_mai_n232_), .Y(mai_mai_n709_));
  NA3        m0681(.A(mai_mai_n709_), .B(mai_mai_n258_), .C(j), .Y(mai_mai_n710_));
  NO3        m0682(.A(mai_mai_n469_), .B(mai_mai_n173_), .C(i), .Y(mai_mai_n711_));
  NA2        m0683(.A(mai_mai_n473_), .B(mai_mai_n80_), .Y(mai_mai_n712_));
  NO4        m0684(.A(mai_mai_n540_), .B(mai_mai_n712_), .C(mai_mai_n128_), .D(mai_mai_n214_), .Y(mai_mai_n713_));
  INV        m0685(.A(mai_mai_n713_), .Y(mai_mai_n714_));
  NA4        m0686(.A(mai_mai_n714_), .B(mai_mai_n710_), .C(mai_mai_n525_), .D(mai_mai_n408_), .Y(mai_mai_n715_));
  NO4        m0687(.A(mai_mai_n715_), .B(mai_mai_n707_), .C(mai_mai_n699_), .D(mai_mai_n684_), .Y(mai_mai_n716_));
  NA4        m0688(.A(mai_mai_n716_), .B(mai_mai_n676_), .C(mai_mai_n629_), .D(mai_mai_n598_), .Y(mai08));
  NO2        m0689(.A(k), .B(h), .Y(mai_mai_n718_));
  AO210      m0690(.A0(mai_mai_n256_), .A1(mai_mai_n459_), .B0(mai_mai_n718_), .Y(mai_mai_n719_));
  NO2        m0691(.A(mai_mai_n719_), .B(mai_mai_n300_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n639_), .B(mai_mai_n80_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n721_), .B(mai_mai_n469_), .Y(mai_mai_n722_));
  AOI210     m0694(.A0(mai_mai_n722_), .A1(mai_mai_n720_), .B0(mai_mai_n501_), .Y(mai_mai_n723_));
  NA2        m0695(.A(mai_mai_n80_), .B(mai_mai_n108_), .Y(mai_mai_n724_));
  NO2        m0696(.A(mai_mai_n724_), .B(mai_mai_n57_), .Y(mai_mai_n725_));
  NO4        m0697(.A(mai_mai_n384_), .B(mai_mai_n110_), .C(j), .D(mai_mai_n215_), .Y(mai_mai_n726_));
  OAI210     m0698(.A0(mai_mai_n594_), .A1(mai_mai_n80_), .B0(mai_mai_n234_), .Y(mai_mai_n727_));
  AOI220     m0699(.A0(mai_mai_n727_), .A1(mai_mai_n351_), .B0(mai_mai_n726_), .B1(mai_mai_n725_), .Y(mai_mai_n728_));
  AOI210     m0700(.A0(mai_mai_n594_), .A1(mai_mai_n155_), .B0(mai_mai_n80_), .Y(mai_mai_n729_));
  NA4        m0701(.A(mai_mai_n217_), .B(mai_mai_n138_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n730_));
  AN2        m0702(.A(l), .B(k), .Y(mai_mai_n731_));
  NA4        m0703(.A(mai_mai_n731_), .B(mai_mai_n106_), .C(mai_mai_n69_), .D(mai_mai_n215_), .Y(mai_mai_n732_));
  OAI210     m0704(.A0(mai_mai_n730_), .A1(m), .B0(mai_mai_n732_), .Y(mai_mai_n733_));
  NA2        m0705(.A(mai_mai_n733_), .B(mai_mai_n729_), .Y(mai_mai_n734_));
  NA4        m0706(.A(mai_mai_n734_), .B(mai_mai_n728_), .C(mai_mai_n723_), .D(mai_mai_n353_), .Y(mai_mai_n735_));
  AN2        m0707(.A(mai_mai_n548_), .B(mai_mai_n92_), .Y(mai_mai_n736_));
  NO4        m0708(.A(mai_mai_n173_), .B(mai_mai_n398_), .C(mai_mai_n110_), .D(m), .Y(mai_mai_n737_));
  AOI210     m0709(.A0(mai_mai_n737_), .A1(mai_mai_n727_), .B0(mai_mai_n532_), .Y(mai_mai_n738_));
  NO2        m0710(.A(mai_mai_n38_), .B(mai_mai_n214_), .Y(mai_mai_n739_));
  AOI220     m0711(.A0(mai_mai_n641_), .A1(mai_mai_n350_), .B0(mai_mai_n739_), .B1(mai_mai_n581_), .Y(mai_mai_n740_));
  NAi31      m0712(.An(mai_mai_n736_), .B(mai_mai_n740_), .C(mai_mai_n738_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n551_), .B(mai_mai_n35_), .Y(mai_mai_n742_));
  OAI210     m0714(.A0(mai_mai_n568_), .A1(mai_mai_n47_), .B0(mai_mai_n672_), .Y(mai_mai_n743_));
  NO2        m0715(.A(mai_mai_n493_), .B(mai_mai_n129_), .Y(mai_mai_n744_));
  AOI210     m0716(.A0(mai_mai_n744_), .A1(mai_mai_n743_), .B0(mai_mai_n742_), .Y(mai_mai_n745_));
  NO3        m0717(.A(mai_mai_n318_), .B(mai_mai_n128_), .C(mai_mai_n41_), .Y(mai_mai_n746_));
  NAi21      m0718(.An(mai_mai_n746_), .B(mai_mai_n732_), .Y(mai_mai_n747_));
  NA2        m0719(.A(mai_mai_n719_), .B(mai_mai_n133_), .Y(mai_mai_n748_));
  AOI220     m0720(.A0(mai_mai_n748_), .A1(mai_mai_n409_), .B0(mai_mai_n747_), .B1(mai_mai_n72_), .Y(mai_mai_n749_));
  OAI210     m0721(.A0(mai_mai_n745_), .A1(mai_mai_n83_), .B0(mai_mai_n749_), .Y(mai_mai_n750_));
  NA2        m0722(.A(mai_mai_n366_), .B(mai_mai_n43_), .Y(mai_mai_n751_));
  NA3        m0723(.A(mai_mai_n709_), .B(mai_mai_n336_), .C(mai_mai_n390_), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n731_), .B(mai_mai_n222_), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n753_), .B(mai_mai_n329_), .Y(mai_mai_n754_));
  AOI210     m0726(.A0(mai_mai_n754_), .A1(mai_mai_n700_), .B0(mai_mai_n500_), .Y(mai_mai_n755_));
  NA3        m0727(.A(m), .B(l), .C(k), .Y(mai_mai_n756_));
  AOI210     m0728(.A0(mai_mai_n681_), .A1(mai_mai_n679_), .B0(mai_mai_n756_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n550_), .B(mai_mai_n274_), .Y(mai_mai_n758_));
  NOi21      m0730(.An(mai_mai_n758_), .B(mai_mai_n544_), .Y(mai_mai_n759_));
  NA4        m0731(.A(mai_mai_n111_), .B(l), .C(k), .D(mai_mai_n83_), .Y(mai_mai_n760_));
  NA3        m0732(.A(mai_mai_n118_), .B(mai_mai_n418_), .C(i), .Y(mai_mai_n761_));
  NO2        m0733(.A(mai_mai_n761_), .B(mai_mai_n760_), .Y(mai_mai_n762_));
  NO3        m0734(.A(mai_mai_n762_), .B(mai_mai_n759_), .C(mai_mai_n757_), .Y(mai_mai_n763_));
  NA4        m0735(.A(mai_mai_n763_), .B(mai_mai_n755_), .C(mai_mai_n752_), .D(mai_mai_n751_), .Y(mai_mai_n764_));
  NO4        m0736(.A(mai_mai_n764_), .B(mai_mai_n750_), .C(mai_mai_n741_), .D(mai_mai_n735_), .Y(mai_mai_n765_));
  NA2        m0737(.A(mai_mai_n641_), .B(mai_mai_n399_), .Y(mai_mai_n766_));
  NOi31      m0738(.An(m), .B(h), .C(f), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n654_), .B(mai_mai_n767_), .Y(mai_mai_n768_));
  AO210      m0740(.A0(mai_mai_n768_), .A1(mai_mai_n608_), .B0(mai_mai_n553_), .Y(mai_mai_n769_));
  NO3        m0741(.A(mai_mai_n403_), .B(mai_mai_n538_), .C(h), .Y(mai_mai_n770_));
  AOI210     m0742(.A0(mai_mai_n770_), .A1(mai_mai_n111_), .B0(mai_mai_n511_), .Y(mai_mai_n771_));
  NA4        m0743(.A(mai_mai_n771_), .B(mai_mai_n769_), .C(mai_mai_n766_), .D(mai_mai_n255_), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n731_), .B(mai_mai_n69_), .Y(mai_mai_n773_));
  NO4        m0745(.A(mai_mai_n708_), .B(mai_mai_n173_), .C(n), .D(i), .Y(mai_mai_n774_));
  NOi21      m0746(.An(h), .B(j), .Y(mai_mai_n775_));
  NA2        m0747(.A(mai_mai_n775_), .B(f), .Y(mai_mai_n776_));
  NO2        m0748(.A(mai_mai_n776_), .B(mai_mai_n249_), .Y(mai_mai_n777_));
  NO3        m0749(.A(mai_mai_n777_), .B(mai_mai_n774_), .C(mai_mai_n711_), .Y(mai_mai_n778_));
  OAI220     m0750(.A0(mai_mai_n778_), .A1(mai_mai_n773_), .B0(mai_mai_n610_), .B1(mai_mai_n62_), .Y(mai_mai_n779_));
  AOI210     m0751(.A0(mai_mai_n772_), .A1(l), .B0(mai_mai_n779_), .Y(mai_mai_n780_));
  NO2        m0752(.A(j), .B(i), .Y(mai_mai_n781_));
  NA3        m0753(.A(mai_mai_n781_), .B(mai_mai_n76_), .C(l), .Y(mai_mai_n782_));
  NA2        m0754(.A(mai_mai_n781_), .B(mai_mai_n33_), .Y(mai_mai_n783_));
  NA2        m0755(.A(mai_mai_n428_), .B(mai_mai_n118_), .Y(mai_mai_n784_));
  OA220      m0756(.A0(mai_mai_n784_), .A1(mai_mai_n783_), .B0(mai_mai_n782_), .B1(mai_mai_n606_), .Y(mai_mai_n785_));
  NO3        m0757(.A(mai_mai_n150_), .B(mai_mai_n49_), .C(mai_mai_n108_), .Y(mai_mai_n786_));
  NO3        m0758(.A(mai_mai_n557_), .B(mai_mai_n148_), .C(mai_mai_n69_), .Y(mai_mai_n787_));
  NO3        m0759(.A(mai_mai_n493_), .B(mai_mai_n447_), .C(j), .Y(mai_mai_n788_));
  OAI210     m0760(.A0(mai_mai_n787_), .A1(mai_mai_n786_), .B0(mai_mai_n788_), .Y(mai_mai_n789_));
  OAI210     m0761(.A0(mai_mai_n768_), .A1(mai_mai_n62_), .B0(mai_mai_n789_), .Y(mai_mai_n790_));
  NA2        m0762(.A(k), .B(j), .Y(mai_mai_n791_));
  NO3        m0763(.A(mai_mai_n300_), .B(mai_mai_n791_), .C(mai_mai_n40_), .Y(mai_mai_n792_));
  AOI210     m0764(.A0(mai_mai_n543_), .A1(n), .B0(mai_mai_n567_), .Y(mai_mai_n793_));
  NA2        m0765(.A(mai_mai_n793_), .B(mai_mai_n570_), .Y(mai_mai_n794_));
  AN3        m0766(.A(mai_mai_n794_), .B(mai_mai_n792_), .C(mai_mai_n95_), .Y(mai_mai_n795_));
  NO3        m0767(.A(mai_mai_n173_), .B(mai_mai_n398_), .C(mai_mai_n110_), .Y(mai_mai_n796_));
  AOI220     m0768(.A0(mai_mai_n796_), .A1(mai_mai_n250_), .B0(mai_mai_n632_), .B1(mai_mai_n311_), .Y(mai_mai_n797_));
  NAi31      m0769(.An(mai_mai_n625_), .B(mai_mai_n89_), .C(mai_mai_n80_), .Y(mai_mai_n798_));
  NA2        m0770(.A(mai_mai_n798_), .B(mai_mai_n797_), .Y(mai_mai_n799_));
  NO2        m0771(.A(mai_mai_n300_), .B(mai_mai_n133_), .Y(mai_mai_n800_));
  AOI220     m0772(.A0(mai_mai_n800_), .A1(mai_mai_n641_), .B0(mai_mai_n746_), .B1(mai_mai_n729_), .Y(mai_mai_n801_));
  NO2        m0773(.A(mai_mai_n756_), .B(mai_mai_n87_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n605_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n607_), .B(mai_mai_n115_), .Y(mai_mai_n804_));
  OAI210     m0776(.A0(mai_mai_n804_), .A1(mai_mai_n788_), .B0(mai_mai_n696_), .Y(mai_mai_n805_));
  NA3        m0777(.A(mai_mai_n805_), .B(mai_mai_n803_), .C(mai_mai_n801_), .Y(mai_mai_n806_));
  OR4        m0778(.A(mai_mai_n806_), .B(mai_mai_n799_), .C(mai_mai_n795_), .D(mai_mai_n790_), .Y(mai_mai_n807_));
  NA3        m0779(.A(mai_mai_n793_), .B(mai_mai_n570_), .C(mai_mai_n569_), .Y(mai_mai_n808_));
  NA4        m0780(.A(mai_mai_n808_), .B(mai_mai_n217_), .C(mai_mai_n459_), .D(mai_mai_n34_), .Y(mai_mai_n809_));
  NO4        m0781(.A(mai_mai_n493_), .B(mai_mai_n442_), .C(j), .D(f), .Y(mai_mai_n810_));
  OAI220     m0782(.A0(mai_mai_n730_), .A1(mai_mai_n721_), .B0(mai_mai_n334_), .B1(mai_mai_n38_), .Y(mai_mai_n811_));
  AOI210     m0783(.A0(mai_mai_n810_), .A1(mai_mai_n262_), .B0(mai_mai_n811_), .Y(mai_mai_n812_));
  NA3        m0784(.A(mai_mai_n560_), .B(mai_mai_n294_), .C(h), .Y(mai_mai_n813_));
  NOi21      m0785(.An(mai_mai_n696_), .B(mai_mai_n813_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n88_), .B(mai_mai_n47_), .Y(mai_mai_n815_));
  OAI220     m0787(.A0(mai_mai_n813_), .A1(mai_mai_n621_), .B0(mai_mai_n782_), .B1(mai_mai_n688_), .Y(mai_mai_n816_));
  AOI210     m0788(.A0(mai_mai_n815_), .A1(mai_mai_n660_), .B0(mai_mai_n816_), .Y(mai_mai_n817_));
  NAi41      m0789(.An(mai_mai_n814_), .B(mai_mai_n817_), .C(mai_mai_n812_), .D(mai_mai_n809_), .Y(mai_mai_n818_));
  OR2        m0790(.A(mai_mai_n802_), .B(mai_mai_n92_), .Y(mai_mai_n819_));
  AOI220     m0791(.A0(mai_mai_n819_), .A1(mai_mai_n240_), .B0(mai_mai_n788_), .B1(mai_mai_n653_), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n680_), .B(mai_mai_n69_), .Y(mai_mai_n821_));
  AOI210     m0793(.A0(mai_mai_n810_), .A1(mai_mai_n821_), .B0(mai_mai_n338_), .Y(mai_mai_n822_));
  OAI210     m0794(.A0(mai_mai_n756_), .A1(mai_mai_n678_), .B0(mai_mai_n531_), .Y(mai_mai_n823_));
  NA3        m0795(.A(mai_mai_n253_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n824_));
  AOI220     m0796(.A0(mai_mai_n620_), .A1(mai_mai_n29_), .B0(mai_mai_n473_), .B1(mai_mai_n80_), .Y(mai_mai_n825_));
  NA2        m0797(.A(mai_mai_n825_), .B(mai_mai_n824_), .Y(mai_mai_n826_));
  NO2        m0798(.A(mai_mai_n813_), .B(mai_mai_n499_), .Y(mai_mai_n827_));
  AOI210     m0799(.A0(mai_mai_n826_), .A1(mai_mai_n823_), .B0(mai_mai_n827_), .Y(mai_mai_n828_));
  NA3        m0800(.A(mai_mai_n828_), .B(mai_mai_n822_), .C(mai_mai_n820_), .Y(mai_mai_n829_));
  NOi41      m0801(.An(mai_mai_n785_), .B(mai_mai_n829_), .C(mai_mai_n818_), .D(mai_mai_n807_), .Y(mai_mai_n830_));
  OR3        m0802(.A(mai_mai_n730_), .B(mai_mai_n234_), .C(m), .Y(mai_mai_n831_));
  NO3        m0803(.A(mai_mai_n344_), .B(mai_mai_n302_), .C(mai_mai_n110_), .Y(mai_mai_n832_));
  NA2        m0804(.A(mai_mai_n832_), .B(mai_mai_n794_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n834_));
  NO3        m0806(.A(mai_mai_n834_), .B(mai_mai_n783_), .C(mai_mai_n280_), .Y(mai_mai_n835_));
  NO3        m0807(.A(mai_mai_n538_), .B(mai_mai_n90_), .C(h), .Y(mai_mai_n836_));
  AOI210     m0808(.A0(mai_mai_n836_), .A1(mai_mai_n725_), .B0(mai_mai_n835_), .Y(mai_mai_n837_));
  NA4        m0809(.A(mai_mai_n837_), .B(mai_mai_n833_), .C(mai_mai_n831_), .D(mai_mai_n411_), .Y(mai_mai_n838_));
  OR2        m0810(.A(mai_mai_n678_), .B(mai_mai_n88_), .Y(mai_mai_n839_));
  NOi31      m0811(.An(b), .B(d), .C(a), .Y(mai_mai_n840_));
  NO2        m0812(.A(mai_mai_n840_), .B(mai_mai_n618_), .Y(mai_mai_n841_));
  NO2        m0813(.A(mai_mai_n841_), .B(n), .Y(mai_mai_n842_));
  NOi21      m0814(.An(mai_mai_n825_), .B(mai_mai_n842_), .Y(mai_mai_n843_));
  OAI220     m0815(.A0(mai_mai_n843_), .A1(mai_mai_n839_), .B0(mai_mai_n813_), .B1(mai_mai_n619_), .Y(mai_mai_n844_));
  NO2        m0816(.A(mai_mai_n568_), .B(mai_mai_n80_), .Y(mai_mai_n845_));
  NO3        m0817(.A(mai_mai_n640_), .B(mai_mai_n329_), .C(mai_mai_n115_), .Y(mai_mai_n846_));
  NOi21      m0818(.An(mai_mai_n846_), .B(mai_mai_n160_), .Y(mai_mai_n847_));
  AOI210     m0819(.A0(mai_mai_n832_), .A1(mai_mai_n845_), .B0(mai_mai_n847_), .Y(mai_mai_n848_));
  OAI210     m0820(.A0(mai_mai_n730_), .A1(mai_mai_n400_), .B0(mai_mai_n848_), .Y(mai_mai_n849_));
  NO2        m0821(.A(mai_mai_n708_), .B(n), .Y(mai_mai_n850_));
  AOI220     m0822(.A0(mai_mai_n800_), .A1(mai_mai_n685_), .B0(mai_mai_n850_), .B1(mai_mai_n720_), .Y(mai_mai_n851_));
  NO2        m0823(.A(mai_mai_n324_), .B(mai_mai_n239_), .Y(mai_mai_n852_));
  OAI210     m0824(.A0(mai_mai_n92_), .A1(mai_mai_n89_), .B0(mai_mai_n852_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n118_), .B(mai_mai_n80_), .Y(mai_mai_n854_));
  AOI210     m0826(.A0(mai_mai_n432_), .A1(mai_mai_n424_), .B0(mai_mai_n854_), .Y(mai_mai_n855_));
  NAi21      m0827(.An(mai_mai_n855_), .B(mai_mai_n853_), .Y(mai_mai_n856_));
  NA2        m0828(.A(mai_mai_n754_), .B(mai_mai_n34_), .Y(mai_mai_n857_));
  NAi21      m0829(.An(mai_mai_n760_), .B(mai_mai_n443_), .Y(mai_mai_n858_));
  NO2        m0830(.A(mai_mai_n274_), .B(i), .Y(mai_mai_n859_));
  NA2        m0831(.A(mai_mai_n737_), .B(mai_mai_n352_), .Y(mai_mai_n860_));
  OAI210     m0832(.A0(mai_mai_n613_), .A1(mai_mai_n612_), .B0(mai_mai_n367_), .Y(mai_mai_n861_));
  AN3        m0833(.A(mai_mai_n861_), .B(mai_mai_n860_), .C(mai_mai_n858_), .Y(mai_mai_n862_));
  NAi41      m0834(.An(mai_mai_n856_), .B(mai_mai_n862_), .C(mai_mai_n857_), .D(mai_mai_n851_), .Y(mai_mai_n863_));
  NO4        m0835(.A(mai_mai_n863_), .B(mai_mai_n849_), .C(mai_mai_n844_), .D(mai_mai_n838_), .Y(mai_mai_n864_));
  NA4        m0836(.A(mai_mai_n864_), .B(mai_mai_n830_), .C(mai_mai_n780_), .D(mai_mai_n765_), .Y(mai09));
  INV        m0837(.A(mai_mai_n119_), .Y(mai_mai_n866_));
  NA2        m0838(.A(f), .B(e), .Y(mai_mai_n867_));
  NO2        m0839(.A(mai_mai_n227_), .B(mai_mai_n110_), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n868_), .B(m), .Y(mai_mai_n869_));
  NO2        m0841(.A(m), .B(mai_mai_n479_), .Y(mai_mai_n870_));
  AOI210     m0842(.A0(mai_mai_n870_), .A1(mai_mai_n869_), .B0(mai_mai_n867_), .Y(mai_mai_n871_));
  NA2        m0843(.A(mai_mai_n453_), .B(e), .Y(mai_mai_n872_));
  NO2        m0844(.A(mai_mai_n872_), .B(mai_mai_n522_), .Y(mai_mai_n873_));
  AOI210     m0845(.A0(mai_mai_n871_), .A1(mai_mai_n866_), .B0(mai_mai_n873_), .Y(mai_mai_n874_));
  NO2        m0846(.A(mai_mai_n204_), .B(mai_mai_n214_), .Y(mai_mai_n875_));
  NA3        m0847(.A(m), .B(l), .C(i), .Y(mai_mai_n876_));
  OAI220     m0848(.A0(mai_mai_n607_), .A1(mai_mai_n876_), .B0(mai_mai_n357_), .B1(mai_mai_n539_), .Y(mai_mai_n877_));
  NA4        m0849(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(m), .D(f), .Y(mai_mai_n878_));
  NAi31      m0850(.An(mai_mai_n877_), .B(mai_mai_n878_), .C(mai_mai_n448_), .Y(mai_mai_n879_));
  OA210      m0851(.A0(mai_mai_n879_), .A1(mai_mai_n875_), .B0(mai_mai_n581_), .Y(mai_mai_n880_));
  NA3        m0852(.A(mai_mai_n839_), .B(mai_mai_n583_), .C(mai_mai_n531_), .Y(mai_mai_n881_));
  OA210      m0853(.A0(mai_mai_n881_), .A1(mai_mai_n880_), .B0(mai_mai_n842_), .Y(mai_mai_n882_));
  INV        m0854(.A(mai_mai_n341_), .Y(mai_mai_n883_));
  NO2        m0855(.A(mai_mai_n124_), .B(mai_mai_n122_), .Y(mai_mai_n884_));
  NOi31      m0856(.An(k), .B(m), .C(l), .Y(mai_mai_n885_));
  NO2        m0857(.A(mai_mai_n343_), .B(mai_mai_n885_), .Y(mai_mai_n886_));
  AOI210     m0858(.A0(mai_mai_n886_), .A1(mai_mai_n884_), .B0(mai_mai_n616_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n824_), .B(mai_mai_n334_), .Y(mai_mai_n888_));
  NA2        m0860(.A(mai_mai_n345_), .B(mai_mai_n347_), .Y(mai_mai_n889_));
  OAI210     m0861(.A0(mai_mai_n204_), .A1(mai_mai_n214_), .B0(mai_mai_n889_), .Y(mai_mai_n890_));
  AOI220     m0862(.A0(mai_mai_n890_), .A1(mai_mai_n888_), .B0(mai_mai_n887_), .B1(mai_mai_n883_), .Y(mai_mai_n891_));
  NA2        m0863(.A(mai_mai_n167_), .B(mai_mai_n112_), .Y(mai_mai_n892_));
  NA3        m0864(.A(mai_mai_n892_), .B(mai_mai_n719_), .C(mai_mai_n133_), .Y(mai_mai_n893_));
  NA3        m0865(.A(mai_mai_n893_), .B(mai_mai_n189_), .C(mai_mai_n31_), .Y(mai_mai_n894_));
  NA4        m0866(.A(mai_mai_n894_), .B(mai_mai_n891_), .C(mai_mai_n642_), .D(mai_mai_n78_), .Y(mai_mai_n895_));
  NO2        m0867(.A(mai_mai_n603_), .B(mai_mai_n507_), .Y(mai_mai_n896_));
  NA2        m0868(.A(mai_mai_n896_), .B(mai_mai_n189_), .Y(mai_mai_n897_));
  NOi21      m0869(.An(f), .B(d), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n898_), .B(m), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n899_), .B(mai_mai_n52_), .Y(mai_mai_n900_));
  NOi32      m0872(.An(m), .Bn(f), .C(d), .Y(mai_mai_n901_));
  NA4        m0873(.A(mai_mai_n901_), .B(mai_mai_n620_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n902_));
  INV        m0874(.A(mai_mai_n902_), .Y(mai_mai_n903_));
  AOI210     m0875(.A0(mai_mai_n900_), .A1(mai_mai_n558_), .B0(mai_mai_n903_), .Y(mai_mai_n904_));
  AN2        m0876(.A(f), .B(d), .Y(mai_mai_n905_));
  NA3        m0877(.A(mai_mai_n484_), .B(mai_mai_n905_), .C(mai_mai_n80_), .Y(mai_mai_n906_));
  NO3        m0878(.A(mai_mai_n906_), .B(mai_mai_n69_), .C(mai_mai_n215_), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n289_), .B(mai_mai_n56_), .Y(mai_mai_n908_));
  INV        m0880(.A(mai_mai_n907_), .Y(mai_mai_n909_));
  NAi41      m0881(.An(mai_mai_n498_), .B(mai_mai_n909_), .C(mai_mai_n904_), .D(mai_mai_n897_), .Y(mai_mai_n910_));
  NO4        m0882(.A(mai_mai_n640_), .B(mai_mai_n129_), .C(mai_mai_n329_), .D(mai_mai_n151_), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n671_), .B(mai_mai_n329_), .Y(mai_mai_n912_));
  AN2        m0884(.A(mai_mai_n912_), .B(mai_mai_n700_), .Y(mai_mai_n913_));
  NO3        m0885(.A(mai_mai_n913_), .B(mai_mai_n911_), .C(mai_mai_n236_), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n618_), .B(mai_mai_n80_), .Y(mai_mai_n915_));
  OAI220     m0887(.A0(mai_mai_n889_), .A1(mai_mai_n915_), .B0(mai_mai_n824_), .B1(mai_mai_n448_), .Y(mai_mai_n916_));
  NA3        m0888(.A(mai_mai_n159_), .B(mai_mai_n106_), .C(mai_mai_n105_), .Y(mai_mai_n917_));
  OAI220     m0889(.A0(mai_mai_n906_), .A1(mai_mai_n437_), .B0(mai_mai_n341_), .B1(mai_mai_n917_), .Y(mai_mai_n918_));
  NOi41      m0890(.An(mai_mai_n225_), .B(mai_mai_n918_), .C(mai_mai_n916_), .D(mai_mai_n309_), .Y(mai_mai_n919_));
  NA2        m0891(.A(c), .B(mai_mai_n114_), .Y(mai_mai_n920_));
  NO2        m0892(.A(mai_mai_n920_), .B(mai_mai_n415_), .Y(mai_mai_n921_));
  NA3        m0893(.A(mai_mai_n921_), .B(mai_mai_n520_), .C(f), .Y(mai_mai_n922_));
  OR2        m0894(.A(mai_mai_n678_), .B(mai_mai_n554_), .Y(mai_mai_n923_));
  INV        m0895(.A(mai_mai_n923_), .Y(mai_mai_n924_));
  NA2        m0896(.A(mai_mai_n841_), .B(mai_mai_n109_), .Y(mai_mai_n925_));
  NA2        m0897(.A(mai_mai_n925_), .B(mai_mai_n924_), .Y(mai_mai_n926_));
  NA4        m0898(.A(mai_mai_n926_), .B(mai_mai_n922_), .C(mai_mai_n919_), .D(mai_mai_n914_), .Y(mai_mai_n927_));
  NO4        m0899(.A(mai_mai_n927_), .B(mai_mai_n910_), .C(mai_mai_n895_), .D(mai_mai_n882_), .Y(mai_mai_n928_));
  OR2        m0900(.A(mai_mai_n906_), .B(mai_mai_n69_), .Y(mai_mai_n929_));
  INV        m0901(.A(mai_mai_n142_), .Y(mai_mai_n930_));
  OAI210     m0902(.A0(mai_mai_n930_), .A1(mai_mai_n868_), .B0(m), .Y(mai_mai_n931_));
  AOI210     m0903(.A0(mai_mai_n931_), .A1(mai_mai_n295_), .B0(mai_mai_n929_), .Y(mai_mai_n932_));
  AOI210     m0904(.A0(mai_mai_n824_), .A1(mai_mai_n334_), .B0(mai_mai_n878_), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n133_), .B(mai_mai_n129_), .Y(mai_mai_n934_));
  NO2        m0906(.A(mai_mai_n232_), .B(mai_mai_n226_), .Y(mai_mai_n935_));
  AOI220     m0907(.A0(mai_mai_n935_), .A1(mai_mai_n229_), .B0(mai_mai_n307_), .B1(mai_mai_n934_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n437_), .B(mai_mai_n867_), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n937_), .B(mai_mai_n575_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n938_), .B(mai_mai_n936_), .Y(mai_mai_n939_));
  NA2        m0911(.A(e), .B(d), .Y(mai_mai_n940_));
  OAI220     m0912(.A0(mai_mai_n940_), .A1(c), .B0(mai_mai_n324_), .B1(d), .Y(mai_mai_n941_));
  NA3        m0913(.A(mai_mai_n941_), .B(mai_mai_n462_), .C(mai_mai_n518_), .Y(mai_mai_n942_));
  AOI210     m0914(.A0(mai_mai_n526_), .A1(mai_mai_n180_), .B0(mai_mai_n232_), .Y(mai_mai_n943_));
  AOI210     m0915(.A0(mai_mai_n641_), .A1(mai_mai_n350_), .B0(mai_mai_n943_), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n907_), .B(mai_mai_n56_), .Y(mai_mai_n945_));
  NA3        m0917(.A(mai_mai_n166_), .B(mai_mai_n81_), .C(mai_mai_n34_), .Y(mai_mai_n946_));
  NA4        m0918(.A(mai_mai_n946_), .B(mai_mai_n945_), .C(mai_mai_n944_), .D(mai_mai_n942_), .Y(mai_mai_n947_));
  NO4        m0919(.A(mai_mai_n947_), .B(mai_mai_n939_), .C(mai_mai_n933_), .D(mai_mai_n932_), .Y(mai_mai_n948_));
  NA2        m0920(.A(mai_mai_n883_), .B(mai_mai_n31_), .Y(mai_mai_n949_));
  AO210      m0921(.A0(mai_mai_n949_), .A1(mai_mai_n721_), .B0(mai_mai_n218_), .Y(mai_mai_n950_));
  OAI220     m0922(.A0(mai_mai_n640_), .A1(mai_mai_n61_), .B0(mai_mai_n302_), .B1(j), .Y(mai_mai_n951_));
  AOI220     m0923(.A0(mai_mai_n951_), .A1(mai_mai_n912_), .B0(mai_mai_n630_), .B1(mai_mai_n639_), .Y(mai_mai_n952_));
  OAI210     m0924(.A0(mai_mai_n872_), .A1(mai_mai_n170_), .B0(mai_mai_n952_), .Y(mai_mai_n953_));
  INV        m0925(.A(mai_mai_n901_), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n954_), .B(mai_mai_n621_), .Y(mai_mai_n955_));
  AOI210     m0927(.A0(mai_mai_n116_), .A1(mai_mai_n115_), .B0(mai_mai_n263_), .Y(mai_mai_n956_));
  NO2        m0928(.A(mai_mai_n956_), .B(mai_mai_n902_), .Y(mai_mai_n957_));
  AO210      m0929(.A0(mai_mai_n888_), .A1(mai_mai_n877_), .B0(mai_mai_n957_), .Y(mai_mai_n958_));
  NOi31      m0930(.An(mai_mai_n558_), .B(mai_mai_n899_), .C(mai_mai_n295_), .Y(mai_mai_n959_));
  NO4        m0931(.A(mai_mai_n959_), .B(mai_mai_n958_), .C(mai_mai_n955_), .D(mai_mai_n953_), .Y(mai_mai_n960_));
  AO220      m0932(.A0(mai_mai_n462_), .A1(mai_mai_n775_), .B0(mai_mai_n175_), .B1(f), .Y(mai_mai_n961_));
  OAI210     m0933(.A0(mai_mai_n961_), .A1(mai_mai_n465_), .B0(mai_mai_n941_), .Y(mai_mai_n962_));
  NO2        m0934(.A(mai_mai_n447_), .B(mai_mai_n66_), .Y(mai_mai_n963_));
  OAI210     m0935(.A0(mai_mai_n881_), .A1(mai_mai_n963_), .B0(mai_mai_n725_), .Y(mai_mai_n964_));
  AN4        m0936(.A(mai_mai_n964_), .B(mai_mai_n962_), .C(mai_mai_n960_), .D(mai_mai_n950_), .Y(mai_mai_n965_));
  NA4        m0937(.A(mai_mai_n965_), .B(mai_mai_n948_), .C(mai_mai_n928_), .D(mai_mai_n874_), .Y(mai12));
  NO2        m0938(.A(mai_mai_n460_), .B(c), .Y(mai_mai_n967_));
  NO4        m0939(.A(mai_mai_n452_), .B(mai_mai_n256_), .C(mai_mai_n599_), .D(mai_mai_n215_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n968_), .B(mai_mai_n967_), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n558_), .B(mai_mai_n963_), .Y(mai_mai_n970_));
  NO3        m0942(.A(mai_mai_n460_), .B(mai_mai_n80_), .C(mai_mai_n114_), .Y(mai_mai_n971_));
  NO2        m0943(.A(mai_mai_n884_), .B(mai_mai_n357_), .Y(mai_mai_n972_));
  NO2        m0944(.A(mai_mai_n678_), .B(mai_mai_n384_), .Y(mai_mai_n973_));
  AOI220     m0945(.A0(mai_mai_n973_), .A1(mai_mai_n556_), .B0(mai_mai_n972_), .B1(mai_mai_n971_), .Y(mai_mai_n974_));
  NA4        m0946(.A(mai_mai_n974_), .B(mai_mai_n970_), .C(mai_mai_n969_), .D(mai_mai_n451_), .Y(mai_mai_n975_));
  AOI210     m0947(.A0(mai_mai_n235_), .A1(mai_mai_n340_), .B0(mai_mai_n201_), .Y(mai_mai_n976_));
  OR2        m0948(.A(mai_mai_n976_), .B(mai_mai_n968_), .Y(mai_mai_n977_));
  AOI210     m0949(.A0(mai_mai_n337_), .A1(mai_mai_n396_), .B0(mai_mai_n215_), .Y(mai_mai_n978_));
  OAI210     m0950(.A0(mai_mai_n978_), .A1(mai_mai_n977_), .B0(mai_mai_n410_), .Y(mai_mai_n979_));
  NO2        m0951(.A(mai_mai_n657_), .B(mai_mai_n265_), .Y(mai_mai_n980_));
  NO2        m0952(.A(mai_mai_n607_), .B(mai_mai_n876_), .Y(mai_mai_n981_));
  AOI220     m0953(.A0(mai_mai_n981_), .A1(mai_mai_n581_), .B0(mai_mai_n852_), .B1(mai_mai_n980_), .Y(mai_mai_n982_));
  NO2        m0954(.A(mai_mai_n150_), .B(mai_mai_n239_), .Y(mai_mai_n983_));
  NA3        m0955(.A(mai_mai_n983_), .B(mai_mai_n242_), .C(i), .Y(mai_mai_n984_));
  NA3        m0956(.A(mai_mai_n984_), .B(mai_mai_n982_), .C(mai_mai_n979_), .Y(mai_mai_n985_));
  OR2        m0957(.A(mai_mai_n325_), .B(mai_mai_n971_), .Y(mai_mai_n986_));
  NA2        m0958(.A(mai_mai_n986_), .B(mai_mai_n358_), .Y(mai_mai_n987_));
  NO3        m0959(.A(mai_mai_n129_), .B(mai_mai_n151_), .C(mai_mai_n215_), .Y(mai_mai_n988_));
  NA2        m0960(.A(mai_mai_n988_), .B(mai_mai_n543_), .Y(mai_mai_n989_));
  NA4        m0961(.A(mai_mai_n453_), .B(mai_mai_n445_), .C(mai_mai_n181_), .D(m), .Y(mai_mai_n990_));
  NA3        m0962(.A(mai_mai_n990_), .B(mai_mai_n989_), .C(mai_mai_n987_), .Y(mai_mai_n991_));
  NO3        m0963(.A(mai_mai_n683_), .B(mai_mai_n88_), .C(mai_mai_n45_), .Y(mai_mai_n992_));
  NO4        m0964(.A(mai_mai_n992_), .B(mai_mai_n991_), .C(mai_mai_n985_), .D(mai_mai_n975_), .Y(mai_mai_n993_));
  NO2        m0965(.A(mai_mai_n374_), .B(mai_mai_n373_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n604_), .B(mai_mai_n68_), .Y(mai_mai_n995_));
  NA2        m0967(.A(mai_mai_n568_), .B(mai_mai_n143_), .Y(mai_mai_n996_));
  NOi21      m0968(.An(mai_mai_n34_), .B(mai_mai_n671_), .Y(mai_mai_n997_));
  AOI220     m0969(.A0(mai_mai_n997_), .A1(mai_mai_n996_), .B0(mai_mai_n995_), .B1(mai_mai_n994_), .Y(mai_mai_n998_));
  OAI210     m0970(.A0(mai_mai_n254_), .A1(mai_mai_n45_), .B0(mai_mai_n998_), .Y(mai_mai_n999_));
  NO3        m0971(.A(mai_mai_n854_), .B(mai_mai_n85_), .C(mai_mai_n415_), .Y(mai_mai_n1000_));
  NAi21      m0972(.An(mai_mai_n1000_), .B(mai_mai_n322_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(mai_mai_n514_), .B(mai_mai_n302_), .Y(mai_mai_n1002_));
  NO2        m0974(.A(mai_mai_n1002_), .B(mai_mai_n370_), .Y(mai_mai_n1003_));
  NO2        m0975(.A(mai_mai_n1003_), .B(mai_mai_n143_), .Y(mai_mai_n1004_));
  INV        m0976(.A(mai_mai_n371_), .Y(mai_mai_n1005_));
  NO4        m0977(.A(mai_mai_n1005_), .B(mai_mai_n1004_), .C(mai_mai_n1001_), .D(mai_mai_n999_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n350_), .B(m), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n162_), .B(i), .Y(mai_mai_n1008_));
  NA2        m0980(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n1009_));
  OAI220     m0981(.A0(mai_mai_n1009_), .A1(mai_mai_n200_), .B0(mai_mai_n1008_), .B1(mai_mai_n88_), .Y(mai_mai_n1010_));
  AOI210     m0982(.A0(mai_mai_n426_), .A1(mai_mai_n37_), .B0(mai_mai_n1010_), .Y(mai_mai_n1011_));
  NO2        m0983(.A(mai_mai_n143_), .B(mai_mai_n80_), .Y(mai_mai_n1012_));
  OR2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n567_), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n568_), .B(mai_mai_n388_), .Y(mai_mai_n1014_));
  AOI210     m0986(.A0(mai_mai_n1014_), .A1(n), .B0(mai_mai_n1013_), .Y(mai_mai_n1015_));
  OAI220     m0987(.A0(mai_mai_n1015_), .A1(mai_mai_n1007_), .B0(mai_mai_n1011_), .B1(mai_mai_n334_), .Y(mai_mai_n1016_));
  NO2        m0988(.A(mai_mai_n678_), .B(mai_mai_n507_), .Y(mai_mai_n1017_));
  NA3        m0989(.A(mai_mai_n345_), .B(j), .C(i), .Y(mai_mai_n1018_));
  INV        m0990(.A(mai_mai_n1018_), .Y(mai_mai_n1019_));
  OAI220     m0991(.A0(mai_mai_n1019_), .A1(mai_mai_n1017_), .B0(mai_mai_n696_), .B1(mai_mai_n787_), .Y(mai_mai_n1020_));
  NA2        m0992(.A(mai_mai_n624_), .B(mai_mai_n111_), .Y(mai_mai_n1021_));
  NA3        m0993(.A(j), .B(mai_mai_n76_), .C(i), .Y(mai_mai_n1022_));
  OR2        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1021_), .Y(mai_mai_n1023_));
  NA3        m0995(.A(mai_mai_n326_), .B(mai_mai_n116_), .C(m), .Y(mai_mai_n1024_));
  AOI210     m0996(.A0(mai_mai_n693_), .A1(mai_mai_n1024_), .B0(m), .Y(mai_mai_n1025_));
  OAI210     m0997(.A0(mai_mai_n1025_), .A1(mai_mai_n972_), .B0(mai_mai_n325_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n712_), .B(mai_mai_n915_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n878_), .B(mai_mai_n448_), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n223_), .B(mai_mai_n73_), .Y(mai_mai_n1029_));
  NA2        m1001(.A(mai_mai_n1029_), .B(mai_mai_n1022_), .Y(mai_mai_n1030_));
  AOI220     m1002(.A0(mai_mai_n1030_), .A1(mai_mai_n262_), .B0(mai_mai_n1028_), .B1(mai_mai_n1027_), .Y(mai_mai_n1031_));
  NA4        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1026_), .C(mai_mai_n1023_), .D(mai_mai_n1020_), .Y(mai_mai_n1032_));
  NO2        m1004(.A(mai_mai_n384_), .B(mai_mai_n87_), .Y(mai_mai_n1033_));
  OAI210     m1005(.A0(mai_mai_n1033_), .A1(mai_mai_n980_), .B0(mai_mai_n240_), .Y(mai_mai_n1034_));
  NA2        m1006(.A(mai_mai_n682_), .B(mai_mai_n84_), .Y(mai_mai_n1035_));
  NO2        m1007(.A(mai_mai_n468_), .B(mai_mai_n215_), .Y(mai_mai_n1036_));
  AOI220     m1008(.A0(mai_mai_n1036_), .A1(mai_mai_n389_), .B0(mai_mai_n986_), .B1(mai_mai_n219_), .Y(mai_mai_n1037_));
  AOI220     m1009(.A0(mai_mai_n973_), .A1(mai_mai_n983_), .B0(mai_mai_n605_), .B1(mai_mai_n86_), .Y(mai_mai_n1038_));
  NA4        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1037_), .C(mai_mai_n1035_), .D(mai_mai_n1034_), .Y(mai_mai_n1039_));
  OAI210     m1011(.A0(mai_mai_n1028_), .A1(mai_mai_n981_), .B0(mai_mai_n556_), .Y(mai_mai_n1040_));
  AOI210     m1012(.A0(mai_mai_n427_), .A1(mai_mai_n419_), .B0(mai_mai_n854_), .Y(mai_mai_n1041_));
  OAI210     m1013(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n107_), .Y(mai_mai_n1042_));
  AOI210     m1014(.A0(mai_mai_n1042_), .A1(mai_mai_n548_), .B0(mai_mai_n1041_), .Y(mai_mai_n1043_));
  NA2        m1015(.A(mai_mai_n1025_), .B(mai_mai_n971_), .Y(mai_mai_n1044_));
  NO3        m1016(.A(mai_mai_n1547_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n1045_));
  AOI220     m1017(.A0(mai_mai_n1045_), .A1(mai_mai_n644_), .B0(mai_mai_n662_), .B1(mai_mai_n543_), .Y(mai_mai_n1046_));
  NA4        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1044_), .C(mai_mai_n1043_), .D(mai_mai_n1040_), .Y(mai_mai_n1047_));
  NO4        m1019(.A(mai_mai_n1047_), .B(mai_mai_n1039_), .C(mai_mai_n1032_), .D(mai_mai_n1016_), .Y(mai_mai_n1048_));
  NAi31      m1020(.An(mai_mai_n139_), .B(mai_mai_n428_), .C(n), .Y(mai_mai_n1049_));
  NO3        m1021(.A(mai_mai_n122_), .B(mai_mai_n343_), .C(mai_mai_n885_), .Y(mai_mai_n1050_));
  NO2        m1022(.A(mai_mai_n1050_), .B(mai_mai_n1049_), .Y(mai_mai_n1051_));
  NO3        m1023(.A(mai_mai_n274_), .B(mai_mai_n139_), .C(mai_mai_n415_), .Y(mai_mai_n1052_));
  AOI210     m1024(.A0(mai_mai_n1052_), .A1(mai_mai_n508_), .B0(mai_mai_n1051_), .Y(mai_mai_n1053_));
  NA2        m1025(.A(mai_mai_n501_), .B(i), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n1054_), .B(mai_mai_n1053_), .Y(mai_mai_n1055_));
  NA2        m1027(.A(mai_mai_n232_), .B(mai_mai_n171_), .Y(mai_mai_n1056_));
  NO3        m1028(.A(mai_mai_n311_), .B(mai_mai_n453_), .C(mai_mai_n175_), .Y(mai_mai_n1057_));
  NOi31      m1029(.An(mai_mai_n1056_), .B(mai_mai_n1057_), .C(mai_mai_n215_), .Y(mai_mai_n1058_));
  NAi21      m1030(.An(mai_mai_n568_), .B(mai_mai_n1036_), .Y(mai_mai_n1059_));
  NA2        m1031(.A(mai_mai_n490_), .B(m), .Y(mai_mai_n1060_));
  NA2        m1032(.A(mai_mai_n1060_), .B(mai_mai_n1059_), .Y(mai_mai_n1061_));
  OAI220     m1033(.A0(mai_mai_n1049_), .A1(mai_mai_n235_), .B0(mai_mai_n1018_), .B1(mai_mai_n619_), .Y(mai_mai_n1062_));
  NO2        m1034(.A(mai_mai_n679_), .B(mai_mai_n384_), .Y(mai_mai_n1063_));
  NA2        m1035(.A(mai_mai_n976_), .B(mai_mai_n967_), .Y(mai_mai_n1064_));
  NO3        m1036(.A(mai_mai_n557_), .B(mai_mai_n148_), .C(mai_mai_n214_), .Y(mai_mai_n1065_));
  OAI210     m1037(.A0(mai_mai_n1065_), .A1(mai_mai_n537_), .B0(mai_mai_n385_), .Y(mai_mai_n1066_));
  OAI220     m1038(.A0(mai_mai_n973_), .A1(mai_mai_n981_), .B0(mai_mai_n558_), .B1(mai_mai_n436_), .Y(mai_mai_n1067_));
  NA4        m1039(.A(mai_mai_n1067_), .B(mai_mai_n1066_), .C(mai_mai_n1064_), .D(mai_mai_n638_), .Y(mai_mai_n1068_));
  OAI210     m1040(.A0(mai_mai_n976_), .A1(mai_mai_n968_), .B0(mai_mai_n1056_), .Y(mai_mai_n1069_));
  NA3        m1041(.A(mai_mai_n1014_), .B(mai_mai_n495_), .C(mai_mai_n46_), .Y(mai_mai_n1070_));
  AOI210     m1042(.A0(mai_mai_n387_), .A1(mai_mai_n385_), .B0(mai_mai_n333_), .Y(mai_mai_n1071_));
  NA4        m1043(.A(mai_mai_n1071_), .B(mai_mai_n1070_), .C(mai_mai_n1069_), .D(mai_mai_n275_), .Y(mai_mai_n1072_));
  OR4        m1044(.A(mai_mai_n1072_), .B(mai_mai_n1068_), .C(mai_mai_n1063_), .D(mai_mai_n1062_), .Y(mai_mai_n1073_));
  NO4        m1045(.A(mai_mai_n1073_), .B(mai_mai_n1061_), .C(mai_mai_n1058_), .D(mai_mai_n1055_), .Y(mai_mai_n1074_));
  NA4        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1048_), .C(mai_mai_n1006_), .D(mai_mai_n993_), .Y(mai13));
  AN2        m1047(.A(c), .B(b), .Y(mai_mai_n1076_));
  NA3        m1048(.A(mai_mai_n253_), .B(mai_mai_n1076_), .C(m), .Y(mai_mai_n1077_));
  NA2        m1049(.A(mai_mai_n505_), .B(f), .Y(mai_mai_n1078_));
  NO4        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1077_), .C(j), .D(mai_mai_n600_), .Y(mai_mai_n1079_));
  INV        m1051(.A(mai_mai_n266_), .Y(mai_mai_n1080_));
  NO4        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1078_), .C(mai_mai_n1008_), .D(a), .Y(mai_mai_n1081_));
  NAi32      m1053(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1082_));
  NA2        m1054(.A(mai_mai_n138_), .B(mai_mai_n45_), .Y(mai_mai_n1083_));
  NO4        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1082_), .C(mai_mai_n607_), .D(mai_mai_n310_), .Y(mai_mai_n1084_));
  NA2        m1056(.A(mai_mai_n418_), .B(mai_mai_n214_), .Y(mai_mai_n1085_));
  AN2        m1057(.A(d), .B(c), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n114_), .Y(mai_mai_n1087_));
  NO4        m1059(.A(mai_mai_n1087_), .B(mai_mai_n1085_), .C(mai_mai_n176_), .D(mai_mai_n167_), .Y(mai_mai_n1088_));
  NA2        m1060(.A(mai_mai_n505_), .B(c), .Y(mai_mai_n1089_));
  NO4        m1061(.A(mai_mai_n1083_), .B(mai_mai_n603_), .C(mai_mai_n1089_), .D(mai_mai_n310_), .Y(mai_mai_n1090_));
  OR2        m1062(.A(mai_mai_n1088_), .B(mai_mai_n1090_), .Y(mai_mai_n1091_));
  OR4        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1084_), .C(mai_mai_n1081_), .D(mai_mai_n1079_), .Y(mai_mai_n1092_));
  NAi32      m1064(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1093_));
  NO2        m1065(.A(mai_mai_n1093_), .B(mai_mai_n145_), .Y(mai_mai_n1094_));
  NA2        m1066(.A(mai_mai_n1094_), .B(m), .Y(mai_mai_n1095_));
  OR3        m1067(.A(mai_mai_n226_), .B(mai_mai_n176_), .C(mai_mai_n167_), .Y(mai_mai_n1096_));
  NO2        m1068(.A(mai_mai_n1096_), .B(mai_mai_n1095_), .Y(mai_mai_n1097_));
  NO2        m1069(.A(mai_mai_n1089_), .B(mai_mai_n310_), .Y(mai_mai_n1098_));
  NO2        m1070(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1099_));
  NA2        m1071(.A(mai_mai_n646_), .B(mai_mai_n1099_), .Y(mai_mai_n1100_));
  NOi21      m1072(.An(mai_mai_n1098_), .B(mai_mai_n1100_), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n791_), .B(mai_mai_n110_), .Y(mai_mai_n1102_));
  NOi41      m1074(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1103_));
  NA2        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1102_), .Y(mai_mai_n1104_));
  NO2        m1076(.A(mai_mai_n1104_), .B(mai_mai_n1095_), .Y(mai_mai_n1105_));
  OR3        m1077(.A(e), .B(d), .C(c), .Y(mai_mai_n1106_));
  NA3        m1078(.A(k), .B(j), .C(i), .Y(mai_mai_n1107_));
  NO3        m1079(.A(mai_mai_n1107_), .B(mai_mai_n310_), .C(mai_mai_n87_), .Y(mai_mai_n1108_));
  NOi21      m1080(.An(mai_mai_n1108_), .B(mai_mai_n1106_), .Y(mai_mai_n1109_));
  OR4        m1081(.A(mai_mai_n1109_), .B(mai_mai_n1105_), .C(mai_mai_n1101_), .D(mai_mai_n1097_), .Y(mai_mai_n1110_));
  NA3        m1082(.A(mai_mai_n476_), .B(mai_mai_n336_), .C(mai_mai_n56_), .Y(mai_mai_n1111_));
  NO2        m1083(.A(mai_mai_n1111_), .B(mai_mai_n1100_), .Y(mai_mai_n1112_));
  NO3        m1084(.A(mai_mai_n1111_), .B(mai_mai_n603_), .C(mai_mai_n459_), .Y(mai_mai_n1113_));
  NO2        m1085(.A(f), .B(c), .Y(mai_mai_n1114_));
  NOi21      m1086(.An(mai_mai_n1114_), .B(mai_mai_n452_), .Y(mai_mai_n1115_));
  NA2        m1087(.A(mai_mai_n1115_), .B(mai_mai_n59_), .Y(mai_mai_n1116_));
  NO3        m1088(.A(i), .B(mai_mai_n246_), .C(l), .Y(mai_mai_n1117_));
  NOi31      m1089(.An(mai_mai_n1117_), .B(mai_mai_n1116_), .C(j), .Y(mai_mai_n1118_));
  OR3        m1090(.A(mai_mai_n1118_), .B(mai_mai_n1113_), .C(mai_mai_n1112_), .Y(mai_mai_n1119_));
  OR3        m1091(.A(mai_mai_n1119_), .B(mai_mai_n1110_), .C(mai_mai_n1092_), .Y(mai02));
  OR3        m1092(.A(h), .B(m), .C(f), .Y(mai_mai_n1121_));
  OR3        m1093(.A(n), .B(m), .C(i), .Y(mai_mai_n1122_));
  NO4        m1094(.A(mai_mai_n1122_), .B(mai_mai_n1121_), .C(l), .D(mai_mai_n1106_), .Y(mai_mai_n1123_));
  NOi31      m1095(.An(e), .B(d), .C(c), .Y(mai_mai_n1124_));
  AOI210     m1096(.A0(mai_mai_n1108_), .A1(mai_mai_n1124_), .B0(mai_mai_n1084_), .Y(mai_mai_n1125_));
  AN3        m1097(.A(m), .B(f), .C(c), .Y(mai_mai_n1126_));
  NA3        m1098(.A(mai_mai_n1126_), .B(mai_mai_n476_), .C(h), .Y(mai_mai_n1127_));
  OR2        m1099(.A(mai_mai_n1107_), .B(mai_mai_n310_), .Y(mai_mai_n1128_));
  OR2        m1100(.A(mai_mai_n1128_), .B(mai_mai_n1127_), .Y(mai_mai_n1129_));
  NO3        m1101(.A(mai_mai_n1111_), .B(mai_mai_n1083_), .C(mai_mai_n603_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n1130_), .B(mai_mai_n1097_), .Y(mai_mai_n1131_));
  NA3        m1103(.A(l), .B(k), .C(j), .Y(mai_mai_n1132_));
  NA2        m1104(.A(i), .B(h), .Y(mai_mai_n1133_));
  NO3        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1132_), .C(mai_mai_n129_), .Y(mai_mai_n1134_));
  NO3        m1106(.A(mai_mai_n140_), .B(mai_mai_n287_), .C(mai_mai_n215_), .Y(mai_mai_n1135_));
  AOI210     m1107(.A0(mai_mai_n1135_), .A1(mai_mai_n1134_), .B0(mai_mai_n1101_), .Y(mai_mai_n1136_));
  NA3        m1108(.A(c), .B(b), .C(a), .Y(mai_mai_n1137_));
  NO3        m1109(.A(mai_mai_n1137_), .B(mai_mai_n940_), .C(mai_mai_n214_), .Y(mai_mai_n1138_));
  NO3        m1110(.A(mai_mai_n1107_), .B(mai_mai_n302_), .C(mai_mai_n49_), .Y(mai_mai_n1139_));
  AOI210     m1111(.A0(mai_mai_n1139_), .A1(mai_mai_n1138_), .B0(mai_mai_n1112_), .Y(mai_mai_n1140_));
  AN4        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1136_), .C(mai_mai_n1131_), .D(mai_mai_n1129_), .Y(mai_mai_n1141_));
  NO2        m1113(.A(mai_mai_n1087_), .B(mai_mai_n1085_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n1104_), .B(mai_mai_n1096_), .Y(mai_mai_n1143_));
  AOI210     m1115(.A0(mai_mai_n1143_), .A1(mai_mai_n1142_), .B0(mai_mai_n1079_), .Y(mai_mai_n1144_));
  NAi41      m1116(.An(mai_mai_n1123_), .B(mai_mai_n1144_), .C(mai_mai_n1141_), .D(mai_mai_n1125_), .Y(mai03));
  NO2        m1117(.A(mai_mai_n539_), .B(mai_mai_n616_), .Y(mai_mai_n1146_));
  NA4        m1118(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(m), .D(mai_mai_n214_), .Y(mai_mai_n1147_));
  NA4        m1119(.A(mai_mai_n591_), .B(m), .C(mai_mai_n110_), .D(mai_mai_n214_), .Y(mai_mai_n1148_));
  NA3        m1120(.A(mai_mai_n1148_), .B(mai_mai_n375_), .C(mai_mai_n1147_), .Y(mai_mai_n1149_));
  NO3        m1121(.A(mai_mai_n1149_), .B(mai_mai_n1146_), .C(mai_mai_n1042_), .Y(mai_mai_n1150_));
  NOi41      m1122(.An(mai_mai_n839_), .B(mai_mai_n890_), .C(mai_mai_n879_), .D(mai_mai_n739_), .Y(mai_mai_n1151_));
  OAI220     m1123(.A0(mai_mai_n1151_), .A1(mai_mai_n712_), .B0(mai_mai_n1150_), .B1(mai_mai_n604_), .Y(mai_mai_n1152_));
  NA4        m1124(.A(i), .B(mai_mai_n1124_), .C(mai_mai_n345_), .D(mai_mai_n336_), .Y(mai_mai_n1153_));
  OAI210     m1125(.A0(mai_mai_n854_), .A1(mai_mai_n429_), .B0(mai_mai_n1153_), .Y(mai_mai_n1154_));
  NOi31      m1126(.An(m), .B(n), .C(f), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n1155_), .B(mai_mai_n51_), .Y(mai_mai_n1156_));
  AN2        m1128(.A(e), .B(c), .Y(mai_mai_n1157_));
  NA2        m1129(.A(mai_mai_n1157_), .B(a), .Y(mai_mai_n1158_));
  OAI220     m1130(.A0(mai_mai_n1158_), .A1(mai_mai_n1156_), .B0(mai_mai_n923_), .B1(mai_mai_n435_), .Y(mai_mai_n1159_));
  NA2        m1131(.A(mai_mai_n518_), .B(l), .Y(mai_mai_n1160_));
  NOi31      m1132(.An(mai_mai_n901_), .B(mai_mai_n1077_), .C(mai_mai_n1160_), .Y(mai_mai_n1161_));
  NO4        m1133(.A(mai_mai_n1161_), .B(mai_mai_n1159_), .C(mai_mai_n1154_), .D(mai_mai_n1041_), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n287_), .B(a), .Y(mai_mai_n1163_));
  INV        m1135(.A(mai_mai_n1084_), .Y(mai_mai_n1164_));
  NO2        m1136(.A(mai_mai_n1133_), .B(mai_mai_n493_), .Y(mai_mai_n1165_));
  NO2        m1137(.A(mai_mai_n83_), .B(m), .Y(mai_mai_n1166_));
  AOI210     m1138(.A0(mai_mai_n1166_), .A1(mai_mai_n1165_), .B0(mai_mai_n1117_), .Y(mai_mai_n1167_));
  OR2        m1139(.A(mai_mai_n1167_), .B(mai_mai_n1116_), .Y(mai_mai_n1168_));
  NA3        m1140(.A(mai_mai_n1168_), .B(mai_mai_n1164_), .C(mai_mai_n1162_), .Y(mai_mai_n1169_));
  NO4        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1152_), .C(mai_mai_n856_), .D(mai_mai_n580_), .Y(mai_mai_n1170_));
  NA2        m1142(.A(c), .B(b), .Y(mai_mai_n1171_));
  NO2        m1143(.A(mai_mai_n724_), .B(mai_mai_n1171_), .Y(mai_mai_n1172_));
  OAI210     m1144(.A0(mai_mai_n899_), .A1(mai_mai_n870_), .B0(mai_mai_n422_), .Y(mai_mai_n1173_));
  OAI210     m1145(.A0(mai_mai_n1173_), .A1(mai_mai_n900_), .B0(mai_mai_n1172_), .Y(mai_mai_n1174_));
  NAi21      m1146(.An(mai_mai_n430_), .B(mai_mai_n1172_), .Y(mai_mai_n1175_));
  NA3        m1147(.A(mai_mai_n436_), .B(mai_mai_n573_), .C(f), .Y(mai_mai_n1176_));
  OAI210     m1148(.A0(mai_mai_n562_), .A1(mai_mai_n39_), .B0(mai_mai_n1163_), .Y(mai_mai_n1177_));
  NA3        m1149(.A(mai_mai_n1177_), .B(mai_mai_n1176_), .C(mai_mai_n1175_), .Y(mai_mai_n1178_));
  INV        m1150(.A(m), .Y(mai_mai_n1179_));
  NAi21      m1151(.An(f), .B(d), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n1180_), .B(mai_mai_n1137_), .Y(mai_mai_n1181_));
  INV        m1153(.A(mai_mai_n1181_), .Y(mai_mai_n1182_));
  AOI210     m1154(.A0(mai_mai_n1179_), .A1(mai_mai_n295_), .B0(mai_mai_n1182_), .Y(mai_mai_n1183_));
  AOI210     m1155(.A0(mai_mai_n1183_), .A1(mai_mai_n111_), .B0(mai_mai_n1178_), .Y(mai_mai_n1184_));
  NA2        m1156(.A(mai_mai_n479_), .B(mai_mai_n478_), .Y(mai_mai_n1185_));
  NO2        m1157(.A(mai_mai_n182_), .B(mai_mai_n239_), .Y(mai_mai_n1186_));
  NA2        m1158(.A(mai_mai_n1186_), .B(m), .Y(mai_mai_n1187_));
  AOI210     m1159(.A0(mai_mai_n1548_), .A1(mai_mai_n1185_), .B0(mai_mai_n1187_), .Y(mai_mai_n1188_));
  NA2        m1160(.A(mai_mai_n575_), .B(mai_mai_n417_), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n456_), .B(mai_mai_n1181_), .Y(mai_mai_n1190_));
  NO2        m1162(.A(mai_mai_n378_), .B(mai_mai_n377_), .Y(mai_mai_n1191_));
  AOI210     m1163(.A0(mai_mai_n1186_), .A1(mai_mai_n438_), .B0(mai_mai_n1000_), .Y(mai_mai_n1192_));
  NAi41      m1164(.An(mai_mai_n1191_), .B(mai_mai_n1192_), .C(mai_mai_n1190_), .D(mai_mai_n1189_), .Y(mai_mai_n1193_));
  NO2        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1188_), .Y(mai_mai_n1194_));
  NA4        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1184_), .C(mai_mai_n1174_), .D(mai_mai_n1170_), .Y(mai00));
  AOI210     m1167(.A0(mai_mai_n301_), .A1(mai_mai_n215_), .B0(mai_mai_n279_), .Y(mai_mai_n1196_));
  NO2        m1168(.A(mai_mai_n1196_), .B(mai_mai_n594_), .Y(mai_mai_n1197_));
  AOI210     m1169(.A0(mai_mai_n937_), .A1(mai_mai_n983_), .B0(mai_mai_n1154_), .Y(mai_mai_n1198_));
  NO3        m1170(.A(mai_mai_n1130_), .B(mai_mai_n1000_), .C(mai_mai_n736_), .Y(mai_mai_n1199_));
  NA3        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1198_), .C(mai_mai_n1043_), .Y(mai_mai_n1200_));
  NA2        m1172(.A(mai_mai_n520_), .B(f), .Y(mai_mai_n1201_));
  OAI210     m1173(.A0(mai_mai_n1050_), .A1(mai_mai_n40_), .B0(mai_mai_n664_), .Y(mai_mai_n1202_));
  NA3        m1174(.A(mai_mai_n1202_), .B(mai_mai_n261_), .C(n), .Y(mai_mai_n1203_));
  AOI210     m1175(.A0(mai_mai_n1203_), .A1(mai_mai_n1201_), .B0(mai_mai_n1087_), .Y(mai_mai_n1204_));
  NO4        m1176(.A(mai_mai_n1204_), .B(mai_mai_n1200_), .C(mai_mai_n1197_), .D(mai_mai_n1110_), .Y(mai_mai_n1205_));
  NA3        m1177(.A(mai_mai_n166_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1206_));
  NA3        m1178(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1207_));
  NOi31      m1179(.An(n), .B(m), .C(i), .Y(mai_mai_n1208_));
  NA3        m1180(.A(mai_mai_n1208_), .B(mai_mai_n667_), .C(mai_mai_n51_), .Y(mai_mai_n1209_));
  OAI210     m1181(.A0(mai_mai_n1207_), .A1(mai_mai_n1206_), .B0(mai_mai_n1209_), .Y(mai_mai_n1210_));
  INV        m1182(.A(mai_mai_n593_), .Y(mai_mai_n1211_));
  NO4        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1210_), .C(mai_mai_n1191_), .D(mai_mai_n959_), .Y(mai_mai_n1212_));
  NO4        m1184(.A(mai_mai_n496_), .B(mai_mai_n360_), .C(mai_mai_n1171_), .D(mai_mai_n59_), .Y(mai_mai_n1213_));
  NA3        m1185(.A(mai_mai_n390_), .B(mai_mai_n222_), .C(m), .Y(mai_mai_n1214_));
  OA220      m1186(.A0(mai_mai_n1214_), .A1(mai_mai_n1207_), .B0(mai_mai_n391_), .B1(mai_mai_n132_), .Y(mai_mai_n1215_));
  NO2        m1187(.A(h), .B(m), .Y(mai_mai_n1216_));
  NA4        m1188(.A(mai_mai_n508_), .B(mai_mai_n476_), .C(mai_mai_n1216_), .D(mai_mai_n1076_), .Y(mai_mai_n1217_));
  OAI220     m1189(.A0(mai_mai_n539_), .A1(mai_mai_n616_), .B0(mai_mai_n88_), .B1(mai_mai_n87_), .Y(mai_mai_n1218_));
  AOI220     m1190(.A0(mai_mai_n1218_), .A1(mai_mai_n548_), .B0(mai_mai_n988_), .B1(mai_mai_n592_), .Y(mai_mai_n1219_));
  AOI220     m1191(.A0(mai_mai_n319_), .A1(mai_mai_n250_), .B0(mai_mai_n177_), .B1(mai_mai_n147_), .Y(mai_mai_n1220_));
  NA4        m1192(.A(mai_mai_n1220_), .B(mai_mai_n1219_), .C(mai_mai_n1217_), .D(mai_mai_n1215_), .Y(mai_mai_n1221_));
  NO3        m1193(.A(mai_mai_n1221_), .B(mai_mai_n1213_), .C(mai_mai_n268_), .Y(mai_mai_n1222_));
  INV        m1194(.A(mai_mai_n323_), .Y(mai_mai_n1223_));
  AOI210     m1195(.A0(mai_mai_n250_), .A1(mai_mai_n350_), .B0(mai_mai_n595_), .Y(mai_mai_n1224_));
  NA3        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1223_), .C(mai_mai_n153_), .Y(mai_mai_n1225_));
  NO2        m1197(.A(mai_mai_n241_), .B(mai_mai_n181_), .Y(mai_mai_n1226_));
  NA2        m1198(.A(mai_mai_n1226_), .B(mai_mai_n436_), .Y(mai_mai_n1227_));
  NA3        m1199(.A(mai_mai_n179_), .B(mai_mai_n110_), .C(m), .Y(mai_mai_n1228_));
  NA3        m1200(.A(mai_mai_n476_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1229_));
  NOi31      m1201(.An(mai_mai_n908_), .B(mai_mai_n1229_), .C(mai_mai_n1228_), .Y(mai_mai_n1230_));
  NAi31      m1202(.An(mai_mai_n185_), .B(mai_mai_n896_), .C(mai_mai_n476_), .Y(mai_mai_n1231_));
  NAi31      m1203(.An(mai_mai_n1230_), .B(mai_mai_n1231_), .C(mai_mai_n1227_), .Y(mai_mai_n1232_));
  NO2        m1204(.A(mai_mai_n278_), .B(mai_mai_n69_), .Y(mai_mai_n1233_));
  NO3        m1205(.A(mai_mai_n435_), .B(mai_mai_n867_), .C(n), .Y(mai_mai_n1234_));
  AOI210     m1206(.A0(mai_mai_n1234_), .A1(mai_mai_n1233_), .B0(mai_mai_n1123_), .Y(mai_mai_n1235_));
  NAi21      m1207(.An(mai_mai_n1090_), .B(mai_mai_n1235_), .Y(mai_mai_n1236_));
  NO4        m1208(.A(mai_mai_n1236_), .B(mai_mai_n1232_), .C(mai_mai_n1225_), .D(mai_mai_n530_), .Y(mai_mai_n1237_));
  AN3        m1209(.A(mai_mai_n1237_), .B(mai_mai_n1222_), .C(mai_mai_n1212_), .Y(mai_mai_n1238_));
  NA2        m1210(.A(mai_mai_n548_), .B(mai_mai_n98_), .Y(mai_mai_n1239_));
  NA3        m1211(.A(mai_mai_n1155_), .B(mai_mai_n624_), .C(mai_mai_n475_), .Y(mai_mai_n1240_));
  NA4        m1212(.A(mai_mai_n1240_), .B(mai_mai_n576_), .C(mai_mai_n1239_), .D(mai_mai_n244_), .Y(mai_mai_n1241_));
  NA2        m1213(.A(mai_mai_n1149_), .B(mai_mai_n548_), .Y(mai_mai_n1242_));
  NA4        m1214(.A(mai_mai_n667_), .B(mai_mai_n206_), .C(mai_mai_n222_), .D(mai_mai_n162_), .Y(mai_mai_n1243_));
  NA3        m1215(.A(mai_mai_n1243_), .B(mai_mai_n1242_), .C(mai_mai_n298_), .Y(mai_mai_n1244_));
  OAI210     m1216(.A0(mai_mai_n474_), .A1(mai_mai_n117_), .B0(mai_mai_n902_), .Y(mai_mai_n1245_));
  AOI210     m1217(.A0(mai_mai_n575_), .A1(mai_mai_n417_), .B0(mai_mai_n1245_), .Y(mai_mai_n1246_));
  OR4        m1218(.A(mai_mai_n1087_), .B(mai_mai_n274_), .C(mai_mai_n224_), .D(e), .Y(mai_mai_n1247_));
  NO2        m1219(.A(mai_mai_n218_), .B(mai_mai_n215_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(n), .B(e), .Y(mai_mai_n1249_));
  NO2        m1221(.A(mai_mai_n1249_), .B(mai_mai_n145_), .Y(mai_mai_n1250_));
  AOI220     m1222(.A0(mai_mai_n1250_), .A1(mai_mai_n276_), .B0(mai_mai_n883_), .B1(mai_mai_n1248_), .Y(mai_mai_n1251_));
  OAI210     m1223(.A0(mai_mai_n361_), .A1(mai_mai_n314_), .B0(mai_mai_n458_), .Y(mai_mai_n1252_));
  NA4        m1224(.A(mai_mai_n1252_), .B(mai_mai_n1251_), .C(mai_mai_n1247_), .D(mai_mai_n1246_), .Y(mai_mai_n1253_));
  AOI210     m1225(.A0(mai_mai_n1250_), .A1(mai_mai_n887_), .B0(mai_mai_n855_), .Y(mai_mai_n1254_));
  AOI220     m1226(.A0(mai_mai_n997_), .A1(mai_mai_n592_), .B0(mai_mai_n667_), .B1(mai_mai_n247_), .Y(mai_mai_n1255_));
  NO2        m1227(.A(mai_mai_n64_), .B(h), .Y(mai_mai_n1256_));
  NO3        m1228(.A(mai_mai_n1087_), .B(mai_mai_n1085_), .C(mai_mai_n753_), .Y(mai_mai_n1257_));
  INV        m1229(.A(mai_mai_n129_), .Y(mai_mai_n1258_));
  AN2        m1230(.A(mai_mai_n1258_), .B(mai_mai_n1135_), .Y(mai_mai_n1259_));
  OAI210     m1231(.A0(mai_mai_n1259_), .A1(mai_mai_n1257_), .B0(mai_mai_n1256_), .Y(mai_mai_n1260_));
  NA4        m1232(.A(mai_mai_n1260_), .B(mai_mai_n1255_), .C(mai_mai_n1254_), .D(mai_mai_n904_), .Y(mai_mai_n1261_));
  NO4        m1233(.A(mai_mai_n1261_), .B(mai_mai_n1253_), .C(mai_mai_n1244_), .D(mai_mai_n1241_), .Y(mai_mai_n1262_));
  NA2        m1234(.A(mai_mai_n871_), .B(mai_mai_n786_), .Y(mai_mai_n1263_));
  NA4        m1235(.A(mai_mai_n1263_), .B(mai_mai_n1262_), .C(mai_mai_n1238_), .D(mai_mai_n1205_), .Y(mai01));
  AN2        m1236(.A(mai_mai_n1066_), .B(mai_mai_n1064_), .Y(mai_mai_n1265_));
  NO4        m1237(.A(mai_mai_n835_), .B(mai_mai_n827_), .C(mai_mai_n487_), .D(mai_mai_n285_), .Y(mai_mai_n1266_));
  NO2        m1238(.A(mai_mai_n609_), .B(mai_mai_n292_), .Y(mai_mai_n1267_));
  OAI210     m1239(.A0(mai_mai_n1267_), .A1(mai_mai_n401_), .B0(i), .Y(mai_mai_n1268_));
  NA3        m1240(.A(mai_mai_n1268_), .B(mai_mai_n1266_), .C(mai_mai_n1265_), .Y(mai_mai_n1269_));
  NA2        m1241(.A(mai_mai_n605_), .B(mai_mai_n86_), .Y(mai_mai_n1270_));
  NA2        m1242(.A(mai_mai_n568_), .B(mai_mai_n273_), .Y(mai_mai_n1271_));
  NA2        m1243(.A(mai_mai_n1002_), .B(mai_mai_n1271_), .Y(mai_mai_n1272_));
  NA4        m1244(.A(mai_mai_n1272_), .B(mai_mai_n1270_), .C(mai_mai_n952_), .D(mai_mai_n335_), .Y(mai_mai_n1273_));
  NA2        m1245(.A(mai_mai_n731_), .B(mai_mai_n93_), .Y(mai_mai_n1274_));
  NO2        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1546_), .Y(mai_mai_n1275_));
  OAI210     m1247(.A0(mai_mai_n813_), .A1(mai_mai_n619_), .B0(mai_mai_n1243_), .Y(mai_mai_n1276_));
  AOI210     m1248(.A0(mai_mai_n1275_), .A1(mai_mai_n653_), .B0(mai_mai_n1276_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n116_), .B(l), .Y(mai_mai_n1278_));
  OA220      m1250(.A0(mai_mai_n1278_), .A1(mai_mai_n602_), .B0(mai_mai_n680_), .B1(mai_mai_n375_), .Y(mai_mai_n1279_));
  NAi41      m1251(.An(mai_mai_n161_), .B(mai_mai_n1279_), .C(mai_mai_n1277_), .D(mai_mai_n936_), .Y(mai_mai_n1280_));
  NO3        m1252(.A(mai_mai_n814_), .B(mai_mai_n695_), .C(mai_mai_n523_), .Y(mai_mai_n1281_));
  NA4        m1253(.A(mai_mai_n731_), .B(mai_mai_n93_), .C(mai_mai_n45_), .D(mai_mai_n214_), .Y(mai_mai_n1282_));
  OA220      m1254(.A0(mai_mai_n1282_), .A1(mai_mai_n688_), .B0(mai_mai_n195_), .B1(mai_mai_n193_), .Y(mai_mai_n1283_));
  NA3        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1281_), .C(mai_mai_n135_), .Y(mai_mai_n1284_));
  NO4        m1256(.A(mai_mai_n1284_), .B(mai_mai_n1280_), .C(mai_mai_n1273_), .D(mai_mai_n1269_), .Y(mai_mai_n1285_));
  NA2        m1257(.A(mai_mai_n1214_), .B(mai_mai_n207_), .Y(mai_mai_n1286_));
  OAI210     m1258(.A0(mai_mai_n1286_), .A1(mai_mai_n304_), .B0(mai_mai_n543_), .Y(mai_mai_n1287_));
  NA2        m1259(.A(mai_mai_n551_), .B(mai_mai_n403_), .Y(mai_mai_n1288_));
  NA2        m1260(.A(mai_mai_n70_), .B(i), .Y(mai_mai_n1289_));
  AOI210     m1261(.A0(mai_mai_n608_), .A1(mai_mai_n602_), .B0(mai_mai_n1289_), .Y(mai_mai_n1290_));
  NOi21      m1262(.An(mai_mai_n577_), .B(mai_mai_n599_), .Y(mai_mai_n1291_));
  AOI210     m1263(.A0(mai_mai_n1291_), .A1(mai_mai_n1288_), .B0(mai_mai_n1290_), .Y(mai_mai_n1292_));
  AOI210     m1264(.A0(mai_mai_n204_), .A1(mai_mai_n85_), .B0(mai_mai_n214_), .Y(mai_mai_n1293_));
  OAI210     m1265(.A0(mai_mai_n842_), .A1(mai_mai_n436_), .B0(mai_mai_n1293_), .Y(mai_mai_n1294_));
  AN3        m1266(.A(m), .B(l), .C(k), .Y(mai_mai_n1295_));
  OAI210     m1267(.A0(mai_mai_n363_), .A1(mai_mai_n34_), .B0(mai_mai_n1295_), .Y(mai_mai_n1296_));
  NA2        m1268(.A(mai_mai_n203_), .B(mai_mai_n34_), .Y(mai_mai_n1297_));
  AO210      m1269(.A0(mai_mai_n1297_), .A1(mai_mai_n1296_), .B0(mai_mai_n334_), .Y(mai_mai_n1298_));
  NA4        m1270(.A(mai_mai_n1298_), .B(mai_mai_n1294_), .C(mai_mai_n1292_), .D(mai_mai_n1287_), .Y(mai_mai_n1299_));
  NA2        m1271(.A(mai_mai_n614_), .B(mai_mai_n116_), .Y(mai_mai_n1300_));
  OAI210     m1272(.A0(mai_mai_n1278_), .A1(mai_mai_n611_), .B0(mai_mai_n1300_), .Y(mai_mai_n1301_));
  NA2        m1273(.A(mai_mai_n284_), .B(mai_mai_n195_), .Y(mai_mai_n1302_));
  OAI210     m1274(.A0(mai_mai_n1302_), .A1(mai_mai_n392_), .B0(mai_mai_n685_), .Y(mai_mai_n1303_));
  NO3        m1275(.A(mai_mai_n854_), .B(mai_mai_n204_), .C(mai_mai_n415_), .Y(mai_mai_n1304_));
  NO2        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1000_), .Y(mai_mai_n1305_));
  OAI210     m1277(.A0(mai_mai_n1275_), .A1(mai_mai_n328_), .B0(mai_mai_n696_), .Y(mai_mai_n1306_));
  NA4        m1278(.A(mai_mai_n1306_), .B(mai_mai_n1305_), .C(mai_mai_n1303_), .D(mai_mai_n817_), .Y(mai_mai_n1307_));
  NO3        m1279(.A(mai_mai_n1307_), .B(mai_mai_n1301_), .C(mai_mai_n1299_), .Y(mai_mai_n1308_));
  NA3        m1280(.A(mai_mai_n620_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n1309_), .B(mai_mai_n204_), .Y(mai_mai_n1310_));
  AOI210     m1282(.A0(mai_mai_n515_), .A1(mai_mai_n58_), .B0(mai_mai_n1310_), .Y(mai_mai_n1311_));
  OR3        m1283(.A(mai_mai_n1274_), .B(mai_mai_n621_), .C(mai_mai_n1546_), .Y(mai_mai_n1312_));
  NA3        m1284(.A(mai_mai_n767_), .B(mai_mai_n70_), .C(i), .Y(mai_mai_n1313_));
  AOI210     m1285(.A0(mai_mai_n1313_), .A1(mai_mai_n1282_), .B0(mai_mai_n1021_), .Y(mai_mai_n1314_));
  NO2        m1286(.A(mai_mai_n207_), .B(mai_mai_n109_), .Y(mai_mai_n1315_));
  NO3        m1287(.A(mai_mai_n1315_), .B(mai_mai_n1314_), .C(mai_mai_n1210_), .Y(mai_mai_n1316_));
  NA4        m1288(.A(mai_mai_n1316_), .B(mai_mai_n1312_), .C(mai_mai_n1311_), .D(mai_mai_n785_), .Y(mai_mai_n1317_));
  NO2        m1289(.A(mai_mai_n1008_), .B(mai_mai_n234_), .Y(mai_mai_n1318_));
  NO2        m1290(.A(mai_mai_n1009_), .B(mai_mai_n570_), .Y(mai_mai_n1319_));
  OAI210     m1291(.A0(mai_mai_n1319_), .A1(mai_mai_n1318_), .B0(mai_mai_n343_), .Y(mai_mai_n1320_));
  NA2        m1292(.A(mai_mai_n587_), .B(mai_mai_n585_), .Y(mai_mai_n1321_));
  NO3        m1293(.A(mai_mai_n75_), .B(mai_mai_n302_), .C(mai_mai_n45_), .Y(mai_mai_n1322_));
  NA2        m1294(.A(mai_mai_n1322_), .B(mai_mai_n567_), .Y(mai_mai_n1323_));
  NA3        m1295(.A(mai_mai_n1323_), .B(mai_mai_n1321_), .C(mai_mai_n690_), .Y(mai_mai_n1324_));
  OR2        m1296(.A(mai_mai_n1214_), .B(mai_mai_n1207_), .Y(mai_mai_n1325_));
  NO2        m1297(.A(mai_mai_n375_), .B(mai_mai_n68_), .Y(mai_mai_n1326_));
  AOI210     m1298(.A0(mai_mai_n758_), .A1(mai_mai_n635_), .B0(mai_mai_n1326_), .Y(mai_mai_n1327_));
  NA2        m1299(.A(mai_mai_n1322_), .B(mai_mai_n845_), .Y(mai_mai_n1328_));
  NA4        m1300(.A(mai_mai_n1328_), .B(mai_mai_n1327_), .C(mai_mai_n1325_), .D(mai_mai_n393_), .Y(mai_mai_n1329_));
  NOi41      m1301(.An(mai_mai_n1320_), .B(mai_mai_n1329_), .C(mai_mai_n1324_), .D(mai_mai_n1317_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n128_), .B(mai_mai_n45_), .Y(mai_mai_n1331_));
  NO2        m1303(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1332_));
  AO220      m1304(.A0(mai_mai_n1332_), .A1(mai_mai_n641_), .B0(mai_mai_n1331_), .B1(mai_mai_n729_), .Y(mai_mai_n1333_));
  NA2        m1305(.A(mai_mai_n1333_), .B(mai_mai_n343_), .Y(mai_mai_n1334_));
  NA2        m1306(.A(mai_mai_n469_), .B(mai_mai_n132_), .Y(mai_mai_n1335_));
  NO3        m1307(.A(mai_mai_n1133_), .B(mai_mai_n176_), .C(mai_mai_n83_), .Y(mai_mai_n1336_));
  AOI220     m1308(.A0(mai_mai_n1336_), .A1(mai_mai_n1335_), .B0(mai_mai_n1322_), .B1(mai_mai_n1012_), .Y(mai_mai_n1337_));
  NA2        m1309(.A(mai_mai_n1337_), .B(mai_mai_n1334_), .Y(mai_mai_n1338_));
  NO2        m1310(.A(mai_mai_n632_), .B(mai_mai_n631_), .Y(mai_mai_n1339_));
  NO4        m1311(.A(mai_mai_n1133_), .B(mai_mai_n1339_), .C(mai_mai_n174_), .D(mai_mai_n83_), .Y(mai_mai_n1340_));
  NO3        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1338_), .C(mai_mai_n656_), .Y(mai_mai_n1341_));
  NA4        m1313(.A(mai_mai_n1341_), .B(mai_mai_n1330_), .C(mai_mai_n1308_), .D(mai_mai_n1285_), .Y(mai06));
  NO2        m1314(.A(mai_mai_n416_), .B(mai_mai_n574_), .Y(mai_mai_n1343_));
  NA2        m1315(.A(mai_mai_n269_), .B(mai_mai_n1343_), .Y(mai_mai_n1344_));
  NO2        m1316(.A(mai_mai_n226_), .B(mai_mai_n100_), .Y(mai_mai_n1345_));
  OAI210     m1317(.A0(mai_mai_n1345_), .A1(mai_mai_n1336_), .B0(mai_mai_n389_), .Y(mai_mai_n1346_));
  NO3        m1318(.A(mai_mai_n617_), .B(mai_mai_n840_), .C(mai_mai_n618_), .Y(mai_mai_n1347_));
  OR2        m1319(.A(mai_mai_n1347_), .B(mai_mai_n923_), .Y(mai_mai_n1348_));
  NA4        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1346_), .C(mai_mai_n1344_), .D(mai_mai_n1320_), .Y(mai_mai_n1349_));
  NO3        m1321(.A(mai_mai_n1349_), .B(mai_mai_n1324_), .C(mai_mai_n260_), .Y(mai_mai_n1350_));
  NO2        m1322(.A(mai_mai_n302_), .B(mai_mai_n45_), .Y(mai_mai_n1351_));
  AOI210     m1323(.A0(mai_mai_n1351_), .A1(mai_mai_n1013_), .B0(mai_mai_n1318_), .Y(mai_mai_n1352_));
  AOI210     m1324(.A0(mai_mai_n1351_), .A1(mai_mai_n571_), .B0(mai_mai_n1333_), .Y(mai_mai_n1353_));
  AOI210     m1325(.A0(mai_mai_n1353_), .A1(mai_mai_n1352_), .B0(mai_mai_n340_), .Y(mai_mai_n1354_));
  OAI210     m1326(.A0(mai_mai_n85_), .A1(mai_mai_n40_), .B0(mai_mai_n694_), .Y(mai_mai_n1355_));
  NA2        m1327(.A(mai_mai_n1355_), .B(mai_mai_n660_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n526_), .B(mai_mai_n171_), .Y(mai_mai_n1357_));
  NOi21      m1329(.An(mai_mai_n134_), .B(mai_mai_n45_), .Y(mai_mai_n1358_));
  AOI210     m1330(.A0(mai_mai_n625_), .A1(mai_mai_n57_), .B0(mai_mai_n1156_), .Y(mai_mai_n1359_));
  OAI210     m1331(.A0(mai_mai_n469_), .A1(mai_mai_n251_), .B0(mai_mai_n946_), .Y(mai_mai_n1360_));
  NO4        m1332(.A(mai_mai_n1360_), .B(mai_mai_n1359_), .C(mai_mai_n1358_), .D(mai_mai_n1357_), .Y(mai_mai_n1361_));
  NO2        m1333(.A(mai_mai_n374_), .B(mai_mai_n133_), .Y(mai_mai_n1362_));
  NA2        m1334(.A(mai_mai_n1362_), .B(mai_mai_n605_), .Y(mai_mai_n1363_));
  NA3        m1335(.A(mai_mai_n1363_), .B(mai_mai_n1361_), .C(mai_mai_n1356_), .Y(mai_mai_n1364_));
  NO2        m1336(.A(mai_mai_n776_), .B(mai_mai_n373_), .Y(mai_mai_n1365_));
  NO3        m1337(.A(mai_mai_n696_), .B(mai_mai_n787_), .C(mai_mai_n653_), .Y(mai_mai_n1366_));
  NOi21      m1338(.An(mai_mai_n1365_), .B(mai_mai_n1366_), .Y(mai_mai_n1367_));
  AN2        m1339(.A(mai_mai_n997_), .B(mai_mai_n663_), .Y(mai_mai_n1368_));
  NO4        m1340(.A(mai_mai_n1368_), .B(mai_mai_n1367_), .C(mai_mai_n1364_), .D(mai_mai_n1354_), .Y(mai_mai_n1369_));
  NO2        m1341(.A(mai_mai_n834_), .B(mai_mai_n280_), .Y(mai_mai_n1370_));
  OAI220     m1342(.A0(mai_mai_n760_), .A1(mai_mai_n47_), .B0(mai_mai_n226_), .B1(mai_mai_n634_), .Y(mai_mai_n1371_));
  OAI210     m1343(.A0(mai_mai_n280_), .A1(c), .B0(mai_mai_n659_), .Y(mai_mai_n1372_));
  AOI220     m1344(.A0(mai_mai_n1372_), .A1(mai_mai_n1371_), .B0(mai_mai_n1370_), .B1(mai_mai_n269_), .Y(mai_mai_n1373_));
  NO3        m1345(.A(mai_mai_n246_), .B(mai_mai_n100_), .C(mai_mai_n287_), .Y(mai_mai_n1374_));
  OAI220     m1346(.A0(mai_mai_n721_), .A1(mai_mai_n251_), .B0(mai_mai_n522_), .B1(mai_mai_n526_), .Y(mai_mai_n1375_));
  OAI210     m1347(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1376_));
  NO3        m1348(.A(mai_mai_n1376_), .B(mai_mai_n616_), .C(j), .Y(mai_mai_n1377_));
  NOi21      m1349(.An(mai_mai_n1377_), .B(mai_mai_n688_), .Y(mai_mai_n1378_));
  NO4        m1350(.A(mai_mai_n1378_), .B(mai_mai_n1375_), .C(mai_mai_n1374_), .D(mai_mai_n1159_), .Y(mai_mai_n1379_));
  NA4        m1351(.A(mai_mai_n825_), .B(mai_mai_n824_), .C(mai_mai_n446_), .D(mai_mai_n915_), .Y(mai_mai_n1380_));
  NAi31      m1352(.An(mai_mai_n776_), .B(mai_mai_n1380_), .C(mai_mai_n203_), .Y(mai_mai_n1381_));
  NA4        m1353(.A(mai_mai_n1381_), .B(mai_mai_n1379_), .C(mai_mai_n1373_), .D(mai_mai_n1255_), .Y(mai_mai_n1382_));
  OR2        m1354(.A(mai_mai_n813_), .B(mai_mai_n554_), .Y(mai_mai_n1383_));
  OR3        m1355(.A(mai_mai_n377_), .B(mai_mai_n226_), .C(mai_mai_n634_), .Y(mai_mai_n1384_));
  AOI210     m1356(.A0(mai_mai_n587_), .A1(mai_mai_n458_), .B0(mai_mai_n379_), .Y(mai_mai_n1385_));
  NA2        m1357(.A(mai_mai_n1377_), .B(mai_mai_n821_), .Y(mai_mai_n1386_));
  NA4        m1358(.A(mai_mai_n1386_), .B(mai_mai_n1385_), .C(mai_mai_n1384_), .D(mai_mai_n1383_), .Y(mai_mai_n1387_));
  AOI220     m1359(.A0(mai_mai_n1365_), .A1(mai_mai_n786_), .B0(mai_mai_n1362_), .B1(mai_mai_n240_), .Y(mai_mai_n1388_));
  AO220      m1360(.A0(mai_mai_n1345_), .A1(mai_mai_n685_), .B0(mai_mai_n968_), .B1(mai_mai_n967_), .Y(mai_mai_n1389_));
  NO4        m1361(.A(mai_mai_n1389_), .B(mai_mai_n913_), .C(mai_mai_n511_), .D(mai_mai_n490_), .Y(mai_mai_n1390_));
  NA3        m1362(.A(mai_mai_n1390_), .B(mai_mai_n1388_), .C(mai_mai_n1328_), .Y(mai_mai_n1391_));
  NAi21      m1363(.An(j), .B(i), .Y(mai_mai_n1392_));
  NO4        m1364(.A(mai_mai_n1339_), .B(mai_mai_n1392_), .C(mai_mai_n452_), .D(mai_mai_n237_), .Y(mai_mai_n1393_));
  NO4        m1365(.A(mai_mai_n1393_), .B(mai_mai_n1391_), .C(mai_mai_n1387_), .D(mai_mai_n1382_), .Y(mai_mai_n1394_));
  NA4        m1366(.A(mai_mai_n1394_), .B(mai_mai_n1369_), .C(mai_mai_n1350_), .D(mai_mai_n1341_), .Y(mai07));
  NOi21      m1367(.An(j), .B(k), .Y(mai_mai_n1396_));
  NA4        m1368(.A(mai_mai_n179_), .B(mai_mai_n106_), .C(mai_mai_n1396_), .D(f), .Y(mai_mai_n1397_));
  NAi32      m1369(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1398_));
  NO3        m1370(.A(mai_mai_n1398_), .B(m), .C(f), .Y(mai_mai_n1399_));
  OAI210     m1371(.A0(i), .A1(mai_mai_n492_), .B0(mai_mai_n1399_), .Y(mai_mai_n1400_));
  NAi21      m1372(.An(f), .B(c), .Y(mai_mai_n1401_));
  OR2        m1373(.A(e), .B(d), .Y(mai_mai_n1402_));
  OAI220     m1374(.A0(mai_mai_n1402_), .A1(mai_mai_n1401_), .B0(mai_mai_n645_), .B1(mai_mai_n324_), .Y(mai_mai_n1403_));
  NA3        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1099_), .C(mai_mai_n179_), .Y(mai_mai_n1404_));
  NOi31      m1376(.An(n), .B(m), .C(b), .Y(mai_mai_n1405_));
  NO3        m1377(.A(mai_mai_n129_), .B(mai_mai_n459_), .C(h), .Y(mai_mai_n1406_));
  NA3        m1378(.A(mai_mai_n1404_), .B(mai_mai_n1400_), .C(mai_mai_n1397_), .Y(mai_mai_n1407_));
  NOi41      m1379(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1408_));
  NO2        m1380(.A(k), .B(i), .Y(mai_mai_n1409_));
  NA3        m1381(.A(mai_mai_n1409_), .B(mai_mai_n935_), .C(mai_mai_n179_), .Y(mai_mai_n1410_));
  NA2        m1382(.A(mai_mai_n83_), .B(mai_mai_n45_), .Y(mai_mai_n1411_));
  NO2        m1383(.A(mai_mai_n1093_), .B(mai_mai_n452_), .Y(mai_mai_n1412_));
  NA3        m1384(.A(mai_mai_n1412_), .B(mai_mai_n1411_), .C(mai_mai_n215_), .Y(mai_mai_n1413_));
  NO2        m1385(.A(mai_mai_n1107_), .B(mai_mai_n310_), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1256_), .B(mai_mai_n293_), .Y(mai_mai_n1415_));
  NA3        m1387(.A(mai_mai_n1415_), .B(mai_mai_n1413_), .C(mai_mai_n1410_), .Y(mai_mai_n1416_));
  NO2        m1388(.A(mai_mai_n1416_), .B(mai_mai_n1407_), .Y(mai_mai_n1417_));
  NO3        m1389(.A(e), .B(d), .C(c), .Y(mai_mai_n1418_));
  OAI210     m1390(.A0(mai_mai_n129_), .A1(mai_mai_n215_), .B0(mai_mai_n622_), .Y(mai_mai_n1419_));
  NA2        m1391(.A(mai_mai_n1419_), .B(mai_mai_n1418_), .Y(mai_mai_n1420_));
  INV        m1392(.A(mai_mai_n1420_), .Y(mai_mai_n1421_));
  NA3        m1393(.A(mai_mai_n718_), .B(mai_mai_n704_), .C(mai_mai_n110_), .Y(mai_mai_n1422_));
  NO2        m1394(.A(mai_mai_n1422_), .B(mai_mai_n45_), .Y(mai_mai_n1423_));
  NO2        m1395(.A(l), .B(k), .Y(mai_mai_n1424_));
  NOi41      m1396(.An(mai_mai_n560_), .B(mai_mai_n1424_), .C(mai_mai_n485_), .D(mai_mai_n452_), .Y(mai_mai_n1425_));
  NO3        m1397(.A(mai_mai_n452_), .B(d), .C(c), .Y(mai_mai_n1426_));
  NO3        m1398(.A(mai_mai_n1425_), .B(mai_mai_n1423_), .C(mai_mai_n1421_), .Y(mai_mai_n1427_));
  NO2        m1399(.A(mai_mai_n146_), .B(h), .Y(mai_mai_n1428_));
  NO2        m1400(.A(m), .B(c), .Y(mai_mai_n1429_));
  NA3        m1401(.A(mai_mai_n1429_), .B(mai_mai_n140_), .C(mai_mai_n186_), .Y(mai_mai_n1430_));
  NO2        m1402(.A(mai_mai_n1430_), .B(mai_mai_n1545_), .Y(mai_mai_n1431_));
  NA2        m1403(.A(mai_mai_n1431_), .B(mai_mai_n179_), .Y(mai_mai_n1432_));
  NO2        m1404(.A(mai_mai_n460_), .B(a), .Y(mai_mai_n1433_));
  NA3        m1405(.A(mai_mai_n1433_), .B(k), .C(mai_mai_n111_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(i), .B(h), .Y(mai_mai_n1435_));
  NA2        m1407(.A(mai_mai_n1180_), .B(h), .Y(mai_mai_n1436_));
  NA2        m1408(.A(mai_mai_n136_), .B(mai_mai_n222_), .Y(mai_mai_n1437_));
  NO2        m1409(.A(mai_mai_n1437_), .B(mai_mai_n1436_), .Y(mai_mai_n1438_));
  NO2        m1410(.A(mai_mai_n783_), .B(mai_mai_n187_), .Y(mai_mai_n1439_));
  NOi31      m1411(.An(m), .B(n), .C(b), .Y(mai_mai_n1440_));
  NOi31      m1412(.An(f), .B(d), .C(c), .Y(mai_mai_n1441_));
  NA2        m1413(.A(mai_mai_n1441_), .B(mai_mai_n1440_), .Y(mai_mai_n1442_));
  INV        m1414(.A(mai_mai_n1442_), .Y(mai_mai_n1443_));
  NO3        m1415(.A(mai_mai_n1443_), .B(mai_mai_n1439_), .C(mai_mai_n1438_), .Y(mai_mai_n1444_));
  NA2        m1416(.A(mai_mai_n1126_), .B(mai_mai_n476_), .Y(mai_mai_n1445_));
  NO4        m1417(.A(mai_mai_n1445_), .B(mai_mai_n1102_), .C(mai_mai_n452_), .D(mai_mai_n45_), .Y(mai_mai_n1446_));
  OAI210     m1418(.A0(mai_mai_n182_), .A1(mai_mai_n538_), .B0(mai_mai_n1103_), .Y(mai_mai_n1447_));
  INV        m1419(.A(mai_mai_n1447_), .Y(mai_mai_n1448_));
  NO2        m1420(.A(mai_mai_n1448_), .B(mai_mai_n1446_), .Y(mai_mai_n1449_));
  AN4        m1421(.A(mai_mai_n1449_), .B(mai_mai_n1444_), .C(mai_mai_n1434_), .D(mai_mai_n1432_), .Y(mai_mai_n1450_));
  NA2        m1422(.A(mai_mai_n1405_), .B(mai_mai_n386_), .Y(mai_mai_n1451_));
  NA2        m1423(.A(mai_mai_n1426_), .B(mai_mai_n216_), .Y(mai_mai_n1452_));
  NA2        m1424(.A(mai_mai_n1134_), .B(mai_mai_n1445_), .Y(mai_mai_n1453_));
  NA2        m1425(.A(mai_mai_n1453_), .B(mai_mai_n1452_), .Y(mai_mai_n1454_));
  NO4        m1426(.A(mai_mai_n129_), .B(m), .C(f), .D(e), .Y(mai_mai_n1455_));
  NA3        m1427(.A(mai_mai_n1409_), .B(mai_mai_n294_), .C(h), .Y(mai_mai_n1456_));
  OR2        m1428(.A(e), .B(a), .Y(mai_mai_n1457_));
  NO2        m1429(.A(mai_mai_n1402_), .B(mai_mai_n1401_), .Y(mai_mai_n1458_));
  AOI210     m1430(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1458_), .Y(mai_mai_n1459_));
  NO2        m1431(.A(mai_mai_n1459_), .B(mai_mai_n1122_), .Y(mai_mai_n1460_));
  NA2        m1432(.A(mai_mai_n1408_), .B(mai_mai_n1424_), .Y(mai_mai_n1461_));
  INV        m1433(.A(mai_mai_n1461_), .Y(mai_mai_n1462_));
  NA2        m1434(.A(mai_mai_n1155_), .B(mai_mai_n415_), .Y(mai_mai_n1463_));
  NO2        m1435(.A(mai_mai_n1463_), .B(mai_mai_n445_), .Y(mai_mai_n1464_));
  AO210      m1436(.A0(mai_mai_n1464_), .A1(mai_mai_n114_), .B0(mai_mai_n1462_), .Y(mai_mai_n1465_));
  NO3        m1437(.A(mai_mai_n1465_), .B(mai_mai_n1460_), .C(mai_mai_n1454_), .Y(mai_mai_n1466_));
  NA4        m1438(.A(mai_mai_n1466_), .B(mai_mai_n1450_), .C(mai_mai_n1427_), .D(mai_mai_n1417_), .Y(mai_mai_n1467_));
  NO2        m1439(.A(mai_mai_n398_), .B(j), .Y(mai_mai_n1468_));
  NAi41      m1440(.An(mai_mai_n1435_), .B(mai_mai_n1115_), .C(mai_mai_n167_), .D(mai_mai_n149_), .Y(mai_mai_n1469_));
  INV        m1441(.A(mai_mai_n1469_), .Y(mai_mai_n1470_));
  NA3        m1442(.A(m), .B(mai_mai_n1468_), .C(mai_mai_n158_), .Y(mai_mai_n1471_));
  INV        m1443(.A(mai_mai_n1471_), .Y(mai_mai_n1472_));
  NO3        m1444(.A(mai_mai_n776_), .B(mai_mai_n174_), .C(mai_mai_n418_), .Y(mai_mai_n1473_));
  NO3        m1445(.A(mai_mai_n1473_), .B(mai_mai_n1472_), .C(mai_mai_n1470_), .Y(mai_mai_n1474_));
  OR2        m1446(.A(n), .B(i), .Y(mai_mai_n1475_));
  OAI210     m1447(.A0(mai_mai_n1475_), .A1(mai_mai_n1114_), .B0(mai_mai_n49_), .Y(mai_mai_n1476_));
  AOI220     m1448(.A0(mai_mai_n1476_), .A1(mai_mai_n1216_), .B0(mai_mai_n859_), .B1(mai_mai_n194_), .Y(mai_mai_n1477_));
  NO3        m1449(.A(mai_mai_n1137_), .B(mai_mai_n1402_), .C(mai_mai_n49_), .Y(mai_mai_n1478_));
  NO2        m1450(.A(mai_mai_n1122_), .B(h), .Y(mai_mai_n1479_));
  NA3        m1451(.A(mai_mai_n1479_), .B(d), .C(mai_mai_n1085_), .Y(mai_mai_n1480_));
  NO2        m1452(.A(mai_mai_n1480_), .B(c), .Y(mai_mai_n1481_));
  NA2        m1453(.A(mai_mai_n179_), .B(mai_mai_n110_), .Y(mai_mai_n1482_));
  NOi21      m1454(.An(d), .B(f), .Y(mai_mai_n1483_));
  INV        m1455(.A(mai_mai_n1481_), .Y(mai_mai_n1484_));
  NA3        m1456(.A(mai_mai_n1484_), .B(mai_mai_n1477_), .C(mai_mai_n1474_), .Y(mai_mai_n1485_));
  NO3        m1457(.A(mai_mai_n1126_), .B(mai_mai_n1114_), .C(mai_mai_n40_), .Y(mai_mai_n1486_));
  NA2        m1458(.A(mai_mai_n1486_), .B(mai_mai_n1414_), .Y(mai_mai_n1487_));
  OAI210     m1459(.A0(mai_mai_n1455_), .A1(mai_mai_n1405_), .B0(mai_mai_n920_), .Y(mai_mai_n1488_));
  NO2        m1460(.A(mai_mai_n1082_), .B(mai_mai_n129_), .Y(mai_mai_n1489_));
  NA2        m1461(.A(mai_mai_n1489_), .B(mai_mai_n640_), .Y(mai_mai_n1490_));
  NA3        m1462(.A(mai_mai_n1490_), .B(mai_mai_n1488_), .C(mai_mai_n1487_), .Y(mai_mai_n1491_));
  NA2        m1463(.A(mai_mai_n1429_), .B(mai_mai_n1483_), .Y(mai_mai_n1492_));
  NO2        m1464(.A(mai_mai_n1492_), .B(m), .Y(mai_mai_n1493_));
  OAI220     m1465(.A0(mai_mai_n150_), .A1(mai_mai_n181_), .B0(mai_mai_n459_), .B1(m), .Y(mai_mai_n1494_));
  OAI210     m1466(.A0(mai_mai_n1494_), .A1(mai_mai_n108_), .B0(mai_mai_n1440_), .Y(mai_mai_n1495_));
  INV        m1467(.A(mai_mai_n1495_), .Y(mai_mai_n1496_));
  NO3        m1468(.A(mai_mai_n1496_), .B(mai_mai_n1493_), .C(mai_mai_n1491_), .Y(mai_mai_n1497_));
  NO2        m1469(.A(mai_mai_n1401_), .B(e), .Y(mai_mai_n1498_));
  NA2        m1470(.A(mai_mai_n1166_), .B(mai_mai_n649_), .Y(mai_mai_n1499_));
  NO2        m1471(.A(mai_mai_n1499_), .B(mai_mai_n454_), .Y(mai_mai_n1500_));
  INV        m1472(.A(mai_mai_n1500_), .Y(mai_mai_n1501_));
  NO2        m1473(.A(mai_mai_n181_), .B(c), .Y(mai_mai_n1502_));
  OAI210     m1474(.A0(mai_mai_n1502_), .A1(mai_mai_n1498_), .B0(mai_mai_n179_), .Y(mai_mai_n1503_));
  AOI220     m1475(.A0(mai_mai_n1503_), .A1(mai_mai_n1116_), .B0(mai_mai_n545_), .B1(mai_mai_n373_), .Y(mai_mai_n1504_));
  NA2        m1476(.A(mai_mai_n553_), .B(m), .Y(mai_mai_n1505_));
  AOI210     m1477(.A0(mai_mai_n1505_), .A1(mai_mai_n1426_), .B0(mai_mai_n1478_), .Y(mai_mai_n1506_));
  NO2        m1478(.A(mai_mai_n1457_), .B(f), .Y(mai_mai_n1507_));
  AOI210     m1479(.A0(mai_mai_n1166_), .A1(a), .B0(mai_mai_n1507_), .Y(mai_mai_n1508_));
  OAI220     m1480(.A0(mai_mai_n1508_), .A1(mai_mai_n65_), .B0(mai_mai_n1506_), .B1(mai_mai_n214_), .Y(mai_mai_n1509_));
  AOI210     m1481(.A0(mai_mai_n940_), .A1(mai_mai_n425_), .B0(mai_mai_n102_), .Y(mai_mai_n1510_));
  OR2        m1482(.A(mai_mai_n1510_), .B(mai_mai_n553_), .Y(mai_mai_n1511_));
  NO2        m1483(.A(mai_mai_n1511_), .B(mai_mai_n174_), .Y(mai_mai_n1512_));
  NA4        m1484(.A(mai_mai_n1135_), .B(mai_mai_n1132_), .C(mai_mai_n222_), .D(mai_mai_n64_), .Y(mai_mai_n1513_));
  NA2        m1485(.A(mai_mai_n1406_), .B(mai_mai_n182_), .Y(mai_mai_n1514_));
  NO2        m1486(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1515_));
  OAI210     m1487(.A0(mai_mai_n1457_), .A1(mai_mai_n898_), .B0(mai_mai_n492_), .Y(mai_mai_n1516_));
  OAI210     m1488(.A0(mai_mai_n1516_), .A1(mai_mai_n1138_), .B0(mai_mai_n1515_), .Y(mai_mai_n1517_));
  NO2        m1489(.A(m), .B(i), .Y(mai_mai_n1518_));
  NA2        m1490(.A(mai_mai_n1518_), .B(mai_mai_n1428_), .Y(mai_mai_n1519_));
  NA4        m1491(.A(mai_mai_n1519_), .B(mai_mai_n1517_), .C(mai_mai_n1514_), .D(mai_mai_n1513_), .Y(mai_mai_n1520_));
  NO4        m1492(.A(mai_mai_n1520_), .B(mai_mai_n1512_), .C(mai_mai_n1509_), .D(mai_mai_n1504_), .Y(mai_mai_n1521_));
  NA3        m1493(.A(mai_mai_n1521_), .B(mai_mai_n1501_), .C(mai_mai_n1497_), .Y(mai_mai_n1522_));
  AO210      m1494(.A0(mai_mai_n130_), .A1(l), .B0(mai_mai_n1451_), .Y(mai_mai_n1523_));
  NO4        m1495(.A(mai_mai_n226_), .B(mai_mai_n185_), .C(mai_mai_n261_), .D(k), .Y(mai_mai_n1524_));
  AOI210     m1496(.A0(mai_mai_n156_), .A1(mai_mai_n56_), .B0(mai_mai_n1498_), .Y(mai_mai_n1525_));
  NO2        m1497(.A(mai_mai_n1525_), .B(mai_mai_n1482_), .Y(mai_mai_n1526_));
  NOi21      m1498(.An(mai_mai_n1406_), .B(e), .Y(mai_mai_n1527_));
  NO3        m1499(.A(mai_mai_n1527_), .B(mai_mai_n1526_), .C(mai_mai_n1524_), .Y(mai_mai_n1528_));
  NA2        m1500(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1529_));
  NO2        m1501(.A(mai_mai_n1463_), .B(mai_mai_n1529_), .Y(mai_mai_n1530_));
  INV        m1502(.A(mai_mai_n1530_), .Y(mai_mai_n1531_));
  NA3        m1503(.A(mai_mai_n1531_), .B(mai_mai_n1528_), .C(mai_mai_n1523_), .Y(mai_mai_n1532_));
  OR4        m1504(.A(mai_mai_n1532_), .B(mai_mai_n1522_), .C(mai_mai_n1485_), .D(mai_mai_n1467_), .Y(mai04));
  NOi31      m1505(.An(mai_mai_n1455_), .B(mai_mai_n1456_), .C(mai_mai_n1087_), .Y(mai_mai_n1534_));
  INV        m1506(.A(mai_mai_n859_), .Y(mai_mai_n1535_));
  NO4        m1507(.A(mai_mai_n1535_), .B(mai_mai_n1077_), .C(mai_mai_n493_), .D(j), .Y(mai_mai_n1536_));
  OR3        m1508(.A(mai_mai_n1536_), .B(mai_mai_n1534_), .C(mai_mai_n1105_), .Y(mai_mai_n1537_));
  NO3        m1509(.A(mai_mai_n1411_), .B(mai_mai_n87_), .C(k), .Y(mai_mai_n1538_));
  AOI210     m1510(.A0(mai_mai_n1538_), .A1(mai_mai_n1098_), .B0(mai_mai_n1230_), .Y(mai_mai_n1539_));
  NA2        m1511(.A(mai_mai_n1539_), .B(mai_mai_n1260_), .Y(mai_mai_n1540_));
  NO4        m1512(.A(mai_mai_n1540_), .B(mai_mai_n1537_), .C(mai_mai_n1113_), .D(mai_mai_n1092_), .Y(mai_mai_n1541_));
  NA4        m1513(.A(mai_mai_n1541_), .B(mai_mai_n1168_), .C(mai_mai_n1153_), .D(mai_mai_n1141_), .Y(mai05));
  INV        m1514(.A(l), .Y(mai_mai_n1545_));
  INV        m1515(.A(f), .Y(mai_mai_n1546_));
  INV        m1516(.A(j), .Y(mai_mai_n1547_));
  INV        m1517(.A(mai_mai_n480_), .Y(mai_mai_n1548_));
  INV        m1518(.A(m), .Y(mai_mai_n1549_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  NA3        u0002(.A(e), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n31_));
  NOi32      u0003(.An(m), .Bn(l), .C(n), .Y(men_men_n32_));
  NOi32      u0004(.An(i), .Bn(u), .C(h), .Y(men_men_n33_));
  NA2        u0005(.A(men_men_n33_), .B(men_men_n32_), .Y(men_men_n34_));
  AN2        u0006(.A(m), .B(l), .Y(men_men_n35_));
  NOi32      u0007(.An(j), .Bn(u), .C(k), .Y(men_men_n36_));
  NA2        u0008(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n37_));
  NO2        u0009(.A(men_men_n37_), .B(n), .Y(men_men_n38_));
  INV        u0010(.A(h), .Y(men_men_n39_));
  NAi21      u0011(.An(j), .B(l), .Y(men_men_n40_));
  NAi32      u0012(.An(n), .Bn(u), .C(m), .Y(men_men_n41_));
  NO3        u0013(.A(men_men_n41_), .B(men_men_n40_), .C(men_men_n39_), .Y(men_men_n42_));
  NAi31      u0014(.An(n), .B(m), .C(l), .Y(men_men_n43_));
  INV        u0015(.A(i), .Y(men_men_n44_));
  AN2        u0016(.A(h), .B(u), .Y(men_men_n45_));
  NA2        u0017(.A(men_men_n45_), .B(men_men_n44_), .Y(men_men_n46_));
  NO2        u0018(.A(men_men_n46_), .B(men_men_n43_), .Y(men_men_n47_));
  NAi21      u0019(.An(n), .B(m), .Y(men_men_n48_));
  NOi32      u0020(.An(k), .Bn(h), .C(l), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(u), .Y(men_men_n50_));
  NO2        u0022(.A(men_men_n50_), .B(men_men_n49_), .Y(men_men_n51_));
  NO4        u0023(.A(men_men_n50_), .B(men_men_n47_), .C(men_men_n42_), .D(men_men_n38_), .Y(men_men_n52_));
  AOI210     u0024(.A0(men_men_n52_), .A1(men_men_n34_), .B0(men_men_n31_), .Y(men_men_n53_));
  INV        u0025(.A(c), .Y(men_men_n54_));
  NA2        u0026(.A(e), .B(b), .Y(men_men_n55_));
  NO2        u0027(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  INV        u0028(.A(d), .Y(men_men_n57_));
  NA2        u0029(.A(u), .B(men_men_n57_), .Y(men_men_n58_));
  NAi21      u0030(.An(i), .B(h), .Y(men_men_n59_));
  NAi31      u0031(.An(i), .B(l), .C(j), .Y(men_men_n60_));
  OAI220     u0032(.A0(men_men_n60_), .A1(men_men_n48_), .B0(men_men_n59_), .B1(men_men_n43_), .Y(men_men_n61_));
  NAi31      u0033(.An(men_men_n58_), .B(men_men_n61_), .C(men_men_n56_), .Y(men_men_n62_));
  NAi41      u0034(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n63_));
  NA2        u0035(.A(u), .B(f), .Y(men_men_n64_));
  NO2        u0036(.A(men_men_n64_), .B(men_men_n63_), .Y(men_men_n65_));
  NAi21      u0037(.An(i), .B(j), .Y(men_men_n66_));
  NAi32      u0038(.An(n), .Bn(k), .C(m), .Y(men_men_n67_));
  NO2        u0039(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n68_));
  NAi31      u0040(.An(l), .B(m), .C(k), .Y(men_men_n69_));
  NAi21      u0041(.An(e), .B(h), .Y(men_men_n70_));
  NAi41      u0042(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n71_));
  NA2        u0043(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n72_));
  INV        u0044(.A(m), .Y(men_men_n73_));
  NOi21      u0045(.An(k), .B(l), .Y(men_men_n74_));
  NA2        u0046(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n75_));
  AN4        u0047(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n76_));
  NA2        u0048(.A(h), .B(men_men_n76_), .Y(men_men_n77_));
  NAi32      u0049(.An(m), .Bn(k), .C(j), .Y(men_men_n78_));
  NOi32      u0050(.An(h), .Bn(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n72_), .B(men_men_n62_), .Y(men_men_n80_));
  INV        u0052(.A(n), .Y(men_men_n81_));
  INV        u0053(.A(j), .Y(men_men_n82_));
  AN3        u0054(.A(m), .B(k), .C(i), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n82_), .C(u), .Y(men_men_n84_));
  NO2        u0056(.A(men_men_n84_), .B(f), .Y(men_men_n85_));
  NAi32      u0057(.An(u), .Bn(f), .C(h), .Y(men_men_n86_));
  NAi31      u0058(.An(j), .B(m), .C(l), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  NA2        u0060(.A(m), .B(l), .Y(men_men_n89_));
  NAi31      u0061(.An(k), .B(j), .C(u), .Y(men_men_n90_));
  NO3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(f), .Y(men_men_n91_));
  AN2        u0063(.A(j), .B(u), .Y(men_men_n92_));
  NOi32      u0064(.An(m), .Bn(l), .C(i), .Y(men_men_n93_));
  NOi21      u0065(.An(u), .B(i), .Y(men_men_n94_));
  NOi32      u0066(.An(m), .Bn(j), .C(k), .Y(men_men_n95_));
  AOI220     u0067(.A0(men_men_n95_), .A1(men_men_n94_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n96_));
  NO2        u0068(.A(men_men_n96_), .B(f), .Y(men_men_n97_));
  NAi41      u0069(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n98_));
  AN2        u0070(.A(e), .B(b), .Y(men_men_n99_));
  NA2        u0071(.A(c), .B(men_men_n99_), .Y(men_men_n100_));
  NOi21      u0072(.An(u), .B(f), .Y(men_men_n101_));
  NOi21      u0073(.An(i), .B(h), .Y(men_men_n102_));
  NA3        u0074(.A(men_men_n102_), .B(men_men_n101_), .C(men_men_n35_), .Y(men_men_n103_));
  INV        u0075(.A(a), .Y(men_men_n104_));
  NA2        u0076(.A(men_men_n99_), .B(men_men_n104_), .Y(men_men_n105_));
  INV        u0077(.A(l), .Y(men_men_n106_));
  NOi21      u0078(.An(m), .B(n), .Y(men_men_n107_));
  AN2        u0079(.A(k), .B(h), .Y(men_men_n108_));
  INV        u0080(.A(b), .Y(men_men_n109_));
  NA2        u0081(.A(l), .B(j), .Y(men_men_n110_));
  AN2        u0082(.A(k), .B(i), .Y(men_men_n111_));
  NA2        u0083(.A(men_men_n111_), .B(men_men_n110_), .Y(men_men_n112_));
  NA2        u0084(.A(u), .B(e), .Y(men_men_n113_));
  NOi32      u0085(.An(c), .Bn(a), .C(d), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n114_), .B(men_men_n107_), .Y(men_men_n115_));
  NO4        u0087(.A(men_men_n115_), .B(men_men_n113_), .C(men_men_n112_), .D(men_men_n109_), .Y(men_men_n116_));
  NOi31      u0088(.An(k), .B(m), .C(j), .Y(men_men_n117_));
  NOi31      u0089(.An(k), .B(m), .C(i), .Y(men_men_n118_));
  NA3        u0090(.A(men_men_n118_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n119_));
  NOi32      u0091(.An(f), .Bn(b), .C(e), .Y(men_men_n120_));
  NAi21      u0092(.An(u), .B(h), .Y(men_men_n121_));
  NAi21      u0093(.An(m), .B(n), .Y(men_men_n122_));
  NO3        u0094(.A(j), .B(men_men_n122_), .C(men_men_n121_), .Y(men_men_n123_));
  NAi31      u0095(.An(j), .B(k), .C(h), .Y(men_men_n124_));
  NA2        u0096(.A(men_men_n123_), .B(men_men_n120_), .Y(men_men_n125_));
  NO2        u0097(.A(k), .B(j), .Y(men_men_n126_));
  INV        u0098(.A(men_men_n122_), .Y(men_men_n127_));
  AN2        u0099(.A(k), .B(j), .Y(men_men_n128_));
  NAi21      u0100(.An(c), .B(b), .Y(men_men_n129_));
  NA2        u0101(.A(f), .B(d), .Y(men_men_n130_));
  NO3        u0102(.A(men_men_n130_), .B(men_men_n129_), .C(men_men_n121_), .Y(men_men_n131_));
  NA2        u0103(.A(men_men_n131_), .B(men_men_n127_), .Y(men_men_n132_));
  NA2        u0104(.A(d), .B(b), .Y(men_men_n133_));
  NAi21      u0105(.An(e), .B(f), .Y(men_men_n134_));
  NO2        u0106(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NA2        u0107(.A(b), .B(a), .Y(men_men_n136_));
  NAi21      u0108(.An(e), .B(u), .Y(men_men_n137_));
  NAi21      u0109(.An(c), .B(d), .Y(men_men_n138_));
  NAi31      u0110(.An(l), .B(k), .C(h), .Y(men_men_n139_));
  NA2        u0111(.A(men_men_n132_), .B(men_men_n125_), .Y(men_men_n140_));
  NAi31      u0112(.An(e), .B(f), .C(b), .Y(men_men_n141_));
  NOi21      u0113(.An(u), .B(d), .Y(men_men_n142_));
  NO2        u0114(.A(men_men_n142_), .B(men_men_n141_), .Y(men_men_n143_));
  NOi21      u0115(.An(h), .B(i), .Y(men_men_n144_));
  NOi21      u0116(.An(k), .B(m), .Y(men_men_n145_));
  NA3        u0117(.A(men_men_n145_), .B(men_men_n144_), .C(n), .Y(men_men_n146_));
  NOi21      u0118(.An(men_men_n143_), .B(men_men_n146_), .Y(men_men_n147_));
  NOi21      u0119(.An(h), .B(u), .Y(men_men_n148_));
  NAi31      u0120(.An(l), .B(j), .C(h), .Y(men_men_n149_));
  NO2        u0121(.A(men_men_n149_), .B(men_men_n48_), .Y(men_men_n150_));
  NA2        u0122(.A(men_men_n150_), .B(men_men_n65_), .Y(men_men_n151_));
  NOi32      u0123(.An(n), .Bn(k), .C(m), .Y(men_men_n152_));
  NA2        u0124(.A(l), .B(i), .Y(men_men_n153_));
  INV        u0125(.A(men_men_n151_), .Y(men_men_n154_));
  NA2        u0126(.A(j), .B(h), .Y(men_men_n155_));
  OR3        u0127(.A(n), .B(m), .C(k), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  NAi32      u0129(.An(m), .Bn(k), .C(n), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n158_), .B(men_men_n155_), .Y(men_men_n159_));
  AOI220     u0131(.A0(men_men_n159_), .A1(men_men_n143_), .B0(men_men_n157_), .B1(f), .Y(men_men_n160_));
  NO2        u0132(.A(n), .B(m), .Y(men_men_n161_));
  NA2        u0133(.A(men_men_n161_), .B(men_men_n49_), .Y(men_men_n162_));
  NAi21      u0134(.An(f), .B(e), .Y(men_men_n163_));
  NA2        u0135(.A(d), .B(c), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NOi21      u0137(.An(men_men_n165_), .B(men_men_n162_), .Y(men_men_n166_));
  NAi21      u0138(.An(d), .B(c), .Y(men_men_n167_));
  NAi31      u0139(.An(m), .B(n), .C(b), .Y(men_men_n168_));
  NA2        u0140(.A(k), .B(i), .Y(men_men_n169_));
  NAi21      u0141(.An(h), .B(f), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NO2        u0143(.A(men_men_n168_), .B(men_men_n138_), .Y(men_men_n172_));
  NA2        u0144(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  NOi32      u0145(.An(f), .Bn(c), .C(d), .Y(men_men_n174_));
  NOi32      u0146(.An(f), .Bn(c), .C(e), .Y(men_men_n175_));
  NO2        u0147(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  NO3        u0148(.A(n), .B(m), .C(j), .Y(men_men_n177_));
  NA2        u0149(.A(men_men_n177_), .B(men_men_n108_), .Y(men_men_n178_));
  AO210      u0150(.A0(men_men_n178_), .A1(men_men_n162_), .B0(men_men_n176_), .Y(men_men_n179_));
  NAi41      u0151(.An(men_men_n166_), .B(men_men_n179_), .C(men_men_n173_), .D(men_men_n160_), .Y(men_men_n180_));
  OR4        u0152(.A(men_men_n180_), .B(men_men_n154_), .C(men_men_n147_), .D(men_men_n140_), .Y(men_men_n181_));
  NO4        u0153(.A(men_men_n181_), .B(men_men_n116_), .C(men_men_n80_), .D(men_men_n53_), .Y(men_men_n182_));
  NA3        u0154(.A(m), .B(men_men_n106_), .C(j), .Y(men_men_n183_));
  NAi31      u0155(.An(n), .B(h), .C(u), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NOi32      u0157(.An(m), .Bn(k), .C(l), .Y(men_men_n186_));
  NA3        u0158(.A(men_men_n186_), .B(men_men_n82_), .C(u), .Y(men_men_n187_));
  NO2        u0159(.A(men_men_n187_), .B(n), .Y(men_men_n188_));
  NOi21      u0160(.An(k), .B(j), .Y(men_men_n189_));
  NA4        u0161(.A(men_men_n189_), .B(men_men_n107_), .C(i), .D(u), .Y(men_men_n190_));
  AN2        u0162(.A(i), .B(u), .Y(men_men_n191_));
  NA3        u0163(.A(men_men_n74_), .B(men_men_n191_), .C(men_men_n107_), .Y(men_men_n192_));
  NA2        u0164(.A(men_men_n192_), .B(men_men_n190_), .Y(men_men_n193_));
  NO3        u0165(.A(men_men_n193_), .B(men_men_n188_), .C(men_men_n185_), .Y(men_men_n194_));
  NAi41      u0166(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n195_));
  INV        u0167(.A(f), .Y(men_men_n196_));
  INV        u0168(.A(u), .Y(men_men_n197_));
  NOi31      u0169(.An(i), .B(j), .C(h), .Y(men_men_n198_));
  NOi21      u0170(.An(l), .B(m), .Y(men_men_n199_));
  NA2        u0171(.A(men_men_n199_), .B(men_men_n198_), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n194_), .B(men_men_n31_), .Y(men_men_n201_));
  NOi21      u0173(.An(n), .B(m), .Y(men_men_n202_));
  NOi32      u0174(.An(l), .Bn(i), .C(j), .Y(men_men_n203_));
  NA2        u0175(.A(men_men_n203_), .B(men_men_n202_), .Y(men_men_n204_));
  OA220      u0176(.A0(men_men_n204_), .A1(men_men_n100_), .B0(men_men_n78_), .B1(men_men_n77_), .Y(men_men_n205_));
  NAi21      u0177(.An(j), .B(h), .Y(men_men_n206_));
  XN2        u0178(.A(i), .B(h), .Y(men_men_n207_));
  NA2        u0179(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NOi31      u0180(.An(k), .B(n), .C(m), .Y(men_men_n209_));
  NOi31      u0181(.An(men_men_n209_), .B(men_men_n164_), .C(men_men_n163_), .Y(men_men_n210_));
  NA2        u0182(.A(men_men_n210_), .B(men_men_n208_), .Y(men_men_n211_));
  NAi31      u0183(.An(f), .B(e), .C(c), .Y(men_men_n212_));
  NO4        u0184(.A(men_men_n212_), .B(men_men_n156_), .C(men_men_n155_), .D(men_men_n57_), .Y(men_men_n213_));
  NA4        u0185(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n214_));
  NAi32      u0186(.An(m), .Bn(i), .C(k), .Y(men_men_n215_));
  NO3        u0187(.A(men_men_n215_), .B(men_men_n86_), .C(men_men_n214_), .Y(men_men_n216_));
  INV        u0188(.A(k), .Y(men_men_n217_));
  NO2        u0189(.A(men_men_n216_), .B(men_men_n213_), .Y(men_men_n218_));
  NAi21      u0190(.An(n), .B(a), .Y(men_men_n219_));
  NO2        u0191(.A(men_men_n219_), .B(men_men_n133_), .Y(men_men_n220_));
  NAi41      u0192(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n221_));
  NO2        u0193(.A(men_men_n221_), .B(e), .Y(men_men_n222_));
  NO3        u0194(.A(men_men_n134_), .B(men_men_n90_), .C(men_men_n89_), .Y(men_men_n223_));
  OAI210     u0195(.A0(men_men_n223_), .A1(men_men_n222_), .B0(men_men_n220_), .Y(men_men_n224_));
  AN4        u0196(.A(men_men_n224_), .B(men_men_n218_), .C(men_men_n211_), .D(men_men_n205_), .Y(men_men_n225_));
  NO2        u0197(.A(h), .B(men_men_n98_), .Y(men_men_n226_));
  NA2        u0198(.A(men_men_n226_), .B(men_men_n120_), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n145_), .B(men_men_n102_), .Y(men_men_n228_));
  NO2        u0200(.A(n), .B(a), .Y(men_men_n229_));
  NAi31      u0201(.An(men_men_n221_), .B(men_men_n229_), .C(men_men_n99_), .Y(men_men_n230_));
  NAi21      u0202(.An(h), .B(i), .Y(men_men_n231_));
  NA2        u0203(.A(men_men_n161_), .B(k), .Y(men_men_n232_));
  NO2        u0204(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  NA2        u0205(.A(men_men_n233_), .B(men_men_n174_), .Y(men_men_n234_));
  NA3        u0206(.A(men_men_n234_), .B(men_men_n230_), .C(men_men_n227_), .Y(men_men_n235_));
  NOi21      u0207(.An(u), .B(e), .Y(men_men_n236_));
  NO2        u0208(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n237_));
  NA2        u0209(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  NOi32      u0210(.An(l), .Bn(j), .C(i), .Y(men_men_n239_));
  AOI210     u0211(.A0(men_men_n74_), .A1(men_men_n82_), .B0(men_men_n239_), .Y(men_men_n240_));
  NO2        u0212(.A(men_men_n231_), .B(men_men_n43_), .Y(men_men_n241_));
  NAi21      u0213(.An(f), .B(u), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n242_), .B(men_men_n63_), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n67_), .B(men_men_n110_), .Y(men_men_n244_));
  AOI220     u0216(.A0(men_men_n244_), .A1(men_men_n243_), .B0(men_men_n241_), .B1(men_men_n65_), .Y(men_men_n245_));
  OAI210     u0217(.A0(men_men_n240_), .A1(men_men_n238_), .B0(men_men_n245_), .Y(men_men_n246_));
  NO3        u0218(.A(j), .B(men_men_n48_), .C(men_men_n44_), .Y(men_men_n247_));
  NOi41      u0219(.An(men_men_n225_), .B(men_men_n246_), .C(men_men_n235_), .D(men_men_n201_), .Y(men_men_n248_));
  NO4        u0220(.A(men_men_n185_), .B(men_men_n47_), .C(men_men_n42_), .D(men_men_n38_), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(men_men_n105_), .Y(men_men_n250_));
  NAi21      u0222(.An(h), .B(u), .Y(men_men_n251_));
  NA2        u0223(.A(men_men_n145_), .B(men_men_n76_), .Y(men_men_n252_));
  NAi31      u0224(.An(u), .B(k), .C(h), .Y(men_men_n253_));
  NO3        u0225(.A(men_men_n122_), .B(men_men_n253_), .C(l), .Y(men_men_n254_));
  NAi31      u0226(.An(e), .B(d), .C(a), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n254_), .B(men_men_n120_), .Y(men_men_n256_));
  NA2        u0228(.A(men_men_n256_), .B(men_men_n252_), .Y(men_men_n257_));
  NA4        u0229(.A(men_men_n145_), .B(men_men_n79_), .C(men_men_n76_), .D(men_men_n110_), .Y(men_men_n258_));
  NA3        u0230(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n81_), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n176_), .Y(men_men_n260_));
  NOi21      u0232(.An(men_men_n258_), .B(men_men_n260_), .Y(men_men_n261_));
  NA3        u0233(.A(e), .B(c), .C(b), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n58_), .B(men_men_n262_), .Y(men_men_n263_));
  NAi32      u0235(.An(k), .Bn(i), .C(j), .Y(men_men_n264_));
  NAi31      u0236(.An(h), .B(l), .C(i), .Y(men_men_n265_));
  NA3        u0237(.A(men_men_n265_), .B(men_men_n264_), .C(men_men_n149_), .Y(men_men_n266_));
  NOi21      u0238(.An(men_men_n266_), .B(men_men_n48_), .Y(men_men_n267_));
  OAI210     u0239(.A0(men_men_n243_), .A1(men_men_n263_), .B0(men_men_n267_), .Y(men_men_n268_));
  NAi21      u0240(.An(l), .B(k), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n269_), .B(men_men_n48_), .Y(men_men_n270_));
  NOi21      u0242(.An(l), .B(j), .Y(men_men_n271_));
  NA2        u0243(.A(men_men_n148_), .B(men_men_n271_), .Y(men_men_n272_));
  NA3        u0244(.A(men_men_n111_), .B(men_men_n110_), .C(u), .Y(men_men_n273_));
  OR3        u0245(.A(men_men_n71_), .B(men_men_n73_), .C(e), .Y(men_men_n274_));
  AOI210     u0246(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n274_), .Y(men_men_n275_));
  INV        u0247(.A(men_men_n275_), .Y(men_men_n276_));
  NAi32      u0248(.An(j), .Bn(h), .C(i), .Y(men_men_n277_));
  NAi21      u0249(.An(m), .B(l), .Y(men_men_n278_));
  NO3        u0250(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n81_), .Y(men_men_n279_));
  NA2        u0251(.A(h), .B(u), .Y(men_men_n280_));
  NA2        u0252(.A(men_men_n279_), .B(b), .Y(men_men_n281_));
  NA4        u0253(.A(men_men_n281_), .B(men_men_n276_), .C(men_men_n268_), .D(men_men_n261_), .Y(men_men_n282_));
  NO2        u0254(.A(men_men_n100_), .B(men_men_n98_), .Y(men_men_n283_));
  NAi32      u0255(.An(n), .Bn(m), .C(l), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n284_), .B(men_men_n277_), .Y(men_men_n285_));
  NA2        u0257(.A(men_men_n285_), .B(men_men_n165_), .Y(men_men_n286_));
  NO2        u0258(.A(men_men_n115_), .B(men_men_n109_), .Y(men_men_n287_));
  NAi31      u0259(.An(k), .B(l), .C(j), .Y(men_men_n288_));
  OAI210     u0260(.A0(men_men_n269_), .A1(j), .B0(men_men_n288_), .Y(men_men_n289_));
  NOi21      u0261(.An(men_men_n289_), .B(men_men_n113_), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n290_), .B(men_men_n287_), .Y(men_men_n291_));
  NA2        u0263(.A(men_men_n291_), .B(men_men_n286_), .Y(men_men_n292_));
  NO4        u0264(.A(men_men_n292_), .B(men_men_n282_), .C(men_men_n257_), .D(men_men_n250_), .Y(men_men_n293_));
  NA2        u0265(.A(men_men_n233_), .B(men_men_n175_), .Y(men_men_n294_));
  NAi21      u0266(.An(m), .B(k), .Y(men_men_n295_));
  NO2        u0267(.A(men_men_n207_), .B(men_men_n295_), .Y(men_men_n296_));
  NAi41      u0268(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n297_), .B(men_men_n137_), .Y(men_men_n298_));
  NA2        u0270(.A(men_men_n298_), .B(men_men_n296_), .Y(men_men_n299_));
  NAi31      u0271(.An(i), .B(l), .C(h), .Y(men_men_n300_));
  NO4        u0272(.A(men_men_n300_), .B(men_men_n137_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n301_));
  NA2        u0273(.A(e), .B(c), .Y(men_men_n302_));
  NOi21      u0274(.An(f), .B(h), .Y(men_men_n303_));
  NA2        u0275(.A(men_men_n303_), .B(men_men_n111_), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n304_), .B(men_men_n197_), .Y(men_men_n305_));
  NAi31      u0277(.An(d), .B(e), .C(b), .Y(men_men_n306_));
  NO2        u0278(.A(men_men_n122_), .B(men_men_n306_), .Y(men_men_n307_));
  NA2        u0279(.A(men_men_n307_), .B(men_men_n305_), .Y(men_men_n308_));
  NAi41      u0280(.An(men_men_n301_), .B(men_men_n308_), .C(men_men_n299_), .D(men_men_n294_), .Y(men_men_n309_));
  NO4        u0281(.A(men_men_n297_), .B(men_men_n78_), .C(men_men_n70_), .D(men_men_n197_), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n229_), .B(men_men_n99_), .Y(men_men_n311_));
  OR2        u0283(.A(men_men_n311_), .B(men_men_n187_), .Y(men_men_n312_));
  NOi31      u0284(.An(l), .B(n), .C(m), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n198_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n314_), .B(men_men_n176_), .Y(men_men_n315_));
  NAi32      u0287(.An(men_men_n315_), .Bn(men_men_n310_), .C(men_men_n312_), .Y(men_men_n316_));
  NAi32      u0288(.An(m), .Bn(j), .C(k), .Y(men_men_n317_));
  NAi41      u0289(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n318_));
  NOi31      u0290(.An(j), .B(m), .C(k), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n117_), .B(men_men_n319_), .Y(men_men_n320_));
  AN3        u0292(.A(h), .B(u), .C(f), .Y(men_men_n321_));
  NAi31      u0293(.An(men_men_n320_), .B(men_men_n321_), .C(b), .Y(men_men_n322_));
  NOi32      u0294(.An(m), .Bn(j), .C(l), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n323_), .B(men_men_n93_), .Y(men_men_n324_));
  NO2        u0296(.A(men_men_n278_), .B(men_men_n277_), .Y(men_men_n325_));
  NO2        u0297(.A(men_men_n200_), .B(u), .Y(men_men_n326_));
  NA2        u0298(.A(f), .B(men_men_n326_), .Y(men_men_n327_));
  INV        u0299(.A(men_men_n215_), .Y(men_men_n328_));
  NA3        u0300(.A(men_men_n328_), .B(men_men_n321_), .C(b), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n329_), .B(men_men_n322_), .Y(men_men_n330_));
  NA3        u0302(.A(h), .B(u), .C(f), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n331_), .B(men_men_n75_), .Y(men_men_n332_));
  NA2        u0304(.A(men_men_n148_), .B(e), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n333_), .B(men_men_n40_), .Y(men_men_n334_));
  AOI220     u0306(.A0(men_men_n334_), .A1(men_men_n287_), .B0(b), .B1(men_men_n332_), .Y(men_men_n335_));
  NOi32      u0307(.An(j), .Bn(u), .C(i), .Y(men_men_n336_));
  NA3        u0308(.A(men_men_n336_), .B(men_men_n269_), .C(men_men_n107_), .Y(men_men_n337_));
  AO210      u0309(.A0(men_men_n105_), .A1(men_men_n31_), .B0(men_men_n337_), .Y(men_men_n338_));
  NOi32      u0310(.An(e), .Bn(b), .C(a), .Y(men_men_n339_));
  AN2        u0311(.A(l), .B(j), .Y(men_men_n340_));
  INV        u0312(.A(men_men_n295_), .Y(men_men_n341_));
  NO3        u0313(.A(men_men_n297_), .B(men_men_n70_), .C(men_men_n197_), .Y(men_men_n342_));
  NA3        u0314(.A(men_men_n192_), .B(men_men_n190_), .C(men_men_n34_), .Y(men_men_n343_));
  AOI220     u0315(.A0(men_men_n343_), .A1(men_men_n339_), .B0(men_men_n342_), .B1(men_men_n341_), .Y(men_men_n344_));
  NA2        u0316(.A(men_men_n191_), .B(k), .Y(men_men_n345_));
  NA3        u0317(.A(m), .B(men_men_n106_), .C(men_men_n196_), .Y(men_men_n346_));
  NA4        u0318(.A(men_men_n186_), .B(men_men_n82_), .C(u), .D(men_men_n196_), .Y(men_men_n347_));
  NAi41      u0319(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n348_));
  NA2        u0320(.A(men_men_n50_), .B(men_men_n107_), .Y(men_men_n349_));
  NO2        u0321(.A(men_men_n349_), .B(men_men_n348_), .Y(men_men_n350_));
  NA2        u0322(.A(men_men_n350_), .B(b), .Y(men_men_n351_));
  NA4        u0323(.A(men_men_n351_), .B(men_men_n344_), .C(men_men_n338_), .D(men_men_n335_), .Y(men_men_n352_));
  NO4        u0324(.A(men_men_n352_), .B(men_men_n330_), .C(men_men_n316_), .D(men_men_n309_), .Y(men_men_n353_));
  NA4        u0325(.A(men_men_n353_), .B(men_men_n293_), .C(men_men_n248_), .D(men_men_n182_), .Y(men10));
  NA3        u0326(.A(m), .B(k), .C(i), .Y(men_men_n355_));
  NO3        u0327(.A(men_men_n355_), .B(j), .C(men_men_n197_), .Y(men_men_n356_));
  NOi21      u0328(.An(e), .B(f), .Y(men_men_n357_));
  NO4        u0329(.A(men_men_n138_), .B(men_men_n357_), .C(n), .D(men_men_n104_), .Y(men_men_n358_));
  NOi32      u0330(.An(k), .Bn(h), .C(j), .Y(men_men_n359_));
  NA2        u0331(.A(men_men_n359_), .B(men_men_n202_), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n146_), .B(men_men_n360_), .Y(men_men_n361_));
  AOI220     u0333(.A0(men_men_n361_), .A1(f), .B0(men_men_n358_), .B1(men_men_n356_), .Y(men_men_n362_));
  AN2        u0334(.A(j), .B(h), .Y(men_men_n363_));
  NO3        u0335(.A(n), .B(m), .C(k), .Y(men_men_n364_));
  NA2        u0336(.A(men_men_n364_), .B(men_men_n363_), .Y(men_men_n365_));
  NO3        u0337(.A(men_men_n365_), .B(men_men_n138_), .C(men_men_n196_), .Y(men_men_n366_));
  NO2        u0338(.A(men_men_n155_), .B(m), .Y(men_men_n367_));
  NA4        u0339(.A(n), .B(f), .C(c), .D(men_men_n109_), .Y(men_men_n368_));
  NOi21      u0340(.An(men_men_n367_), .B(men_men_n368_), .Y(men_men_n369_));
  NOi32      u0341(.An(d), .Bn(a), .C(c), .Y(men_men_n370_));
  NA2        u0342(.A(men_men_n370_), .B(men_men_n163_), .Y(men_men_n371_));
  NAi21      u0343(.An(i), .B(u), .Y(men_men_n372_));
  NAi31      u0344(.An(k), .B(m), .C(j), .Y(men_men_n373_));
  NO3        u0345(.A(men_men_n373_), .B(men_men_n372_), .C(n), .Y(men_men_n374_));
  NOi21      u0346(.An(men_men_n374_), .B(men_men_n371_), .Y(men_men_n375_));
  NO3        u0347(.A(men_men_n375_), .B(men_men_n369_), .C(men_men_n366_), .Y(men_men_n376_));
  NA2        u0348(.A(f), .B(men_men_n285_), .Y(men_men_n377_));
  NA3        u0349(.A(men_men_n377_), .B(men_men_n376_), .C(men_men_n362_), .Y(men_men_n378_));
  NO2        u0350(.A(men_men_n57_), .B(men_men_n109_), .Y(men_men_n379_));
  NA2        u0351(.A(men_men_n229_), .B(men_men_n379_), .Y(men_men_n380_));
  INV        u0352(.A(e), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n45_), .B(e), .Y(men_men_n382_));
  OAI220     u0354(.A0(men_men_n382_), .A1(men_men_n183_), .B0(men_men_n187_), .B1(men_men_n381_), .Y(men_men_n383_));
  AN2        u0355(.A(u), .B(e), .Y(men_men_n384_));
  NA3        u0356(.A(men_men_n384_), .B(men_men_n186_), .C(i), .Y(men_men_n385_));
  OAI210     u0357(.A0(men_men_n84_), .A1(men_men_n381_), .B0(men_men_n385_), .Y(men_men_n386_));
  NO2        u0358(.A(men_men_n96_), .B(men_men_n381_), .Y(men_men_n387_));
  NO3        u0359(.A(men_men_n387_), .B(men_men_n386_), .C(men_men_n383_), .Y(men_men_n388_));
  NOi32      u0360(.An(h), .Bn(e), .C(u), .Y(men_men_n389_));
  NA3        u0361(.A(men_men_n389_), .B(men_men_n271_), .C(m), .Y(men_men_n390_));
  NOi21      u0362(.An(u), .B(h), .Y(men_men_n391_));
  AN3        u0363(.A(m), .B(l), .C(i), .Y(men_men_n392_));
  NA3        u0364(.A(men_men_n392_), .B(men_men_n391_), .C(e), .Y(men_men_n393_));
  AN3        u0365(.A(h), .B(u), .C(e), .Y(men_men_n394_));
  NA2        u0366(.A(men_men_n394_), .B(men_men_n93_), .Y(men_men_n395_));
  AN3        u0367(.A(men_men_n395_), .B(men_men_n393_), .C(men_men_n390_), .Y(men_men_n396_));
  AOI210     u0368(.A0(men_men_n396_), .A1(men_men_n388_), .B0(men_men_n380_), .Y(men_men_n397_));
  NA3        u0369(.A(men_men_n36_), .B(men_men_n35_), .C(e), .Y(men_men_n398_));
  NO2        u0370(.A(men_men_n398_), .B(men_men_n380_), .Y(men_men_n399_));
  NA3        u0371(.A(men_men_n370_), .B(men_men_n163_), .C(men_men_n81_), .Y(men_men_n400_));
  NAi31      u0372(.An(b), .B(c), .C(a), .Y(men_men_n401_));
  NO2        u0373(.A(men_men_n401_), .B(n), .Y(men_men_n402_));
  OAI210     u0374(.A0(men_men_n50_), .A1(men_men_n49_), .B0(m), .Y(men_men_n403_));
  NO2        u0375(.A(men_men_n403_), .B(men_men_n134_), .Y(men_men_n404_));
  NA2        u0376(.A(men_men_n404_), .B(men_men_n402_), .Y(men_men_n405_));
  INV        u0377(.A(men_men_n405_), .Y(men_men_n406_));
  NO4        u0378(.A(men_men_n406_), .B(men_men_n399_), .C(men_men_n397_), .D(men_men_n378_), .Y(men_men_n407_));
  NA2        u0379(.A(i), .B(u), .Y(men_men_n408_));
  NO3        u0380(.A(men_men_n255_), .B(men_men_n408_), .C(c), .Y(men_men_n409_));
  NOi21      u0381(.An(a), .B(n), .Y(men_men_n410_));
  NOi21      u0382(.An(d), .B(c), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n411_), .B(men_men_n410_), .Y(men_men_n412_));
  NA3        u0384(.A(i), .B(u), .C(f), .Y(men_men_n413_));
  OR2        u0385(.A(men_men_n413_), .B(men_men_n69_), .Y(men_men_n414_));
  NA3        u0386(.A(men_men_n392_), .B(men_men_n391_), .C(men_men_n163_), .Y(men_men_n415_));
  AOI210     u0387(.A0(men_men_n415_), .A1(men_men_n414_), .B0(men_men_n412_), .Y(men_men_n416_));
  AOI210     u0388(.A0(men_men_n409_), .A1(men_men_n270_), .B0(men_men_n416_), .Y(men_men_n417_));
  OR2        u0389(.A(n), .B(m), .Y(men_men_n418_));
  NO2        u0390(.A(men_men_n418_), .B(men_men_n139_), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n164_), .B(men_men_n134_), .Y(men_men_n420_));
  OAI210     u0392(.A0(men_men_n419_), .A1(men_men_n157_), .B0(men_men_n420_), .Y(men_men_n421_));
  INV        u0393(.A(men_men_n349_), .Y(men_men_n422_));
  NA3        u0394(.A(men_men_n422_), .B(men_men_n339_), .C(d), .Y(men_men_n423_));
  NO2        u0395(.A(men_men_n401_), .B(men_men_n48_), .Y(men_men_n424_));
  NO3        u0396(.A(men_men_n64_), .B(men_men_n106_), .C(e), .Y(men_men_n425_));
  NAi21      u0397(.An(k), .B(j), .Y(men_men_n426_));
  NA2        u0398(.A(men_men_n231_), .B(men_men_n426_), .Y(men_men_n427_));
  NA3        u0399(.A(men_men_n427_), .B(men_men_n425_), .C(men_men_n424_), .Y(men_men_n428_));
  NAi21      u0400(.An(e), .B(d), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n232_), .B(men_men_n196_), .Y(men_men_n430_));
  NA3        u0402(.A(men_men_n430_), .B(d), .C(men_men_n208_), .Y(men_men_n431_));
  NA4        u0403(.A(men_men_n431_), .B(men_men_n428_), .C(men_men_n423_), .D(men_men_n421_), .Y(men_men_n432_));
  NO2        u0404(.A(men_men_n314_), .B(men_men_n196_), .Y(men_men_n433_));
  NOi31      u0405(.An(n), .B(m), .C(k), .Y(men_men_n434_));
  AOI220     u0406(.A0(men_men_n434_), .A1(men_men_n363_), .B0(men_men_n202_), .B1(men_men_n49_), .Y(men_men_n435_));
  NAi31      u0407(.An(u), .B(f), .C(c), .Y(men_men_n436_));
  OR3        u0408(.A(men_men_n436_), .B(men_men_n435_), .C(e), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n437_), .B(men_men_n286_), .Y(men_men_n438_));
  NOi41      u0410(.An(men_men_n417_), .B(men_men_n438_), .C(men_men_n432_), .D(men_men_n246_), .Y(men_men_n439_));
  NOi32      u0411(.An(c), .Bn(a), .C(b), .Y(men_men_n440_));
  NA2        u0412(.A(men_men_n440_), .B(men_men_n107_), .Y(men_men_n441_));
  INV        u0413(.A(men_men_n253_), .Y(men_men_n442_));
  AN2        u0414(.A(e), .B(d), .Y(men_men_n443_));
  NA2        u0415(.A(men_men_n443_), .B(men_men_n442_), .Y(men_men_n444_));
  INV        u0416(.A(men_men_n134_), .Y(men_men_n445_));
  NO2        u0417(.A(men_men_n121_), .B(men_men_n40_), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n64_), .B(e), .Y(men_men_n447_));
  NOi31      u0419(.An(j), .B(k), .C(i), .Y(men_men_n448_));
  NOi21      u0420(.An(men_men_n149_), .B(men_men_n448_), .Y(men_men_n449_));
  NA4        u0421(.A(men_men_n300_), .B(men_men_n449_), .C(men_men_n240_), .D(men_men_n112_), .Y(men_men_n450_));
  AOI220     u0422(.A0(men_men_n450_), .A1(men_men_n447_), .B0(men_men_n446_), .B1(men_men_n445_), .Y(men_men_n451_));
  AOI210     u0423(.A0(men_men_n451_), .A1(men_men_n444_), .B0(men_men_n441_), .Y(men_men_n452_));
  NO2        u0424(.A(men_men_n193_), .B(men_men_n188_), .Y(men_men_n453_));
  NOi21      u0425(.An(a), .B(b), .Y(men_men_n454_));
  NA3        u0426(.A(e), .B(d), .C(c), .Y(men_men_n455_));
  NAi21      u0427(.An(men_men_n455_), .B(men_men_n454_), .Y(men_men_n456_));
  NO2        u0428(.A(men_men_n400_), .B(men_men_n187_), .Y(men_men_n457_));
  NOi21      u0429(.An(men_men_n456_), .B(men_men_n457_), .Y(men_men_n458_));
  AOI210     u0430(.A0(men_men_n249_), .A1(men_men_n453_), .B0(men_men_n458_), .Y(men_men_n459_));
  OR2        u0431(.A(k), .B(j), .Y(men_men_n460_));
  NA2        u0432(.A(l), .B(k), .Y(men_men_n461_));
  NA2        u0433(.A(men_men_n215_), .B(men_men_n317_), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n258_), .B(men_men_n119_), .Y(men_men_n463_));
  NA2        u0435(.A(men_men_n370_), .B(men_men_n107_), .Y(men_men_n464_));
  NO4        u0436(.A(men_men_n464_), .B(men_men_n90_), .C(men_men_n106_), .D(e), .Y(men_men_n465_));
  NO3        u0437(.A(men_men_n400_), .B(men_men_n87_), .C(men_men_n121_), .Y(men_men_n466_));
  NO4        u0438(.A(men_men_n466_), .B(men_men_n465_), .C(men_men_n463_), .D(men_men_n301_), .Y(men_men_n467_));
  INV        u0439(.A(men_men_n467_), .Y(men_men_n468_));
  NO3        u0440(.A(men_men_n468_), .B(men_men_n459_), .C(men_men_n452_), .Y(men_men_n469_));
  NA2        u0441(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n470_));
  NO2        u0442(.A(men_men_n170_), .B(men_men_n54_), .Y(men_men_n471_));
  NAi31      u0443(.An(j), .B(l), .C(i), .Y(men_men_n472_));
  OAI210     u0444(.A0(men_men_n472_), .A1(men_men_n122_), .B0(men_men_n98_), .Y(men_men_n473_));
  NA2        u0445(.A(men_men_n473_), .B(men_men_n471_), .Y(men_men_n474_));
  NO3        u0446(.A(men_men_n371_), .B(men_men_n324_), .C(men_men_n184_), .Y(men_men_n475_));
  NO2        u0447(.A(men_men_n371_), .B(men_men_n349_), .Y(men_men_n476_));
  NO4        u0448(.A(men_men_n476_), .B(men_men_n475_), .C(men_men_n166_), .D(men_men_n283_), .Y(men_men_n477_));
  NA4        u0449(.A(men_men_n477_), .B(men_men_n474_), .C(men_men_n470_), .D(men_men_n225_), .Y(men_men_n478_));
  OAI210     u0450(.A0(men_men_n118_), .A1(men_men_n117_), .B0(n), .Y(men_men_n479_));
  NO2        u0451(.A(men_men_n479_), .B(men_men_n121_), .Y(men_men_n480_));
  XO2        u0452(.A(i), .B(h), .Y(men_men_n481_));
  NA3        u0453(.A(men_men_n481_), .B(men_men_n145_), .C(n), .Y(men_men_n482_));
  NAi41      u0454(.An(men_men_n279_), .B(men_men_n482_), .C(men_men_n435_), .D(men_men_n360_), .Y(men_men_n483_));
  AN2        u0455(.A(men_men_n483_), .B(men_men_n447_), .Y(men_men_n484_));
  NAi31      u0456(.An(c), .B(f), .C(d), .Y(men_men_n485_));
  NA3        u0457(.A(men_men_n358_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n486_));
  NA2        u0458(.A(men_men_n209_), .B(men_men_n102_), .Y(men_men_n487_));
  AOI210     u0459(.A0(men_men_n487_), .A1(men_men_n162_), .B0(men_men_n485_), .Y(men_men_n488_));
  AOI210     u0460(.A0(men_men_n337_), .A1(men_men_n34_), .B0(men_men_n456_), .Y(men_men_n489_));
  NOi31      u0461(.An(men_men_n486_), .B(men_men_n489_), .C(men_men_n488_), .Y(men_men_n490_));
  AO220      u0462(.A0(men_men_n267_), .A1(men_men_n243_), .B0(men_men_n150_), .B1(men_men_n65_), .Y(men_men_n491_));
  NA3        u0463(.A(men_men_n36_), .B(men_men_n35_), .C(f), .Y(men_men_n492_));
  NO2        u0464(.A(men_men_n492_), .B(men_men_n412_), .Y(men_men_n493_));
  NO2        u0465(.A(men_men_n493_), .B(men_men_n275_), .Y(men_men_n494_));
  NAi31      u0466(.An(men_men_n491_), .B(men_men_n494_), .C(men_men_n490_), .Y(men_men_n495_));
  NO3        u0467(.A(men_men_n495_), .B(men_men_n484_), .C(men_men_n478_), .Y(men_men_n496_));
  NA4        u0468(.A(men_men_n496_), .B(men_men_n469_), .C(men_men_n439_), .D(men_men_n407_), .Y(men11));
  NO2        u0469(.A(men_men_n71_), .B(f), .Y(men_men_n498_));
  NA2        u0470(.A(j), .B(u), .Y(men_men_n499_));
  NAi31      u0471(.An(i), .B(m), .C(l), .Y(men_men_n500_));
  NA3        u0472(.A(m), .B(k), .C(j), .Y(men_men_n501_));
  OAI220     u0473(.A0(men_men_n501_), .A1(men_men_n121_), .B0(men_men_n500_), .B1(men_men_n499_), .Y(men_men_n502_));
  NA2        u0474(.A(men_men_n502_), .B(men_men_n498_), .Y(men_men_n503_));
  NOi32      u0475(.An(e), .Bn(b), .C(f), .Y(men_men_n504_));
  NA2        u0476(.A(men_men_n239_), .B(men_men_n107_), .Y(men_men_n505_));
  NA2        u0477(.A(men_men_n45_), .B(j), .Y(men_men_n506_));
  NAi31      u0478(.An(d), .B(e), .C(a), .Y(men_men_n507_));
  NO2        u0479(.A(men_men_n507_), .B(n), .Y(men_men_n508_));
  NA2        u0480(.A(men_men_n508_), .B(men_men_n97_), .Y(men_men_n509_));
  NAi41      u0481(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n510_));
  BUFFER     u0482(.A(men_men_n510_), .Y(men_men_n511_));
  NA2        u0483(.A(j), .B(i), .Y(men_men_n512_));
  NAi31      u0484(.An(n), .B(m), .C(k), .Y(men_men_n513_));
  NO3        u0485(.A(men_men_n513_), .B(men_men_n512_), .C(men_men_n106_), .Y(men_men_n514_));
  OR2        u0486(.A(n), .B(c), .Y(men_men_n515_));
  NO2        u0487(.A(men_men_n515_), .B(men_men_n136_), .Y(men_men_n516_));
  NOi32      u0488(.An(u), .Bn(f), .C(i), .Y(men_men_n517_));
  AOI220     u0489(.A0(men_men_n517_), .A1(men_men_n95_), .B0(men_men_n502_), .B1(f), .Y(men_men_n518_));
  NO2        u0490(.A(men_men_n253_), .B(men_men_n48_), .Y(men_men_n519_));
  NO2        u0491(.A(men_men_n518_), .B(n), .Y(men_men_n520_));
  INV        u0492(.A(men_men_n520_), .Y(men_men_n521_));
  NA2        u0493(.A(men_men_n128_), .B(men_men_n33_), .Y(men_men_n522_));
  OAI220     u0494(.A0(men_men_n522_), .A1(m), .B0(men_men_n506_), .B1(men_men_n215_), .Y(men_men_n523_));
  OAI220     u0495(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n500_), .B1(men_men_n499_), .Y(men_men_n524_));
  NAi31      u0496(.An(d), .B(c), .C(a), .Y(men_men_n525_));
  NO2        u0497(.A(men_men_n525_), .B(n), .Y(men_men_n526_));
  NA3        u0498(.A(men_men_n526_), .B(men_men_n524_), .C(e), .Y(men_men_n527_));
  NO3        u0499(.A(men_men_n60_), .B(men_men_n48_), .C(men_men_n197_), .Y(men_men_n528_));
  NO2        u0500(.A(men_men_n212_), .B(men_men_n104_), .Y(men_men_n529_));
  OAI210     u0501(.A0(men_men_n528_), .A1(men_men_n374_), .B0(men_men_n529_), .Y(men_men_n530_));
  NA2        u0502(.A(men_men_n530_), .B(men_men_n527_), .Y(men_men_n531_));
  NA2        u0503(.A(men_men_n524_), .B(f), .Y(men_men_n532_));
  NO2        u0504(.A(d), .B(men_men_n48_), .Y(men_men_n533_));
  NA2        u0505(.A(h), .B(f), .Y(men_men_n534_));
  NO2        u0506(.A(men_men_n534_), .B(men_men_n90_), .Y(men_men_n535_));
  NO3        u0507(.A(men_men_n158_), .B(men_men_n155_), .C(u), .Y(men_men_n536_));
  AOI220     u0508(.A0(men_men_n536_), .A1(men_men_n56_), .B0(men_men_n535_), .B1(men_men_n533_), .Y(men_men_n537_));
  INV        u0509(.A(men_men_n537_), .Y(men_men_n538_));
  AN3        u0510(.A(j), .B(h), .C(u), .Y(men_men_n539_));
  NA3        u0511(.A(d), .B(men_men_n539_), .C(men_men_n434_), .Y(men_men_n540_));
  NA3        u0512(.A(f), .B(d), .C(b), .Y(men_men_n541_));
  NO4        u0513(.A(men_men_n541_), .B(men_men_n158_), .C(men_men_n155_), .D(u), .Y(men_men_n542_));
  NO4        u0514(.A(men_men_n542_), .B(men_men_n538_), .C(men_men_n531_), .D(men_men_n523_), .Y(men_men_n543_));
  AN4        u0515(.A(men_men_n543_), .B(men_men_n521_), .C(men_men_n509_), .D(men_men_n503_), .Y(men_men_n544_));
  INV        u0516(.A(k), .Y(men_men_n545_));
  NA3        u0517(.A(l), .B(men_men_n545_), .C(i), .Y(men_men_n546_));
  INV        u0518(.A(men_men_n546_), .Y(men_men_n547_));
  NA4        u0519(.A(men_men_n370_), .B(men_men_n391_), .C(men_men_n163_), .D(men_men_n107_), .Y(men_men_n548_));
  NAi32      u0520(.An(h), .Bn(f), .C(u), .Y(men_men_n549_));
  NAi41      u0521(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n550_));
  OAI210     u0522(.A0(men_men_n507_), .A1(n), .B0(men_men_n550_), .Y(men_men_n551_));
  NA2        u0523(.A(men_men_n551_), .B(m), .Y(men_men_n552_));
  NAi31      u0524(.An(h), .B(u), .C(f), .Y(men_men_n553_));
  OR3        u0525(.A(men_men_n553_), .B(men_men_n255_), .C(men_men_n48_), .Y(men_men_n554_));
  OA210      u0526(.A0(men_men_n552_), .A1(men_men_n549_), .B0(men_men_n554_), .Y(men_men_n555_));
  NO3        u0527(.A(men_men_n549_), .B(men_men_n71_), .C(men_men_n73_), .Y(men_men_n556_));
  NAi31      u0528(.An(men_men_n556_), .B(men_men_n555_), .C(men_men_n548_), .Y(men_men_n557_));
  NAi31      u0529(.An(f), .B(h), .C(u), .Y(men_men_n558_));
  NO4        u0530(.A(men_men_n288_), .B(men_men_n558_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n559_));
  NOi32      u0531(.An(b), .Bn(a), .C(c), .Y(men_men_n560_));
  NOi32      u0532(.An(d), .Bn(a), .C(e), .Y(men_men_n561_));
  NO2        u0533(.A(n), .B(c), .Y(men_men_n562_));
  NOi32      u0534(.An(e), .Bn(a), .C(d), .Y(men_men_n563_));
  AOI210     u0535(.A0(men_men_n29_), .A1(d), .B0(men_men_n563_), .Y(men_men_n564_));
  INV        u0536(.A(men_men_n522_), .Y(men_men_n565_));
  AOI210     u0537(.A0(men_men_n565_), .A1(men_men_n107_), .B0(men_men_n559_), .Y(men_men_n566_));
  INV        u0538(.A(men_men_n566_), .Y(men_men_n567_));
  AOI210     u0539(.A0(men_men_n557_), .A1(men_men_n547_), .B0(men_men_n567_), .Y(men_men_n568_));
  NO3        u0540(.A(men_men_n295_), .B(men_men_n59_), .C(n), .Y(men_men_n569_));
  INV        u0541(.A(men_men_n212_), .Y(men_men_n570_));
  NA2        u0542(.A(men_men_n74_), .B(men_men_n107_), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n1312_), .B(men_men_n82_), .Y(men_men_n572_));
  NA2        u0544(.A(men_men_n319_), .B(men_men_n45_), .Y(men_men_n573_));
  NOi32      u0545(.An(e), .Bn(c), .C(f), .Y(men_men_n574_));
  INV        u0546(.A(men_men_n195_), .Y(men_men_n575_));
  AOI220     u0547(.A0(men_men_n575_), .A1(men_men_n367_), .B0(men_men_n574_), .B1(men_men_n157_), .Y(men_men_n576_));
  NA3        u0548(.A(men_men_n576_), .B(men_men_n573_), .C(men_men_n160_), .Y(men_men_n577_));
  AOI210     u0549(.A0(men_men_n511_), .A1(men_men_n371_), .B0(men_men_n280_), .Y(men_men_n578_));
  NA2        u0550(.A(men_men_n578_), .B(men_men_n244_), .Y(men_men_n579_));
  NOi21      u0551(.An(j), .B(l), .Y(men_men_n580_));
  NAi21      u0552(.An(k), .B(h), .Y(men_men_n581_));
  NO2        u0553(.A(men_men_n581_), .B(men_men_n242_), .Y(men_men_n582_));
  NA2        u0554(.A(men_men_n582_), .B(men_men_n580_), .Y(men_men_n583_));
  OR2        u0555(.A(men_men_n583_), .B(men_men_n552_), .Y(men_men_n584_));
  NOi31      u0556(.An(m), .B(n), .C(k), .Y(men_men_n585_));
  NA2        u0557(.A(men_men_n580_), .B(men_men_n585_), .Y(men_men_n586_));
  NO2        u0558(.A(men_men_n371_), .B(men_men_n280_), .Y(men_men_n587_));
  NAi21      u0559(.An(men_men_n586_), .B(men_men_n587_), .Y(men_men_n588_));
  NO2        u0560(.A(men_men_n255_), .B(men_men_n48_), .Y(men_men_n589_));
  NO2        u0561(.A(men_men_n288_), .B(men_men_n558_), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n507_), .B(men_men_n48_), .Y(men_men_n591_));
  AOI220     u0563(.A0(men_men_n591_), .A1(men_men_n590_), .B0(men_men_n589_), .B1(men_men_n535_), .Y(men_men_n592_));
  NA4        u0564(.A(men_men_n592_), .B(men_men_n588_), .C(men_men_n584_), .D(men_men_n579_), .Y(men_men_n593_));
  NA2        u0565(.A(men_men_n102_), .B(men_men_n35_), .Y(men_men_n594_));
  NO2        u0566(.A(k), .B(men_men_n197_), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n504_), .B(men_men_n339_), .Y(men_men_n596_));
  NO2        u0568(.A(men_men_n596_), .B(n), .Y(men_men_n597_));
  NAi31      u0569(.An(men_men_n594_), .B(men_men_n597_), .C(men_men_n595_), .Y(men_men_n598_));
  AN3        u0570(.A(f), .B(d), .C(b), .Y(men_men_n599_));
  NA3        u0571(.A(men_men_n481_), .B(men_men_n145_), .C(men_men_n197_), .Y(men_men_n600_));
  AOI210     u0572(.A0(men_men_n1313_), .A1(men_men_n214_), .B0(men_men_n600_), .Y(men_men_n601_));
  NAi31      u0573(.An(m), .B(n), .C(k), .Y(men_men_n602_));
  INV        u0574(.A(men_men_n230_), .Y(men_men_n603_));
  OAI210     u0575(.A0(men_men_n603_), .A1(men_men_n601_), .B0(j), .Y(men_men_n604_));
  NA2        u0576(.A(men_men_n604_), .B(men_men_n598_), .Y(men_men_n605_));
  NO4        u0577(.A(men_men_n605_), .B(men_men_n593_), .C(men_men_n577_), .D(men_men_n572_), .Y(men_men_n606_));
  NA2        u0578(.A(men_men_n358_), .B(men_men_n148_), .Y(men_men_n607_));
  NAi31      u0579(.An(u), .B(h), .C(f), .Y(men_men_n608_));
  OA210      u0580(.A0(men_men_n507_), .A1(n), .B0(men_men_n550_), .Y(men_men_n609_));
  NO2        u0581(.A(men_men_n609_), .B(men_men_n86_), .Y(men_men_n610_));
  INV        u0582(.A(men_men_n610_), .Y(men_men_n611_));
  AOI210     u0583(.A0(men_men_n611_), .A1(men_men_n607_), .B0(men_men_n501_), .Y(men_men_n612_));
  NAi21      u0584(.An(h), .B(j), .Y(men_men_n613_));
  OR2        u0585(.A(men_men_n583_), .B(men_men_n71_), .Y(men_men_n614_));
  NA3        u0586(.A(men_men_n498_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n615_));
  NA2        u0587(.A(h), .B(men_men_n36_), .Y(men_men_n616_));
  NA2        u0588(.A(men_men_n95_), .B(men_men_n45_), .Y(men_men_n617_));
  OAI220     u0589(.A0(men_men_n617_), .A1(men_men_n311_), .B0(men_men_n616_), .B1(men_men_n441_), .Y(men_men_n618_));
  AOI210     u0590(.A0(d), .A1(men_men_n401_), .B0(men_men_n48_), .Y(men_men_n619_));
  OAI220     u0591(.A0(men_men_n553_), .A1(men_men_n546_), .B0(men_men_n304_), .B1(men_men_n499_), .Y(men_men_n620_));
  AOI210     u0592(.A0(men_men_n620_), .A1(men_men_n619_), .B0(men_men_n618_), .Y(men_men_n621_));
  NA3        u0593(.A(men_men_n621_), .B(men_men_n615_), .C(men_men_n614_), .Y(men_men_n622_));
  NA2        u0594(.A(men_men_n307_), .B(men_men_n128_), .Y(men_men_n623_));
  NA2        u0595(.A(men_men_n122_), .B(men_men_n48_), .Y(men_men_n624_));
  OR2        u0596(.A(men_men_n337_), .B(men_men_n105_), .Y(men_men_n625_));
  NA2        u0597(.A(men_men_n623_), .B(men_men_n625_), .Y(men_men_n626_));
  INV        u0598(.A(men_men_n212_), .Y(men_men_n627_));
  NA3        u0599(.A(men_men_n627_), .B(men_men_n233_), .C(j), .Y(men_men_n628_));
  NA2        u0600(.A(men_men_n440_), .B(men_men_n81_), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n628_), .B(men_men_n486_), .C(men_men_n376_), .Y(men_men_n630_));
  NO4        u0602(.A(men_men_n630_), .B(men_men_n626_), .C(men_men_n622_), .D(men_men_n612_), .Y(men_men_n631_));
  NA4        u0603(.A(men_men_n631_), .B(men_men_n606_), .C(men_men_n568_), .D(men_men_n544_), .Y(men08));
  NO2        u0604(.A(k), .B(h), .Y(men_men_n633_));
  AO210      u0605(.A0(men_men_n231_), .A1(men_men_n426_), .B0(men_men_n633_), .Y(men_men_n634_));
  NO2        u0606(.A(men_men_n634_), .B(men_men_n278_), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n574_), .B(men_men_n81_), .Y(men_men_n636_));
  AOI210     u0608(.A0(men_men_n574_), .A1(men_men_n635_), .B0(men_men_n466_), .Y(men_men_n637_));
  NO2        u0609(.A(n), .B(men_men_n55_), .Y(men_men_n638_));
  NO4        u0610(.A(men_men_n355_), .B(men_men_n106_), .C(j), .D(men_men_n197_), .Y(men_men_n639_));
  INV        u0611(.A(men_men_n214_), .Y(men_men_n640_));
  AOI220     u0612(.A0(men_men_n640_), .A1(men_men_n326_), .B0(men_men_n639_), .B1(men_men_n638_), .Y(men_men_n641_));
  NA4        u0613(.A(men_men_n199_), .B(men_men_n128_), .C(men_men_n44_), .D(h), .Y(men_men_n642_));
  AN2        u0614(.A(l), .B(k), .Y(men_men_n643_));
  NA3        u0615(.A(men_men_n641_), .B(men_men_n637_), .C(men_men_n327_), .Y(men_men_n644_));
  AN2        u0616(.A(men_men_n508_), .B(men_men_n91_), .Y(men_men_n645_));
  NO4        u0617(.A(men_men_n155_), .B(m), .C(men_men_n106_), .D(u), .Y(men_men_n646_));
  AOI210     u0618(.A0(men_men_n646_), .A1(men_men_n640_), .B0(men_men_n493_), .Y(men_men_n647_));
  NO2        u0619(.A(men_men_n37_), .B(men_men_n196_), .Y(men_men_n648_));
  NA2        u0620(.A(men_men_n575_), .B(men_men_n325_), .Y(men_men_n649_));
  NA2        u0621(.A(men_men_n649_), .B(men_men_n647_), .Y(men_men_n650_));
  NA2        u0622(.A(men_men_n1314_), .B(men_men_n76_), .Y(men_men_n651_));
  OAI210     u0623(.A0(men_men_n34_), .A1(men_men_n82_), .B0(men_men_n651_), .Y(men_men_n652_));
  NA2        u0624(.A(men_men_n339_), .B(men_men_n42_), .Y(men_men_n653_));
  NA3        u0625(.A(men_men_n627_), .B(men_men_n313_), .C(men_men_n359_), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n643_), .B(men_men_n202_), .Y(men_men_n655_));
  NO2        u0627(.A(men_men_n655_), .B(men_men_n306_), .Y(men_men_n656_));
  AOI210     u0628(.A0(men_men_n656_), .A1(i), .B0(men_men_n465_), .Y(men_men_n657_));
  NA3        u0629(.A(m), .B(l), .C(k), .Y(men_men_n658_));
  NO2        u0630(.A(men_men_n510_), .B(men_men_n251_), .Y(men_men_n659_));
  NOi21      u0631(.An(men_men_n659_), .B(men_men_n505_), .Y(men_men_n660_));
  NA4        u0632(.A(men_men_n107_), .B(l), .C(k), .D(men_men_n82_), .Y(men_men_n661_));
  INV        u0633(.A(men_men_n660_), .Y(men_men_n662_));
  NA4        u0634(.A(men_men_n662_), .B(men_men_n657_), .C(men_men_n654_), .D(men_men_n653_), .Y(men_men_n663_));
  NO4        u0635(.A(men_men_n663_), .B(men_men_n652_), .C(men_men_n650_), .D(men_men_n644_), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n575_), .B(men_men_n367_), .Y(men_men_n665_));
  NA2        u0637(.A(men_men_n591_), .B(u), .Y(men_men_n666_));
  NO3        u0638(.A(men_men_n371_), .B(men_men_n499_), .C(h), .Y(men_men_n667_));
  AOI210     u0639(.A0(men_men_n667_), .A1(men_men_n107_), .B0(men_men_n476_), .Y(men_men_n668_));
  NA4        u0640(.A(men_men_n668_), .B(men_men_n666_), .C(men_men_n665_), .D(men_men_n230_), .Y(men_men_n669_));
  NOi21      u0641(.An(h), .B(j), .Y(men_men_n670_));
  NA2        u0642(.A(men_men_n670_), .B(f), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n554_), .B(men_men_n60_), .Y(men_men_n672_));
  AOI210     u0644(.A0(men_men_n669_), .A1(l), .B0(men_men_n672_), .Y(men_men_n673_));
  NO2        u0645(.A(j), .B(i), .Y(men_men_n674_));
  NA3        u0646(.A(men_men_n674_), .B(men_men_n79_), .C(l), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n674_), .B(men_men_n32_), .Y(men_men_n676_));
  OR2        u0648(.A(men_men_n675_), .B(men_men_n552_), .Y(men_men_n677_));
  NO3        u0649(.A(men_men_n138_), .B(men_men_n48_), .C(men_men_n104_), .Y(men_men_n678_));
  NO3        u0650(.A(men_men_n461_), .B(men_men_n413_), .C(j), .Y(men_men_n679_));
  NA2        u0651(.A(men_men_n678_), .B(men_men_n679_), .Y(men_men_n680_));
  INV        u0652(.A(men_men_n680_), .Y(men_men_n681_));
  NA2        u0653(.A(k), .B(j), .Y(men_men_n682_));
  NA2        u0654(.A(men_men_n570_), .B(men_men_n285_), .Y(men_men_n683_));
  NAi31      u0655(.An(men_men_n564_), .B(men_men_n88_), .C(men_men_n81_), .Y(men_men_n684_));
  NA2        u0656(.A(men_men_n684_), .B(men_men_n683_), .Y(men_men_n685_));
  NO2        u0657(.A(men_men_n278_), .B(men_men_n124_), .Y(men_men_n686_));
  NA2        u0658(.A(men_men_n686_), .B(men_men_n575_), .Y(men_men_n687_));
  NO2        u0659(.A(men_men_n658_), .B(men_men_n86_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n688_), .B(men_men_n551_), .Y(men_men_n689_));
  NO2        u0661(.A(men_men_n553_), .B(men_men_n110_), .Y(men_men_n690_));
  OAI210     u0662(.A0(men_men_n690_), .A1(men_men_n679_), .B0(men_men_n619_), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n691_), .B(men_men_n689_), .C(men_men_n687_), .Y(men_men_n692_));
  OR3        u0664(.A(men_men_n692_), .B(men_men_n685_), .C(men_men_n681_), .Y(men_men_n693_));
  NA3        u0665(.A(men_men_n199_), .B(men_men_n426_), .C(men_men_n33_), .Y(men_men_n694_));
  NO4        u0666(.A(men_men_n461_), .B(men_men_n408_), .C(j), .D(f), .Y(men_men_n695_));
  NO2        u0667(.A(men_men_n311_), .B(men_men_n37_), .Y(men_men_n696_));
  AOI210     u0668(.A0(men_men_n695_), .A1(men_men_n237_), .B0(men_men_n696_), .Y(men_men_n697_));
  NA3        u0669(.A(men_men_n517_), .B(men_men_n271_), .C(h), .Y(men_men_n698_));
  NO2        u0670(.A(men_men_n87_), .B(men_men_n46_), .Y(men_men_n699_));
  NO2        u0671(.A(men_men_n675_), .B(men_men_n71_), .Y(men_men_n700_));
  AOI210     u0672(.A0(men_men_n699_), .A1(men_men_n597_), .B0(men_men_n700_), .Y(men_men_n701_));
  NA3        u0673(.A(men_men_n701_), .B(men_men_n697_), .C(men_men_n694_), .Y(men_men_n702_));
  OR2        u0674(.A(men_men_n688_), .B(men_men_n91_), .Y(men_men_n703_));
  AOI220     u0675(.A0(men_men_n703_), .A1(men_men_n220_), .B0(men_men_n679_), .B1(men_men_n589_), .Y(men_men_n704_));
  NO2        u0676(.A(men_men_n609_), .B(men_men_n73_), .Y(men_men_n705_));
  AOI210     u0677(.A0(men_men_n695_), .A1(men_men_n705_), .B0(men_men_n315_), .Y(men_men_n706_));
  OAI210     u0678(.A0(men_men_n658_), .A1(men_men_n608_), .B0(men_men_n492_), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n81_), .B(men_men_n707_), .Y(men_men_n708_));
  NA3        u0680(.A(men_men_n708_), .B(men_men_n706_), .C(men_men_n704_), .Y(men_men_n709_));
  NOi41      u0681(.An(men_men_n677_), .B(men_men_n709_), .C(men_men_n702_), .D(men_men_n693_), .Y(men_men_n710_));
  BUFFER     u0682(.A(men_men_n642_), .Y(men_men_n711_));
  NO3        u0683(.A(men_men_n320_), .B(men_men_n280_), .C(men_men_n106_), .Y(men_men_n712_));
  INV        u0684(.A(men_men_n712_), .Y(men_men_n713_));
  NA2        u0685(.A(men_men_n45_), .B(men_men_n54_), .Y(men_men_n714_));
  NO3        u0686(.A(men_men_n714_), .B(men_men_n676_), .C(men_men_n255_), .Y(men_men_n715_));
  NO3        u0687(.A(men_men_n499_), .B(men_men_n89_), .C(h), .Y(men_men_n716_));
  AOI210     u0688(.A0(men_men_n716_), .A1(men_men_n638_), .B0(men_men_n715_), .Y(men_men_n717_));
  NA4        u0689(.A(men_men_n717_), .B(men_men_n713_), .C(men_men_n711_), .D(men_men_n377_), .Y(men_men_n718_));
  OR2        u0690(.A(men_men_n608_), .B(men_men_n87_), .Y(men_men_n719_));
  NOi31      u0691(.An(b), .B(d), .C(a), .Y(men_men_n720_));
  OAI220     u0692(.A0(n), .A1(men_men_n719_), .B0(men_men_n698_), .B1(n), .Y(men_men_n721_));
  AOI220     u0693(.A0(men_men_n686_), .A1(f), .B0(f), .B1(men_men_n635_), .Y(men_men_n722_));
  NO2        u0694(.A(men_men_n302_), .B(men_men_n219_), .Y(men_men_n723_));
  OAI210     u0695(.A0(men_men_n91_), .A1(men_men_n88_), .B0(men_men_n723_), .Y(men_men_n724_));
  NA2        u0696(.A(men_men_n114_), .B(men_men_n81_), .Y(men_men_n725_));
  AOI210     u0697(.A0(men_men_n398_), .A1(men_men_n390_), .B0(men_men_n725_), .Y(men_men_n726_));
  INV        u0698(.A(men_men_n724_), .Y(men_men_n727_));
  NAi21      u0699(.An(men_men_n661_), .B(men_men_n409_), .Y(men_men_n728_));
  NO2        u0700(.A(men_men_n251_), .B(i), .Y(men_men_n729_));
  NA2        u0701(.A(men_men_n556_), .B(men_men_n340_), .Y(men_men_n730_));
  AN2        u0702(.A(men_men_n730_), .B(men_men_n728_), .Y(men_men_n731_));
  NAi31      u0703(.An(men_men_n727_), .B(men_men_n731_), .C(men_men_n722_), .Y(men_men_n732_));
  NO3        u0704(.A(men_men_n732_), .B(men_men_n721_), .C(men_men_n718_), .Y(men_men_n733_));
  NA4        u0705(.A(men_men_n733_), .B(men_men_n710_), .C(men_men_n673_), .D(men_men_n664_), .Y(men09));
  NA2        u0706(.A(f), .B(e), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n207_), .B(men_men_n106_), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n736_), .B(u), .Y(men_men_n737_));
  NA4        u0709(.A(men_men_n288_), .B(men_men_n449_), .C(men_men_n240_), .D(men_men_n112_), .Y(men_men_n738_));
  AOI210     u0710(.A0(men_men_n738_), .A1(u), .B0(men_men_n446_), .Y(men_men_n739_));
  AOI210     u0711(.A0(men_men_n739_), .A1(men_men_n737_), .B0(men_men_n735_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n419_), .B(e), .Y(men_men_n741_));
  NO2        u0713(.A(men_men_n187_), .B(men_men_n196_), .Y(men_men_n742_));
  NA3        u0714(.A(m), .B(l), .C(i), .Y(men_men_n743_));
  OAI220     u0715(.A0(men_men_n553_), .A1(men_men_n743_), .B0(men_men_n331_), .B1(men_men_n500_), .Y(men_men_n744_));
  NA4        u0716(.A(men_men_n83_), .B(men_men_n82_), .C(u), .D(f), .Y(men_men_n745_));
  NAi31      u0717(.An(men_men_n744_), .B(men_men_n745_), .C(men_men_n414_), .Y(men_men_n746_));
  OR2        u0718(.A(men_men_n746_), .B(men_men_n742_), .Y(men_men_n747_));
  NA3        u0719(.A(men_men_n719_), .B(men_men_n532_), .C(men_men_n492_), .Y(men_men_n748_));
  OA210      u0720(.A0(men_men_n748_), .A1(men_men_n747_), .B0(men_men_n1309_), .Y(men_men_n749_));
  INV        u0721(.A(men_men_n318_), .Y(men_men_n750_));
  NO2        u0722(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n751_));
  NO2        u0723(.A(m), .B(men_men_n558_), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n321_), .B(men_men_n323_), .Y(men_men_n753_));
  OAI210     u0725(.A0(men_men_n187_), .A1(men_men_n196_), .B0(men_men_n753_), .Y(men_men_n754_));
  NA2        u0726(.A(men_men_n752_), .B(men_men_n750_), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n755_), .B(men_men_n576_), .Y(men_men_n756_));
  NA2        u0728(.A(f), .B(m), .Y(men_men_n757_));
  NO2        u0729(.A(men_men_n757_), .B(men_men_n51_), .Y(men_men_n758_));
  NOi32      u0730(.An(u), .Bn(f), .C(d), .Y(men_men_n759_));
  NA4        u0731(.A(men_men_n759_), .B(men_men_n562_), .C(men_men_n29_), .D(m), .Y(men_men_n760_));
  NOi21      u0732(.An(men_men_n289_), .B(men_men_n760_), .Y(men_men_n761_));
  AOI210     u0733(.A0(men_men_n758_), .A1(men_men_n516_), .B0(men_men_n761_), .Y(men_men_n762_));
  AN2        u0734(.A(f), .B(d), .Y(men_men_n763_));
  NO2        u0735(.A(men_men_n602_), .B(men_men_n306_), .Y(men_men_n764_));
  NO2        u0736(.A(men_men_n764_), .B(men_men_n216_), .Y(men_men_n765_));
  NO2        u0737(.A(men_men_n753_), .B(n), .Y(men_men_n766_));
  NA3        u0738(.A(men_men_n145_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n767_));
  NO2        u0739(.A(men_men_n318_), .B(men_men_n767_), .Y(men_men_n768_));
  NOi41      u0740(.An(men_men_n205_), .B(men_men_n768_), .C(men_men_n766_), .D(men_men_n283_), .Y(men_men_n769_));
  NA2        u0741(.A(c), .B(men_men_n109_), .Y(men_men_n770_));
  NA3        u0742(.A(e), .B(men_men_n483_), .C(f), .Y(men_men_n771_));
  OR2        u0743(.A(men_men_n608_), .B(men_men_n513_), .Y(men_men_n772_));
  NA4        u0744(.A(men_men_n772_), .B(men_men_n771_), .C(men_men_n769_), .D(men_men_n765_), .Y(men_men_n773_));
  NO4        u0745(.A(men_men_n773_), .B(men_men_n463_), .C(men_men_n756_), .D(men_men_n749_), .Y(men_men_n774_));
  NO2        u0746(.A(men_men_n212_), .B(men_men_n206_), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n775_), .B(men_men_n209_), .Y(men_men_n776_));
  NO2        u0748(.A(men_men_n403_), .B(men_men_n735_), .Y(men_men_n777_));
  NA2        u0749(.A(e), .B(d), .Y(men_men_n778_));
  NA3        u0750(.A(e), .B(men_men_n430_), .C(men_men_n481_), .Y(men_men_n779_));
  AOI210     u0751(.A0(men_men_n487_), .A1(men_men_n162_), .B0(men_men_n212_), .Y(men_men_n780_));
  AOI210     u0752(.A0(men_men_n575_), .A1(men_men_n325_), .B0(men_men_n780_), .Y(men_men_n781_));
  NA2        u0753(.A(men_men_n781_), .B(men_men_n779_), .Y(men_men_n782_));
  NO2        u0754(.A(men_men_n782_), .B(men_men_n1307_), .Y(men_men_n783_));
  AO210      u0755(.A0(men_men_n318_), .A1(men_men_n636_), .B0(men_men_n200_), .Y(men_men_n784_));
  AOI220     u0756(.A0(h), .A1(men_men_n764_), .B0(men_men_n569_), .B1(men_men_n574_), .Y(men_men_n785_));
  AOI210     u0757(.A0(men_men_n111_), .A1(men_men_n110_), .B0(men_men_n239_), .Y(men_men_n786_));
  NOi31      u0758(.An(men_men_n516_), .B(men_men_n757_), .C(men_men_n272_), .Y(men_men_n787_));
  AO220      u0759(.A0(men_men_n430_), .A1(men_men_n670_), .B0(men_men_n157_), .B1(f), .Y(men_men_n788_));
  OAI210     u0760(.A0(men_men_n788_), .A1(men_men_n433_), .B0(e), .Y(men_men_n789_));
  AN3        u0761(.A(men_men_n789_), .B(men_men_n785_), .C(men_men_n784_), .Y(men_men_n790_));
  NA4        u0762(.A(men_men_n790_), .B(men_men_n783_), .C(men_men_n774_), .D(men_men_n741_), .Y(men12));
  NO4        u0763(.A(men_men_n418_), .B(men_men_n231_), .C(men_men_n545_), .D(men_men_n197_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n792_), .B(d), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n751_), .B(men_men_n331_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n608_), .B(men_men_n355_), .Y(men_men_n795_));
  AOI210     u0767(.A0(men_men_n795_), .A1(men_men_n1308_), .B0(men_men_n794_), .Y(men_men_n796_));
  NA3        u0768(.A(men_men_n796_), .B(men_men_n793_), .C(men_men_n417_), .Y(men_men_n797_));
  AOI210     u0769(.A0(men_men_n215_), .A1(men_men_n317_), .B0(men_men_n184_), .Y(men_men_n798_));
  NO2        u0770(.A(men_men_n594_), .B(men_men_n242_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n553_), .B(men_men_n743_), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n723_), .B(men_men_n799_), .Y(men_men_n801_));
  NO2        u0773(.A(men_men_n138_), .B(men_men_n219_), .Y(men_men_n802_));
  NA3        u0774(.A(men_men_n802_), .B(men_men_n222_), .C(i), .Y(men_men_n803_));
  NA2        u0775(.A(men_men_n803_), .B(men_men_n801_), .Y(men_men_n804_));
  NO3        u0776(.A(men_men_n122_), .B(men_men_n139_), .C(men_men_n197_), .Y(men_men_n805_));
  NO3        u0777(.A(men_men_n611_), .B(men_men_n87_), .C(men_men_n44_), .Y(men_men_n806_));
  NO4        u0778(.A(men_men_n806_), .B(men_men_n805_), .C(men_men_n804_), .D(men_men_n797_), .Y(men_men_n807_));
  NO2        u0779(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n808_));
  NA2        u0780(.A(men_men_n550_), .B(men_men_n71_), .Y(men_men_n809_));
  NOi21      u0781(.An(men_men_n33_), .B(men_men_n602_), .Y(men_men_n810_));
  AOI220     u0782(.A0(men_men_n810_), .A1(c), .B0(men_men_n809_), .B1(men_men_n808_), .Y(men_men_n811_));
  OAI210     u0783(.A0(men_men_n230_), .A1(men_men_n44_), .B0(men_men_n811_), .Y(men_men_n812_));
  NA2        u0784(.A(men_men_n409_), .B(men_men_n244_), .Y(men_men_n813_));
  NO3        u0785(.A(men_men_n725_), .B(men_men_n84_), .C(men_men_n381_), .Y(men_men_n814_));
  NA2        u0786(.A(men_men_n813_), .B(men_men_n299_), .Y(men_men_n815_));
  NO2        u0787(.A(men_men_n48_), .B(men_men_n44_), .Y(men_men_n816_));
  NA2        u0788(.A(men_men_n585_), .B(men_men_n340_), .Y(men_men_n817_));
  INV        u0789(.A(men_men_n344_), .Y(men_men_n818_));
  NO3        u0790(.A(men_men_n818_), .B(men_men_n815_), .C(men_men_n812_), .Y(men_men_n819_));
  NA2        u0791(.A(men_men_n325_), .B(u), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n148_), .B(i), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n45_), .B(i), .Y(men_men_n822_));
  OAI220     u0794(.A0(men_men_n822_), .A1(men_men_n183_), .B0(men_men_n821_), .B1(men_men_n87_), .Y(men_men_n823_));
  AOI210     u0795(.A0(men_men_n392_), .A1(men_men_n36_), .B0(men_men_n823_), .Y(men_men_n824_));
  OAI210     u0796(.A0(men_men_n824_), .A1(men_men_n311_), .B0(men_men_n820_), .Y(men_men_n825_));
  NO2        u0797(.A(men_men_n608_), .B(men_men_n472_), .Y(men_men_n826_));
  NA3        u0798(.A(men_men_n321_), .B(men_men_n580_), .C(i), .Y(men_men_n827_));
  NO2        u0799(.A(men_men_n413_), .B(men_men_n288_), .Y(men_men_n828_));
  OAI210     u0800(.A0(men_men_n828_), .A1(men_men_n826_), .B0(men_men_n619_), .Y(men_men_n829_));
  NA2        u0801(.A(men_men_n563_), .B(men_men_n107_), .Y(men_men_n830_));
  OR3        u0802(.A(men_men_n288_), .B(men_men_n408_), .C(f), .Y(men_men_n831_));
  NA3        u0803(.A(men_men_n580_), .B(men_men_n79_), .C(i), .Y(men_men_n832_));
  OA220      u0804(.A0(men_men_n832_), .A1(men_men_n830_), .B0(men_men_n831_), .B1(men_men_n552_), .Y(men_men_n833_));
  NA3        u0805(.A(men_men_n303_), .B(men_men_n111_), .C(u), .Y(men_men_n834_));
  AOI210     u0806(.A0(men_men_n616_), .A1(men_men_n834_), .B0(m), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n745_), .B(men_men_n414_), .Y(men_men_n836_));
  NA2        u0808(.A(men_men_n203_), .B(h), .Y(men_men_n837_));
  NA3        u0809(.A(men_men_n837_), .B(men_men_n832_), .C(men_men_n831_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n838_), .B(men_men_n237_), .Y(men_men_n839_));
  NA3        u0811(.A(men_men_n839_), .B(men_men_n833_), .C(men_men_n829_), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n355_), .B(men_men_n86_), .Y(men_men_n841_));
  OAI210     u0813(.A0(men_men_n841_), .A1(men_men_n799_), .B0(men_men_n220_), .Y(men_men_n842_));
  NA2        u0814(.A(men_men_n610_), .B(men_men_n83_), .Y(men_men_n843_));
  NA2        u0815(.A(men_men_n551_), .B(men_men_n85_), .Y(men_men_n844_));
  NA3        u0816(.A(men_men_n844_), .B(men_men_n843_), .C(men_men_n842_), .Y(men_men_n845_));
  OAI210     u0817(.A0(men_men_n836_), .A1(men_men_n800_), .B0(men_men_n1308_), .Y(men_men_n846_));
  AOI210     u0818(.A0(men_men_n393_), .A1(men_men_n385_), .B0(men_men_n725_), .Y(men_men_n847_));
  OAI210     u0819(.A0(men_men_n346_), .A1(men_men_n345_), .B0(men_men_n103_), .Y(men_men_n848_));
  AOI210     u0820(.A0(men_men_n848_), .A1(men_men_n508_), .B0(men_men_n847_), .Y(men_men_n849_));
  INV        u0821(.A(men_men_n835_), .Y(men_men_n850_));
  NO3        u0822(.A(l), .B(men_men_n48_), .C(men_men_n44_), .Y(men_men_n851_));
  NA2        u0823(.A(men_men_n851_), .B(men_men_n578_), .Y(men_men_n852_));
  NA4        u0824(.A(men_men_n852_), .B(men_men_n850_), .C(men_men_n849_), .D(men_men_n846_), .Y(men_men_n853_));
  NO4        u0825(.A(men_men_n853_), .B(men_men_n845_), .C(men_men_n840_), .D(men_men_n825_), .Y(men_men_n854_));
  NAi31      u0826(.An(men_men_n129_), .B(men_men_n394_), .C(n), .Y(men_men_n855_));
  NO2        u0827(.A(m), .B(men_men_n855_), .Y(men_men_n856_));
  NO2        u0828(.A(men_men_n251_), .B(men_men_n381_), .Y(men_men_n857_));
  AOI210     u0829(.A0(men_men_n857_), .A1(men_men_n473_), .B0(men_men_n856_), .Y(men_men_n858_));
  NA2        u0830(.A(men_men_n466_), .B(i), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n859_), .B(men_men_n858_), .Y(men_men_n860_));
  NO3        u0832(.A(men_men_n285_), .B(men_men_n419_), .C(men_men_n157_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n861_), .B(men_men_n197_), .Y(men_men_n862_));
  NO3        u0834(.A(men_men_n413_), .B(men_men_n288_), .C(men_men_n73_), .Y(men_men_n863_));
  NA2        u0835(.A(men_men_n863_), .B(men_men_n410_), .Y(men_men_n864_));
  INV        u0836(.A(men_men_n864_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n827_), .B(n), .Y(men_men_n866_));
  NA2        u0838(.A(men_men_n798_), .B(d), .Y(men_men_n867_));
  NA2        u0839(.A(men_men_n498_), .B(men_men_n356_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n792_), .B(c), .Y(men_men_n869_));
  NA3        u0841(.A(c), .B(men_men_n462_), .C(men_men_n45_), .Y(men_men_n870_));
  AOI210     u0842(.A0(men_men_n358_), .A1(men_men_n356_), .B0(men_men_n310_), .Y(men_men_n871_));
  NA3        u0843(.A(men_men_n871_), .B(men_men_n870_), .C(men_men_n869_), .Y(men_men_n872_));
  OR3        u0844(.A(men_men_n872_), .B(men_men_n798_), .C(men_men_n866_), .Y(men_men_n873_));
  NO4        u0845(.A(men_men_n873_), .B(men_men_n865_), .C(men_men_n862_), .D(men_men_n860_), .Y(men_men_n874_));
  NA4        u0846(.A(men_men_n874_), .B(men_men_n854_), .C(men_men_n819_), .D(men_men_n807_), .Y(men13));
  NA2        u0847(.A(men_men_n45_), .B(men_men_n82_), .Y(men_men_n876_));
  AN2        u0848(.A(c), .B(b), .Y(men_men_n877_));
  NA3        u0849(.A(men_men_n229_), .B(men_men_n877_), .C(m), .Y(men_men_n878_));
  NO4        u0850(.A(e), .B(men_men_n878_), .C(men_men_n876_), .D(men_men_n546_), .Y(men_men_n879_));
  NA2        u0851(.A(men_men_n244_), .B(men_men_n877_), .Y(men_men_n880_));
  NO4        u0852(.A(men_men_n880_), .B(e), .C(men_men_n821_), .D(a), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n128_), .B(men_men_n44_), .Y(men_men_n882_));
  NO4        u0854(.A(men_men_n882_), .B(d), .C(men_men_n553_), .D(men_men_n284_), .Y(men_men_n883_));
  NA2        u0855(.A(men_men_n613_), .B(men_men_n206_), .Y(men_men_n884_));
  AN2        u0856(.A(d), .B(c), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n885_), .B(men_men_n109_), .Y(men_men_n886_));
  NO3        u0858(.A(men_men_n886_), .B(men_men_n158_), .C(men_men_n153_), .Y(men_men_n887_));
  NA2        u0859(.A(d), .B(c), .Y(men_men_n888_));
  NO4        u0860(.A(men_men_n882_), .B(men_men_n549_), .C(men_men_n888_), .D(men_men_n284_), .Y(men_men_n889_));
  AO210      u0861(.A0(men_men_n887_), .A1(men_men_n884_), .B0(men_men_n889_), .Y(men_men_n890_));
  OR4        u0862(.A(men_men_n890_), .B(men_men_n883_), .C(men_men_n881_), .D(men_men_n879_), .Y(men_men_n891_));
  NAi32      u0863(.An(f), .Bn(e), .C(c), .Y(men_men_n892_));
  OR3        u0864(.A(men_men_n206_), .B(men_men_n158_), .C(men_men_n153_), .Y(men_men_n893_));
  NO2        u0865(.A(men_men_n893_), .B(men_men_n892_), .Y(men_men_n894_));
  NO2        u0866(.A(men_men_n888_), .B(men_men_n284_), .Y(men_men_n895_));
  NA2        u0867(.A(men_men_n582_), .B(men_men_n1305_), .Y(men_men_n896_));
  NOi21      u0868(.An(men_men_n895_), .B(men_men_n896_), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n682_), .B(men_men_n106_), .Y(men_men_n898_));
  NOi41      u0870(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n899_));
  NA2        u0871(.A(men_men_n899_), .B(men_men_n898_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n900_), .B(men_men_n892_), .Y(men_men_n901_));
  NA3        u0873(.A(k), .B(j), .C(i), .Y(men_men_n902_));
  NO3        u0874(.A(men_men_n902_), .B(men_men_n284_), .C(men_men_n86_), .Y(men_men_n903_));
  OR4        u0875(.A(men_men_n903_), .B(men_men_n901_), .C(men_men_n897_), .D(men_men_n894_), .Y(men_men_n904_));
  NA3        u0876(.A(men_men_n443_), .B(men_men_n313_), .C(men_men_n54_), .Y(men_men_n905_));
  NO2        u0877(.A(men_men_n905_), .B(men_men_n896_), .Y(men_men_n906_));
  NO3        u0878(.A(men_men_n905_), .B(men_men_n549_), .C(men_men_n44_), .Y(men_men_n907_));
  NO2        u0879(.A(f), .B(c), .Y(men_men_n908_));
  NOi21      u0880(.An(men_men_n908_), .B(men_men_n418_), .Y(men_men_n909_));
  NA2        u0881(.A(men_men_n909_), .B(men_men_n57_), .Y(men_men_n910_));
  NO3        u0882(.A(k), .B(h), .C(l), .Y(men_men_n911_));
  NOi31      u0883(.An(men_men_n911_), .B(men_men_n910_), .C(j), .Y(men_men_n912_));
  OR3        u0884(.A(men_men_n912_), .B(men_men_n907_), .C(men_men_n906_), .Y(men_men_n913_));
  OR3        u0885(.A(men_men_n913_), .B(men_men_n904_), .C(men_men_n891_), .Y(men02));
  OR2        u0886(.A(l), .B(k), .Y(men_men_n915_));
  OR3        u0887(.A(h), .B(u), .C(f), .Y(men_men_n916_));
  OR3        u0888(.A(n), .B(m), .C(i), .Y(men_men_n917_));
  NO4        u0889(.A(men_men_n917_), .B(men_men_n916_), .C(men_men_n915_), .D(e), .Y(men_men_n918_));
  AOI210     u0890(.A0(men_men_n903_), .A1(e), .B0(men_men_n883_), .Y(men_men_n919_));
  AN3        u0891(.A(u), .B(f), .C(c), .Y(men_men_n920_));
  NA3        u0892(.A(men_men_n920_), .B(men_men_n443_), .C(h), .Y(men_men_n921_));
  OR2        u0893(.A(men_men_n284_), .B(men_men_n921_), .Y(men_men_n922_));
  NO3        u0894(.A(men_men_n905_), .B(men_men_n882_), .C(men_men_n549_), .Y(men_men_n923_));
  NO2        u0895(.A(men_men_n923_), .B(men_men_n894_), .Y(men_men_n924_));
  NA2        u0896(.A(i), .B(h), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n925_), .B(men_men_n122_), .Y(men_men_n926_));
  NO3        u0898(.A(men_men_n130_), .B(men_men_n262_), .C(men_men_n197_), .Y(men_men_n927_));
  AOI210     u0899(.A0(men_men_n927_), .A1(men_men_n926_), .B0(men_men_n897_), .Y(men_men_n928_));
  NA3        u0900(.A(c), .B(b), .C(a), .Y(men_men_n929_));
  NO3        u0901(.A(men_men_n929_), .B(men_men_n778_), .C(men_men_n196_), .Y(men_men_n930_));
  NO3        u0902(.A(men_men_n902_), .B(men_men_n48_), .C(men_men_n106_), .Y(men_men_n931_));
  AOI210     u0903(.A0(men_men_n931_), .A1(men_men_n930_), .B0(men_men_n906_), .Y(men_men_n932_));
  AN4        u0904(.A(men_men_n932_), .B(men_men_n928_), .C(men_men_n924_), .D(men_men_n922_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n900_), .B(men_men_n893_), .Y(men_men_n934_));
  AOI210     u0906(.A0(men_men_n934_), .A1(men_men_n885_), .B0(men_men_n879_), .Y(men_men_n935_));
  NAi41      u0907(.An(men_men_n918_), .B(men_men_n935_), .C(men_men_n933_), .D(men_men_n919_), .Y(men03));
  NO2        u0908(.A(men_men_n500_), .B(men_men_n558_), .Y(men_men_n937_));
  NA4        u0909(.A(men_men_n83_), .B(men_men_n82_), .C(u), .D(men_men_n196_), .Y(men_men_n938_));
  NA4        u0910(.A(men_men_n539_), .B(m), .C(men_men_n106_), .D(men_men_n196_), .Y(men_men_n939_));
  NA3        u0911(.A(men_men_n939_), .B(men_men_n347_), .C(men_men_n938_), .Y(men_men_n940_));
  NO3        u0912(.A(men_men_n940_), .B(men_men_n937_), .C(men_men_n848_), .Y(men_men_n941_));
  NOi41      u0913(.An(men_men_n719_), .B(men_men_n754_), .C(men_men_n746_), .D(men_men_n648_), .Y(men_men_n942_));
  OAI220     u0914(.A0(men_men_n942_), .A1(men_men_n629_), .B0(men_men_n941_), .B1(men_men_n550_), .Y(men_men_n943_));
  NOi31      u0915(.An(i), .B(k), .C(j), .Y(men_men_n944_));
  NA4        u0916(.A(men_men_n944_), .B(e), .C(men_men_n321_), .D(men_men_n313_), .Y(men_men_n945_));
  OAI210     u0917(.A0(men_men_n725_), .A1(men_men_n395_), .B0(men_men_n945_), .Y(men_men_n946_));
  NOi31      u0918(.An(m), .B(n), .C(f), .Y(men_men_n947_));
  NA2        u0919(.A(men_men_n947_), .B(men_men_n50_), .Y(men_men_n948_));
  AN2        u0920(.A(e), .B(c), .Y(men_men_n949_));
  NA2        u0921(.A(men_men_n949_), .B(a), .Y(men_men_n950_));
  OAI220     u0922(.A0(men_men_n950_), .A1(men_men_n948_), .B0(men_men_n772_), .B1(men_men_n401_), .Y(men_men_n951_));
  NA2        u0923(.A(men_men_n481_), .B(l), .Y(men_men_n952_));
  NOi31      u0924(.An(men_men_n759_), .B(men_men_n878_), .C(men_men_n952_), .Y(men_men_n953_));
  NO3        u0925(.A(men_men_n953_), .B(men_men_n951_), .C(men_men_n946_), .Y(men_men_n954_));
  NO2        u0926(.A(men_men_n262_), .B(a), .Y(men_men_n955_));
  INV        u0927(.A(men_men_n883_), .Y(men_men_n956_));
  NO2        u0928(.A(men_men_n82_), .B(u), .Y(men_men_n957_));
  AOI210     u0929(.A0(men_men_n957_), .A1(h), .B0(men_men_n911_), .Y(men_men_n958_));
  OR2        u0930(.A(men_men_n958_), .B(men_men_n910_), .Y(men_men_n959_));
  NA3        u0931(.A(men_men_n959_), .B(men_men_n956_), .C(men_men_n954_), .Y(men_men_n960_));
  NO4        u0932(.A(men_men_n960_), .B(men_men_n943_), .C(men_men_n727_), .D(men_men_n531_), .Y(men_men_n961_));
  NA2        u0933(.A(c), .B(b), .Y(men_men_n962_));
  NO2        u0934(.A(n), .B(men_men_n962_), .Y(men_men_n963_));
  OAI210     u0935(.A0(men_men_n757_), .A1(men_men_n739_), .B0(men_men_n388_), .Y(men_men_n964_));
  OAI210     u0936(.A0(men_men_n964_), .A1(men_men_n758_), .B0(men_men_n963_), .Y(men_men_n965_));
  NAi21      u0937(.An(men_men_n396_), .B(men_men_n963_), .Y(men_men_n966_));
  NA3        u0938(.A(men_men_n402_), .B(men_men_n524_), .C(f), .Y(men_men_n967_));
  OAI210     u0939(.A0(men_men_n519_), .A1(men_men_n38_), .B0(men_men_n955_), .Y(men_men_n968_));
  NA3        u0940(.A(men_men_n968_), .B(men_men_n967_), .C(men_men_n966_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n240_), .B(men_men_n112_), .Y(men_men_n970_));
  OAI210     u0942(.A0(men_men_n970_), .A1(men_men_n266_), .B0(u), .Y(men_men_n971_));
  NO2        u0943(.A(f), .B(men_men_n929_), .Y(men_men_n972_));
  AOI210     u0944(.A0(men_men_n971_), .A1(men_men_n272_), .B0(men_men_n929_), .Y(men_men_n973_));
  AOI210     u0945(.A0(men_men_n973_), .A1(men_men_n107_), .B0(men_men_n969_), .Y(men_men_n974_));
  NO2        u0946(.A(men_men_n164_), .B(men_men_n219_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n975_), .B(m), .Y(men_men_n976_));
  NA3        u0948(.A(men_men_n786_), .B(men_men_n952_), .C(men_men_n449_), .Y(men_men_n977_));
  OAI210     u0949(.A0(men_men_n977_), .A1(men_men_n289_), .B0(men_men_n447_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n978_), .B(men_men_n976_), .Y(men_men_n979_));
  NA2        u0951(.A(men_men_n144_), .B(men_men_n32_), .Y(men_men_n980_));
  AOI210     u0952(.A0(men_men_n817_), .A1(men_men_n980_), .B0(men_men_n197_), .Y(men_men_n981_));
  OAI210     u0953(.A0(men_men_n981_), .A1(men_men_n422_), .B0(men_men_n972_), .Y(men_men_n982_));
  NO2        u0954(.A(men_men_n349_), .B(men_men_n348_), .Y(men_men_n983_));
  INV        u0955(.A(men_men_n982_), .Y(men_men_n984_));
  NO2        u0956(.A(men_men_n984_), .B(men_men_n979_), .Y(men_men_n985_));
  NA4        u0957(.A(men_men_n985_), .B(men_men_n974_), .C(men_men_n965_), .D(men_men_n961_), .Y(men00));
  NO2        u0958(.A(men_men_n279_), .B(men_men_n254_), .Y(men_men_n987_));
  NO2        u0959(.A(men_men_n987_), .B(men_men_n541_), .Y(men_men_n988_));
  AOI210     u0960(.A0(men_men_n777_), .A1(men_men_n802_), .B0(men_men_n946_), .Y(men_men_n989_));
  NO3        u0961(.A(men_men_n923_), .B(men_men_n814_), .C(men_men_n645_), .Y(men_men_n990_));
  NA3        u0962(.A(men_men_n990_), .B(men_men_n989_), .C(men_men_n849_), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n483_), .B(f), .Y(men_men_n992_));
  NO2        u0964(.A(men_men_n992_), .B(men_men_n886_), .Y(men_men_n993_));
  NO4        u0965(.A(men_men_n993_), .B(men_men_n991_), .C(men_men_n988_), .D(men_men_n904_), .Y(men_men_n994_));
  NA3        u0966(.A(men_men_n152_), .B(men_men_n45_), .C(men_men_n44_), .Y(men_men_n995_));
  NOi31      u0967(.An(n), .B(m), .C(i), .Y(men_men_n996_));
  NA3        u0968(.A(men_men_n996_), .B(men_men_n599_), .C(men_men_n50_), .Y(men_men_n997_));
  OAI210     u0969(.A0(men_men_n1311_), .A1(men_men_n995_), .B0(men_men_n997_), .Y(men_men_n998_));
  INV        u0970(.A(men_men_n540_), .Y(men_men_n999_));
  NO4        u0971(.A(men_men_n999_), .B(men_men_n998_), .C(men_men_n983_), .D(men_men_n787_), .Y(men_men_n1000_));
  NO4        u0972(.A(men_men_n1306_), .B(men_men_n333_), .C(men_men_n962_), .D(men_men_n57_), .Y(men_men_n1001_));
  NA3        u0973(.A(men_men_n359_), .B(men_men_n202_), .C(u), .Y(men_men_n1002_));
  OR2        u0974(.A(men_men_n1002_), .B(men_men_n1311_), .Y(men_men_n1003_));
  NO2        u0975(.A(h), .B(u), .Y(men_men_n1004_));
  NA3        u0976(.A(men_men_n473_), .B(men_men_n443_), .C(men_men_n877_), .Y(men_men_n1005_));
  OAI220     u0977(.A0(men_men_n500_), .A1(men_men_n558_), .B0(men_men_n87_), .B1(men_men_n86_), .Y(men_men_n1006_));
  AOI220     u0978(.A0(men_men_n1006_), .A1(men_men_n508_), .B0(men_men_n805_), .B1(d), .Y(men_men_n1007_));
  NA3        u0979(.A(men_men_n1007_), .B(men_men_n1005_), .C(men_men_n1003_), .Y(men_men_n1008_));
  NO3        u0980(.A(men_men_n1008_), .B(men_men_n1001_), .C(men_men_n246_), .Y(men_men_n1009_));
  INV        u0981(.A(men_men_n301_), .Y(men_men_n1010_));
  INV        u0982(.A(men_men_n542_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n1011_), .B(men_men_n1010_), .Y(men_men_n1012_));
  NO2        u0984(.A(men_men_n221_), .B(men_men_n163_), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n1013_), .B(men_men_n402_), .Y(men_men_n1014_));
  NA3        u0986(.A(men_men_n161_), .B(men_men_n106_), .C(u), .Y(men_men_n1015_));
  NA3        u0987(.A(men_men_n443_), .B(men_men_n39_), .C(f), .Y(men_men_n1016_));
  NOi31      u0988(.An(j), .B(men_men_n1016_), .C(men_men_n1015_), .Y(men_men_n1017_));
  NAi21      u0989(.An(men_men_n1017_), .B(men_men_n1014_), .Y(men_men_n1018_));
  NO2        u0990(.A(men_men_n253_), .B(men_men_n73_), .Y(men_men_n1019_));
  NO3        u0991(.A(men_men_n401_), .B(men_men_n735_), .C(n), .Y(men_men_n1020_));
  AOI210     u0992(.A0(men_men_n1020_), .A1(men_men_n1019_), .B0(men_men_n918_), .Y(men_men_n1021_));
  NAi31      u0993(.An(men_men_n889_), .B(men_men_n1021_), .C(men_men_n72_), .Y(men_men_n1022_));
  NO4        u0994(.A(men_men_n1022_), .B(men_men_n1018_), .C(men_men_n1012_), .D(men_men_n491_), .Y(men_men_n1023_));
  AN3        u0995(.A(men_men_n1023_), .B(men_men_n1009_), .C(men_men_n1000_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n508_), .B(men_men_n97_), .Y(men_men_n1025_));
  NA3        u0997(.A(men_men_n947_), .B(men_men_n563_), .C(men_men_n442_), .Y(men_men_n1026_));
  NA4        u0998(.A(men_men_n1026_), .B(men_men_n527_), .C(men_men_n1025_), .D(men_men_n224_), .Y(men_men_n1027_));
  NA2        u0999(.A(men_men_n940_), .B(men_men_n508_), .Y(men_men_n1028_));
  NA4        u1000(.A(men_men_n599_), .B(men_men_n189_), .C(men_men_n202_), .D(men_men_n148_), .Y(men_men_n1029_));
  NA3        u1001(.A(men_men_n1029_), .B(men_men_n1028_), .C(men_men_n276_), .Y(men_men_n1030_));
  OAI210     u1002(.A0(men_men_n441_), .A1(men_men_n113_), .B0(men_men_n760_), .Y(men_men_n1031_));
  AOI220     u1003(.A0(men_men_n1031_), .A1(men_men_n977_), .B0(men_men_n526_), .B1(men_men_n383_), .Y(men_men_n1032_));
  OR3        u1004(.A(men_men_n886_), .B(men_men_n204_), .C(e), .Y(men_men_n1033_));
  NO2        u1005(.A(men_men_n200_), .B(men_men_n197_), .Y(men_men_n1034_));
  NA2        u1006(.A(men_men_n750_), .B(men_men_n1034_), .Y(men_men_n1035_));
  OAI210     u1007(.A0(men_men_n334_), .A1(men_men_n290_), .B0(men_men_n424_), .Y(men_men_n1036_));
  NA4        u1008(.A(men_men_n1036_), .B(men_men_n1035_), .C(men_men_n1033_), .D(men_men_n1032_), .Y(men_men_n1037_));
  INV        u1009(.A(men_men_n726_), .Y(men_men_n1038_));
  AOI220     u1010(.A0(men_men_n810_), .A1(d), .B0(men_men_n599_), .B1(men_men_n226_), .Y(men_men_n1039_));
  NO2        u1011(.A(men_men_n66_), .B(h), .Y(men_men_n1040_));
  NO2        u1012(.A(men_men_n886_), .B(men_men_n655_), .Y(men_men_n1041_));
  NO2        u1013(.A(men_men_n915_), .B(men_men_n122_), .Y(men_men_n1042_));
  AN2        u1014(.A(men_men_n1042_), .B(men_men_n927_), .Y(men_men_n1043_));
  OAI210     u1015(.A0(men_men_n1043_), .A1(men_men_n1041_), .B0(men_men_n1040_), .Y(men_men_n1044_));
  NA4        u1016(.A(men_men_n1044_), .B(men_men_n1039_), .C(men_men_n1038_), .D(men_men_n762_), .Y(men_men_n1045_));
  NO4        u1017(.A(men_men_n1045_), .B(men_men_n1037_), .C(men_men_n1030_), .D(men_men_n1027_), .Y(men_men_n1046_));
  NA2        u1018(.A(men_men_n740_), .B(men_men_n678_), .Y(men_men_n1047_));
  NA4        u1019(.A(men_men_n1047_), .B(men_men_n1046_), .C(men_men_n1024_), .D(men_men_n994_), .Y(men01));
  AN2        u1020(.A(men_men_n868_), .B(men_men_n867_), .Y(men_men_n1049_));
  NO3        u1021(.A(men_men_n715_), .B(men_men_n457_), .C(men_men_n260_), .Y(men_men_n1050_));
  NA2        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .Y(men_men_n1051_));
  NA2        u1023(.A(men_men_n551_), .B(men_men_n85_), .Y(men_men_n1052_));
  NA3        u1024(.A(men_men_n1052_), .B(men_men_n785_), .C(men_men_n312_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n643_), .B(men_men_n92_), .Y(men_men_n1054_));
  NO2        u1026(.A(men_men_n1054_), .B(i), .Y(men_men_n1055_));
  OAI210     u1027(.A0(men_men_n698_), .A1(n), .B0(men_men_n1029_), .Y(men_men_n1056_));
  AOI210     u1028(.A0(men_men_n1055_), .A1(men_men_n589_), .B0(men_men_n1056_), .Y(men_men_n1057_));
  OA220      u1029(.A0(men_men_n1310_), .A1(men_men_n548_), .B0(men_men_n609_), .B1(men_men_n347_), .Y(men_men_n1058_));
  NAi41      u1030(.An(men_men_n147_), .B(men_men_n1058_), .C(men_men_n1057_), .D(men_men_n776_), .Y(men_men_n1059_));
  NO4        u1031(.A(men_men_n618_), .B(men_men_n1059_), .C(men_men_n1053_), .D(men_men_n1051_), .Y(men_men_n1060_));
  INV        u1032(.A(men_men_n190_), .Y(men_men_n1061_));
  NA2        u1033(.A(men_men_n1061_), .B(men_men_n504_), .Y(men_men_n1062_));
  NA2        u1034(.A(men_men_n528_), .B(a), .Y(men_men_n1063_));
  AOI210     u1035(.A0(men_men_n187_), .A1(men_men_n84_), .B0(men_men_n196_), .Y(men_men_n1064_));
  OAI210     u1036(.A0(men_men_n1309_), .A1(men_men_n402_), .B0(men_men_n1064_), .Y(men_men_n1065_));
  OAI210     u1037(.A0(men_men_n336_), .A1(men_men_n33_), .B0(k), .Y(men_men_n1066_));
  OR2        u1038(.A(men_men_n1066_), .B(men_men_n311_), .Y(men_men_n1067_));
  NA4        u1039(.A(men_men_n1067_), .B(men_men_n1065_), .C(men_men_n1063_), .D(men_men_n1062_), .Y(men_men_n1068_));
  AOI210     u1040(.A0(men_men_n556_), .A1(men_men_n111_), .B0(men_men_n559_), .Y(men_men_n1069_));
  OAI210     u1041(.A0(men_men_n1310_), .A1(men_men_n555_), .B0(men_men_n1069_), .Y(men_men_n1070_));
  NA2        u1042(.A(men_men_n259_), .B(men_men_n178_), .Y(men_men_n1071_));
  OAI210     u1043(.A0(men_men_n1071_), .A1(men_men_n361_), .B0(f), .Y(men_men_n1072_));
  OAI210     u1044(.A0(men_men_n1055_), .A1(men_men_n305_), .B0(men_men_n619_), .Y(men_men_n1073_));
  NA3        u1045(.A(men_men_n1073_), .B(men_men_n1072_), .C(men_men_n701_), .Y(men_men_n1074_));
  NO3        u1046(.A(men_men_n1074_), .B(men_men_n1070_), .C(men_men_n1068_), .Y(men_men_n1075_));
  NA2        u1047(.A(men_men_n480_), .B(men_men_n56_), .Y(men_men_n1076_));
  NA3        u1048(.A(men_men_n995_), .B(men_men_n1076_), .C(men_men_n677_), .Y(men_men_n1077_));
  INV        u1049(.A(men_men_n214_), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n535_), .B(men_men_n533_), .Y(men_men_n1079_));
  NO3        u1051(.A(men_men_n78_), .B(men_men_n280_), .C(men_men_n44_), .Y(men_men_n1080_));
  INV        u1052(.A(men_men_n1080_), .Y(men_men_n1081_));
  NA3        u1053(.A(men_men_n1081_), .B(men_men_n1079_), .C(men_men_n614_), .Y(men_men_n1082_));
  BUFFER     u1054(.A(men_men_n1002_), .Y(men_men_n1083_));
  NO2        u1055(.A(men_men_n347_), .B(men_men_n71_), .Y(men_men_n1084_));
  INV        u1056(.A(men_men_n1084_), .Y(men_men_n1085_));
  NA3        u1057(.A(men_men_n1085_), .B(men_men_n1083_), .C(men_men_n362_), .Y(men_men_n1086_));
  NO3        u1058(.A(men_men_n1086_), .B(men_men_n1082_), .C(men_men_n1077_), .Y(men_men_n1087_));
  AN2        u1059(.A(i), .B(f), .Y(men_men_n1088_));
  NO3        u1060(.A(men_men_n925_), .B(men_men_n158_), .C(men_men_n82_), .Y(men_men_n1089_));
  NO2        u1061(.A(men_men_n570_), .B(f), .Y(men_men_n1090_));
  NO4        u1062(.A(men_men_n925_), .B(men_men_n1090_), .C(men_men_n156_), .D(men_men_n82_), .Y(men_men_n1091_));
  NO3        u1063(.A(men_men_n1091_), .B(men_men_n1089_), .C(men_men_n593_), .Y(men_men_n1092_));
  NA4        u1064(.A(men_men_n1092_), .B(men_men_n1087_), .C(men_men_n1075_), .D(men_men_n1060_), .Y(men06));
  NO2        u1065(.A(men_men_n382_), .B(men_men_n525_), .Y(men_men_n1094_));
  OAI210     u1066(.A0(men_men_n107_), .A1(men_men_n247_), .B0(men_men_n1094_), .Y(men_men_n1095_));
  NO3        u1067(.A(men_men_n560_), .B(men_men_n720_), .C(men_men_n561_), .Y(men_men_n1096_));
  BUFFER     u1068(.A(men_men_n772_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n1097_), .B(men_men_n1095_), .Y(men_men_n1098_));
  NO3        u1070(.A(men_men_n1098_), .B(men_men_n1082_), .C(men_men_n235_), .Y(men_men_n1099_));
  NO2        u1071(.A(men_men_n280_), .B(men_men_n44_), .Y(men_men_n1100_));
  NO2        u1072(.A(men_men_n1100_), .B(men_men_n1078_), .Y(men_men_n1101_));
  INV        u1073(.A(men_men_n1088_), .Y(men_men_n1102_));
  AOI210     u1074(.A0(men_men_n1102_), .A1(men_men_n1101_), .B0(men_men_n317_), .Y(men_men_n1103_));
  OAI210     u1075(.A0(men_men_n84_), .A1(men_men_n39_), .B0(men_men_n617_), .Y(men_men_n1104_));
  NA2        u1076(.A(men_men_n1104_), .B(men_men_n597_), .Y(men_men_n1105_));
  NO2        u1077(.A(men_men_n564_), .B(men_men_n948_), .Y(men_men_n1106_));
  NO2        u1078(.A(men_men_n436_), .B(men_men_n228_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n1107_), .B(men_men_n1106_), .Y(men_men_n1108_));
  INV        u1080(.A(men_men_n559_), .Y(men_men_n1109_));
  NA3        u1081(.A(men_men_n1109_), .B(men_men_n1108_), .C(men_men_n1105_), .Y(men_men_n1110_));
  NO2        u1082(.A(men_men_n671_), .B(men_men_n345_), .Y(men_men_n1111_));
  NOi21      u1083(.An(men_men_n1111_), .B(men_men_n48_), .Y(men_men_n1112_));
  NO4        u1084(.A(men_men_n810_), .B(men_men_n1112_), .C(men_men_n1110_), .D(men_men_n1103_), .Y(men_men_n1113_));
  NO2        u1085(.A(men_men_n714_), .B(men_men_n255_), .Y(men_men_n1114_));
  OAI220     u1086(.A0(men_men_n661_), .A1(men_men_n46_), .B0(men_men_n206_), .B1(men_men_n571_), .Y(men_men_n1115_));
  OAI210     u1087(.A0(men_men_n255_), .A1(c), .B0(men_men_n596_), .Y(men_men_n1116_));
  AOI220     u1088(.A0(men_men_n1116_), .A1(men_men_n1115_), .B0(men_men_n1114_), .B1(men_men_n247_), .Y(men_men_n1117_));
  NO3        u1089(.A(h), .B(men_men_n98_), .C(men_men_n262_), .Y(men_men_n1118_));
  OAI220     u1090(.A0(men_men_n636_), .A1(men_men_n228_), .B0(men_men_n485_), .B1(men_men_n487_), .Y(men_men_n1119_));
  NO2        u1091(.A(men_men_n558_), .B(j), .Y(men_men_n1120_));
  NOi21      u1092(.An(men_men_n1120_), .B(men_men_n71_), .Y(men_men_n1121_));
  NO4        u1093(.A(men_men_n1121_), .B(men_men_n1119_), .C(men_men_n1118_), .D(men_men_n951_), .Y(men_men_n1122_));
  NAi31      u1094(.An(men_men_n671_), .B(men_men_n81_), .C(men_men_n186_), .Y(men_men_n1123_));
  NA4        u1095(.A(men_men_n1123_), .B(men_men_n1122_), .C(men_men_n1117_), .D(men_men_n1039_), .Y(men_men_n1124_));
  NOi31      u1096(.An(men_men_n1096_), .B(men_men_n440_), .C(men_men_n370_), .Y(men_men_n1125_));
  OR3        u1097(.A(men_men_n1125_), .B(men_men_n698_), .C(men_men_n513_), .Y(men_men_n1126_));
  NA2        u1098(.A(men_men_n535_), .B(men_men_n424_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n1120_), .B(men_men_n705_), .Y(men_men_n1128_));
  NA3        u1100(.A(men_men_n1128_), .B(men_men_n1127_), .C(men_men_n1126_), .Y(men_men_n1129_));
  NO3        u1101(.A(men_men_n792_), .B(men_men_n764_), .C(men_men_n476_), .Y(men_men_n1130_));
  INV        u1102(.A(men_men_n1130_), .Y(men_men_n1131_));
  NAi21      u1103(.An(j), .B(i), .Y(men_men_n1132_));
  NO4        u1104(.A(men_men_n1090_), .B(men_men_n1132_), .C(men_men_n418_), .D(men_men_n217_), .Y(men_men_n1133_));
  NO4        u1105(.A(men_men_n1133_), .B(men_men_n1131_), .C(men_men_n1129_), .D(men_men_n1124_), .Y(men_men_n1134_));
  NA4        u1106(.A(men_men_n1134_), .B(men_men_n1113_), .C(men_men_n1099_), .D(men_men_n1092_), .Y(men07));
  NOi21      u1107(.An(j), .B(k), .Y(men_men_n1136_));
  NAi32      u1108(.An(m), .Bn(b), .C(n), .Y(men_men_n1137_));
  NAi21      u1109(.An(f), .B(c), .Y(men_men_n1138_));
  OR2        u1110(.A(e), .B(d), .Y(men_men_n1139_));
  NOi31      u1111(.An(n), .B(m), .C(b), .Y(men_men_n1140_));
  NOi41      u1112(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1141_));
  NA3        u1113(.A(men_men_n1141_), .B(men_men_n763_), .C(men_men_n384_), .Y(men_men_n1142_));
  NO2        u1114(.A(men_men_n1142_), .B(men_men_n54_), .Y(men_men_n1143_));
  NA2        u1115(.A(men_men_n927_), .B(men_men_n202_), .Y(men_men_n1144_));
  NO2        u1116(.A(men_men_n1144_), .B(men_men_n59_), .Y(men_men_n1145_));
  NO2        u1117(.A(k), .B(i), .Y(men_men_n1146_));
  NA2        u1118(.A(men_men_n82_), .B(men_men_n44_), .Y(men_men_n1147_));
  NO2        u1119(.A(men_men_n892_), .B(men_men_n418_), .Y(men_men_n1148_));
  NA3        u1120(.A(men_men_n1148_), .B(men_men_n1147_), .C(men_men_n197_), .Y(men_men_n1149_));
  NO2        u1121(.A(men_men_n902_), .B(men_men_n284_), .Y(men_men_n1150_));
  NA2        u1122(.A(men_men_n514_), .B(men_men_n79_), .Y(men_men_n1151_));
  NA2        u1123(.A(men_men_n1151_), .B(men_men_n1149_), .Y(men_men_n1152_));
  NO3        u1124(.A(men_men_n1152_), .B(men_men_n1145_), .C(men_men_n1143_), .Y(men_men_n1153_));
  OR2        u1125(.A(h), .B(f), .Y(men_men_n1154_));
  NO3        u1126(.A(n), .B(m), .C(i), .Y(men_men_n1155_));
  OAI210     u1127(.A0(men_men_n949_), .A1(men_men_n142_), .B0(men_men_n1155_), .Y(men_men_n1156_));
  NO2        u1128(.A(i), .B(u), .Y(men_men_n1157_));
  OR3        u1129(.A(men_men_n1157_), .B(men_men_n1137_), .C(men_men_n70_), .Y(men_men_n1158_));
  OAI220     u1130(.A0(men_men_n1158_), .A1(men_men_n460_), .B0(men_men_n1156_), .B1(men_men_n1154_), .Y(men_men_n1159_));
  NA3        u1131(.A(men_men_n633_), .B(men_men_n624_), .C(men_men_n106_), .Y(men_men_n1160_));
  NA3        u1132(.A(men_men_n1140_), .B(men_men_n898_), .C(h), .Y(men_men_n1161_));
  AOI210     u1133(.A0(men_men_n1161_), .A1(men_men_n1160_), .B0(men_men_n44_), .Y(men_men_n1162_));
  NA2        u1134(.A(men_men_n1155_), .B(men_men_n595_), .Y(men_men_n1163_));
  NO2        u1135(.A(l), .B(k), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n1162_), .B(men_men_n1159_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n134_), .B(h), .Y(men_men_n1166_));
  NO2        u1138(.A(u), .B(c), .Y(men_men_n1167_));
  NO2        u1139(.A(men_men_n429_), .B(a), .Y(men_men_n1168_));
  NA3        u1140(.A(men_men_n1168_), .B(men_men_n1304_), .C(men_men_n107_), .Y(men_men_n1169_));
  NO2        u1141(.A(i), .B(h), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n1170_), .B(men_men_n202_), .Y(men_men_n1171_));
  AOI210     u1143(.A0(men_men_n236_), .A1(men_men_n109_), .B0(men_men_n504_), .Y(men_men_n1172_));
  NO2        u1144(.A(men_men_n1172_), .B(men_men_n1171_), .Y(men_men_n1173_));
  NOi31      u1145(.An(m), .B(n), .C(b), .Y(men_men_n1174_));
  NOi31      u1146(.An(f), .B(d), .C(c), .Y(men_men_n1175_));
  INV        u1147(.A(men_men_n1173_), .Y(men_men_n1176_));
  OAI210     u1148(.A0(men_men_n164_), .A1(men_men_n499_), .B0(men_men_n899_), .Y(men_men_n1177_));
  NO3        u1149(.A(men_men_n40_), .B(i), .C(h), .Y(men_men_n1178_));
  AN3        u1150(.A(men_men_n1177_), .B(men_men_n1176_), .C(men_men_n1169_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n1140_), .B(men_men_n357_), .Y(men_men_n1180_));
  NO2        u1152(.A(men_men_n1180_), .B(men_men_n884_), .Y(men_men_n1181_));
  NO2        u1153(.A(men_men_n170_), .B(b), .Y(men_men_n1182_));
  NA2        u1154(.A(men_men_n996_), .B(men_men_n1182_), .Y(men_men_n1183_));
  NO2        u1155(.A(i), .B(men_men_n196_), .Y(men_men_n1184_));
  NA4        u1156(.A(men_men_n975_), .B(men_men_n1184_), .C(men_men_n99_), .D(m), .Y(men_men_n1185_));
  NAi31      u1157(.An(men_men_n1181_), .B(men_men_n1185_), .C(men_men_n1183_), .Y(men_men_n1186_));
  NO4        u1158(.A(men_men_n122_), .B(u), .C(f), .D(e), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n177_), .B(men_men_n94_), .Y(men_men_n1188_));
  OR2        u1160(.A(e), .B(a), .Y(men_men_n1189_));
  NOi41      u1161(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n1190_), .B(men_men_n107_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n1141_), .B(men_men_n1164_), .Y(men_men_n1192_));
  NA2        u1164(.A(men_men_n1192_), .B(men_men_n1191_), .Y(men_men_n1193_));
  OR3        u1165(.A(men_men_n513_), .B(men_men_n512_), .C(men_men_n106_), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n947_), .B(men_men_n381_), .Y(men_men_n1195_));
  OAI220     u1167(.A0(men_men_n1195_), .A1(men_men_n411_), .B0(men_men_n1194_), .B1(men_men_n280_), .Y(men_men_n1196_));
  AO210      u1168(.A0(men_men_n1196_), .A1(men_men_n109_), .B0(men_men_n1193_), .Y(men_men_n1197_));
  NO2        u1169(.A(men_men_n1197_), .B(men_men_n1186_), .Y(men_men_n1198_));
  NA4        u1170(.A(men_men_n1198_), .B(men_men_n1179_), .C(men_men_n1165_), .D(men_men_n1153_), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n962_), .B(men_men_n104_), .Y(men_men_n1200_));
  NA2        u1172(.A(men_men_n357_), .B(men_men_n54_), .Y(men_men_n1201_));
  AOI210     u1173(.A0(men_men_n1201_), .A1(men_men_n892_), .B0(men_men_n1163_), .Y(men_men_n1202_));
  NA2        u1174(.A(men_men_n198_), .B(men_men_n161_), .Y(men_men_n1203_));
  AOI210     u1175(.A0(men_men_n1203_), .A1(men_men_n1015_), .B0(men_men_n1201_), .Y(men_men_n1204_));
  NO2        u1176(.A(men_men_n921_), .B(men_men_n917_), .Y(men_men_n1205_));
  NO3        u1177(.A(men_men_n1205_), .B(men_men_n1204_), .C(men_men_n1202_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n1178_), .B(men_men_n1139_), .C(men_men_n947_), .Y(men_men_n1207_));
  NO3        u1179(.A(men_men_n917_), .B(men_men_n545_), .C(u), .Y(men_men_n1208_));
  NOi21      u1180(.An(men_men_n1203_), .B(men_men_n1208_), .Y(men_men_n1209_));
  AOI210     u1181(.A0(men_men_n1209_), .A1(men_men_n1188_), .B0(men_men_n892_), .Y(men_men_n1210_));
  INV        u1182(.A(men_men_n48_), .Y(men_men_n1211_));
  AOI220     u1183(.A0(men_men_n1211_), .A1(men_men_n1004_), .B0(men_men_n729_), .B1(men_men_n177_), .Y(men_men_n1212_));
  INV        u1184(.A(men_men_n1212_), .Y(men_men_n1213_));
  OAI220     u1185(.A0(men_men_n613_), .A1(u), .B0(men_men_n206_), .B1(c), .Y(men_men_n1214_));
  AOI210     u1186(.A0(men_men_n1182_), .A1(men_men_n40_), .B0(men_men_n1214_), .Y(men_men_n1215_));
  NO2        u1187(.A(men_men_n122_), .B(l), .Y(men_men_n1216_));
  NO2        u1188(.A(men_men_n206_), .B(k), .Y(men_men_n1217_));
  OAI210     u1189(.A0(men_men_n1217_), .A1(men_men_n1170_), .B0(men_men_n1216_), .Y(men_men_n1218_));
  OAI220     u1190(.A0(men_men_n1218_), .A1(e), .B0(men_men_n1215_), .B1(men_men_n158_), .Y(men_men_n1219_));
  NO3        u1191(.A(men_men_n1194_), .B(men_men_n443_), .C(men_men_n331_), .Y(men_men_n1220_));
  NO4        u1192(.A(men_men_n1220_), .B(men_men_n1219_), .C(men_men_n1213_), .D(men_men_n1210_), .Y(men_men_n1221_));
  NO2        u1193(.A(men_men_n48_), .B(men_men_n545_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n930_), .B(men_men_n1222_), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n917_), .B(h), .Y(men_men_n1224_));
  NO2        u1196(.A(men_men_n1223_), .B(j), .Y(men_men_n1225_));
  NA3        u1197(.A(men_men_n1200_), .B(men_men_n443_), .C(f), .Y(men_men_n1226_));
  NO2        u1198(.A(men_men_n1136_), .B(men_men_n41_), .Y(men_men_n1227_));
  AOI210     u1199(.A0(men_men_n107_), .A1(men_men_n39_), .B0(men_men_n1227_), .Y(men_men_n1228_));
  NO2        u1200(.A(men_men_n1228_), .B(men_men_n1226_), .Y(men_men_n1229_));
  AOI210     u1201(.A0(men_men_n499_), .A1(h), .B0(men_men_n67_), .Y(men_men_n1230_));
  NA2        u1202(.A(men_men_n1230_), .B(men_men_n1168_), .Y(men_men_n1231_));
  NO2        u1203(.A(men_men_n1132_), .B(men_men_n156_), .Y(men_men_n1232_));
  NOi21      u1204(.An(d), .B(f), .Y(men_men_n1233_));
  NO3        u1205(.A(men_men_n1175_), .B(men_men_n1233_), .C(men_men_n39_), .Y(men_men_n1234_));
  NA2        u1206(.A(men_men_n1234_), .B(men_men_n1232_), .Y(men_men_n1235_));
  NO2        u1207(.A(men_men_n1139_), .B(f), .Y(men_men_n1236_));
  NA2        u1208(.A(men_men_n1168_), .B(men_men_n1227_), .Y(men_men_n1237_));
  NO2        u1209(.A(men_men_n280_), .B(c), .Y(men_men_n1238_));
  NA2        u1210(.A(men_men_n1238_), .B(men_men_n514_), .Y(men_men_n1239_));
  NA4        u1211(.A(men_men_n1239_), .B(men_men_n1237_), .C(men_men_n1235_), .D(men_men_n1231_), .Y(men_men_n1240_));
  NO3        u1212(.A(men_men_n1240_), .B(men_men_n1229_), .C(men_men_n1225_), .Y(men_men_n1241_));
  NA4        u1213(.A(men_men_n1241_), .B(men_men_n1221_), .C(men_men_n1207_), .D(men_men_n1206_), .Y(men_men_n1242_));
  OAI220     u1214(.A0(men_men_n443_), .A1(men_men_n280_), .B0(men_men_n121_), .B1(men_men_n57_), .Y(men_men_n1243_));
  NA2        u1215(.A(men_men_n1243_), .B(men_men_n1150_), .Y(men_men_n1244_));
  OAI210     u1216(.A0(men_men_n1187_), .A1(men_men_n1140_), .B0(men_men_n770_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n1245_), .B(men_men_n1244_), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n1167_), .B(men_men_n1233_), .Y(men_men_n1247_));
  NO2        u1219(.A(men_men_n1247_), .B(m), .Y(men_men_n1248_));
  NA3        u1220(.A(men_men_n927_), .B(men_men_n102_), .C(men_men_n202_), .Y(men_men_n1249_));
  NA2        u1221(.A(men_men_n104_), .B(men_men_n1174_), .Y(men_men_n1250_));
  NA2        u1222(.A(men_men_n1250_), .B(men_men_n1249_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n1251_), .B(men_men_n1248_), .C(men_men_n1246_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n1138_), .B(e), .Y(men_men_n1253_));
  NA2        u1225(.A(men_men_n1253_), .B(men_men_n379_), .Y(men_men_n1254_));
  NA2        u1226(.A(men_men_n957_), .B(men_men_n585_), .Y(men_men_n1255_));
  OR3        u1227(.A(men_men_n1217_), .B(men_men_n1040_), .C(men_men_n122_), .Y(men_men_n1256_));
  OAI220     u1228(.A0(men_men_n1256_), .A1(men_men_n1254_), .B0(men_men_n1255_), .B1(men_men_n420_), .Y(men_men_n1257_));
  NO3        u1229(.A(men_men_n1194_), .B(men_men_n331_), .C(a), .Y(men_men_n1258_));
  NO2        u1230(.A(men_men_n1258_), .B(men_men_n1257_), .Y(men_men_n1259_));
  NO2        u1231(.A(men_men_n1189_), .B(f), .Y(men_men_n1260_));
  NA2        u1232(.A(men_men_n1260_), .B(men_men_n1147_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n1261_), .B(men_men_n48_), .Y(men_men_n1262_));
  NO2        u1234(.A(men_men_n48_), .B(l), .Y(men_men_n1263_));
  INV        u1235(.A(men_men_n460_), .Y(men_men_n1264_));
  OAI210     u1236(.A0(men_men_n1264_), .A1(men_men_n930_), .B0(men_men_n1263_), .Y(men_men_n1265_));
  NO2        u1237(.A(men_men_n231_), .B(u), .Y(men_men_n1266_));
  NO2        u1238(.A(m), .B(i), .Y(men_men_n1267_));
  AOI220     u1239(.A0(men_men_n1267_), .A1(men_men_n1166_), .B0(men_men_n909_), .B1(men_men_n1266_), .Y(men_men_n1268_));
  NA2        u1240(.A(men_men_n1268_), .B(men_men_n1265_), .Y(men_men_n1269_));
  NO2        u1241(.A(men_men_n1269_), .B(men_men_n1262_), .Y(men_men_n1270_));
  NA3        u1242(.A(men_men_n1270_), .B(men_men_n1259_), .C(men_men_n1252_), .Y(men_men_n1271_));
  NA3        u1243(.A(men_men_n816_), .B(men_men_n126_), .C(men_men_n45_), .Y(men_men_n1272_));
  AOI210     u1244(.A0(men_men_n135_), .A1(c), .B0(men_men_n1272_), .Y(men_men_n1273_));
  OAI210     u1245(.A0(men_men_n545_), .A1(u), .B0(men_men_n167_), .Y(men_men_n1274_));
  NA2        u1246(.A(men_men_n1274_), .B(men_men_n1224_), .Y(men_men_n1275_));
  NO2        u1247(.A(men_men_n70_), .B(c), .Y(men_men_n1276_));
  NO4        u1248(.A(men_men_n1154_), .B(men_men_n168_), .C(men_men_n426_), .D(men_men_n44_), .Y(men_men_n1277_));
  AOI210     u1249(.A0(men_men_n1232_), .A1(men_men_n1276_), .B0(men_men_n1277_), .Y(men_men_n1278_));
  NA2        u1250(.A(men_men_n1278_), .B(men_men_n1275_), .Y(men_men_n1279_));
  NO2        u1251(.A(men_men_n1279_), .B(men_men_n1273_), .Y(men_men_n1280_));
  NO2        u1252(.A(men_men_n1272_), .B(men_men_n104_), .Y(men_men_n1281_));
  INV        u1253(.A(men_men_n1281_), .Y(men_men_n1282_));
  AN2        u1254(.A(men_men_n927_), .B(men_men_n915_), .Y(men_men_n1283_));
  AOI220     u1255(.A0(men_men_n1267_), .A1(men_men_n595_), .B0(men_men_n1305_), .B1(men_men_n145_), .Y(men_men_n1284_));
  NOi31      u1256(.An(men_men_n30_), .B(men_men_n1284_), .C(n), .Y(men_men_n1285_));
  AOI210     u1257(.A0(men_men_n1283_), .A1(men_men_n996_), .B0(men_men_n1285_), .Y(men_men_n1286_));
  NO2        u1258(.A(men_men_n1226_), .B(men_men_n67_), .Y(men_men_n1287_));
  NO2        u1259(.A(men_men_n1146_), .B(men_men_n111_), .Y(men_men_n1288_));
  NO2        u1260(.A(men_men_n1288_), .B(men_men_n1180_), .Y(men_men_n1289_));
  NO2        u1261(.A(men_men_n1289_), .B(men_men_n1287_), .Y(men_men_n1290_));
  NA4        u1262(.A(men_men_n1290_), .B(men_men_n1286_), .C(men_men_n1282_), .D(men_men_n1280_), .Y(men_men_n1291_));
  OR4        u1263(.A(men_men_n1291_), .B(men_men_n1271_), .C(men_men_n1242_), .D(men_men_n1199_), .Y(men04));
  NOi21      u1264(.An(men_men_n1187_), .B(men_men_n886_), .Y(men_men_n1293_));
  NA2        u1265(.A(men_men_n1236_), .B(men_men_n729_), .Y(men_men_n1294_));
  NO4        u1266(.A(men_men_n1294_), .B(men_men_n878_), .C(men_men_n461_), .D(j), .Y(men_men_n1295_));
  OR3        u1267(.A(men_men_n1295_), .B(men_men_n1293_), .C(men_men_n901_), .Y(men_men_n1296_));
  NO3        u1268(.A(men_men_n1147_), .B(men_men_n86_), .C(k), .Y(men_men_n1297_));
  AOI210     u1269(.A0(men_men_n1297_), .A1(men_men_n895_), .B0(men_men_n1017_), .Y(men_men_n1298_));
  NA2        u1270(.A(men_men_n1298_), .B(men_men_n1044_), .Y(men_men_n1299_));
  NO4        u1271(.A(men_men_n1299_), .B(men_men_n1296_), .C(men_men_n907_), .D(men_men_n891_), .Y(men_men_n1300_));
  NA4        u1272(.A(men_men_n1300_), .B(men_men_n959_), .C(men_men_n945_), .D(men_men_n933_), .Y(men05));
  INV        u1273(.A(i), .Y(men_men_n1304_));
  INV        u1274(.A(j), .Y(men_men_n1305_));
  INV        u1275(.A(men_men_n202_), .Y(men_men_n1306_));
  INV        u1276(.A(men_men_n776_), .Y(men_men_n1307_));
  INV        u1277(.A(n), .Y(men_men_n1308_));
  INV        u1278(.A(n), .Y(men_men_n1309_));
  INV        u1279(.A(k), .Y(men_men_n1310_));
  INV        u1280(.A(d), .Y(men_men_n1311_));
  INV        u1281(.A(men_men_n569_), .Y(men_men_n1312_));
  INV        u1282(.A(f), .Y(men_men_n1313_));
  INV        u1283(.A(men_men_n295_), .Y(men_men_n1314_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule