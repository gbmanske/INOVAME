library verilog;
use verilog.vl_types.all;
entity tb_lzc_4bit is
end tb_lzc_4bit;
