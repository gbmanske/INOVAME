// Benchmark "top" written by ABC on Thu Jun 20 14:59:12 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n136_, new_new_n137_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n352_, new_new_n353_,
    new_new_n354_, new_new_n355_, new_new_n356_, new_new_n357_,
    new_new_n358_, new_new_n359_, new_new_n360_, new_new_n361_,
    new_new_n362_, new_new_n363_, new_new_n364_, new_new_n365_,
    new_new_n366_, new_new_n367_, new_new_n368_, new_new_n369_,
    new_new_n370_, new_new_n371_, new_new_n372_, new_new_n373_,
    new_new_n374_, new_new_n375_, new_new_n376_, new_new_n377_,
    new_new_n378_, new_new_n379_, new_new_n380_, new_new_n381_,
    new_new_n382_, new_new_n383_, new_new_n384_, new_new_n385_,
    new_new_n386_, new_new_n387_, new_new_n388_, new_new_n389_,
    new_new_n390_, new_new_n391_, new_new_n392_, new_new_n393_,
    new_new_n394_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n460_, new_new_n461_, new_new_n462_,
    new_new_n463_, new_new_n464_, new_new_n465_, new_new_n466_,
    new_new_n467_, new_new_n468_, new_new_n469_, new_new_n470_,
    new_new_n471_, new_new_n472_, new_new_n473_, new_new_n474_,
    new_new_n475_, new_new_n476_, new_new_n477_, new_new_n478_,
    new_new_n479_, new_new_n480_, new_new_n481_, new_new_n482_,
    new_new_n483_, new_new_n484_, new_new_n485_, new_new_n486_,
    new_new_n487_, new_new_n488_, new_new_n489_, new_new_n490_,
    new_new_n491_, new_new_n492_, new_new_n493_, new_new_n494_,
    new_new_n495_, new_new_n496_, new_new_n497_, new_new_n498_,
    new_new_n499_, new_new_n500_, new_new_n501_, new_new_n502_,
    new_new_n503_, new_new_n504_, new_new_n505_, new_new_n506_,
    new_new_n508_, new_new_n509_, new_new_n510_, new_new_n511_,
    new_new_n512_, new_new_n513_, new_new_n514_, new_new_n515_,
    new_new_n516_, new_new_n517_, new_new_n518_, new_new_n519_,
    new_new_n520_, new_new_n521_, new_new_n522_, new_new_n523_,
    new_new_n524_, new_new_n525_, new_new_n526_, new_new_n527_,
    new_new_n528_, new_new_n529_, new_new_n530_, new_new_n531_,
    new_new_n532_, new_new_n533_, new_new_n534_, new_new_n535_,
    new_new_n536_, new_new_n537_, new_new_n538_, new_new_n539_,
    new_new_n540_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n645_, new_new_n646_, new_new_n647_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  NO2        g036(.A(new_new_n58_), .B(new_new_n57_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA3        g041(.A(new_new_n63_), .B(new_new_n61_), .C(new_new_n31_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_10_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(i_6_), .Y(new_new_n66_));
  NAi31      g044(.An(new_new_n66_), .B(new_new_n64_), .C(new_new_n60_), .Y(new_new_n67_));
  NA2        g045(.A(new_new_n50_), .B(i_2_), .Y(new_new_n68_));
  AOI210     g046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n69_));
  NA2        g047(.A(i_1_), .B(i_6_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n25_), .Y(new_new_n71_));
  INV        g049(.A(i_0_), .Y(new_new_n72_));
  NAi21      g050(.An(i_5_), .B(i_10_), .Y(new_new_n73_));
  NA2        g051(.A(i_5_), .B(i_9_), .Y(new_new_n74_));
  AOI210     g052(.A0(new_new_n74_), .A1(new_new_n73_), .B0(new_new_n72_), .Y(new_new_n75_));
  NO2        g053(.A(new_new_n75_), .B(new_new_n71_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n76_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n77_), .A1(new_new_n67_), .B0(i_0_), .Y(new_new_n78_));
  NA2        g056(.A(i_12_), .B(i_5_), .Y(new_new_n79_));
  NA2        g057(.A(i_2_), .B(i_8_), .Y(new_new_n80_));
  NO2        g058(.A(new_new_n80_), .B(new_new_n57_), .Y(new_new_n81_));
  NO2        g059(.A(i_3_), .B(i_9_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_7_), .Y(new_new_n83_));
  NO2        g061(.A(new_new_n82_), .B(new_new_n62_), .Y(new_new_n84_));
  INV        g062(.A(i_6_), .Y(new_new_n85_));
  NO2        g063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  INV        g064(.A(new_new_n86_), .Y(new_new_n87_));
  OAI210     g065(.A0(new_new_n84_), .A1(new_new_n81_), .B0(new_new_n87_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n62_), .Y(new_new_n91_));
  NA2        g069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  INV        g070(.A(new_new_n91_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n88_), .B0(new_new_n79_), .Y(new_new_n94_));
  AN3        g072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n95_));
  NAi21      g073(.An(i_6_), .B(i_11_), .Y(new_new_n96_));
  NO2        g074(.A(i_5_), .B(i_8_), .Y(new_new_n97_));
  NOi21      g075(.An(new_new_n97_), .B(new_new_n96_), .Y(new_new_n98_));
  AOI220     g076(.A0(new_new_n98_), .A1(new_new_n61_), .B0(new_new_n95_), .B1(new_new_n32_), .Y(new_new_n99_));
  INV        g077(.A(i_7_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n46_), .B(new_new_n100_), .Y(new_new_n101_));
  NO2        g079(.A(i_0_), .B(i_5_), .Y(new_new_n102_));
  NO2        g080(.A(new_new_n102_), .B(new_new_n85_), .Y(new_new_n103_));
  NA2        g081(.A(i_12_), .B(i_3_), .Y(new_new_n104_));
  INV        g082(.A(new_new_n104_), .Y(new_new_n105_));
  NA3        g083(.A(new_new_n105_), .B(new_new_n103_), .C(new_new_n101_), .Y(new_new_n106_));
  NAi21      g084(.An(i_7_), .B(i_11_), .Y(new_new_n107_));
  AN2        g085(.A(i_2_), .B(i_10_), .Y(new_new_n108_));
  NO2        g086(.A(new_new_n108_), .B(i_7_), .Y(new_new_n109_));
  OR2        g087(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n110_));
  NO2        g088(.A(i_8_), .B(new_new_n100_), .Y(new_new_n111_));
  NO3        g089(.A(new_new_n111_), .B(new_new_n110_), .C(new_new_n109_), .Y(new_new_n112_));
  NA2        g090(.A(i_12_), .B(i_7_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n114_));
  NA2        g092(.A(i_11_), .B(i_12_), .Y(new_new_n115_));
  INV        g093(.A(new_new_n115_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n116_), .B(new_new_n112_), .Y(new_new_n117_));
  NA3        g095(.A(new_new_n117_), .B(new_new_n106_), .C(new_new_n99_), .Y(new_new_n118_));
  NOi21      g096(.An(i_1_), .B(i_5_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_11_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n100_), .B(new_new_n37_), .Y(new_new_n121_));
  NA2        g099(.A(i_7_), .B(new_new_n25_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n122_), .B(new_new_n121_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n123_), .B(new_new_n46_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n125_));
  NAi21      g103(.An(i_3_), .B(i_8_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n61_), .Y(new_new_n127_));
  NOi31      g105(.An(new_new_n127_), .B(new_new_n125_), .C(new_new_n124_), .Y(new_new_n128_));
  NO2        g106(.A(i_1_), .B(new_new_n85_), .Y(new_new_n129_));
  NO2        g107(.A(i_6_), .B(i_5_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(i_3_), .Y(new_new_n131_));
  AO210      g109(.A0(new_new_n131_), .A1(new_new_n47_), .B0(new_new_n129_), .Y(new_new_n132_));
  OAI220     g110(.A0(new_new_n132_), .A1(new_new_n107_), .B0(new_new_n128_), .B1(new_new_n120_), .Y(new_new_n133_));
  NO3        g111(.A(new_new_n133_), .B(new_new_n118_), .C(new_new_n94_), .Y(new_new_n134_));
  NA3        g112(.A(new_new_n134_), .B(new_new_n78_), .C(new_new_n56_), .Y(ori2));
  NO2        g113(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n646_), .B(new_new_n136_), .Y(new_new_n137_));
  NA4        g115(.A(new_new_n137_), .B(new_new_n76_), .C(new_new_n68_), .D(new_new_n30_), .Y(ori0));
  AN2        g116(.A(i_8_), .B(i_7_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(i_6_), .Y(new_new_n140_));
  NO2        g118(.A(i_12_), .B(i_13_), .Y(new_new_n141_));
  NAi21      g119(.An(i_5_), .B(i_11_), .Y(new_new_n142_));
  NO2        g120(.A(i_0_), .B(i_1_), .Y(new_new_n143_));
  NA2        g121(.A(i_2_), .B(i_3_), .Y(new_new_n144_));
  NO2        g122(.A(new_new_n144_), .B(i_4_), .Y(new_new_n145_));
  AN2        g123(.A(new_new_n141_), .B(new_new_n82_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  OR2        g125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NO3        g126(.A(new_new_n148_), .B(new_new_n79_), .C(i_13_), .Y(new_new_n149_));
  NAi32      g127(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n150_));
  NAi21      g128(.An(new_new_n150_), .B(new_new_n149_), .Y(new_new_n151_));
  NOi21      g129(.An(i_4_), .B(i_10_), .Y(new_new_n152_));
  NA2        g130(.A(new_new_n152_), .B(new_new_n40_), .Y(new_new_n153_));
  NOi21      g131(.An(i_4_), .B(i_9_), .Y(new_new_n154_));
  NOi21      g132(.An(i_11_), .B(i_13_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n72_), .B(new_new_n62_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n72_), .B(i_5_), .Y(new_new_n158_));
  NO2        g136(.A(i_2_), .B(i_1_), .Y(new_new_n159_));
  NAi21      g137(.An(i_4_), .B(i_12_), .Y(new_new_n160_));
  INV        g138(.A(i_8_), .Y(new_new_n161_));
  NO2        g139(.A(i_3_), .B(i_8_), .Y(new_new_n162_));
  NO3        g140(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n102_), .B(new_new_n57_), .Y(new_new_n164_));
  NO2        g142(.A(i_13_), .B(i_9_), .Y(new_new_n165_));
  NAi21      g143(.An(i_12_), .B(i_3_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n44_), .B(i_5_), .Y(new_new_n167_));
  NAi21      g145(.An(i_12_), .B(i_7_), .Y(new_new_n168_));
  NA3        g146(.A(i_13_), .B(new_new_n161_), .C(i_10_), .Y(new_new_n169_));
  NA2        g147(.A(i_0_), .B(i_5_), .Y(new_new_n170_));
  NAi31      g148(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n171_));
  INV        g149(.A(i_13_), .Y(new_new_n172_));
  NO2        g150(.A(i_12_), .B(new_new_n172_), .Y(new_new_n173_));
  NO2        g151(.A(i_12_), .B(new_new_n37_), .Y(new_new_n174_));
  OR2        g152(.A(i_8_), .B(i_7_), .Y(new_new_n175_));
  INV        g153(.A(i_12_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n44_), .B(new_new_n176_), .Y(new_new_n177_));
  NO3        g155(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n178_));
  NA2        g156(.A(i_2_), .B(i_1_), .Y(new_new_n179_));
  NO3        g157(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n180_));
  NAi21      g158(.An(i_4_), .B(i_3_), .Y(new_new_n181_));
  NO2        g159(.A(i_0_), .B(i_6_), .Y(new_new_n182_));
  NOi41      g160(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n183_));
  NO2        g161(.A(i_11_), .B(new_new_n172_), .Y(new_new_n184_));
  NOi21      g162(.An(i_1_), .B(i_6_), .Y(new_new_n185_));
  NAi21      g163(.An(i_3_), .B(i_7_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n176_), .B(i_9_), .Y(new_new_n187_));
  OR4        g165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n185_), .D(new_new_n158_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n72_), .B(i_5_), .Y(new_new_n189_));
  NA2        g167(.A(i_3_), .B(i_9_), .Y(new_new_n190_));
  NAi21      g168(.An(i_7_), .B(i_10_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n191_), .B(new_new_n190_), .Y(new_new_n192_));
  NA3        g170(.A(new_new_n192_), .B(new_new_n189_), .C(new_new_n63_), .Y(new_new_n193_));
  NA2        g171(.A(new_new_n193_), .B(new_new_n188_), .Y(new_new_n194_));
  INV        g172(.A(new_new_n140_), .Y(new_new_n195_));
  NA2        g173(.A(new_new_n176_), .B(i_13_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n196_), .B(new_new_n74_), .Y(new_new_n197_));
  AOI220     g175(.A0(new_new_n197_), .A1(new_new_n195_), .B0(new_new_n194_), .B1(new_new_n184_), .Y(new_new_n198_));
  NA2        g176(.A(i_12_), .B(i_6_), .Y(new_new_n199_));
  OR2        g177(.A(i_13_), .B(i_9_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n181_), .B(i_2_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n184_), .B(i_9_), .Y(new_new_n202_));
  NO3        g180(.A(i_11_), .B(new_new_n172_), .C(new_new_n25_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n186_), .B(i_8_), .Y(new_new_n204_));
  NO3        g182(.A(i_12_), .B(new_new_n172_), .C(new_new_n37_), .Y(new_new_n205_));
  NO2        g183(.A(i_2_), .B(new_new_n100_), .Y(new_new_n206_));
  AN2        g184(.A(i_3_), .B(i_10_), .Y(new_new_n207_));
  NO2        g185(.A(i_5_), .B(new_new_n37_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n209_));
  NO3        g187(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n210_));
  NO2        g188(.A(i_2_), .B(i_3_), .Y(new_new_n211_));
  OR2        g189(.A(i_0_), .B(i_5_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(i_10_), .Y(new_new_n213_));
  NOi21      g191(.An(i_5_), .B(i_0_), .Y(new_new_n214_));
  NO2        g192(.A(i_1_), .B(i_7_), .Y(new_new_n215_));
  NOi21      g193(.An(new_new_n147_), .B(new_new_n103_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n216_), .B(new_new_n122_), .Y(new_new_n217_));
  NA2        g195(.A(new_new_n217_), .B(i_3_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n161_), .B(i_9_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n219_), .B(new_new_n164_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n220_), .B(new_new_n46_), .Y(new_new_n221_));
  INV        g199(.A(new_new_n221_), .Y(new_new_n222_));
  AOI210     g200(.A0(new_new_n222_), .A1(new_new_n218_), .B0(new_new_n153_), .Y(new_new_n223_));
  INV        g201(.A(new_new_n223_), .Y(new_new_n224_));
  NOi32      g202(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n225_));
  INV        g203(.A(new_new_n225_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n150_), .B(new_new_n148_), .Y(new_new_n227_));
  NOi32      g205(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n228_));
  NAi21      g206(.An(i_6_), .B(i_1_), .Y(new_new_n229_));
  NO2        g207(.A(i_1_), .B(new_new_n100_), .Y(new_new_n230_));
  NAi21      g208(.An(i_3_), .B(i_4_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n231_), .B(i_9_), .Y(new_new_n232_));
  AN2        g210(.A(i_6_), .B(i_7_), .Y(new_new_n233_));
  OAI210     g211(.A0(new_new_n233_), .A1(new_new_n230_), .B0(new_new_n232_), .Y(new_new_n234_));
  NA2        g212(.A(i_2_), .B(i_7_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n231_), .B(i_10_), .Y(new_new_n236_));
  NA3        g214(.A(new_new_n236_), .B(new_new_n235_), .C(new_new_n182_), .Y(new_new_n237_));
  AOI210     g215(.A0(new_new_n237_), .A1(new_new_n234_), .B0(new_new_n158_), .Y(new_new_n238_));
  AOI210     g216(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n239_));
  OAI210     g217(.A0(new_new_n239_), .A1(new_new_n159_), .B0(new_new_n236_), .Y(new_new_n240_));
  AOI220     g218(.A0(new_new_n236_), .A1(new_new_n215_), .B0(new_new_n178_), .B1(new_new_n159_), .Y(new_new_n241_));
  AOI210     g219(.A0(new_new_n241_), .A1(new_new_n240_), .B0(i_5_), .Y(new_new_n242_));
  NO3        g220(.A(new_new_n242_), .B(new_new_n238_), .C(new_new_n227_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n243_), .B(new_new_n226_), .Y(new_new_n244_));
  AN2        g222(.A(i_12_), .B(i_5_), .Y(new_new_n245_));
  NO2        g223(.A(i_11_), .B(i_6_), .Y(new_new_n246_));
  NO2        g224(.A(i_5_), .B(i_10_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n248_));
  NO3        g226(.A(new_new_n85_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n249_));
  NO2        g227(.A(i_11_), .B(i_12_), .Y(new_new_n250_));
  NAi21      g228(.An(i_13_), .B(i_0_), .Y(new_new_n251_));
  NO3        g229(.A(i_1_), .B(i_12_), .C(new_new_n85_), .Y(new_new_n252_));
  NO2        g230(.A(i_0_), .B(i_11_), .Y(new_new_n253_));
  AN2        g231(.A(i_1_), .B(i_6_), .Y(new_new_n254_));
  NOi21      g232(.An(i_2_), .B(i_12_), .Y(new_new_n255_));
  NAi21      g233(.An(i_9_), .B(i_4_), .Y(new_new_n256_));
  OR2        g234(.A(i_13_), .B(i_10_), .Y(new_new_n257_));
  NO3        g235(.A(new_new_n257_), .B(new_new_n115_), .C(new_new_n256_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n156_), .B(new_new_n121_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n100_), .B(new_new_n25_), .Y(new_new_n260_));
  NA2        g238(.A(new_new_n205_), .B(new_new_n260_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n261_), .B(new_new_n216_), .Y(new_new_n262_));
  INV        g240(.A(new_new_n262_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n263_), .B(new_new_n26_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n161_), .B(i_10_), .Y(new_new_n265_));
  NA3        g243(.A(new_new_n189_), .B(new_new_n63_), .C(i_2_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n266_), .B(new_new_n265_), .Y(new_new_n267_));
  INV        g245(.A(new_new_n267_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n268_), .B(new_new_n202_), .Y(new_new_n269_));
  NO3        g247(.A(new_new_n269_), .B(new_new_n264_), .C(new_new_n244_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n72_), .B(i_13_), .Y(new_new_n271_));
  NO2        g249(.A(i_10_), .B(i_9_), .Y(new_new_n272_));
  NAi21      g250(.An(i_12_), .B(i_8_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(i_3_), .Y(new_new_n274_));
  NO3        g252(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n199_), .B(new_new_n96_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n276_), .B(new_new_n275_), .Y(new_new_n277_));
  NA2        g255(.A(i_8_), .B(i_9_), .Y(new_new_n278_));
  AOI210     g256(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n279_));
  OR2        g257(.A(new_new_n279_), .B(new_new_n278_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n205_), .B(new_new_n164_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n281_), .B(new_new_n280_), .Y(new_new_n282_));
  NA2        g260(.A(new_new_n184_), .B(new_new_n208_), .Y(new_new_n283_));
  NO3        g261(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n284_));
  INV        g262(.A(new_new_n284_), .Y(new_new_n285_));
  NA3        g263(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n286_));
  NA4        g264(.A(new_new_n142_), .B(new_new_n114_), .C(new_new_n79_), .D(new_new_n23_), .Y(new_new_n287_));
  OAI220     g265(.A0(new_new_n287_), .A1(new_new_n286_), .B0(new_new_n285_), .B1(new_new_n283_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n288_), .B(new_new_n282_), .Y(new_new_n289_));
  NA2        g267(.A(new_new_n95_), .B(i_13_), .Y(new_new_n290_));
  NO2        g268(.A(i_11_), .B(i_1_), .Y(new_new_n291_));
  NOi21      g269(.An(i_2_), .B(i_7_), .Y(new_new_n292_));
  NO2        g270(.A(i_6_), .B(i_10_), .Y(new_new_n293_));
  NA3        g271(.A(new_new_n183_), .B(new_new_n155_), .C(new_new_n130_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n148_), .B(i_3_), .Y(new_new_n296_));
  NAi31      g274(.An(new_new_n295_), .B(new_new_n296_), .C(new_new_n173_), .Y(new_new_n297_));
  NA3        g275(.A(new_new_n248_), .B(new_new_n157_), .C(new_new_n145_), .Y(new_new_n298_));
  NA3        g276(.A(new_new_n298_), .B(new_new_n297_), .C(new_new_n294_), .Y(new_new_n299_));
  INV        g277(.A(new_new_n299_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n275_), .B(new_new_n245_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n284_), .B(new_new_n247_), .Y(new_new_n302_));
  NAi21      g280(.An(new_new_n169_), .B(new_new_n250_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n27_), .B(i_10_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n210_), .B(new_new_n178_), .Y(new_new_n305_));
  OAI220     g283(.A0(new_new_n305_), .A1(new_new_n266_), .B0(new_new_n304_), .B1(new_new_n290_), .Y(new_new_n306_));
  INV        g284(.A(new_new_n306_), .Y(new_new_n307_));
  NA3        g285(.A(new_new_n307_), .B(new_new_n300_), .C(new_new_n289_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n245_), .B(new_new_n172_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n233_), .B(new_new_n228_), .Y(new_new_n310_));
  OR2        g288(.A(new_new_n309_), .B(new_new_n310_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n36_), .B(i_8_), .Y(new_new_n312_));
  AOI210     g290(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n258_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n313_), .B(new_new_n311_), .Y(new_new_n314_));
  INV        g292(.A(new_new_n314_), .Y(new_new_n315_));
  INV        g293(.A(new_new_n132_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n259_), .Y(new_new_n317_));
  NA2        g295(.A(new_new_n317_), .B(new_new_n315_), .Y(new_new_n318_));
  NO2        g296(.A(i_12_), .B(new_new_n161_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n44_), .B(i_10_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(i_6_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n148_), .B(i_5_), .Y(new_new_n322_));
  NA3        g300(.A(new_new_n170_), .B(new_new_n70_), .C(new_new_n44_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n205_), .B(new_new_n83_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n323_), .B(new_new_n324_), .Y(new_new_n325_));
  AOI210     g303(.A0(new_new_n229_), .A1(new_new_n46_), .B0(new_new_n230_), .Y(new_new_n326_));
  NA2        g304(.A(i_0_), .B(new_new_n48_), .Y(new_new_n327_));
  NA3        g305(.A(new_new_n319_), .B(new_new_n203_), .C(new_new_n327_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n326_), .B(new_new_n328_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n329_), .B(new_new_n325_), .Y(new_new_n330_));
  NO3        g308(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n257_), .B(i_1_), .Y(new_new_n332_));
  NOi31      g310(.An(new_new_n332_), .B(new_new_n276_), .C(new_new_n72_), .Y(new_new_n333_));
  NOi21      g311(.An(i_10_), .B(i_6_), .Y(new_new_n334_));
  NO2        g312(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n113_), .B(new_new_n23_), .Y(new_new_n336_));
  NO2        g314(.A(i_12_), .B(new_new_n85_), .Y(new_new_n337_));
  OR2        g315(.A(i_2_), .B(i_5_), .Y(new_new_n338_));
  OR2        g316(.A(new_new_n338_), .B(new_new_n254_), .Y(new_new_n339_));
  NA2        g317(.A(new_new_n235_), .B(new_new_n182_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n340_), .A1(new_new_n339_), .B0(new_new_n303_), .Y(new_new_n341_));
  INV        g319(.A(new_new_n341_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n330_), .Y(new_new_n343_));
  NO3        g321(.A(new_new_n343_), .B(new_new_n318_), .C(new_new_n308_), .Y(new_new_n344_));
  NA4        g322(.A(new_new_n344_), .B(new_new_n270_), .C(new_new_n224_), .D(new_new_n198_), .Y(ori7));
  NO2        g323(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n293_), .B(new_new_n83_), .Y(new_new_n347_));
  NA2        g325(.A(i_11_), .B(new_new_n161_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n141_), .B(new_new_n348_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(new_new_n347_), .Y(new_new_n350_));
  NA3        g328(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n176_), .B(i_4_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n352_), .B(i_8_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n104_), .B(new_new_n351_), .Y(new_new_n354_));
  NA2        g332(.A(i_2_), .B(new_new_n85_), .Y(new_new_n355_));
  OAI210     g333(.A0(new_new_n86_), .A1(new_new_n162_), .B0(new_new_n163_), .Y(new_new_n356_));
  NO2        g334(.A(i_7_), .B(new_new_n37_), .Y(new_new_n357_));
  NA2        g335(.A(i_4_), .B(i_8_), .Y(new_new_n358_));
  AOI210     g336(.A0(new_new_n358_), .A1(new_new_n207_), .B0(new_new_n357_), .Y(new_new_n359_));
  OAI220     g337(.A0(new_new_n359_), .A1(new_new_n355_), .B0(new_new_n356_), .B1(i_13_), .Y(new_new_n360_));
  NO4        g338(.A(new_new_n360_), .B(new_new_n354_), .C(new_new_n350_), .D(new_new_n346_), .Y(new_new_n361_));
  AOI210     g339(.A0(new_new_n126_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n362_));
  AOI210     g340(.A0(new_new_n362_), .A1(new_new_n176_), .B0(new_new_n152_), .Y(new_new_n363_));
  OR2        g341(.A(i_6_), .B(i_10_), .Y(new_new_n364_));
  OR3        g342(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n365_));
  OR2        g343(.A(new_new_n363_), .B(new_new_n200_), .Y(new_new_n366_));
  AOI210     g344(.A0(new_new_n366_), .A1(new_new_n361_), .B0(new_new_n62_), .Y(new_new_n367_));
  NOi21      g345(.An(i_11_), .B(i_7_), .Y(new_new_n368_));
  AO210      g346(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n370_), .B(new_new_n165_), .Y(new_new_n371_));
  NA3        g349(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n372_));
  NO2        g350(.A(new_new_n371_), .B(new_new_n62_), .Y(new_new_n373_));
  OR2        g351(.A(new_new_n241_), .B(new_new_n41_), .Y(new_new_n374_));
  NA2        g352(.A(new_new_n173_), .B(new_new_n62_), .Y(new_new_n375_));
  OR2        g353(.A(new_new_n166_), .B(new_new_n107_), .Y(new_new_n376_));
  NO2        g354(.A(i_1_), .B(i_12_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n375_), .B(new_new_n374_), .Y(new_new_n378_));
  OAI210     g356(.A0(new_new_n378_), .A1(new_new_n373_), .B0(i_6_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n372_), .B(new_new_n107_), .Y(new_new_n380_));
  NA2        g358(.A(new_new_n380_), .B(new_new_n337_), .Y(new_new_n381_));
  NO2        g359(.A(i_6_), .B(i_11_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n381_), .B(new_new_n277_), .Y(new_new_n383_));
  NO3        g361(.A(new_new_n364_), .B(new_new_n175_), .C(new_new_n23_), .Y(new_new_n384_));
  AOI210     g362(.A0(i_1_), .A1(new_new_n192_), .B0(new_new_n384_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n385_), .B(new_new_n44_), .Y(new_new_n386_));
  INV        g364(.A(i_2_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n136_), .B(i_9_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n46_), .B(i_1_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n388_), .B(new_new_n387_), .Y(new_new_n390_));
  AOI210     g368(.A0(new_new_n291_), .A1(new_new_n260_), .B0(new_new_n180_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n391_), .B(new_new_n355_), .Y(new_new_n392_));
  NO2        g370(.A(i_11_), .B(new_new_n37_), .Y(new_new_n393_));
  OR2        g371(.A(new_new_n392_), .B(new_new_n390_), .Y(new_new_n394_));
  NO3        g372(.A(new_new_n394_), .B(new_new_n386_), .C(new_new_n383_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n176_), .B(new_new_n100_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n396_), .B(new_new_n368_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n397_), .B(i_1_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n365_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n256_), .B(new_new_n85_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n399_), .B(new_new_n46_), .Y(new_new_n401_));
  NA2        g379(.A(i_3_), .B(new_new_n161_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(new_new_n113_), .Y(new_new_n403_));
  AN2        g381(.A(new_new_n403_), .B(new_new_n321_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n175_), .B(new_new_n44_), .Y(new_new_n405_));
  NO3        g383(.A(new_new_n405_), .B(new_new_n209_), .C(new_new_n177_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n115_), .B(new_new_n37_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n407_), .B(i_6_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n85_), .B(i_9_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n62_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n410_), .B(new_new_n377_), .Y(new_new_n411_));
  NO4        g389(.A(new_new_n411_), .B(new_new_n408_), .C(new_new_n406_), .D(i_4_), .Y(new_new_n412_));
  NA2        g390(.A(i_1_), .B(i_3_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n278_), .B(new_new_n92_), .Y(new_new_n414_));
  AOI210     g392(.A0(new_new_n405_), .A1(new_new_n334_), .B0(new_new_n414_), .Y(new_new_n415_));
  NO2        g393(.A(new_new_n415_), .B(new_new_n413_), .Y(new_new_n416_));
  NO3        g394(.A(new_new_n416_), .B(new_new_n412_), .C(new_new_n404_), .Y(new_new_n417_));
  NA4        g395(.A(new_new_n417_), .B(new_new_n401_), .C(new_new_n395_), .D(new_new_n379_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n419_));
  INV        g397(.A(new_new_n419_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n420_), .B(i_1_), .Y(new_new_n421_));
  AOI210     g399(.A0(new_new_n199_), .A1(new_new_n96_), .B0(i_1_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n231_), .B(i_2_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n423_), .B(new_new_n422_), .Y(new_new_n424_));
  AOI210     g402(.A0(new_new_n424_), .A1(new_new_n421_), .B0(i_13_), .Y(new_new_n425_));
  OR2        g403(.A(i_11_), .B(i_7_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n54_), .B(i_12_), .Y(new_new_n427_));
  NO2        g405(.A(new_new_n292_), .B(new_new_n24_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n428_), .B(new_new_n400_), .Y(new_new_n429_));
  OAI220     g407(.A0(new_new_n429_), .A1(new_new_n41_), .B0(new_new_n645_), .B1(new_new_n92_), .Y(new_new_n430_));
  INV        g408(.A(new_new_n430_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n246_), .B(new_new_n389_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n432_), .B(new_new_n181_), .Y(new_new_n433_));
  AOI210     g411(.A0(new_new_n273_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n434_));
  NOi31      g412(.An(new_new_n434_), .B(new_new_n347_), .C(new_new_n44_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n125_), .B(i_13_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n422_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n26_), .B(new_new_n161_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(i_7_), .Y(new_new_n439_));
  AOI220     g417(.A0(new_new_n246_), .A1(new_new_n389_), .B0(new_new_n91_), .B1(new_new_n101_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n440_), .B(new_new_n353_), .Y(new_new_n441_));
  NO4        g419(.A(new_new_n441_), .B(new_new_n437_), .C(new_new_n435_), .D(new_new_n433_), .Y(new_new_n442_));
  OR2        g420(.A(i_11_), .B(i_6_), .Y(new_new_n443_));
  NA3        g421(.A(new_new_n352_), .B(new_new_n438_), .C(i_7_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n444_), .B(new_new_n443_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n255_), .B(new_new_n357_), .C(new_new_n96_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n382_), .B(i_13_), .Y(new_new_n447_));
  NAi21      g425(.An(i_11_), .B(i_12_), .Y(new_new_n448_));
  NOi41      g426(.An(new_new_n109_), .B(new_new_n448_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n449_), .B(new_new_n46_), .Y(new_new_n450_));
  NA3        g428(.A(new_new_n450_), .B(new_new_n447_), .C(new_new_n446_), .Y(new_new_n451_));
  OAI210     g429(.A0(new_new_n451_), .A1(new_new_n445_), .B0(new_new_n62_), .Y(new_new_n452_));
  NO2        g430(.A(i_2_), .B(i_12_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n230_), .B(new_new_n453_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n232_), .B(new_new_n230_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n456_), .B(new_new_n45_), .C(new_new_n172_), .Y(new_new_n457_));
  NA4        g435(.A(new_new_n457_), .B(new_new_n452_), .C(new_new_n442_), .D(new_new_n431_), .Y(new_new_n458_));
  OR4        g436(.A(new_new_n458_), .B(new_new_n425_), .C(new_new_n418_), .D(new_new_n367_), .Y(ori5));
  NA2        g437(.A(new_new_n397_), .B(new_new_n201_), .Y(new_new_n460_));
  AN2        g438(.A(new_new_n24_), .B(i_10_), .Y(new_new_n461_));
  NA3        g439(.A(new_new_n461_), .B(new_new_n453_), .C(new_new_n107_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n353_), .B(i_11_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n86_), .B(new_new_n463_), .Y(new_new_n464_));
  NA3        g442(.A(new_new_n464_), .B(new_new_n462_), .C(new_new_n460_), .Y(new_new_n465_));
  NO3        g443(.A(i_11_), .B(new_new_n176_), .C(i_13_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n122_), .B(new_new_n23_), .Y(new_new_n467_));
  NA2        g445(.A(i_12_), .B(i_8_), .Y(new_new_n468_));
  OAI210     g446(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n468_), .Y(new_new_n469_));
  INV        g447(.A(new_new_n272_), .Y(new_new_n470_));
  AOI220     g448(.A0(new_new_n211_), .A1(new_new_n336_), .B0(new_new_n469_), .B1(new_new_n467_), .Y(new_new_n471_));
  INV        g449(.A(new_new_n471_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n465_), .Y(new_new_n473_));
  INV        g451(.A(new_new_n155_), .Y(new_new_n474_));
  INV        g452(.A(new_new_n183_), .Y(new_new_n475_));
  OAI210     g453(.A0(new_new_n423_), .A1(new_new_n274_), .B0(new_new_n109_), .Y(new_new_n476_));
  AOI210     g454(.A0(new_new_n476_), .A1(new_new_n475_), .B0(new_new_n474_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n278_), .B(new_new_n26_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n478_), .B(new_new_n260_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(i_2_), .Y(new_new_n480_));
  INV        g458(.A(new_new_n480_), .Y(new_new_n481_));
  AOI210     g459(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n257_), .Y(new_new_n482_));
  AOI210     g460(.A0(new_new_n482_), .A1(new_new_n481_), .B0(new_new_n477_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n160_), .B(new_new_n123_), .Y(new_new_n484_));
  OAI210     g462(.A0(new_new_n484_), .A1(new_new_n467_), .B0(i_2_), .Y(new_new_n485_));
  INV        g463(.A(new_new_n156_), .Y(new_new_n486_));
  NO3        g464(.A(new_new_n369_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n486_), .A1(new_new_n86_), .B0(new_new_n487_), .Y(new_new_n488_));
  AOI210     g466(.A0(new_new_n488_), .A1(new_new_n485_), .B0(new_new_n161_), .Y(new_new_n489_));
  OA210      g467(.A0(new_new_n370_), .A1(new_new_n124_), .B0(i_13_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n146_), .B(new_new_n348_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n491_), .B(new_new_n235_), .Y(new_new_n492_));
  AOI210     g470(.A0(new_new_n166_), .A1(new_new_n144_), .B0(new_new_n312_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n260_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n101_), .B(new_new_n44_), .Y(new_new_n495_));
  INV        g473(.A(new_new_n206_), .Y(new_new_n496_));
  NA4        g474(.A(new_new_n496_), .B(new_new_n207_), .C(new_new_n122_), .D(new_new_n42_), .Y(new_new_n497_));
  OAI210     g475(.A0(new_new_n497_), .A1(new_new_n495_), .B0(new_new_n494_), .Y(new_new_n498_));
  NO4        g476(.A(new_new_n498_), .B(new_new_n492_), .C(new_new_n490_), .D(new_new_n489_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n336_), .B(new_new_n28_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n466_), .B(new_new_n204_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n501_), .B(new_new_n500_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n61_), .B(i_12_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(new_new_n124_), .Y(new_new_n504_));
  NO2        g482(.A(new_new_n504_), .B(new_new_n348_), .Y(new_new_n505_));
  AOI220     g483(.A0(new_new_n505_), .A1(new_new_n36_), .B0(new_new_n502_), .B1(new_new_n46_), .Y(new_new_n506_));
  NA4        g484(.A(new_new_n506_), .B(new_new_n499_), .C(new_new_n483_), .D(new_new_n473_), .Y(ori6));
  NO2        g485(.A(new_new_n171_), .B(new_new_n295_), .Y(new_new_n508_));
  OR2        g486(.A(new_new_n647_), .B(i_12_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n337_), .B(new_new_n62_), .Y(new_new_n510_));
  INV        g488(.A(new_new_n510_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n72_), .Y(new_new_n512_));
  INV        g490(.A(new_new_n213_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n74_), .B(new_new_n129_), .Y(new_new_n514_));
  INV        g492(.A(new_new_n122_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n515_), .B(new_new_n46_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n516_), .A1(new_new_n514_), .B0(new_new_n513_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n185_), .B(i_9_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n518_), .B(new_new_n503_), .Y(new_new_n519_));
  AOI210     g497(.A0(new_new_n519_), .A1(new_new_n310_), .B0(new_new_n158_), .Y(new_new_n520_));
  NAi32      g498(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n443_), .B(new_new_n521_), .Y(new_new_n522_));
  OR3        g500(.A(new_new_n522_), .B(new_new_n520_), .C(new_new_n517_), .Y(new_new_n523_));
  NO2        g501(.A(new_new_n426_), .B(i_2_), .Y(new_new_n524_));
  BUFFER     g502(.A(new_new_n370_), .Y(new_new_n525_));
  NA3        g503(.A(new_new_n525_), .B(new_new_n143_), .C(new_new_n68_), .Y(new_new_n526_));
  AO210      g504(.A0(new_new_n302_), .A1(new_new_n470_), .B0(new_new_n36_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n527_), .B(new_new_n526_), .Y(new_new_n528_));
  NO2        g506(.A(i_6_), .B(i_11_), .Y(new_new_n529_));
  AOI220     g507(.A0(new_new_n529_), .A1(new_new_n331_), .B0(new_new_n508_), .B1(new_new_n439_), .Y(new_new_n530_));
  NA3        g508(.A(new_new_n235_), .B(new_new_n178_), .C(new_new_n143_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n249_), .B(new_new_n69_), .Y(new_new_n532_));
  NA4        g510(.A(new_new_n532_), .B(new_new_n531_), .C(new_new_n530_), .D(new_new_n356_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n274_), .B(new_new_n272_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n364_), .B(new_new_n101_), .Y(new_new_n535_));
  OAI210     g513(.A0(new_new_n535_), .A1(new_new_n110_), .B0(new_new_n253_), .Y(new_new_n536_));
  INV        g514(.A(new_new_n339_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n537_), .B(new_new_n213_), .C(i_7_), .Y(new_new_n538_));
  NA3        g516(.A(new_new_n538_), .B(new_new_n536_), .C(new_new_n534_), .Y(new_new_n539_));
  NO4        g517(.A(new_new_n539_), .B(new_new_n533_), .C(new_new_n528_), .D(new_new_n523_), .Y(new_new_n540_));
  NA4        g518(.A(new_new_n540_), .B(new_new_n512_), .C(new_new_n509_), .D(new_new_n243_), .Y(ori3));
  NA2        g519(.A(i_12_), .B(i_10_), .Y(new_new_n542_));
  NO2        g520(.A(i_11_), .B(new_new_n176_), .Y(new_new_n543_));
  NA3        g521(.A(new_new_n531_), .B(new_new_n356_), .C(new_new_n234_), .Y(new_new_n544_));
  NA2        g522(.A(new_new_n544_), .B(new_new_n40_), .Y(new_new_n545_));
  NOi21      g523(.An(new_new_n95_), .B(new_new_n479_), .Y(new_new_n546_));
  NO3        g524(.A(new_new_n376_), .B(new_new_n278_), .C(new_new_n129_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n255_), .B(new_new_n45_), .Y(new_new_n548_));
  AN2        g526(.A(new_new_n276_), .B(new_new_n55_), .Y(new_new_n549_));
  NO3        g527(.A(new_new_n549_), .B(new_new_n547_), .C(new_new_n546_), .Y(new_new_n550_));
  AOI210     g528(.A0(new_new_n550_), .A1(new_new_n545_), .B0(new_new_n48_), .Y(new_new_n551_));
  NO4        g529(.A(new_new_n239_), .B(new_new_n245_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n552_));
  NA2        g530(.A(new_new_n158_), .B(new_new_n334_), .Y(new_new_n553_));
  NOi21      g531(.An(new_new_n553_), .B(new_new_n552_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n554_), .B(new_new_n62_), .Y(new_new_n555_));
  NOi21      g533(.An(i_5_), .B(i_9_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n556_), .B(new_new_n271_), .Y(new_new_n557_));
  BUFFER     g535(.A(new_new_n199_), .Y(new_new_n558_));
  NA2        g536(.A(new_new_n558_), .B(new_new_n291_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n559_), .B(new_new_n557_), .Y(new_new_n560_));
  NO3        g538(.A(new_new_n560_), .B(new_new_n555_), .C(new_new_n551_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n335_), .B(i_0_), .Y(new_new_n562_));
  NO4        g540(.A(new_new_n338_), .B(new_new_n168_), .C(new_new_n257_), .D(new_new_n254_), .Y(new_new_n563_));
  NA2        g541(.A(new_new_n563_), .B(i_11_), .Y(new_new_n564_));
  NA2        g542(.A(new_new_n466_), .B(new_new_n214_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n293_), .A1(new_new_n86_), .B0(new_new_n57_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n566_), .B(new_new_n565_), .Y(new_new_n567_));
  NO2        g545(.A(new_new_n187_), .B(new_new_n147_), .Y(new_new_n568_));
  NA2        g546(.A(i_0_), .B(i_10_), .Y(new_new_n569_));
  INV        g547(.A(new_new_n320_), .Y(new_new_n570_));
  NO4        g548(.A(new_new_n113_), .B(new_new_n57_), .C(new_new_n402_), .D(i_5_), .Y(new_new_n571_));
  AO220      g549(.A0(new_new_n571_), .A1(new_new_n570_), .B0(new_new_n568_), .B1(i_6_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n572_), .B(new_new_n567_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n573_), .B(new_new_n564_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n575_));
  NA2        g553(.A(i_11_), .B(i_9_), .Y(new_new_n576_));
  NO3        g554(.A(i_12_), .B(new_new_n576_), .C(new_new_n355_), .Y(new_new_n577_));
  AN2        g555(.A(new_new_n577_), .B(new_new_n575_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n248_), .B(new_new_n157_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n579_), .B(new_new_n151_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n576_), .B(new_new_n72_), .Y(new_new_n581_));
  INV        g559(.A(new_new_n252_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n582_), .B(new_new_n557_), .Y(new_new_n583_));
  NO3        g561(.A(new_new_n583_), .B(new_new_n580_), .C(new_new_n578_), .Y(new_new_n584_));
  NA2        g562(.A(new_new_n393_), .B(new_new_n119_), .Y(new_new_n585_));
  NO2        g563(.A(i_6_), .B(new_new_n585_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n155_), .B(new_new_n102_), .Y(new_new_n587_));
  INV        g565(.A(new_new_n586_), .Y(new_new_n588_));
  INV        g566(.A(new_new_n212_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n588_), .B(new_new_n584_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n542_), .B(new_new_n211_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n581_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n428_), .B(new_new_n322_), .Y(new_new_n593_));
  NAi21      g571(.An(i_9_), .B(i_5_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n594_), .B(new_new_n251_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n595_), .B(new_new_n370_), .Y(new_new_n596_));
  OAI220     g574(.A0(new_new_n596_), .A1(new_new_n85_), .B0(new_new_n593_), .B1(new_new_n156_), .Y(new_new_n597_));
  NO2        g575(.A(new_new_n597_), .B(new_new_n314_), .Y(new_new_n598_));
  NA2        g576(.A(new_new_n598_), .B(new_new_n592_), .Y(new_new_n599_));
  NO3        g577(.A(new_new_n599_), .B(new_new_n590_), .C(new_new_n574_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n510_), .A1(new_new_n419_), .B0(new_new_n587_), .Y(new_new_n601_));
  INV        g579(.A(new_new_n601_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n182_), .B(new_new_n174_), .Y(new_new_n603_));
  AOI210     g581(.A0(new_new_n603_), .A1(new_new_n562_), .B0(new_new_n147_), .Y(new_new_n604_));
  INV        g582(.A(new_new_n604_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n605_), .B(new_new_n602_), .Y(new_new_n606_));
  NO3        g584(.A(new_new_n569_), .B(new_new_n556_), .C(new_new_n160_), .Y(new_new_n607_));
  AOI220     g585(.A0(new_new_n607_), .A1(i_11_), .B0(new_new_n333_), .B1(new_new_n74_), .Y(new_new_n608_));
  NO3        g586(.A(new_new_n167_), .B(new_new_n245_), .C(i_0_), .Y(new_new_n609_));
  OAI210     g587(.A0(new_new_n609_), .A1(new_new_n75_), .B0(i_13_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(new_new_n608_), .Y(new_new_n611_));
  NO3        g589(.A(new_new_n548_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n612_));
  NA2        g590(.A(new_new_n301_), .B(new_new_n294_), .Y(new_new_n613_));
  NO2        g591(.A(new_new_n613_), .B(new_new_n612_), .Y(new_new_n614_));
  NA3        g592(.A(new_new_n247_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n615_));
  INV        g593(.A(new_new_n615_), .Y(new_new_n616_));
  NO3        g594(.A(new_new_n576_), .B(new_new_n170_), .C(new_new_n160_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n617_), .B(new_new_n616_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n618_), .B(new_new_n614_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n85_), .B(i_5_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n543_), .B(new_new_n108_), .C(new_new_n122_), .Y(new_new_n621_));
  INV        g599(.A(new_new_n621_), .Y(new_new_n622_));
  NA2        g600(.A(new_new_n622_), .B(new_new_n620_), .Y(new_new_n623_));
  NAi21      g601(.An(new_new_n180_), .B(new_new_n181_), .Y(new_new_n624_));
  NO4        g602(.A(new_new_n179_), .B(new_new_n167_), .C(i_0_), .D(i_12_), .Y(new_new_n625_));
  NA2        g603(.A(new_new_n625_), .B(new_new_n624_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n626_), .B(new_new_n623_), .Y(new_new_n627_));
  NO4        g605(.A(new_new_n627_), .B(new_new_n619_), .C(new_new_n611_), .D(new_new_n606_), .Y(new_new_n628_));
  NA2        g606(.A(new_new_n524_), .B(new_new_n37_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n629_), .B(new_new_n363_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n630_), .B(new_new_n165_), .Y(new_new_n631_));
  NAi31      g609(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n69_), .B(new_new_n632_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n633_), .A1(new_new_n48_), .B0(new_new_n563_), .Y(new_new_n634_));
  AOI210     g612(.A0(new_new_n634_), .A1(new_new_n631_), .B0(new_new_n72_), .Y(new_new_n635_));
  INV        g613(.A(new_new_n242_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n636_), .B(new_new_n474_), .Y(new_new_n637_));
  NO3        g615(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n638_));
  OAI210     g616(.A0(new_new_n589_), .A1(new_new_n208_), .B0(new_new_n638_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n639_), .B(new_new_n448_), .Y(new_new_n640_));
  NO3        g618(.A(new_new_n640_), .B(new_new_n637_), .C(new_new_n635_), .Y(new_new_n641_));
  NA4        g619(.A(new_new_n641_), .B(new_new_n628_), .C(new_new_n600_), .D(new_new_n561_), .Y(ori4));
  INV        g620(.A(new_new_n427_), .Y(new_new_n645_));
  INV        g621(.A(i_6_), .Y(new_new_n646_));
  INV        g622(.A(new_new_n214_), .Y(new_new_n647_));
endmodule


