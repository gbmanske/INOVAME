// Benchmark "top" written by ABC on Thu Jun 20 14:59:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n781_,
    new_new_n782_, new_new_n783_, new_new_n784_, new_new_n785_,
    new_new_n786_, new_new_n787_, new_new_n788_, new_new_n789_,
    new_new_n790_, new_new_n791_, new_new_n792_, new_new_n793_,
    new_new_n794_, new_new_n795_, new_new_n796_, new_new_n797_,
    new_new_n798_, new_new_n799_, new_new_n800_, new_new_n801_,
    new_new_n802_, new_new_n803_, new_new_n804_, new_new_n805_,
    new_new_n806_, new_new_n807_, new_new_n808_, new_new_n809_,
    new_new_n810_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n827_, new_new_n828_, new_new_n829_, new_new_n830_,
    new_new_n831_, new_new_n832_, new_new_n833_, new_new_n834_,
    new_new_n835_, new_new_n836_, new_new_n837_, new_new_n838_,
    new_new_n839_, new_new_n840_, new_new_n841_, new_new_n842_,
    new_new_n843_, new_new_n844_, new_new_n845_, new_new_n846_,
    new_new_n847_, new_new_n848_, new_new_n849_, new_new_n850_,
    new_new_n851_, new_new_n852_, new_new_n853_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n881_, new_new_n882_, new_new_n883_,
    new_new_n884_, new_new_n885_, new_new_n886_, new_new_n887_,
    new_new_n888_, new_new_n889_, new_new_n890_, new_new_n891_,
    new_new_n892_, new_new_n893_, new_new_n894_, new_new_n895_,
    new_new_n896_, new_new_n897_, new_new_n898_, new_new_n899_,
    new_new_n900_, new_new_n901_, new_new_n902_, new_new_n903_,
    new_new_n904_, new_new_n905_, new_new_n906_, new_new_n907_,
    new_new_n908_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1107_, new_new_n1108_,
    new_new_n1109_, new_new_n1110_, new_new_n1111_, new_new_n1112_,
    new_new_n1113_, new_new_n1114_, new_new_n1115_, new_new_n1116_,
    new_new_n1117_, new_new_n1118_, new_new_n1119_, new_new_n1120_,
    new_new_n1121_, new_new_n1122_, new_new_n1123_, new_new_n1124_,
    new_new_n1125_, new_new_n1126_, new_new_n1127_, new_new_n1128_,
    new_new_n1129_, new_new_n1130_, new_new_n1131_, new_new_n1132_,
    new_new_n1133_, new_new_n1134_, new_new_n1135_, new_new_n1136_,
    new_new_n1137_, new_new_n1138_, new_new_n1139_, new_new_n1140_,
    new_new_n1141_, new_new_n1142_, new_new_n1146_, new_new_n1147_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NO2        g0028(.A(new_new_n50_), .B(i_3_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  OR4        g0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g0066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  OAI210     g0067(.A0(new_new_n85_), .A1(new_new_n82_), .B0(i_2_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_10_), .Y(new_new_n91_));
  NA2        g0069(.A(i_6_), .B(i_9_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n91_), .B0(new_new_n63_), .Y(new_new_n93_));
  NA2        g0071(.A(i_2_), .B(i_6_), .Y(new_new_n94_));
  NO3        g0072(.A(new_new_n94_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n95_));
  NO2        g0073(.A(new_new_n95_), .B(new_new_n93_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n90_), .B0(new_new_n80_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n101_), .B(new_new_n62_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n46_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n86_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  NO3        g0088(.A(new_new_n110_), .B(new_new_n91_), .C(new_new_n53_), .Y(new_new_n111_));
  AN2        g0089(.A(i_2_), .B(i_10_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n112_), .B(i_7_), .Y(new_new_n113_));
  OR2        g0091(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n114_));
  NO2        g0092(.A(i_8_), .B(new_new_n103_), .Y(new_new_n115_));
  NO3        g0093(.A(new_new_n115_), .B(new_new_n114_), .C(new_new_n113_), .Y(new_new_n116_));
  NA2        g0094(.A(i_12_), .B(i_7_), .Y(new_new_n117_));
  NO2        g0095(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n118_));
  INV        g0096(.A(new_new_n118_), .Y(new_new_n119_));
  NA2        g0097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  OAI210     g0098(.A0(new_new_n119_), .A1(new_new_n117_), .B0(new_new_n120_), .Y(new_new_n121_));
  NO2        g0099(.A(new_new_n121_), .B(new_new_n116_), .Y(new_new_n122_));
  NA3        g0100(.A(new_new_n122_), .B(new_new_n109_), .C(new_new_n102_), .Y(new_new_n123_));
  NOi21      g0101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g0104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g0106(.A(new_new_n128_), .B(new_new_n46_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n92_), .B(new_new_n91_), .Y(new_new_n130_));
  NAi21      g0108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(new_new_n62_), .Y(new_new_n132_));
  NOi31      g0110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g0111(.A(i_1_), .B(new_new_n86_), .Y(new_new_n134_));
  NO2        g0112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g0113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g0114(.A0(new_new_n136_), .A1(new_new_n47_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g0115(.A0(new_new_n137_), .A1(new_new_n110_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g0116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n97_), .Y(new_new_n139_));
  NA3        g0117(.A(new_new_n139_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0118(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g0119(.A(i_6_), .B(new_new_n25_), .Y(new_new_n142_));
  NA3        g0120(.A(new_new_n77_), .B(new_new_n69_), .C(new_new_n30_), .Y(men0));
  AN2        g0121(.A(i_8_), .B(i_7_), .Y(new_new_n144_));
  NA2        g0122(.A(new_new_n144_), .B(i_6_), .Y(new_new_n145_));
  NO2        g0123(.A(i_12_), .B(i_13_), .Y(new_new_n146_));
  NAi21      g0124(.An(i_5_), .B(i_11_), .Y(new_new_n147_));
  NOi21      g0125(.An(new_new_n146_), .B(new_new_n147_), .Y(new_new_n148_));
  NO2        g0126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NA2        g0127(.A(i_2_), .B(i_3_), .Y(new_new_n150_));
  NO2        g0128(.A(new_new_n150_), .B(i_4_), .Y(new_new_n151_));
  NA3        g0129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  OR2        g0130(.A(new_new_n152_), .B(new_new_n25_), .Y(new_new_n153_));
  AN2        g0131(.A(new_new_n146_), .B(new_new_n83_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n154_), .B(new_new_n27_), .Y(new_new_n155_));
  NA2        g0133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  NO2        g0134(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n36_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n156_), .C(new_new_n155_), .Y(new_new_n159_));
  OR2        g0137(.A(i_0_), .B(i_1_), .Y(new_new_n160_));
  NO3        g0138(.A(new_new_n160_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n161_));
  NAi32      g0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n162_));
  NAi21      g0140(.An(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NOi21      g0141(.An(i_4_), .B(i_10_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n39_), .Y(new_new_n165_));
  NO2        g0143(.A(i_3_), .B(i_5_), .Y(new_new_n166_));
  NO3        g0144(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n167_));
  NA2        g0145(.A(new_new_n167_), .B(new_new_n166_), .Y(new_new_n168_));
  OAI210     g0146(.A0(new_new_n168_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n169_));
  NO2        g0147(.A(new_new_n169_), .B(new_new_n159_), .Y(new_new_n170_));
  AOI210     g0148(.A0(new_new_n170_), .A1(new_new_n153_), .B0(new_new_n145_), .Y(new_new_n171_));
  NA3        g0149(.A(new_new_n73_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n172_));
  NA2        g0150(.A(i_3_), .B(new_new_n48_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_4_), .B(i_9_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_11_), .B(i_13_), .Y(new_new_n175_));
  NA2        g0153(.A(new_new_n175_), .B(new_new_n174_), .Y(new_new_n176_));
  OR2        g0154(.A(new_new_n176_), .B(new_new_n173_), .Y(new_new_n177_));
  NO2        g0155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g0156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n83_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n172_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n183_), .B(new_new_n46_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n36_), .B(i_5_), .Y(new_new_n185_));
  NAi31      g0163(.An(new_new_n185_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n186_));
  NA2        g0164(.A(i_3_), .B(i_5_), .Y(new_new_n187_));
  OR2        g0165(.A(new_new_n187_), .B(new_new_n176_), .Y(new_new_n188_));
  AOI210     g0166(.A0(new_new_n188_), .A1(new_new_n186_), .B0(new_new_n184_), .Y(new_new_n189_));
  NO2        g0167(.A(new_new_n73_), .B(i_5_), .Y(new_new_n190_));
  NO2        g0168(.A(i_13_), .B(i_10_), .Y(new_new_n191_));
  NA3        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n44_), .Y(new_new_n192_));
  NO2        g0170(.A(i_2_), .B(i_1_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_3_), .Y(new_new_n194_));
  NAi21      g0172(.An(i_4_), .B(i_12_), .Y(new_new_n195_));
  NO4        g0173(.A(new_new_n195_), .B(new_new_n194_), .C(new_new_n192_), .D(new_new_n25_), .Y(new_new_n196_));
  NO3        g0174(.A(new_new_n196_), .B(new_new_n189_), .C(new_new_n182_), .Y(new_new_n197_));
  INV        g0175(.A(i_8_), .Y(new_new_n198_));
  NO2        g0176(.A(new_new_n198_), .B(i_7_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(i_6_), .Y(new_new_n200_));
  NO3        g0178(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n201_));
  NA2        g0179(.A(new_new_n201_), .B(new_new_n115_), .Y(new_new_n202_));
  NO3        g0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n205_));
  OAI210     g0183(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n205_), .Y(new_new_n206_));
  AOI210     g0184(.A0(new_new_n206_), .A1(new_new_n204_), .B0(new_new_n202_), .Y(new_new_n207_));
  NO2        g0185(.A(i_3_), .B(i_8_), .Y(new_new_n208_));
  NO3        g0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(new_new_n208_), .C(new_new_n39_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n105_), .B(new_new_n58_), .Y(new_new_n211_));
  INV        g0189(.A(new_new_n211_), .Y(new_new_n212_));
  NO2        g0190(.A(i_13_), .B(i_9_), .Y(new_new_n213_));
  NA3        g0191(.A(new_new_n213_), .B(i_6_), .C(new_new_n198_), .Y(new_new_n214_));
  NAi21      g0192(.An(i_12_), .B(i_3_), .Y(new_new_n215_));
  OR2        g0193(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n44_), .B(i_5_), .Y(new_new_n217_));
  NO3        g0195(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n218_));
  NA3        g0196(.A(new_new_n218_), .B(new_new_n217_), .C(i_10_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n219_), .A1(new_new_n216_), .B0(new_new_n212_), .B1(new_new_n210_), .Y(new_new_n220_));
  AOI210     g0198(.A0(new_new_n220_), .A1(i_7_), .B0(new_new_n207_), .Y(new_new_n221_));
  OAI220     g0199(.A0(new_new_n221_), .A1(i_4_), .B0(new_new_n200_), .B1(new_new_n197_), .Y(new_new_n222_));
  NAi21      g0200(.An(i_12_), .B(i_7_), .Y(new_new_n223_));
  NA3        g0201(.A(i_13_), .B(new_new_n198_), .C(i_10_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  NA2        g0203(.A(i_0_), .B(i_5_), .Y(new_new_n226_));
  NA2        g0204(.A(new_new_n226_), .B(new_new_n106_), .Y(new_new_n227_));
  OAI220     g0205(.A0(new_new_n227_), .A1(new_new_n194_), .B0(new_new_n184_), .B1(new_new_n136_), .Y(new_new_n228_));
  NAi31      g0206(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n36_), .B(i_13_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n232_));
  NA3        g0210(.A(new_new_n232_), .B(new_new_n231_), .C(new_new_n230_), .Y(new_new_n233_));
  INV        g0211(.A(i_13_), .Y(new_new_n234_));
  NO2        g0212(.A(i_12_), .B(new_new_n234_), .Y(new_new_n235_));
  NA3        g0213(.A(new_new_n235_), .B(new_new_n203_), .C(new_new_n201_), .Y(new_new_n236_));
  OAI210     g0214(.A0(new_new_n233_), .A1(new_new_n229_), .B0(new_new_n236_), .Y(new_new_n237_));
  AOI220     g0215(.A0(new_new_n237_), .A1(new_new_n144_), .B0(new_new_n228_), .B1(new_new_n225_), .Y(new_new_n238_));
  NO2        g0216(.A(i_12_), .B(new_new_n37_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n187_), .B(i_4_), .Y(new_new_n240_));
  NA2        g0218(.A(new_new_n240_), .B(new_new_n239_), .Y(new_new_n241_));
  OR2        g0219(.A(i_8_), .B(i_7_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n242_), .B(new_new_n86_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n53_), .B(i_1_), .Y(new_new_n244_));
  NA2        g0222(.A(new_new_n244_), .B(new_new_n243_), .Y(new_new_n245_));
  INV        g0223(.A(i_12_), .Y(new_new_n246_));
  NO2        g0224(.A(new_new_n44_), .B(new_new_n246_), .Y(new_new_n247_));
  NO3        g0225(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n248_));
  NA2        g0226(.A(i_2_), .B(i_1_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n245_), .B(new_new_n241_), .Y(new_new_n250_));
  NO3        g0228(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n251_));
  NAi21      g0229(.An(i_4_), .B(i_3_), .Y(new_new_n252_));
  NO2        g0230(.A(new_new_n252_), .B(new_new_n75_), .Y(new_new_n253_));
  NO2        g0231(.A(i_0_), .B(i_6_), .Y(new_new_n254_));
  NOi41      g0232(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n255_));
  NA2        g0233(.A(new_new_n255_), .B(new_new_n254_), .Y(new_new_n256_));
  NO2        g0234(.A(new_new_n249_), .B(new_new_n187_), .Y(new_new_n257_));
  NAi21      g0235(.An(new_new_n256_), .B(new_new_n257_), .Y(new_new_n258_));
  INV        g0236(.A(new_new_n258_), .Y(new_new_n259_));
  AOI220     g0237(.A0(new_new_n259_), .A1(new_new_n39_), .B0(new_new_n250_), .B1(new_new_n213_), .Y(new_new_n260_));
  NO2        g0238(.A(i_11_), .B(new_new_n234_), .Y(new_new_n261_));
  NOi21      g0239(.An(i_1_), .B(i_6_), .Y(new_new_n262_));
  NAi21      g0240(.An(i_3_), .B(i_7_), .Y(new_new_n263_));
  NA2        g0241(.A(new_new_n246_), .B(i_9_), .Y(new_new_n264_));
  OR4        g0242(.A(new_new_n264_), .B(new_new_n263_), .C(new_new_n262_), .D(new_new_n190_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n266_));
  NO2        g0244(.A(i_12_), .B(i_3_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n73_), .B(i_5_), .Y(new_new_n268_));
  NA2        g0246(.A(i_3_), .B(i_9_), .Y(new_new_n269_));
  NAi21      g0247(.An(i_7_), .B(i_10_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n270_), .B(new_new_n269_), .Y(new_new_n271_));
  NA3        g0249(.A(new_new_n271_), .B(new_new_n268_), .C(new_new_n64_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n272_), .B(new_new_n265_), .Y(new_new_n273_));
  NA3        g0251(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n274_));
  INV        g0252(.A(new_new_n145_), .Y(new_new_n275_));
  NA2        g0253(.A(new_new_n246_), .B(i_13_), .Y(new_new_n276_));
  NO2        g0254(.A(new_new_n276_), .B(new_new_n75_), .Y(new_new_n277_));
  AOI220     g0255(.A0(new_new_n277_), .A1(new_new_n275_), .B0(new_new_n273_), .B1(new_new_n261_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n242_), .B(new_new_n37_), .Y(new_new_n279_));
  NA2        g0257(.A(i_12_), .B(i_6_), .Y(new_new_n280_));
  OR2        g0258(.A(i_13_), .B(i_9_), .Y(new_new_n281_));
  NO3        g0259(.A(new_new_n281_), .B(new_new_n280_), .C(new_new_n48_), .Y(new_new_n282_));
  NO2        g0260(.A(new_new_n252_), .B(i_2_), .Y(new_new_n283_));
  NA3        g0261(.A(new_new_n283_), .B(new_new_n282_), .C(new_new_n44_), .Y(new_new_n284_));
  NA2        g0262(.A(new_new_n261_), .B(i_9_), .Y(new_new_n285_));
  NA2        g0263(.A(new_new_n268_), .B(new_new_n64_), .Y(new_new_n286_));
  OAI210     g0264(.A0(new_new_n286_), .A1(new_new_n285_), .B0(new_new_n284_), .Y(new_new_n287_));
  NA2        g0265(.A(new_new_n157_), .B(new_new_n63_), .Y(new_new_n288_));
  NO3        g0266(.A(i_11_), .B(new_new_n234_), .C(new_new_n25_), .Y(new_new_n289_));
  NO2        g0267(.A(new_new_n263_), .B(i_8_), .Y(new_new_n290_));
  NO2        g0268(.A(i_6_), .B(new_new_n48_), .Y(new_new_n291_));
  NA3        g0269(.A(new_new_n291_), .B(new_new_n290_), .C(new_new_n289_), .Y(new_new_n292_));
  NO3        g0270(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n293_));
  NA3        g0271(.A(new_new_n293_), .B(new_new_n279_), .C(new_new_n235_), .Y(new_new_n294_));
  AOI210     g0272(.A0(new_new_n294_), .A1(new_new_n292_), .B0(new_new_n288_), .Y(new_new_n295_));
  AOI210     g0273(.A0(new_new_n287_), .A1(new_new_n279_), .B0(new_new_n295_), .Y(new_new_n296_));
  NA4        g0274(.A(new_new_n296_), .B(new_new_n278_), .C(new_new_n260_), .D(new_new_n238_), .Y(new_new_n297_));
  NO3        g0275(.A(i_12_), .B(new_new_n234_), .C(new_new_n37_), .Y(new_new_n298_));
  INV        g0276(.A(new_new_n298_), .Y(new_new_n299_));
  NA2        g0277(.A(i_8_), .B(new_new_n103_), .Y(new_new_n300_));
  NOi21      g0278(.An(new_new_n166_), .B(new_new_n86_), .Y(new_new_n301_));
  NO3        g0279(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n302_));
  AOI220     g0280(.A0(new_new_n302_), .A1(new_new_n201_), .B0(new_new_n301_), .B1(new_new_n244_), .Y(new_new_n303_));
  NO2        g0281(.A(new_new_n303_), .B(new_new_n300_), .Y(new_new_n304_));
  NO3        g0282(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n305_));
  NO2        g0283(.A(new_new_n249_), .B(i_0_), .Y(new_new_n306_));
  AOI220     g0284(.A0(new_new_n306_), .A1(new_new_n199_), .B0(new_new_n305_), .B1(new_new_n144_), .Y(new_new_n307_));
  NA2        g0285(.A(new_new_n291_), .B(new_new_n26_), .Y(new_new_n308_));
  NO2        g0286(.A(new_new_n308_), .B(new_new_n307_), .Y(new_new_n309_));
  NA2        g0287(.A(i_0_), .B(i_1_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n310_), .B(i_2_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n59_), .B(i_6_), .Y(new_new_n312_));
  NA3        g0290(.A(new_new_n312_), .B(new_new_n311_), .C(new_new_n166_), .Y(new_new_n313_));
  OAI210     g0291(.A0(new_new_n168_), .A1(new_new_n145_), .B0(new_new_n313_), .Y(new_new_n314_));
  NO3        g0292(.A(new_new_n314_), .B(new_new_n309_), .C(new_new_n304_), .Y(new_new_n315_));
  NO2        g0293(.A(i_3_), .B(i_10_), .Y(new_new_n316_));
  NA3        g0294(.A(new_new_n316_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n317_));
  NO2        g0295(.A(i_2_), .B(new_new_n103_), .Y(new_new_n318_));
  NA2        g0296(.A(i_1_), .B(new_new_n36_), .Y(new_new_n319_));
  NO2        g0297(.A(new_new_n319_), .B(i_8_), .Y(new_new_n320_));
  NOi21      g0298(.An(new_new_n226_), .B(new_new_n105_), .Y(new_new_n321_));
  NA3        g0299(.A(new_new_n321_), .B(new_new_n320_), .C(new_new_n318_), .Y(new_new_n322_));
  AN2        g0300(.A(i_3_), .B(i_10_), .Y(new_new_n323_));
  NA4        g0301(.A(new_new_n323_), .B(new_new_n203_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n324_));
  NO2        g0302(.A(i_5_), .B(new_new_n37_), .Y(new_new_n325_));
  NO2        g0303(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n326_));
  OR2        g0304(.A(new_new_n322_), .B(new_new_n317_), .Y(new_new_n327_));
  OAI220     g0305(.A0(new_new_n327_), .A1(i_6_), .B0(new_new_n315_), .B1(new_new_n299_), .Y(new_new_n328_));
  NO4        g0306(.A(new_new_n328_), .B(new_new_n297_), .C(new_new_n222_), .D(new_new_n171_), .Y(new_new_n329_));
  NO3        g0307(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n330_));
  NO2        g0308(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n331_));
  NA2        g0309(.A(new_new_n306_), .B(new_new_n331_), .Y(new_new_n332_));
  NO3        g0310(.A(i_6_), .B(new_new_n198_), .C(i_7_), .Y(new_new_n333_));
  NA2        g0311(.A(new_new_n333_), .B(new_new_n203_), .Y(new_new_n334_));
  AOI210     g0312(.A0(new_new_n334_), .A1(new_new_n332_), .B0(new_new_n173_), .Y(new_new_n335_));
  NO2        g0313(.A(i_2_), .B(i_3_), .Y(new_new_n336_));
  OR2        g0314(.A(i_0_), .B(i_5_), .Y(new_new_n337_));
  NA2        g0315(.A(new_new_n226_), .B(new_new_n337_), .Y(new_new_n338_));
  NA4        g0316(.A(new_new_n338_), .B(new_new_n243_), .C(new_new_n336_), .D(i_1_), .Y(new_new_n339_));
  NA3        g0317(.A(new_new_n306_), .B(new_new_n301_), .C(new_new_n115_), .Y(new_new_n340_));
  NAi21      g0318(.An(i_8_), .B(i_7_), .Y(new_new_n341_));
  NO2        g0319(.A(new_new_n341_), .B(i_6_), .Y(new_new_n342_));
  NO2        g0320(.A(new_new_n160_), .B(new_new_n46_), .Y(new_new_n343_));
  NA3        g0321(.A(new_new_n343_), .B(new_new_n342_), .C(new_new_n166_), .Y(new_new_n344_));
  NA3        g0322(.A(new_new_n344_), .B(new_new_n340_), .C(new_new_n339_), .Y(new_new_n345_));
  OAI210     g0323(.A0(new_new_n345_), .A1(new_new_n335_), .B0(i_4_), .Y(new_new_n346_));
  NO2        g0324(.A(i_12_), .B(i_10_), .Y(new_new_n347_));
  NOi21      g0325(.An(i_5_), .B(i_0_), .Y(new_new_n348_));
  AOI210     g0326(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n103_), .Y(new_new_n349_));
  NO4        g0327(.A(new_new_n349_), .B(new_new_n319_), .C(new_new_n348_), .D(new_new_n131_), .Y(new_new_n350_));
  NA4        g0328(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n351_));
  NA2        g0329(.A(new_new_n350_), .B(new_new_n347_), .Y(new_new_n352_));
  NO2        g0330(.A(i_6_), .B(i_8_), .Y(new_new_n353_));
  NOi21      g0331(.An(i_0_), .B(i_2_), .Y(new_new_n354_));
  AN2        g0332(.A(new_new_n354_), .B(new_new_n353_), .Y(new_new_n355_));
  NO2        g0333(.A(i_1_), .B(i_7_), .Y(new_new_n356_));
  AO220      g0334(.A0(new_new_n356_), .A1(new_new_n355_), .B0(new_new_n342_), .B1(new_new_n244_), .Y(new_new_n357_));
  NA3        g0335(.A(new_new_n357_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n358_));
  NA3        g0336(.A(new_new_n358_), .B(new_new_n352_), .C(new_new_n346_), .Y(new_new_n359_));
  NO3        g0337(.A(new_new_n242_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n360_));
  NO3        g0338(.A(new_new_n341_), .B(i_2_), .C(i_1_), .Y(new_new_n361_));
  OAI210     g0339(.A0(new_new_n361_), .A1(new_new_n360_), .B0(i_6_), .Y(new_new_n362_));
  NA3        g0340(.A(new_new_n262_), .B(new_new_n318_), .C(new_new_n198_), .Y(new_new_n363_));
  AOI210     g0341(.A0(new_new_n363_), .A1(new_new_n362_), .B0(new_new_n338_), .Y(new_new_n364_));
  NOi21      g0342(.An(new_new_n156_), .B(new_new_n106_), .Y(new_new_n365_));
  NO2        g0343(.A(new_new_n365_), .B(new_new_n127_), .Y(new_new_n366_));
  OAI210     g0344(.A0(new_new_n366_), .A1(new_new_n364_), .B0(i_3_), .Y(new_new_n367_));
  INV        g0345(.A(new_new_n84_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n310_), .B(new_new_n81_), .Y(new_new_n369_));
  NA2        g0347(.A(new_new_n369_), .B(new_new_n135_), .Y(new_new_n370_));
  NO2        g0348(.A(new_new_n94_), .B(new_new_n198_), .Y(new_new_n371_));
  NA3        g0349(.A(new_new_n321_), .B(new_new_n371_), .C(new_new_n63_), .Y(new_new_n372_));
  AOI210     g0350(.A0(new_new_n372_), .A1(new_new_n370_), .B0(new_new_n368_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n198_), .B(i_9_), .Y(new_new_n374_));
  NA2        g0352(.A(new_new_n374_), .B(new_new_n211_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n375_), .B(new_new_n46_), .Y(new_new_n376_));
  NO3        g0354(.A(new_new_n376_), .B(new_new_n373_), .C(new_new_n309_), .Y(new_new_n377_));
  AOI210     g0355(.A0(new_new_n377_), .A1(new_new_n367_), .B0(new_new_n165_), .Y(new_new_n378_));
  AOI210     g0356(.A0(new_new_n359_), .A1(new_new_n330_), .B0(new_new_n378_), .Y(new_new_n379_));
  NOi32      g0357(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n380_));
  INV        g0358(.A(new_new_n380_), .Y(new_new_n381_));
  NAi21      g0359(.An(i_0_), .B(i_6_), .Y(new_new_n382_));
  NAi21      g0360(.An(i_1_), .B(i_5_), .Y(new_new_n383_));
  NA2        g0361(.A(new_new_n383_), .B(new_new_n382_), .Y(new_new_n384_));
  NA2        g0362(.A(new_new_n384_), .B(new_new_n25_), .Y(new_new_n385_));
  OAI210     g0363(.A0(new_new_n385_), .A1(new_new_n162_), .B0(new_new_n256_), .Y(new_new_n386_));
  NAi41      g0364(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n387_));
  OAI220     g0365(.A0(new_new_n387_), .A1(new_new_n383_), .B0(new_new_n229_), .B1(new_new_n162_), .Y(new_new_n388_));
  AOI210     g0366(.A0(new_new_n387_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n389_));
  NOi32      g0367(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n390_));
  NAi21      g0368(.An(i_6_), .B(i_1_), .Y(new_new_n391_));
  NA3        g0369(.A(new_new_n391_), .B(new_new_n390_), .C(new_new_n46_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n392_), .B(i_0_), .Y(new_new_n393_));
  OR3        g0371(.A(new_new_n393_), .B(new_new_n389_), .C(new_new_n388_), .Y(new_new_n394_));
  NO2        g0372(.A(i_1_), .B(new_new_n103_), .Y(new_new_n395_));
  NAi21      g0373(.An(i_3_), .B(i_4_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n396_), .B(i_9_), .Y(new_new_n397_));
  AN2        g0375(.A(i_6_), .B(i_7_), .Y(new_new_n398_));
  OAI210     g0376(.A0(new_new_n398_), .A1(new_new_n395_), .B0(new_new_n397_), .Y(new_new_n399_));
  NA2        g0377(.A(i_2_), .B(i_7_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n396_), .B(i_10_), .Y(new_new_n401_));
  NA3        g0379(.A(new_new_n401_), .B(new_new_n400_), .C(new_new_n254_), .Y(new_new_n402_));
  AOI210     g0380(.A0(new_new_n402_), .A1(new_new_n399_), .B0(new_new_n190_), .Y(new_new_n403_));
  AOI210     g0381(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n404_));
  OAI210     g0382(.A0(new_new_n404_), .A1(new_new_n193_), .B0(new_new_n401_), .Y(new_new_n405_));
  AOI220     g0383(.A0(new_new_n401_), .A1(new_new_n356_), .B0(new_new_n248_), .B1(new_new_n193_), .Y(new_new_n406_));
  AOI210     g0384(.A0(new_new_n406_), .A1(new_new_n405_), .B0(i_5_), .Y(new_new_n407_));
  NO4        g0385(.A(new_new_n407_), .B(new_new_n403_), .C(new_new_n394_), .D(new_new_n386_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n408_), .B(new_new_n381_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n410_));
  AN2        g0388(.A(i_12_), .B(i_5_), .Y(new_new_n411_));
  NO2        g0389(.A(i_4_), .B(new_new_n26_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n412_), .B(new_new_n411_), .Y(new_new_n413_));
  NO2        g0391(.A(i_11_), .B(i_6_), .Y(new_new_n414_));
  NA3        g0392(.A(new_new_n414_), .B(new_new_n343_), .C(new_new_n234_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n415_), .B(new_new_n413_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n252_), .B(i_5_), .Y(new_new_n417_));
  NO2        g0395(.A(i_5_), .B(i_10_), .Y(new_new_n418_));
  AOI220     g0396(.A0(new_new_n418_), .A1(new_new_n283_), .B0(new_new_n417_), .B1(new_new_n203_), .Y(new_new_n419_));
  NA2        g0397(.A(new_new_n146_), .B(new_new_n45_), .Y(new_new_n420_));
  NO2        g0398(.A(new_new_n420_), .B(new_new_n419_), .Y(new_new_n421_));
  OAI210     g0399(.A0(new_new_n421_), .A1(new_new_n416_), .B0(new_new_n410_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n152_), .B(new_new_n86_), .Y(new_new_n424_));
  OAI210     g0402(.A0(new_new_n424_), .A1(new_new_n416_), .B0(new_new_n423_), .Y(new_new_n425_));
  NO3        g0403(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n426_));
  NO2        g0404(.A(i_3_), .B(new_new_n103_), .Y(new_new_n427_));
  NA3        g0405(.A(new_new_n316_), .B(new_new_n75_), .C(new_new_n54_), .Y(new_new_n428_));
  NO2        g0406(.A(i_11_), .B(i_12_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n429_), .B(new_new_n36_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n428_), .B(new_new_n430_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n418_), .B(new_new_n246_), .Y(new_new_n432_));
  NA3        g0410(.A(new_new_n115_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n433_), .B(new_new_n229_), .Y(new_new_n434_));
  NAi21      g0412(.An(i_13_), .B(i_0_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n435_), .B(new_new_n249_), .Y(new_new_n436_));
  OAI210     g0414(.A0(new_new_n434_), .A1(new_new_n431_), .B0(new_new_n436_), .Y(new_new_n437_));
  NA3        g0415(.A(new_new_n437_), .B(new_new_n425_), .C(new_new_n422_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n44_), .B(new_new_n234_), .Y(new_new_n439_));
  NO3        g0417(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n440_));
  NO2        g0418(.A(i_0_), .B(i_11_), .Y(new_new_n441_));
  AN2        g0419(.A(i_1_), .B(i_6_), .Y(new_new_n442_));
  NOi21      g0420(.An(i_2_), .B(i_12_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n443_), .B(new_new_n442_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(new_new_n1147_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n144_), .B(i_9_), .Y(new_new_n446_));
  NO2        g0424(.A(new_new_n446_), .B(i_4_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n445_), .B(new_new_n447_), .Y(new_new_n448_));
  NAi21      g0426(.An(i_9_), .B(i_4_), .Y(new_new_n449_));
  OR2        g0427(.A(i_13_), .B(i_10_), .Y(new_new_n450_));
  NO3        g0428(.A(new_new_n450_), .B(new_new_n120_), .C(new_new_n449_), .Y(new_new_n451_));
  NO2        g0429(.A(new_new_n176_), .B(new_new_n126_), .Y(new_new_n452_));
  OR2        g0430(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n298_), .B(new_new_n454_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n291_), .B(new_new_n218_), .Y(new_new_n456_));
  OAI220     g0434(.A0(new_new_n456_), .A1(new_new_n453_), .B0(new_new_n455_), .B1(new_new_n365_), .Y(new_new_n457_));
  INV        g0435(.A(new_new_n457_), .Y(new_new_n458_));
  AOI210     g0436(.A0(new_new_n458_), .A1(new_new_n448_), .B0(new_new_n26_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n340_), .B(new_new_n339_), .Y(new_new_n460_));
  AOI220     g0438(.A0(new_new_n312_), .A1(new_new_n302_), .B0(new_new_n306_), .B1(new_new_n331_), .Y(new_new_n461_));
  NO2        g0439(.A(new_new_n461_), .B(new_new_n173_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n187_), .B(new_new_n86_), .Y(new_new_n463_));
  AOI220     g0441(.A0(new_new_n463_), .A1(new_new_n311_), .B0(new_new_n293_), .B1(new_new_n218_), .Y(new_new_n464_));
  NO2        g0442(.A(new_new_n464_), .B(new_new_n300_), .Y(new_new_n465_));
  NO3        g0443(.A(new_new_n465_), .B(new_new_n462_), .C(new_new_n460_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n201_), .B(new_new_n98_), .Y(new_new_n467_));
  NA3        g0445(.A(new_new_n343_), .B(new_new_n166_), .C(new_new_n86_), .Y(new_new_n468_));
  AOI210     g0446(.A0(new_new_n468_), .A1(new_new_n467_), .B0(new_new_n341_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n198_), .B(i_10_), .Y(new_new_n470_));
  NA3        g0448(.A(new_new_n268_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n312_), .B(new_new_n244_), .Y(new_new_n472_));
  OAI220     g0450(.A0(new_new_n472_), .A1(new_new_n187_), .B0(new_new_n471_), .B1(new_new_n470_), .Y(new_new_n473_));
  NO2        g0451(.A(i_3_), .B(new_new_n48_), .Y(new_new_n474_));
  NA3        g0452(.A(new_new_n356_), .B(new_new_n355_), .C(new_new_n474_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n333_), .B(new_new_n338_), .Y(new_new_n476_));
  OAI210     g0454(.A0(new_new_n476_), .A1(new_new_n194_), .B0(new_new_n475_), .Y(new_new_n477_));
  NO3        g0455(.A(new_new_n477_), .B(new_new_n473_), .C(new_new_n469_), .Y(new_new_n478_));
  AOI210     g0456(.A0(new_new_n478_), .A1(new_new_n466_), .B0(new_new_n285_), .Y(new_new_n479_));
  NO4        g0457(.A(new_new_n479_), .B(new_new_n459_), .C(new_new_n438_), .D(new_new_n409_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n63_), .B(i_4_), .Y(new_new_n481_));
  NO2        g0459(.A(i_10_), .B(i_9_), .Y(new_new_n482_));
  NAi21      g0460(.An(i_12_), .B(i_8_), .Y(new_new_n483_));
  NO2        g0461(.A(new_new_n483_), .B(i_3_), .Y(new_new_n484_));
  NO2        g0462(.A(new_new_n46_), .B(i_4_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n485_), .B(new_new_n106_), .Y(new_new_n486_));
  NO2        g0464(.A(new_new_n486_), .B(new_new_n210_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n326_), .B(i_0_), .Y(new_new_n488_));
  NO3        g0466(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n280_), .B(new_new_n99_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n490_), .B(new_new_n489_), .Y(new_new_n491_));
  NA2        g0469(.A(i_8_), .B(i_9_), .Y(new_new_n492_));
  AOI210     g0470(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n493_));
  OR2        g0471(.A(new_new_n493_), .B(new_new_n492_), .Y(new_new_n494_));
  NA2        g0472(.A(new_new_n298_), .B(new_new_n211_), .Y(new_new_n495_));
  OAI220     g0473(.A0(new_new_n495_), .A1(new_new_n494_), .B0(new_new_n491_), .B1(new_new_n488_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n261_), .B(new_new_n325_), .Y(new_new_n497_));
  NO3        g0475(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n498_));
  INV        g0476(.A(new_new_n498_), .Y(new_new_n499_));
  NA3        g0477(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n500_));
  NA4        g0478(.A(new_new_n147_), .B(new_new_n118_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n501_));
  OAI220     g0479(.A0(new_new_n501_), .A1(new_new_n500_), .B0(new_new_n499_), .B1(new_new_n497_), .Y(new_new_n502_));
  NO3        g0480(.A(new_new_n502_), .B(new_new_n496_), .C(new_new_n487_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n311_), .B(new_new_n110_), .Y(new_new_n504_));
  OR2        g0482(.A(new_new_n504_), .B(new_new_n214_), .Y(new_new_n505_));
  OA210      g0483(.A0(new_new_n375_), .A1(new_new_n103_), .B0(new_new_n313_), .Y(new_new_n506_));
  OA220      g0484(.A0(new_new_n506_), .A1(new_new_n165_), .B0(new_new_n505_), .B1(new_new_n241_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n98_), .B(i_13_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n463_), .B(new_new_n410_), .Y(new_new_n509_));
  NO2        g0487(.A(i_2_), .B(i_13_), .Y(new_new_n510_));
  NA3        g0488(.A(new_new_n510_), .B(new_new_n164_), .C(new_new_n101_), .Y(new_new_n511_));
  OAI220     g0489(.A0(new_new_n511_), .A1(new_new_n246_), .B0(new_new_n509_), .B1(new_new_n508_), .Y(new_new_n512_));
  NO3        g0490(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n513_));
  NO2        g0491(.A(i_6_), .B(i_7_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n514_), .B(new_new_n513_), .Y(new_new_n515_));
  NO2        g0493(.A(i_11_), .B(i_1_), .Y(new_new_n516_));
  NO2        g0494(.A(new_new_n73_), .B(i_3_), .Y(new_new_n517_));
  OR2        g0495(.A(i_11_), .B(i_8_), .Y(new_new_n518_));
  NOi21      g0496(.An(i_2_), .B(i_7_), .Y(new_new_n519_));
  NAi31      g0497(.An(new_new_n518_), .B(new_new_n519_), .C(new_new_n517_), .Y(new_new_n520_));
  NO2        g0498(.A(new_new_n450_), .B(i_6_), .Y(new_new_n521_));
  NA3        g0499(.A(new_new_n521_), .B(new_new_n481_), .C(new_new_n75_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n522_), .B(new_new_n520_), .Y(new_new_n523_));
  NO2        g0501(.A(i_3_), .B(new_new_n198_), .Y(new_new_n524_));
  NO2        g0502(.A(i_6_), .B(i_10_), .Y(new_new_n525_));
  NA4        g0503(.A(new_new_n525_), .B(new_new_n330_), .C(new_new_n524_), .D(new_new_n246_), .Y(new_new_n526_));
  NO2        g0504(.A(new_new_n526_), .B(new_new_n158_), .Y(new_new_n527_));
  NA3        g0505(.A(new_new_n255_), .B(new_new_n175_), .C(new_new_n135_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n160_), .B(i_3_), .Y(new_new_n530_));
  NAi31      g0508(.An(new_new_n529_), .B(new_new_n530_), .C(new_new_n235_), .Y(new_new_n531_));
  NA3        g0509(.A(new_new_n423_), .B(new_new_n183_), .C(new_new_n151_), .Y(new_new_n532_));
  NA3        g0510(.A(new_new_n532_), .B(new_new_n531_), .C(new_new_n528_), .Y(new_new_n533_));
  NO4        g0511(.A(new_new_n533_), .B(new_new_n527_), .C(new_new_n523_), .D(new_new_n512_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n489_), .B(new_new_n411_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n498_), .B(new_new_n418_), .Y(new_new_n536_));
  NO2        g0514(.A(new_new_n536_), .B(new_new_n233_), .Y(new_new_n537_));
  NAi21      g0515(.An(new_new_n224_), .B(new_new_n429_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n356_), .B(new_new_n226_), .Y(new_new_n539_));
  NO2        g0517(.A(new_new_n26_), .B(i_5_), .Y(new_new_n540_));
  NO2        g0518(.A(i_0_), .B(new_new_n86_), .Y(new_new_n541_));
  NA3        g0519(.A(new_new_n541_), .B(new_new_n540_), .C(new_new_n144_), .Y(new_new_n542_));
  OR3        g0520(.A(new_new_n319_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n543_));
  OAI220     g0521(.A0(new_new_n543_), .A1(new_new_n542_), .B0(new_new_n539_), .B1(new_new_n538_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n27_), .B(i_10_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n330_), .B(new_new_n248_), .Y(new_new_n546_));
  OAI220     g0524(.A0(new_new_n546_), .A1(new_new_n471_), .B0(new_new_n545_), .B1(new_new_n508_), .Y(new_new_n547_));
  NA4        g0525(.A(new_new_n323_), .B(new_new_n232_), .C(new_new_n73_), .D(new_new_n246_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n548_), .B(new_new_n515_), .Y(new_new_n549_));
  NO4        g0527(.A(new_new_n549_), .B(new_new_n547_), .C(new_new_n544_), .D(new_new_n537_), .Y(new_new_n550_));
  NA4        g0528(.A(new_new_n550_), .B(new_new_n534_), .C(new_new_n507_), .D(new_new_n503_), .Y(new_new_n551_));
  NA3        g0529(.A(new_new_n323_), .B(new_new_n180_), .C(new_new_n178_), .Y(new_new_n552_));
  OAI210     g0530(.A0(new_new_n317_), .A1(new_new_n185_), .B0(new_new_n552_), .Y(new_new_n553_));
  AN2        g0531(.A(new_new_n302_), .B(new_new_n243_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n553_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n125_), .B(new_new_n114_), .Y(new_new_n556_));
  AO220      g0534(.A0(new_new_n556_), .A1(new_new_n489_), .B0(new_new_n451_), .B1(i_6_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n330_), .B(new_new_n167_), .Y(new_new_n558_));
  OAI210     g0536(.A0(new_new_n558_), .A1(new_new_n241_), .B0(new_new_n324_), .Y(new_new_n559_));
  AOI220     g0537(.A0(new_new_n559_), .A1(new_new_n342_), .B0(new_new_n557_), .B1(new_new_n326_), .Y(new_new_n560_));
  NA2        g0538(.A(new_new_n411_), .B(new_new_n234_), .Y(new_new_n561_));
  NA2        g0539(.A(new_new_n380_), .B(new_new_n73_), .Y(new_new_n562_));
  NA2        g0540(.A(new_new_n398_), .B(new_new_n390_), .Y(new_new_n563_));
  AO210      g0541(.A0(new_new_n562_), .A1(new_new_n561_), .B0(new_new_n563_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n36_), .B(i_8_), .Y(new_new_n565_));
  INV        g0543(.A(new_new_n451_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n566_), .B(new_new_n564_), .Y(new_new_n567_));
  INV        g0545(.A(new_new_n567_), .Y(new_new_n568_));
  NA2        g0546(.A(new_new_n268_), .B(new_new_n64_), .Y(new_new_n569_));
  OAI210     g0547(.A0(i_8_), .A1(new_new_n569_), .B0(new_new_n137_), .Y(new_new_n570_));
  AOI210     g0548(.A0(new_new_n199_), .A1(i_9_), .B0(new_new_n279_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n571_), .B(new_new_n204_), .Y(new_new_n572_));
  OR2        g0550(.A(new_new_n187_), .B(i_4_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n573_), .B(new_new_n86_), .Y(new_new_n574_));
  AOI220     g0552(.A0(new_new_n574_), .A1(new_new_n572_), .B0(new_new_n570_), .B1(new_new_n452_), .Y(new_new_n575_));
  NA4        g0553(.A(new_new_n575_), .B(new_new_n568_), .C(new_new_n560_), .D(new_new_n555_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n417_), .B(new_new_n311_), .Y(new_new_n577_));
  OAI210     g0555(.A0(new_new_n413_), .A1(new_new_n172_), .B0(new_new_n577_), .Y(new_new_n578_));
  NO2        g0556(.A(i_12_), .B(new_new_n198_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n579_), .B(new_new_n234_), .Y(new_new_n580_));
  NA3        g0558(.A(new_new_n525_), .B(new_new_n178_), .C(new_new_n27_), .Y(new_new_n581_));
  NO3        g0559(.A(new_new_n581_), .B(new_new_n580_), .C(new_new_n504_), .Y(new_new_n582_));
  NOi31      g0560(.An(new_new_n333_), .B(new_new_n450_), .C(new_new_n38_), .Y(new_new_n583_));
  OAI210     g0561(.A0(new_new_n583_), .A1(new_new_n582_), .B0(new_new_n578_), .Y(new_new_n584_));
  NO2        g0562(.A(i_8_), .B(i_7_), .Y(new_new_n585_));
  OAI210     g0563(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n586_));
  NA2        g0564(.A(new_new_n586_), .B(new_new_n232_), .Y(new_new_n587_));
  AOI220     g0565(.A0(new_new_n343_), .A1(new_new_n39_), .B0(new_new_n244_), .B1(new_new_n213_), .Y(new_new_n588_));
  OAI220     g0566(.A0(new_new_n588_), .A1(new_new_n573_), .B0(new_new_n587_), .B1(new_new_n252_), .Y(new_new_n589_));
  NA2        g0567(.A(new_new_n44_), .B(i_10_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n590_), .B(i_6_), .Y(new_new_n591_));
  NA3        g0569(.A(new_new_n591_), .B(new_new_n589_), .C(new_new_n585_), .Y(new_new_n592_));
  AOI220     g0570(.A0(new_new_n463_), .A1(new_new_n343_), .B0(new_new_n257_), .B1(new_new_n254_), .Y(new_new_n593_));
  OAI220     g0571(.A0(new_new_n593_), .A1(new_new_n276_), .B0(new_new_n508_), .B1(new_new_n136_), .Y(new_new_n594_));
  NA2        g0572(.A(new_new_n594_), .B(new_new_n279_), .Y(new_new_n595_));
  NOi31      g0573(.An(new_new_n306_), .B(new_new_n317_), .C(new_new_n185_), .Y(new_new_n596_));
  NA3        g0574(.A(new_new_n323_), .B(new_new_n178_), .C(new_new_n98_), .Y(new_new_n597_));
  NO2        g0575(.A(new_new_n230_), .B(new_new_n44_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n160_), .B(i_5_), .Y(new_new_n599_));
  NA3        g0577(.A(new_new_n599_), .B(new_new_n439_), .C(new_new_n336_), .Y(new_new_n600_));
  OAI210     g0578(.A0(new_new_n600_), .A1(new_new_n598_), .B0(new_new_n597_), .Y(new_new_n601_));
  OAI210     g0579(.A0(new_new_n601_), .A1(new_new_n596_), .B0(new_new_n498_), .Y(new_new_n602_));
  NA4        g0580(.A(new_new_n602_), .B(new_new_n595_), .C(new_new_n592_), .D(new_new_n584_), .Y(new_new_n603_));
  NA3        g0581(.A(new_new_n226_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n604_));
  NA2        g0582(.A(new_new_n298_), .B(new_new_n84_), .Y(new_new_n605_));
  AOI210     g0583(.A0(new_new_n604_), .A1(new_new_n370_), .B0(new_new_n605_), .Y(new_new_n606_));
  NA2        g0584(.A(new_new_n312_), .B(new_new_n302_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n607_), .B(new_new_n177_), .Y(new_new_n608_));
  NA2        g0586(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n609_));
  NA2        g0587(.A(new_new_n482_), .B(new_new_n230_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n609_), .B(new_new_n610_), .Y(new_new_n611_));
  AOI210     g0589(.A0(new_new_n391_), .A1(new_new_n46_), .B0(new_new_n395_), .Y(new_new_n612_));
  NA2        g0590(.A(i_0_), .B(new_new_n48_), .Y(new_new_n613_));
  NA3        g0591(.A(new_new_n579_), .B(new_new_n289_), .C(new_new_n613_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n612_), .B(new_new_n614_), .Y(new_new_n615_));
  NO4        g0593(.A(new_new_n615_), .B(new_new_n611_), .C(new_new_n608_), .D(new_new_n606_), .Y(new_new_n616_));
  NO4        g0594(.A(new_new_n262_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n617_));
  NO3        g0595(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n242_), .B(new_new_n36_), .Y(new_new_n619_));
  AN2        g0597(.A(new_new_n619_), .B(new_new_n618_), .Y(new_new_n620_));
  OA210      g0598(.A0(new_new_n620_), .A1(new_new_n617_), .B0(new_new_n380_), .Y(new_new_n621_));
  NO2        g0599(.A(new_new_n450_), .B(i_1_), .Y(new_new_n622_));
  NOi31      g0600(.An(new_new_n622_), .B(new_new_n490_), .C(new_new_n73_), .Y(new_new_n623_));
  AN4        g0601(.A(new_new_n623_), .B(new_new_n447_), .C(new_new_n540_), .D(i_2_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n461_), .B(new_new_n181_), .Y(new_new_n625_));
  NO3        g0603(.A(new_new_n625_), .B(new_new_n624_), .C(new_new_n621_), .Y(new_new_n626_));
  NOi21      g0604(.An(i_10_), .B(i_6_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n628_));
  AOI220     g0606(.A0(new_new_n298_), .A1(new_new_n628_), .B0(new_new_n289_), .B1(new_new_n627_), .Y(new_new_n629_));
  NO2        g0607(.A(new_new_n629_), .B(new_new_n488_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n631_));
  NA2        g0609(.A(new_new_n333_), .B(new_new_n167_), .Y(new_new_n632_));
  AOI220     g0610(.A0(new_new_n632_), .A1(new_new_n472_), .B0(new_new_n188_), .B1(new_new_n186_), .Y(new_new_n633_));
  NO2        g0611(.A(new_new_n203_), .B(new_new_n37_), .Y(new_new_n634_));
  NOi31      g0612(.An(new_new_n148_), .B(new_new_n634_), .C(new_new_n351_), .Y(new_new_n635_));
  NO3        g0613(.A(new_new_n635_), .B(new_new_n633_), .C(new_new_n630_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n562_), .B(new_new_n406_), .Y(new_new_n637_));
  INV        g0615(.A(new_new_n336_), .Y(new_new_n638_));
  NO2        g0616(.A(i_12_), .B(new_new_n86_), .Y(new_new_n639_));
  NA3        g0617(.A(new_new_n639_), .B(new_new_n289_), .C(new_new_n613_), .Y(new_new_n640_));
  NA3        g0618(.A(new_new_n414_), .B(new_new_n298_), .C(new_new_n226_), .Y(new_new_n641_));
  AOI210     g0619(.A0(new_new_n641_), .A1(new_new_n640_), .B0(new_new_n638_), .Y(new_new_n642_));
  NA2        g0620(.A(new_new_n178_), .B(i_0_), .Y(new_new_n643_));
  NO3        g0621(.A(new_new_n643_), .B(new_new_n362_), .C(new_new_n317_), .Y(new_new_n644_));
  OR2        g0622(.A(i_2_), .B(i_5_), .Y(new_new_n645_));
  OR2        g0623(.A(new_new_n645_), .B(new_new_n442_), .Y(new_new_n646_));
  AOI210     g0624(.A0(new_new_n400_), .A1(new_new_n254_), .B0(new_new_n203_), .Y(new_new_n647_));
  AOI210     g0625(.A0(new_new_n647_), .A1(new_new_n646_), .B0(new_new_n538_), .Y(new_new_n648_));
  NO4        g0626(.A(new_new_n648_), .B(new_new_n644_), .C(new_new_n642_), .D(new_new_n637_), .Y(new_new_n649_));
  NA4        g0627(.A(new_new_n649_), .B(new_new_n636_), .C(new_new_n626_), .D(new_new_n616_), .Y(new_new_n650_));
  NO4        g0628(.A(new_new_n650_), .B(new_new_n603_), .C(new_new_n576_), .D(new_new_n551_), .Y(new_new_n651_));
  NA4        g0629(.A(new_new_n651_), .B(new_new_n480_), .C(new_new_n379_), .D(new_new_n329_), .Y(men7));
  NO2        g0630(.A(new_new_n94_), .B(new_new_n54_), .Y(new_new_n653_));
  NO2        g0631(.A(new_new_n110_), .B(new_new_n91_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n412_), .B(new_new_n654_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n525_), .B(new_new_n84_), .Y(new_new_n656_));
  NA2        g0634(.A(i_11_), .B(new_new_n198_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n146_), .B(new_new_n657_), .Y(new_new_n658_));
  OAI210     g0636(.A0(new_new_n658_), .A1(new_new_n656_), .B0(new_new_n655_), .Y(new_new_n659_));
  NA3        g0637(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n246_), .B(i_4_), .Y(new_new_n661_));
  NA2        g0639(.A(new_new_n661_), .B(i_8_), .Y(new_new_n662_));
  AOI210     g0640(.A0(new_new_n662_), .A1(new_new_n107_), .B0(new_new_n660_), .Y(new_new_n663_));
  NA2        g0641(.A(i_2_), .B(new_new_n86_), .Y(new_new_n664_));
  OAI210     g0642(.A0(new_new_n89_), .A1(new_new_n208_), .B0(new_new_n209_), .Y(new_new_n665_));
  NO2        g0643(.A(i_7_), .B(new_new_n37_), .Y(new_new_n666_));
  NA2        g0644(.A(i_4_), .B(i_8_), .Y(new_new_n667_));
  AOI210     g0645(.A0(new_new_n667_), .A1(new_new_n323_), .B0(new_new_n666_), .Y(new_new_n668_));
  OAI220     g0646(.A0(new_new_n668_), .A1(new_new_n664_), .B0(new_new_n665_), .B1(i_13_), .Y(new_new_n669_));
  NO4        g0647(.A(new_new_n669_), .B(new_new_n663_), .C(new_new_n659_), .D(new_new_n653_), .Y(new_new_n670_));
  AOI210     g0648(.A0(new_new_n131_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n671_));
  AOI210     g0649(.A0(new_new_n671_), .A1(new_new_n246_), .B0(new_new_n164_), .Y(new_new_n672_));
  OR2        g0650(.A(i_6_), .B(i_10_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n673_), .B(new_new_n23_), .Y(new_new_n674_));
  OR3        g0652(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n675_));
  NO3        g0653(.A(new_new_n675_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n676_));
  INV        g0654(.A(new_new_n205_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n676_), .B(new_new_n674_), .Y(new_new_n678_));
  OA220      g0656(.A0(new_new_n678_), .A1(new_new_n638_), .B0(new_new_n672_), .B1(new_new_n281_), .Y(new_new_n679_));
  AOI210     g0657(.A0(new_new_n679_), .A1(new_new_n670_), .B0(new_new_n63_), .Y(new_new_n680_));
  NOi21      g0658(.An(i_11_), .B(i_7_), .Y(new_new_n681_));
  AO210      g0659(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n682_), .B(new_new_n681_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n683_), .B(new_new_n213_), .Y(new_new_n684_));
  NA3        g0662(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n685_));
  NAi31      g0663(.An(new_new_n685_), .B(new_new_n223_), .C(i_11_), .Y(new_new_n686_));
  AOI210     g0664(.A0(new_new_n686_), .A1(new_new_n684_), .B0(new_new_n63_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n688_));
  AO210      g0666(.A0(new_new_n688_), .A1(new_new_n406_), .B0(new_new_n40_), .Y(new_new_n689_));
  NO3        g0667(.A(new_new_n270_), .B(new_new_n215_), .C(new_new_n657_), .Y(new_new_n690_));
  NA2        g0668(.A(new_new_n690_), .B(new_new_n63_), .Y(new_new_n691_));
  NA2        g0669(.A(new_new_n443_), .B(new_new_n31_), .Y(new_new_n692_));
  OR2        g0670(.A(new_new_n215_), .B(new_new_n110_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n693_), .B(new_new_n692_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n63_), .B(i_9_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(i_4_), .Y(new_new_n696_));
  NA2        g0674(.A(new_new_n696_), .B(new_new_n694_), .Y(new_new_n697_));
  NO2        g0675(.A(i_1_), .B(i_12_), .Y(new_new_n698_));
  NA3        g0676(.A(new_new_n698_), .B(new_new_n112_), .C(new_new_n24_), .Y(new_new_n699_));
  NA4        g0677(.A(new_new_n699_), .B(new_new_n697_), .C(new_new_n691_), .D(new_new_n689_), .Y(new_new_n700_));
  OAI210     g0678(.A0(new_new_n700_), .A1(new_new_n687_), .B0(i_6_), .Y(new_new_n701_));
  OAI210     g0679(.A0(new_new_n685_), .A1(new_new_n110_), .B0(new_new_n500_), .Y(new_new_n702_));
  NA2        g0680(.A(new_new_n702_), .B(new_new_n639_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n246_), .B(new_new_n86_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n703_), .B(new_new_n491_), .Y(new_new_n705_));
  NO4        g0683(.A(new_new_n223_), .B(new_new_n131_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n706_), .B(new_new_n695_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n246_), .B(i_6_), .Y(new_new_n708_));
  NO3        g0686(.A(new_new_n673_), .B(new_new_n242_), .C(new_new_n23_), .Y(new_new_n709_));
  AOI210     g0687(.A0(i_1_), .A1(new_new_n271_), .B0(new_new_n709_), .Y(new_new_n710_));
  OAI210     g0688(.A0(new_new_n710_), .A1(new_new_n44_), .B0(new_new_n707_), .Y(new_new_n711_));
  NA3        g0689(.A(new_new_n585_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n712_));
  NA3        g0690(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n46_), .B(i_1_), .Y(new_new_n714_));
  NA3        g0692(.A(new_new_n714_), .B(new_new_n280_), .C(new_new_n44_), .Y(new_new_n715_));
  NO2        g0693(.A(new_new_n715_), .B(new_new_n713_), .Y(new_new_n716_));
  NA3        g0694(.A(new_new_n695_), .B(new_new_n336_), .C(i_6_), .Y(new_new_n717_));
  NO2        g0695(.A(new_new_n717_), .B(new_new_n23_), .Y(new_new_n718_));
  NAi21      g0696(.An(new_new_n712_), .B(new_new_n93_), .Y(new_new_n719_));
  NA2        g0697(.A(new_new_n714_), .B(new_new_n280_), .Y(new_new_n720_));
  NO2        g0698(.A(i_11_), .B(new_new_n37_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n721_), .B(new_new_n24_), .Y(new_new_n722_));
  OAI210     g0700(.A0(new_new_n722_), .A1(new_new_n720_), .B0(new_new_n719_), .Y(new_new_n723_));
  OR3        g0701(.A(new_new_n723_), .B(new_new_n718_), .C(new_new_n716_), .Y(new_new_n724_));
  NO3        g0702(.A(new_new_n724_), .B(new_new_n711_), .C(new_new_n705_), .Y(new_new_n725_));
  NO2        g0703(.A(new_new_n246_), .B(new_new_n103_), .Y(new_new_n726_));
  NO2        g0704(.A(new_new_n726_), .B(new_new_n681_), .Y(new_new_n727_));
  NA2        g0705(.A(new_new_n727_), .B(i_1_), .Y(new_new_n728_));
  NO2        g0706(.A(new_new_n728_), .B(new_new_n675_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n449_), .B(new_new_n86_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n729_), .B(new_new_n46_), .Y(new_new_n731_));
  NA2        g0709(.A(i_3_), .B(new_new_n198_), .Y(new_new_n732_));
  NO2        g0710(.A(new_new_n732_), .B(new_new_n117_), .Y(new_new_n733_));
  AN2        g0711(.A(new_new_n733_), .B(new_new_n591_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n242_), .B(new_new_n44_), .Y(new_new_n735_));
  NO3        g0713(.A(new_new_n735_), .B(new_new_n326_), .C(new_new_n247_), .Y(new_new_n736_));
  NO2        g0714(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n737_));
  NO2        g0715(.A(new_new_n737_), .B(i_6_), .Y(new_new_n738_));
  NO2        g0716(.A(new_new_n86_), .B(i_9_), .Y(new_new_n739_));
  NO2        g0717(.A(new_new_n739_), .B(new_new_n63_), .Y(new_new_n740_));
  NO2        g0718(.A(new_new_n740_), .B(new_new_n698_), .Y(new_new_n741_));
  NO4        g0719(.A(new_new_n741_), .B(new_new_n738_), .C(new_new_n736_), .D(i_4_), .Y(new_new_n742_));
  NA2        g0720(.A(i_1_), .B(i_3_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n492_), .B(new_new_n94_), .Y(new_new_n744_));
  AOI210     g0722(.A0(new_new_n735_), .A1(new_new_n627_), .B0(new_new_n744_), .Y(new_new_n745_));
  NO2        g0723(.A(new_new_n745_), .B(new_new_n743_), .Y(new_new_n746_));
  NO3        g0724(.A(new_new_n746_), .B(new_new_n742_), .C(new_new_n734_), .Y(new_new_n747_));
  NA4        g0725(.A(new_new_n747_), .B(new_new_n731_), .C(new_new_n725_), .D(new_new_n701_), .Y(new_new_n748_));
  NO3        g0726(.A(new_new_n518_), .B(i_3_), .C(i_7_), .Y(new_new_n749_));
  NOi21      g0727(.An(new_new_n749_), .B(i_10_), .Y(new_new_n750_));
  OA210      g0728(.A0(new_new_n750_), .A1(new_new_n255_), .B0(new_new_n86_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n398_), .B(new_new_n397_), .Y(new_new_n752_));
  NA3        g0730(.A(new_new_n525_), .B(new_new_n565_), .C(new_new_n46_), .Y(new_new_n753_));
  NO3        g0731(.A(new_new_n519_), .B(new_new_n667_), .C(new_new_n86_), .Y(new_new_n754_));
  NA2        g0732(.A(new_new_n754_), .B(new_new_n25_), .Y(new_new_n755_));
  NA3        g0733(.A(new_new_n164_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n756_));
  NA4        g0734(.A(new_new_n756_), .B(new_new_n755_), .C(new_new_n753_), .D(new_new_n752_), .Y(new_new_n757_));
  OAI210     g0735(.A0(new_new_n757_), .A1(new_new_n751_), .B0(i_1_), .Y(new_new_n758_));
  AOI210     g0736(.A0(new_new_n280_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n396_), .B(i_2_), .Y(new_new_n760_));
  NA2        g0738(.A(new_new_n760_), .B(new_new_n759_), .Y(new_new_n761_));
  OAI210     g0739(.A0(new_new_n717_), .A1(new_new_n483_), .B0(new_new_n761_), .Y(new_new_n762_));
  INV        g0740(.A(new_new_n762_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n763_), .B(new_new_n758_), .Y(new_new_n764_));
  OR2        g0742(.A(i_11_), .B(i_7_), .Y(new_new_n765_));
  NA3        g0743(.A(new_new_n765_), .B(new_new_n108_), .C(new_new_n141_), .Y(new_new_n766_));
  AOI220     g0744(.A0(new_new_n510_), .A1(new_new_n164_), .B0(new_new_n485_), .B1(new_new_n141_), .Y(new_new_n767_));
  OAI210     g0745(.A0(new_new_n767_), .A1(new_new_n44_), .B0(new_new_n766_), .Y(new_new_n768_));
  AOI210     g0746(.A0(new_new_n713_), .A1(new_new_n54_), .B0(i_12_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n519_), .B(new_new_n24_), .Y(new_new_n770_));
  AOI220     g0748(.A0(new_new_n770_), .A1(new_new_n730_), .B0(new_new_n255_), .B1(new_new_n134_), .Y(new_new_n771_));
  OAI220     g0749(.A0(new_new_n771_), .A1(new_new_n40_), .B0(new_new_n1146_), .B1(new_new_n94_), .Y(new_new_n772_));
  AOI210     g0750(.A0(new_new_n768_), .A1(new_new_n353_), .B0(new_new_n772_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n117_), .B(new_new_n110_), .Y(new_new_n774_));
  AOI220     g0752(.A0(new_new_n774_), .A1(new_new_n72_), .B0(new_new_n414_), .B1(new_new_n714_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n775_), .B(new_new_n252_), .Y(new_new_n776_));
  AOI210     g0754(.A0(new_new_n483_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n777_));
  NOi31      g0755(.An(new_new_n777_), .B(new_new_n656_), .C(new_new_n44_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n713_), .B(new_new_n117_), .Y(new_new_n779_));
  INV        g0757(.A(new_new_n779_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n780_), .B(new_new_n71_), .Y(new_new_n781_));
  NO3        g0759(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n103_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n26_), .B(new_new_n198_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(i_7_), .Y(new_new_n784_));
  NO3        g0762(.A(new_new_n519_), .B(new_new_n246_), .C(new_new_n86_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n785_), .A1(new_new_n784_), .B0(new_new_n782_), .Y(new_new_n786_));
  AOI220     g0764(.A0(new_new_n414_), .A1(new_new_n714_), .B0(new_new_n93_), .B1(new_new_n104_), .Y(new_new_n787_));
  OAI220     g0765(.A0(new_new_n787_), .A1(new_new_n662_), .B0(new_new_n786_), .B1(new_new_n677_), .Y(new_new_n788_));
  NO4        g0766(.A(new_new_n788_), .B(new_new_n781_), .C(new_new_n778_), .D(new_new_n776_), .Y(new_new_n789_));
  OR2        g0767(.A(i_11_), .B(i_6_), .Y(new_new_n790_));
  NA3        g0768(.A(new_new_n661_), .B(new_new_n783_), .C(i_7_), .Y(new_new_n791_));
  AOI210     g0769(.A0(new_new_n791_), .A1(new_new_n780_), .B0(new_new_n790_), .Y(new_new_n792_));
  NA3        g0770(.A(new_new_n443_), .B(new_new_n666_), .C(new_new_n99_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n104_), .B(new_new_n783_), .Y(new_new_n794_));
  NAi21      g0772(.An(i_11_), .B(i_12_), .Y(new_new_n795_));
  NOi41      g0773(.An(new_new_n113_), .B(new_new_n795_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n796_));
  NO3        g0774(.A(new_new_n519_), .B(new_new_n639_), .C(new_new_n667_), .Y(new_new_n797_));
  AOI220     g0775(.A0(new_new_n797_), .A1(new_new_n330_), .B0(new_new_n796_), .B1(new_new_n794_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n798_), .B(new_new_n793_), .Y(new_new_n799_));
  OAI210     g0777(.A0(new_new_n799_), .A1(new_new_n792_), .B0(new_new_n63_), .Y(new_new_n800_));
  NO2        g0778(.A(i_2_), .B(i_12_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n395_), .B(new_new_n801_), .Y(new_new_n802_));
  NA2        g0780(.A(i_8_), .B(new_new_n25_), .Y(new_new_n803_));
  NO3        g0781(.A(new_new_n803_), .B(new_new_n412_), .C(new_new_n661_), .Y(new_new_n804_));
  OAI210     g0782(.A0(new_new_n804_), .A1(new_new_n397_), .B0(new_new_n395_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n131_), .B(i_2_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n806_), .B(new_new_n698_), .Y(new_new_n807_));
  NA3        g0785(.A(new_new_n807_), .B(new_new_n805_), .C(new_new_n802_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n808_), .B(new_new_n45_), .Y(new_new_n809_));
  NA4        g0787(.A(new_new_n809_), .B(new_new_n800_), .C(new_new_n789_), .D(new_new_n773_), .Y(new_new_n810_));
  OR4        g0788(.A(new_new_n810_), .B(new_new_n764_), .C(new_new_n748_), .D(new_new_n680_), .Y(men5));
  AOI210     g0789(.A0(new_new_n727_), .A1(new_new_n283_), .B0(new_new_n452_), .Y(new_new_n812_));
  NA3        g0790(.A(new_new_n24_), .B(new_new_n801_), .C(new_new_n110_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n89_), .B(new_new_n661_), .Y(new_new_n814_));
  NA3        g0792(.A(new_new_n814_), .B(new_new_n813_), .C(new_new_n812_), .Y(new_new_n815_));
  NO3        g0793(.A(i_11_), .B(new_new_n246_), .C(i_13_), .Y(new_new_n816_));
  NO2        g0794(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n817_));
  NA2        g0795(.A(i_12_), .B(i_8_), .Y(new_new_n818_));
  OAI210     g0796(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n818_), .Y(new_new_n819_));
  AOI220     g0797(.A0(new_new_n336_), .A1(new_new_n631_), .B0(new_new_n819_), .B1(new_new_n817_), .Y(new_new_n820_));
  INV        g0798(.A(new_new_n820_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n821_), .B(new_new_n815_), .Y(new_new_n822_));
  INV        g0800(.A(new_new_n175_), .Y(new_new_n823_));
  INV        g0801(.A(new_new_n255_), .Y(new_new_n824_));
  OAI210     g0802(.A0(new_new_n760_), .A1(new_new_n484_), .B0(new_new_n113_), .Y(new_new_n825_));
  AOI210     g0803(.A0(new_new_n825_), .A1(new_new_n824_), .B0(new_new_n823_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n492_), .B(new_new_n26_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n827_), .B(new_new_n454_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n828_), .B(i_2_), .Y(new_new_n829_));
  INV        g0807(.A(new_new_n829_), .Y(new_new_n830_));
  AOI210     g0808(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n450_), .Y(new_new_n831_));
  AOI210     g0809(.A0(new_new_n831_), .A1(new_new_n830_), .B0(new_new_n826_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n195_), .B(new_new_n128_), .Y(new_new_n833_));
  OAI210     g0811(.A0(new_new_n833_), .A1(new_new_n817_), .B0(i_2_), .Y(new_new_n834_));
  INV        g0812(.A(new_new_n176_), .Y(new_new_n835_));
  NO3        g0813(.A(new_new_n682_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n836_));
  AOI210     g0814(.A0(new_new_n835_), .A1(new_new_n89_), .B0(new_new_n836_), .Y(new_new_n837_));
  AOI210     g0815(.A0(new_new_n837_), .A1(new_new_n834_), .B0(new_new_n198_), .Y(new_new_n838_));
  NA2        g0816(.A(new_new_n205_), .B(new_new_n208_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n154_), .B(new_new_n657_), .Y(new_new_n840_));
  AOI210     g0818(.A0(new_new_n840_), .A1(new_new_n839_), .B0(new_new_n400_), .Y(new_new_n841_));
  AOI210     g0819(.A0(new_new_n215_), .A1(new_new_n150_), .B0(new_new_n565_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n842_), .B(new_new_n454_), .Y(new_new_n843_));
  NA3        g0821(.A(new_new_n103_), .B(new_new_n323_), .C(new_new_n42_), .Y(new_new_n844_));
  OAI210     g0822(.A0(new_new_n844_), .A1(i_11_), .B0(new_new_n843_), .Y(new_new_n845_));
  NO3        g0823(.A(new_new_n845_), .B(new_new_n841_), .C(new_new_n838_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n631_), .B(new_new_n28_), .Y(new_new_n847_));
  INV        g0825(.A(new_new_n290_), .Y(new_new_n848_));
  NA2        g0826(.A(new_new_n848_), .B(new_new_n847_), .Y(new_new_n849_));
  NO2        g0827(.A(new_new_n62_), .B(i_12_), .Y(new_new_n850_));
  INV        g0828(.A(new_new_n129_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n851_), .B(new_new_n657_), .Y(new_new_n852_));
  AOI220     g0830(.A0(new_new_n852_), .A1(new_new_n36_), .B0(new_new_n849_), .B1(new_new_n46_), .Y(new_new_n853_));
  NA4        g0831(.A(new_new_n853_), .B(new_new_n846_), .C(new_new_n832_), .D(new_new_n822_), .Y(men6));
  NO2        g0832(.A(new_new_n325_), .B(i_1_), .Y(new_new_n855_));
  NO2        g0833(.A(new_new_n190_), .B(new_new_n142_), .Y(new_new_n856_));
  OAI210     g0834(.A0(new_new_n856_), .A1(new_new_n855_), .B0(new_new_n806_), .Y(new_new_n857_));
  NA4        g0835(.A(new_new_n418_), .B(new_new_n524_), .C(new_new_n71_), .D(new_new_n103_), .Y(new_new_n858_));
  INV        g0836(.A(new_new_n858_), .Y(new_new_n859_));
  NO2        g0837(.A(new_new_n229_), .B(new_new_n529_), .Y(new_new_n860_));
  NO2        g0838(.A(i_11_), .B(i_9_), .Y(new_new_n861_));
  AO210      g0839(.A0(new_new_n858_), .A1(new_new_n857_), .B0(i_12_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n401_), .B(new_new_n356_), .Y(new_new_n863_));
  NA2        g0841(.A(new_new_n639_), .B(new_new_n63_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n750_), .B(new_new_n71_), .Y(new_new_n865_));
  NA4        g0843(.A(new_new_n688_), .B(new_new_n865_), .C(new_new_n864_), .D(new_new_n863_), .Y(new_new_n866_));
  INV        g0844(.A(new_new_n202_), .Y(new_new_n867_));
  AOI220     g0845(.A0(new_new_n867_), .A1(new_new_n861_), .B0(new_new_n866_), .B1(new_new_n73_), .Y(new_new_n868_));
  INV        g0846(.A(new_new_n347_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n75_), .B(new_new_n134_), .Y(new_new_n870_));
  INV        g0848(.A(new_new_n127_), .Y(new_new_n871_));
  NA2        g0849(.A(new_new_n871_), .B(new_new_n46_), .Y(new_new_n872_));
  AOI210     g0850(.A0(new_new_n872_), .A1(new_new_n870_), .B0(new_new_n869_), .Y(new_new_n873_));
  NO3        g0851(.A(new_new_n262_), .B(new_new_n135_), .C(i_9_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n874_), .B(new_new_n850_), .Y(new_new_n875_));
  AOI210     g0853(.A0(new_new_n875_), .A1(new_new_n563_), .B0(new_new_n190_), .Y(new_new_n876_));
  NO2        g0854(.A(new_new_n32_), .B(i_11_), .Y(new_new_n877_));
  NA3        g0855(.A(new_new_n877_), .B(new_new_n514_), .C(new_new_n418_), .Y(new_new_n878_));
  NAi32      g0856(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n879_));
  AOI210     g0857(.A0(new_new_n790_), .A1(new_new_n87_), .B0(new_new_n879_), .Y(new_new_n880_));
  OAI210     g0858(.A0(new_new_n749_), .A1(new_new_n619_), .B0(new_new_n618_), .Y(new_new_n881_));
  NAi31      g0859(.An(new_new_n880_), .B(new_new_n881_), .C(new_new_n878_), .Y(new_new_n882_));
  OR3        g0860(.A(new_new_n882_), .B(new_new_n876_), .C(new_new_n873_), .Y(new_new_n883_));
  NO2        g0861(.A(new_new_n765_), .B(i_2_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n885_));
  OAI210     g0863(.A0(new_new_n885_), .A1(new_new_n442_), .B0(new_new_n385_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n886_), .B(new_new_n884_), .Y(new_new_n887_));
  AO220      g0865(.A0(new_new_n384_), .A1(new_new_n374_), .B0(new_new_n426_), .B1(new_new_n657_), .Y(new_new_n888_));
  NA3        g0866(.A(new_new_n888_), .B(new_new_n267_), .C(i_7_), .Y(new_new_n889_));
  OR2        g0867(.A(new_new_n683_), .B(new_new_n484_), .Y(new_new_n890_));
  NA3        g0868(.A(new_new_n890_), .B(new_new_n149_), .C(new_new_n69_), .Y(new_new_n891_));
  OR2        g0869(.A(new_new_n536_), .B(new_new_n36_), .Y(new_new_n892_));
  NA4        g0870(.A(new_new_n892_), .B(new_new_n891_), .C(new_new_n889_), .D(new_new_n887_), .Y(new_new_n893_));
  OAI210     g0871(.A0(new_new_n704_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n894_));
  AOI220     g0872(.A0(new_new_n894_), .A1(new_new_n618_), .B0(new_new_n860_), .B1(new_new_n784_), .Y(new_new_n895_));
  NA3        g0873(.A(new_new_n400_), .B(new_new_n248_), .C(new_new_n149_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n426_), .B(new_new_n70_), .Y(new_new_n897_));
  NA4        g0875(.A(new_new_n897_), .B(new_new_n896_), .C(new_new_n895_), .D(new_new_n665_), .Y(new_new_n898_));
  AO210      g0876(.A0(new_new_n565_), .A1(new_new_n46_), .B0(new_new_n88_), .Y(new_new_n899_));
  NA2        g0877(.A(new_new_n899_), .B(new_new_n525_), .Y(new_new_n900_));
  AOI210     g0878(.A0(new_new_n484_), .A1(new_new_n482_), .B0(new_new_n617_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n673_), .B(new_new_n104_), .Y(new_new_n902_));
  OAI210     g0880(.A0(new_new_n902_), .A1(new_new_n114_), .B0(new_new_n441_), .Y(new_new_n903_));
  NA2        g0881(.A(new_new_n254_), .B(new_new_n46_), .Y(new_new_n904_));
  INV        g0882(.A(new_new_n646_), .Y(new_new_n905_));
  NA3        g0883(.A(new_new_n905_), .B(new_new_n347_), .C(i_7_), .Y(new_new_n906_));
  NA4        g0884(.A(new_new_n906_), .B(new_new_n903_), .C(new_new_n901_), .D(new_new_n900_), .Y(new_new_n907_));
  NO4        g0885(.A(new_new_n907_), .B(new_new_n898_), .C(new_new_n893_), .D(new_new_n883_), .Y(new_new_n908_));
  NA4        g0886(.A(new_new_n908_), .B(new_new_n868_), .C(new_new_n862_), .D(new_new_n408_), .Y(men3));
  NA2        g0887(.A(i_12_), .B(i_10_), .Y(new_new_n910_));
  NA2        g0888(.A(i_6_), .B(i_7_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n911_), .B(i_0_), .Y(new_new_n912_));
  NO2        g0890(.A(i_11_), .B(new_new_n246_), .Y(new_new_n913_));
  OAI210     g0891(.A0(new_new_n912_), .A1(new_new_n306_), .B0(new_new_n913_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n914_), .B(new_new_n198_), .Y(new_new_n915_));
  NO3        g0893(.A(new_new_n488_), .B(new_new_n91_), .C(new_new_n44_), .Y(new_new_n916_));
  OA210      g0894(.A0(new_new_n916_), .A1(new_new_n915_), .B0(new_new_n178_), .Y(new_new_n917_));
  NA3        g0895(.A(new_new_n896_), .B(new_new_n665_), .C(new_new_n399_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n918_), .B(new_new_n39_), .Y(new_new_n919_));
  NOi21      g0897(.An(new_new_n98_), .B(new_new_n828_), .Y(new_new_n920_));
  NO3        g0898(.A(new_new_n693_), .B(new_new_n492_), .C(new_new_n134_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n443_), .B(new_new_n45_), .Y(new_new_n922_));
  AN2        g0900(.A(new_new_n490_), .B(new_new_n55_), .Y(new_new_n923_));
  NO3        g0901(.A(new_new_n923_), .B(new_new_n921_), .C(new_new_n920_), .Y(new_new_n924_));
  AOI210     g0902(.A0(new_new_n924_), .A1(new_new_n919_), .B0(new_new_n48_), .Y(new_new_n925_));
  NO4        g0903(.A(new_new_n404_), .B(new_new_n411_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n190_), .B(new_new_n627_), .Y(new_new_n927_));
  NOi21      g0905(.An(new_new_n927_), .B(new_new_n926_), .Y(new_new_n928_));
  NA2        g0906(.A(new_new_n777_), .B(new_new_n739_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n354_), .B(new_new_n474_), .Y(new_new_n930_));
  OAI220     g0908(.A0(new_new_n930_), .A1(new_new_n929_), .B0(new_new_n928_), .B1(new_new_n63_), .Y(new_new_n931_));
  NOi21      g0909(.An(i_5_), .B(i_9_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n932_), .B(i_0_), .Y(new_new_n933_));
  AOI210     g0911(.A0(new_new_n280_), .A1(new_new_n516_), .B0(new_new_n754_), .Y(new_new_n934_));
  NO3        g0912(.A(new_new_n446_), .B(new_new_n280_), .C(new_new_n73_), .Y(new_new_n935_));
  NO2        g0913(.A(new_new_n179_), .B(new_new_n150_), .Y(new_new_n936_));
  AOI210     g0914(.A0(new_new_n936_), .A1(new_new_n254_), .B0(new_new_n935_), .Y(new_new_n937_));
  OAI220     g0915(.A0(new_new_n937_), .A1(new_new_n185_), .B0(new_new_n934_), .B1(new_new_n933_), .Y(new_new_n938_));
  NO4        g0916(.A(new_new_n938_), .B(new_new_n931_), .C(new_new_n925_), .D(new_new_n917_), .Y(new_new_n939_));
  NA2        g0917(.A(new_new_n190_), .B(new_new_n24_), .Y(new_new_n940_));
  NO2        g0918(.A(new_new_n737_), .B(new_new_n654_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n941_), .B(new_new_n940_), .Y(new_new_n942_));
  NA2        g0920(.A(new_new_n330_), .B(new_new_n132_), .Y(new_new_n943_));
  NAi21      g0921(.An(new_new_n165_), .B(new_new_n474_), .Y(new_new_n944_));
  OAI220     g0922(.A0(new_new_n944_), .A1(new_new_n904_), .B0(new_new_n943_), .B1(new_new_n432_), .Y(new_new_n945_));
  NO2        g0923(.A(new_new_n945_), .B(new_new_n942_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n418_), .B(new_new_n310_), .Y(new_new_n947_));
  NA2        g0925(.A(new_new_n947_), .B(new_new_n779_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n628_), .B(i_0_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n949_), .B(new_new_n413_), .C(new_new_n89_), .Y(new_new_n950_));
  NO4        g0928(.A(new_new_n645_), .B(new_new_n223_), .C(new_new_n450_), .D(new_new_n442_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n951_), .A1(i_11_), .B0(new_new_n950_), .Y(new_new_n952_));
  INV        g0930(.A(new_new_n514_), .Y(new_new_n953_));
  AN2        g0931(.A(new_new_n98_), .B(new_new_n253_), .Y(new_new_n954_));
  NA2        g0932(.A(new_new_n816_), .B(new_new_n348_), .Y(new_new_n955_));
  AOI210     g0933(.A0(new_new_n525_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n956_));
  OAI220     g0934(.A0(new_new_n956_), .A1(new_new_n955_), .B0(new_new_n722_), .B1(new_new_n587_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n264_), .B(new_new_n156_), .Y(new_new_n958_));
  NA2        g0936(.A(i_0_), .B(i_10_), .Y(new_new_n959_));
  NO4        g0937(.A(new_new_n117_), .B(new_new_n58_), .C(new_new_n732_), .D(i_5_), .Y(new_new_n960_));
  AO220      g0938(.A0(new_new_n960_), .A1(i_10_), .B0(new_new_n958_), .B1(i_6_), .Y(new_new_n961_));
  AOI220     g0939(.A0(new_new_n354_), .A1(new_new_n100_), .B0(new_new_n190_), .B1(new_new_n84_), .Y(new_new_n962_));
  NA2        g0940(.A(new_new_n622_), .B(i_4_), .Y(new_new_n963_));
  NA2        g0941(.A(new_new_n193_), .B(new_new_n208_), .Y(new_new_n964_));
  OAI220     g0942(.A0(new_new_n964_), .A1(new_new_n955_), .B0(new_new_n963_), .B1(new_new_n962_), .Y(new_new_n965_));
  NO4        g0943(.A(new_new_n965_), .B(new_new_n961_), .C(new_new_n957_), .D(new_new_n954_), .Y(new_new_n966_));
  NA4        g0944(.A(new_new_n966_), .B(new_new_n952_), .C(new_new_n948_), .D(new_new_n946_), .Y(new_new_n967_));
  NO2        g0945(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n968_));
  NA2        g0946(.A(i_11_), .B(i_9_), .Y(new_new_n969_));
  NO3        g0947(.A(i_12_), .B(new_new_n969_), .C(new_new_n664_), .Y(new_new_n970_));
  AO220      g0948(.A0(new_new_n970_), .A1(new_new_n968_), .B0(new_new_n282_), .B1(new_new_n88_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n48_), .B(i_7_), .Y(new_new_n972_));
  NAi31      g0950(.An(new_new_n277_), .B(new_new_n497_), .C(new_new_n163_), .Y(new_new_n973_));
  NO2        g0951(.A(new_new_n969_), .B(new_new_n73_), .Y(new_new_n974_));
  NO2        g0952(.A(new_new_n179_), .B(i_0_), .Y(new_new_n975_));
  INV        g0953(.A(new_new_n975_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n514_), .B(new_new_n240_), .Y(new_new_n977_));
  AOI210     g0955(.A0(new_new_n398_), .A1(new_new_n41_), .B0(new_new_n440_), .Y(new_new_n978_));
  OAI220     g0956(.A0(new_new_n978_), .A1(new_new_n933_), .B0(new_new_n977_), .B1(new_new_n976_), .Y(new_new_n979_));
  NO3        g0957(.A(new_new_n979_), .B(new_new_n973_), .C(new_new_n971_), .Y(new_new_n980_));
  AOI210     g0958(.A0(new_new_n483_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n175_), .B(new_new_n105_), .Y(new_new_n982_));
  NOi32      g0960(.An(new_new_n981_), .Bn(new_new_n193_), .C(new_new_n982_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n666_), .A1(new_new_n348_), .B0(new_new_n253_), .Y(new_new_n984_));
  NO2        g0962(.A(new_new_n984_), .B(new_new_n922_), .Y(new_new_n985_));
  NO2        g0963(.A(new_new_n985_), .B(new_new_n983_), .Y(new_new_n986_));
  NOi21      g0964(.An(i_7_), .B(i_5_), .Y(new_new_n987_));
  NOi31      g0965(.An(new_new_n987_), .B(i_0_), .C(new_new_n795_), .Y(new_new_n988_));
  NA3        g0966(.A(new_new_n988_), .B(new_new_n412_), .C(i_6_), .Y(new_new_n989_));
  OA210      g0967(.A0(new_new_n982_), .A1(new_new_n563_), .B0(new_new_n989_), .Y(new_new_n990_));
  NO3        g0968(.A(new_new_n435_), .B(new_new_n387_), .C(new_new_n383_), .Y(new_new_n991_));
  NO2        g0969(.A(new_new_n274_), .B(new_new_n337_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n795_), .B(new_new_n269_), .Y(new_new_n993_));
  AOI210     g0971(.A0(new_new_n993_), .A1(new_new_n992_), .B0(new_new_n991_), .Y(new_new_n994_));
  NA4        g0972(.A(new_new_n994_), .B(new_new_n990_), .C(new_new_n986_), .D(new_new_n980_), .Y(new_new_n995_));
  NO2        g0973(.A(new_new_n940_), .B(new_new_n249_), .Y(new_new_n996_));
  AN2        g0974(.A(new_new_n353_), .B(new_new_n348_), .Y(new_new_n997_));
  AO220      g0975(.A0(new_new_n997_), .A1(new_new_n936_), .B0(new_new_n369_), .B1(new_new_n27_), .Y(new_new_n998_));
  OAI210     g0976(.A0(new_new_n998_), .A1(new_new_n996_), .B0(i_10_), .Y(new_new_n999_));
  NO2        g0977(.A(new_new_n910_), .B(new_new_n336_), .Y(new_new_n1000_));
  OA210      g0978(.A0(new_new_n514_), .A1(new_new_n232_), .B0(new_new_n513_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n1000_), .B(new_new_n974_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n513_), .B(new_new_n443_), .C(new_new_n45_), .Y(new_new_n1003_));
  OAI210     g0981(.A0(new_new_n944_), .A1(new_new_n953_), .B0(new_new_n1003_), .Y(new_new_n1004_));
  NO2        g0982(.A(new_new_n267_), .B(new_new_n46_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n974_), .B(new_new_n323_), .Y(new_new_n1006_));
  OAI210     g0984(.A0(new_new_n1005_), .A1(new_new_n192_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  AOI220     g0985(.A0(new_new_n1007_), .A1(new_new_n514_), .B0(new_new_n1004_), .B1(new_new_n73_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n885_), .B(new_new_n410_), .C(new_new_n704_), .Y(new_new_n1009_));
  NA2        g0987(.A(new_new_n94_), .B(new_new_n44_), .Y(new_new_n1010_));
  NO2        g0988(.A(new_new_n75_), .B(new_new_n818_), .Y(new_new_n1011_));
  AOI220     g0989(.A0(new_new_n1011_), .A1(new_new_n1010_), .B0(new_new_n178_), .B1(new_new_n654_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1012_), .A1(new_new_n1009_), .B0(new_new_n47_), .Y(new_new_n1013_));
  NO3        g0991(.A(new_new_n645_), .B(new_new_n382_), .C(new_new_n24_), .Y(new_new_n1014_));
  AOI210     g0992(.A0(new_new_n770_), .A1(new_new_n599_), .B0(new_new_n1014_), .Y(new_new_n1015_));
  NAi21      g0993(.An(i_9_), .B(i_5_), .Y(new_new_n1016_));
  NO2        g0994(.A(new_new_n1016_), .B(new_new_n435_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n660_), .B(new_new_n107_), .Y(new_new_n1018_));
  AOI220     g0996(.A0(new_new_n1018_), .A1(i_0_), .B0(new_new_n1017_), .B1(new_new_n683_), .Y(new_new_n1019_));
  OAI220     g0997(.A0(new_new_n1019_), .A1(new_new_n86_), .B0(new_new_n1015_), .B1(new_new_n176_), .Y(new_new_n1020_));
  NO3        g0998(.A(new_new_n1020_), .B(new_new_n1013_), .C(new_new_n567_), .Y(new_new_n1021_));
  NA4        g0999(.A(new_new_n1021_), .B(new_new_n1008_), .C(new_new_n1002_), .D(new_new_n999_), .Y(new_new_n1022_));
  NO3        g1000(.A(new_new_n1022_), .B(new_new_n995_), .C(new_new_n967_), .Y(new_new_n1023_));
  NO2        g1001(.A(i_0_), .B(new_new_n795_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n73_), .B(new_new_n44_), .Y(new_new_n1025_));
  NA2        g1003(.A(new_new_n959_), .B(new_new_n1025_), .Y(new_new_n1026_));
  NO3        g1004(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n1027_));
  AO220      g1005(.A0(new_new_n1027_), .A1(new_new_n1026_), .B0(new_new_n1024_), .B1(new_new_n178_), .Y(new_new_n1028_));
  AOI210     g1006(.A0(new_new_n864_), .A1(new_new_n752_), .B0(new_new_n982_), .Y(new_new_n1029_));
  AOI210     g1007(.A0(new_new_n1028_), .A1(new_new_n371_), .B0(new_new_n1029_), .Y(new_new_n1030_));
  NA2        g1008(.A(new_new_n806_), .B(new_new_n148_), .Y(new_new_n1031_));
  INV        g1009(.A(new_new_n1031_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n1032_), .B(new_new_n739_), .C(new_new_n73_), .Y(new_new_n1033_));
  NO2        g1011(.A(new_new_n881_), .B(new_new_n435_), .Y(new_new_n1034_));
  NA3        g1012(.A(new_new_n912_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n1035_));
  NA2        g1013(.A(new_new_n913_), .B(i_9_), .Y(new_new_n1036_));
  AOI210     g1014(.A0(new_new_n1035_), .A1(new_new_n542_), .B0(new_new_n1036_), .Y(new_new_n1037_));
  OAI210     g1015(.A0(new_new_n254_), .A1(i_9_), .B0(new_new_n239_), .Y(new_new_n1038_));
  AOI210     g1016(.A0(new_new_n1038_), .A1(new_new_n949_), .B0(new_new_n156_), .Y(new_new_n1039_));
  NO3        g1017(.A(new_new_n1039_), .B(new_new_n1037_), .C(new_new_n1034_), .Y(new_new_n1040_));
  NA3        g1018(.A(new_new_n1040_), .B(new_new_n1033_), .C(new_new_n1030_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n997_), .B(new_new_n400_), .Y(new_new_n1042_));
  AOI210     g1020(.A0(new_new_n317_), .A1(new_new_n165_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  NA3        g1021(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n1044_));
  NA2        g1022(.A(new_new_n972_), .B(new_new_n530_), .Y(new_new_n1045_));
  AOI210     g1023(.A0(new_new_n1044_), .A1(new_new_n165_), .B0(new_new_n1045_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n1046_), .B(new_new_n1043_), .Y(new_new_n1047_));
  NO2        g1025(.A(new_new_n959_), .B(new_new_n195_), .Y(new_new_n1048_));
  AOI220     g1026(.A0(new_new_n1048_), .A1(i_11_), .B0(new_new_n623_), .B1(new_new_n75_), .Y(new_new_n1049_));
  INV        g1027(.A(new_new_n226_), .Y(new_new_n1050_));
  OAI220     g1028(.A0(new_new_n580_), .A1(new_new_n142_), .B0(new_new_n708_), .B1(new_new_n677_), .Y(new_new_n1051_));
  NA3        g1029(.A(new_new_n1051_), .B(new_new_n427_), .C(new_new_n1050_), .Y(new_new_n1052_));
  NA3        g1030(.A(new_new_n1052_), .B(new_new_n1049_), .C(new_new_n1047_), .Y(new_new_n1053_));
  NO2        g1031(.A(new_new_n252_), .B(new_new_n94_), .Y(new_new_n1054_));
  AOI210     g1032(.A0(new_new_n1054_), .A1(new_new_n1024_), .B0(new_new_n111_), .Y(new_new_n1055_));
  AOI220     g1033(.A0(new_new_n987_), .A1(new_new_n530_), .B0(new_new_n912_), .B1(new_new_n166_), .Y(new_new_n1056_));
  NA2        g1034(.A(new_new_n374_), .B(new_new_n180_), .Y(new_new_n1057_));
  OA220      g1035(.A0(new_new_n1057_), .A1(new_new_n1056_), .B0(new_new_n1055_), .B1(i_5_), .Y(new_new_n1058_));
  AOI210     g1036(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n1059_));
  NA2        g1037(.A(new_new_n1059_), .B(new_new_n1001_), .Y(new_new_n1060_));
  NA3        g1038(.A(new_new_n674_), .B(new_new_n190_), .C(new_new_n84_), .Y(new_new_n1061_));
  NA2        g1039(.A(new_new_n1061_), .B(new_new_n597_), .Y(new_new_n1062_));
  NO3        g1040(.A(new_new_n922_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n1063_));
  NA3        g1041(.A(new_new_n535_), .B(new_new_n528_), .C(new_new_n511_), .Y(new_new_n1064_));
  NO3        g1042(.A(new_new_n1064_), .B(new_new_n1063_), .C(new_new_n1062_), .Y(new_new_n1065_));
  NA3        g1043(.A(new_new_n418_), .B(new_new_n175_), .C(new_new_n174_), .Y(new_new_n1066_));
  NA3        g1044(.A(new_new_n972_), .B(new_new_n306_), .C(new_new_n239_), .Y(new_new_n1067_));
  NA2        g1045(.A(new_new_n1067_), .B(new_new_n1066_), .Y(new_new_n1068_));
  NA3        g1046(.A(new_new_n418_), .B(new_new_n355_), .C(new_new_n230_), .Y(new_new_n1069_));
  INV        g1047(.A(new_new_n1069_), .Y(new_new_n1070_));
  NOi31      g1048(.An(new_new_n417_), .B(new_new_n1025_), .C(new_new_n249_), .Y(new_new_n1071_));
  NO2        g1049(.A(new_new_n969_), .B(new_new_n195_), .Y(new_new_n1072_));
  NO4        g1050(.A(new_new_n1072_), .B(new_new_n1071_), .C(new_new_n1070_), .D(new_new_n1068_), .Y(new_new_n1073_));
  NA4        g1051(.A(new_new_n1073_), .B(new_new_n1065_), .C(new_new_n1060_), .D(new_new_n1058_), .Y(new_new_n1074_));
  AOI210     g1052(.A0(new_new_n622_), .A1(new_new_n579_), .B0(new_new_n676_), .Y(new_new_n1075_));
  NO3        g1053(.A(new_new_n1075_), .B(new_new_n613_), .C(new_new_n368_), .Y(new_new_n1076_));
  NO2        g1054(.A(new_new_n86_), .B(i_5_), .Y(new_new_n1077_));
  NA3        g1055(.A(new_new_n913_), .B(new_new_n112_), .C(new_new_n127_), .Y(new_new_n1078_));
  INV        g1056(.A(new_new_n1078_), .Y(new_new_n1079_));
  AOI210     g1057(.A0(new_new_n1079_), .A1(new_new_n1077_), .B0(new_new_n1076_), .Y(new_new_n1080_));
  NA3        g1058(.A(new_new_n323_), .B(i_5_), .C(new_new_n198_), .Y(new_new_n1081_));
  NAi31      g1059(.An(new_new_n251_), .B(new_new_n1081_), .C(new_new_n252_), .Y(new_new_n1082_));
  NO4        g1060(.A(new_new_n249_), .B(new_new_n217_), .C(i_0_), .D(i_12_), .Y(new_new_n1083_));
  AOI220     g1061(.A0(new_new_n1083_), .A1(new_new_n1082_), .B0(new_new_n859_), .B1(new_new_n180_), .Y(new_new_n1084_));
  AN2        g1062(.A(new_new_n959_), .B(new_new_n156_), .Y(new_new_n1085_));
  NO4        g1063(.A(new_new_n1085_), .B(i_12_), .C(new_new_n712_), .D(new_new_n134_), .Y(new_new_n1086_));
  NA2        g1064(.A(new_new_n1086_), .B(new_new_n226_), .Y(new_new_n1087_));
  NA3        g1065(.A(new_new_n100_), .B(new_new_n627_), .C(i_11_), .Y(new_new_n1088_));
  NO2        g1066(.A(new_new_n1088_), .B(new_new_n158_), .Y(new_new_n1089_));
  NA2        g1067(.A(new_new_n987_), .B(new_new_n510_), .Y(new_new_n1090_));
  NA2        g1068(.A(new_new_n64_), .B(new_new_n103_), .Y(new_new_n1091_));
  OAI220     g1069(.A0(new_new_n1091_), .A1(new_new_n1081_), .B0(new_new_n1090_), .B1(new_new_n740_), .Y(new_new_n1092_));
  AOI210     g1070(.A0(new_new_n1092_), .A1(new_new_n975_), .B0(new_new_n1089_), .Y(new_new_n1093_));
  NA4        g1071(.A(new_new_n1093_), .B(new_new_n1087_), .C(new_new_n1084_), .D(new_new_n1080_), .Y(new_new_n1094_));
  NO4        g1072(.A(new_new_n1094_), .B(new_new_n1074_), .C(new_new_n1053_), .D(new_new_n1041_), .Y(new_new_n1095_));
  OAI210     g1073(.A0(new_new_n884_), .A1(new_new_n877_), .B0(new_new_n37_), .Y(new_new_n1096_));
  NA3        g1074(.A(new_new_n981_), .B(new_new_n395_), .C(i_5_), .Y(new_new_n1097_));
  NA3        g1075(.A(new_new_n1097_), .B(new_new_n1096_), .C(new_new_n672_), .Y(new_new_n1098_));
  NA2        g1076(.A(new_new_n1098_), .B(new_new_n213_), .Y(new_new_n1099_));
  AN2        g1077(.A(new_new_n765_), .B(new_new_n396_), .Y(new_new_n1100_));
  NA2        g1078(.A(new_new_n191_), .B(new_new_n193_), .Y(new_new_n1101_));
  AO210      g1079(.A0(new_new_n1100_), .A1(new_new_n33_), .B0(new_new_n1101_), .Y(new_new_n1102_));
  OAI210     g1080(.A0(new_new_n676_), .A1(new_new_n674_), .B0(new_new_n336_), .Y(new_new_n1103_));
  NAi31      g1081(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1104_));
  NO2        g1082(.A(new_new_n70_), .B(new_new_n1104_), .Y(new_new_n1105_));
  NO2        g1083(.A(new_new_n1105_), .B(new_new_n709_), .Y(new_new_n1106_));
  NA3        g1084(.A(new_new_n1106_), .B(new_new_n1103_), .C(new_new_n1102_), .Y(new_new_n1107_));
  NO2        g1085(.A(new_new_n500_), .B(new_new_n280_), .Y(new_new_n1108_));
  NO4        g1086(.A(new_new_n242_), .B(new_new_n147_), .C(new_new_n743_), .D(new_new_n37_), .Y(new_new_n1109_));
  NO3        g1087(.A(new_new_n1109_), .B(new_new_n1108_), .C(new_new_n951_), .Y(new_new_n1110_));
  OAI210     g1088(.A0(new_new_n1088_), .A1(new_new_n150_), .B0(new_new_n1110_), .Y(new_new_n1111_));
  AOI210     g1089(.A0(new_new_n1107_), .A1(new_new_n48_), .B0(new_new_n1111_), .Y(new_new_n1112_));
  AOI210     g1090(.A0(new_new_n1112_), .A1(new_new_n1099_), .B0(new_new_n73_), .Y(new_new_n1113_));
  NO2        g1091(.A(new_new_n620_), .B(new_new_n407_), .Y(new_new_n1114_));
  NO2        g1092(.A(new_new_n1114_), .B(new_new_n823_), .Y(new_new_n1115_));
  OAI210     g1093(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n110_), .Y(new_new_n1116_));
  NA2        g1094(.A(new_new_n1116_), .B(new_new_n76_), .Y(new_new_n1117_));
  AOI210     g1095(.A0(new_new_n1059_), .A1(new_new_n972_), .B0(new_new_n988_), .Y(new_new_n1118_));
  AOI210     g1096(.A0(new_new_n1118_), .A1(new_new_n1117_), .B0(new_new_n743_), .Y(new_new_n1119_));
  NA2        g1097(.A(new_new_n274_), .B(new_new_n57_), .Y(new_new_n1120_));
  AOI220     g1098(.A0(new_new_n1120_), .A1(new_new_n76_), .B0(new_new_n369_), .B1(new_new_n266_), .Y(new_new_n1121_));
  NO2        g1099(.A(new_new_n1121_), .B(new_new_n246_), .Y(new_new_n1122_));
  NA3        g1100(.A(new_new_n98_), .B(new_new_n325_), .C(new_new_n31_), .Y(new_new_n1123_));
  INV        g1101(.A(new_new_n1123_), .Y(new_new_n1124_));
  NO3        g1102(.A(new_new_n1124_), .B(new_new_n1122_), .C(new_new_n1119_), .Y(new_new_n1125_));
  OAI210     g1103(.A0(new_new_n282_), .A1(new_new_n161_), .B0(new_new_n89_), .Y(new_new_n1126_));
  NA3        g1104(.A(new_new_n827_), .B(new_new_n306_), .C(new_new_n80_), .Y(new_new_n1127_));
  AOI210     g1105(.A0(new_new_n1127_), .A1(new_new_n1126_), .B0(i_11_), .Y(new_new_n1128_));
  NA2        g1106(.A(new_new_n667_), .B(new_new_n223_), .Y(new_new_n1129_));
  OAI210     g1107(.A0(new_new_n1129_), .A1(new_new_n981_), .B0(new_new_n213_), .Y(new_new_n1130_));
  NA2        g1108(.A(new_new_n167_), .B(i_5_), .Y(new_new_n1131_));
  AOI210     g1109(.A0(new_new_n1130_), .A1(new_new_n839_), .B0(new_new_n1131_), .Y(new_new_n1132_));
  NO3        g1110(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1133_));
  OAI210     g1111(.A0(new_new_n992_), .A1(new_new_n325_), .B0(new_new_n1133_), .Y(new_new_n1134_));
  NO2        g1112(.A(new_new_n1134_), .B(new_new_n795_), .Y(new_new_n1135_));
  NO4        g1113(.A(new_new_n1016_), .B(new_new_n518_), .C(new_new_n263_), .D(new_new_n262_), .Y(new_new_n1136_));
  NO2        g1114(.A(new_new_n1136_), .B(new_new_n617_), .Y(new_new_n1137_));
  NO2        g1115(.A(new_new_n880_), .B(new_new_n388_), .Y(new_new_n1138_));
  AOI210     g1116(.A0(new_new_n1138_), .A1(new_new_n1137_), .B0(new_new_n40_), .Y(new_new_n1139_));
  NO4        g1117(.A(new_new_n1139_), .B(new_new_n1135_), .C(new_new_n1132_), .D(new_new_n1128_), .Y(new_new_n1140_));
  OAI210     g1118(.A0(new_new_n1125_), .A1(i_4_), .B0(new_new_n1140_), .Y(new_new_n1141_));
  NO3        g1119(.A(new_new_n1141_), .B(new_new_n1115_), .C(new_new_n1113_), .Y(new_new_n1142_));
  NA4        g1120(.A(new_new_n1142_), .B(new_new_n1095_), .C(new_new_n1023_), .D(new_new_n939_), .Y(men4));
  INV        g1121(.A(new_new_n769_), .Y(new_new_n1146_));
  INV        g1122(.A(i_5_), .Y(new_new_n1147_));
endmodule


