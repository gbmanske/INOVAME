//Benchmark atmr_intb_466_0.0156

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n363_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n421_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n383_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n387_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n458_, men_men_n459_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  INV        o039(.A(ori_ori_n59_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(ori_ori_n24_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .Y(ori_ori_n65_));
  NA2        o043(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n66_));
  OAI210     o044(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n66_), .Y(ori_ori_n67_));
  AOI220     o045(.A0(ori_ori_n67_), .A1(ori_ori_n59_), .B0(ori_ori_n65_), .B1(ori_ori_n31_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n61_), .B(ori_ori_n23_), .Y(ori_ori_n70_));
  NA2        o048(.A(x09), .B(x05), .Y(ori_ori_n71_));
  NA2        o049(.A(x10), .B(x06), .Y(ori_ori_n72_));
  NA3        o050(.A(ori_ori_n72_), .B(ori_ori_n71_), .C(ori_ori_n28_), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n73_), .A1(ori_ori_n70_), .B0(x03), .Y(ori_ori_n75_));
  NOi31      o053(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n76_));
  INV        o054(.A(x07), .Y(ori_ori_n77_));
  NO2        o055(.A(ori_ori_n77_), .B(ori_ori_n24_), .Y(ori_ori_n78_));
  NO2        o056(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n36_), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n79_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n81_));
  AOI210     o059(.A0(ori_ori_n80_), .A1(ori_ori_n48_), .B0(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n83_));
  NO2        o061(.A(x08), .B(x01), .Y(ori_ori_n84_));
  OAI210     o062(.A0(ori_ori_n84_), .A1(ori_ori_n83_), .B0(ori_ori_n35_), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n86_));
  NO3        o064(.A(ori_ori_n85_), .B(ori_ori_n82_), .C(ori_ori_n78_), .Y(ori_ori_n87_));
  AN2        o065(.A(ori_ori_n87_), .B(ori_ori_n75_), .Y(ori_ori_n88_));
  INV        o066(.A(ori_ori_n85_), .Y(ori_ori_n89_));
  NO2        o067(.A(x06), .B(x05), .Y(ori_ori_n90_));
  NA2        o068(.A(x11), .B(x00), .Y(ori_ori_n91_));
  NO2        o069(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n92_));
  NOi21      o070(.An(ori_ori_n91_), .B(ori_ori_n92_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NOi21      o072(.An(x01), .B(x10), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n96_));
  NO3        o074(.A(ori_ori_n96_), .B(ori_ori_n95_), .C(x06), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n97_), .B(ori_ori_n27_), .Y(ori_ori_n98_));
  OAI210     o076(.A0(ori_ori_n94_), .A1(x07), .B0(ori_ori_n98_), .Y(ori_ori_n99_));
  NO3        o077(.A(ori_ori_n99_), .B(ori_ori_n88_), .C(ori_ori_n69_), .Y(ori01));
  INV        o078(.A(x12), .Y(ori_ori_n101_));
  INV        o079(.A(x13), .Y(ori_ori_n102_));
  NA2        o080(.A(x08), .B(x04), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n95_), .B(ori_ori_n28_), .Y(ori_ori_n104_));
  NO2        o082(.A(x10), .B(x01), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n105_), .Y(ori_ori_n107_));
  NA2        o085(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n109_));
  NOi21      o087(.An(ori_ori_n109_), .B(ori_ori_n58_), .Y(ori_ori_n110_));
  INV        o088(.A(x13), .Y(ori_ori_n111_));
  NA2        o089(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n112_));
  NA2        o090(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(x05), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n115_));
  AOI210     o093(.A0(ori_ori_n57_), .A1(ori_ori_n80_), .B0(ori_ori_n110_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n72_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n118_));
  NA2        o096(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n122_));
  NA3        o100(.A(ori_ori_n122_), .B(ori_ori_n121_), .C(x13), .Y(ori_ori_n123_));
  NO2        o101(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n124_));
  NOi31      o102(.An(ori_ori_n123_), .B(ori_ori_n124_), .C(ori_ori_n120_), .Y(ori_ori_n125_));
  NO3        o103(.A(ori_ori_n125_), .B(x06), .C(x03), .Y(ori_ori_n126_));
  NO2        o104(.A(ori_ori_n126_), .B(ori_ori_n117_), .Y(ori_ori_n127_));
  NA2        o105(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n128_));
  OAI210     o106(.A0(ori_ori_n84_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  NO2        o108(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n132_));
  AOI210     o110(.A0(ori_ori_n132_), .A1(ori_ori_n49_), .B0(ori_ori_n131_), .Y(ori_ori_n133_));
  AN2        o111(.A(ori_ori_n133_), .B(ori_ori_n130_), .Y(ori_ori_n134_));
  NO2        o112(.A(x09), .B(x05), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n135_), .B(ori_ori_n47_), .Y(ori_ori_n136_));
  AOI210     o114(.A0(ori_ori_n136_), .A1(ori_ori_n107_), .B0(ori_ori_n49_), .Y(ori_ori_n137_));
  NA2        o115(.A(x09), .B(x00), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n109_), .B(ori_ori_n138_), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n139_), .B(ori_ori_n132_), .Y(ori_ori_n140_));
  NO3        o118(.A(ori_ori_n140_), .B(ori_ori_n137_), .C(ori_ori_n134_), .Y(ori_ori_n141_));
  NO2        o119(.A(x03), .B(x02), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n85_), .B(ori_ori_n102_), .Y(ori_ori_n143_));
  OAI210     o121(.A0(ori_ori_n143_), .A1(ori_ori_n110_), .B0(ori_ori_n142_), .Y(ori_ori_n144_));
  OA210      o122(.A0(ori_ori_n141_), .A1(x11), .B0(ori_ori_n144_), .Y(ori_ori_n145_));
  OAI210     o123(.A0(ori_ori_n127_), .A1(ori_ori_n23_), .B0(ori_ori_n145_), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n107_), .B(ori_ori_n40_), .Y(ori_ori_n147_));
  NAi21      o125(.An(x06), .B(x10), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n147_), .B(ori_ori_n41_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n150_));
  NA2        o128(.A(ori_ori_n102_), .B(x01), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n151_), .B(x08), .Y(ori_ori_n152_));
  OAI210     o130(.A0(x05), .A1(ori_ori_n152_), .B0(ori_ori_n51_), .Y(ori_ori_n153_));
  AOI210     o131(.A0(ori_ori_n153_), .A1(ori_ori_n150_), .B0(ori_ori_n48_), .Y(ori_ori_n154_));
  AOI210     o132(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n155_));
  OAI210     o133(.A0(ori_ori_n154_), .A1(ori_ori_n149_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o134(.A(x04), .B(x02), .Y(ori_ori_n157_));
  NA2        o135(.A(x10), .B(x05), .Y(ori_ori_n158_));
  NO2        o136(.A(x09), .B(x01), .Y(ori_ori_n159_));
  NO3        o137(.A(ori_ori_n159_), .B(ori_ori_n105_), .C(ori_ori_n31_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(x00), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n109_), .B(x08), .Y(ori_ori_n162_));
  INV        o140(.A(ori_ori_n161_), .Y(ori_ori_n163_));
  NAi21      o141(.An(ori_ori_n157_), .B(ori_ori_n163_), .Y(ori_ori_n164_));
  INV        o142(.A(ori_ori_n25_), .Y(ori_ori_n165_));
  NAi21      o143(.An(x13), .B(x00), .Y(ori_ori_n166_));
  AOI210     o144(.A0(ori_ori_n29_), .A1(ori_ori_n48_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  AOI220     o145(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(ori_ori_n168_));
  OAI210     o146(.A0(ori_ori_n158_), .A1(ori_ori_n35_), .B0(ori_ori_n168_), .Y(ori_ori_n169_));
  AN2        o147(.A(ori_ori_n169_), .B(ori_ori_n167_), .Y(ori_ori_n170_));
  AN2        o148(.A(ori_ori_n72_), .B(ori_ori_n71_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n96_), .B(x06), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n166_), .B(ori_ori_n36_), .Y(ori_ori_n173_));
  INV        o151(.A(ori_ori_n173_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n172_), .B(ori_ori_n171_), .Y(ori_ori_n175_));
  OAI210     o153(.A0(ori_ori_n175_), .A1(ori_ori_n170_), .B0(ori_ori_n165_), .Y(ori_ori_n176_));
  NOi21      o154(.An(x09), .B(x00), .Y(ori_ori_n177_));
  NO3        o155(.A(ori_ori_n83_), .B(ori_ori_n177_), .C(ori_ori_n47_), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n178_), .B(ori_ori_n119_), .Y(ori_ori_n179_));
  NA2        o157(.A(x10), .B(x08), .Y(ori_ori_n180_));
  INV        o158(.A(ori_ori_n180_), .Y(ori_ori_n181_));
  NA2        o159(.A(x06), .B(x05), .Y(ori_ori_n182_));
  OAI210     o160(.A0(ori_ori_n182_), .A1(ori_ori_n35_), .B0(ori_ori_n101_), .Y(ori_ori_n183_));
  AOI210     o161(.A0(ori_ori_n181_), .A1(ori_ori_n58_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n184_), .B(ori_ori_n179_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n102_), .B(x12), .Y(ori_ori_n186_));
  AOI210     o164(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n186_), .Y(ori_ori_n187_));
  NA2        o165(.A(ori_ori_n95_), .B(ori_ori_n51_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n189_), .B(x02), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n187_), .B(ori_ori_n185_), .Y(ori_ori_n191_));
  NA4        o169(.A(ori_ori_n191_), .B(ori_ori_n176_), .C(ori_ori_n164_), .D(ori_ori_n156_), .Y(ori_ori_n192_));
  AOI210     o170(.A0(ori_ori_n146_), .A1(ori_ori_n101_), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  INV        o171(.A(ori_ori_n73_), .Y(ori_ori_n194_));
  NA2        o172(.A(ori_ori_n194_), .B(ori_ori_n130_), .Y(ori_ori_n195_));
  NA2        o173(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n196_), .B(ori_ori_n129_), .Y(ori_ori_n197_));
  AOI210     o175(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n118_), .B(x06), .Y(ori_ori_n199_));
  AOI210     o177(.A0(ori_ori_n198_), .A1(ori_ori_n197_), .B0(ori_ori_n199_), .Y(ori_ori_n200_));
  AOI210     o178(.A0(ori_ori_n200_), .A1(ori_ori_n195_), .B0(x12), .Y(ori_ori_n201_));
  INV        o179(.A(ori_ori_n76_), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n95_), .B(x06), .Y(ori_ori_n203_));
  AOI210     o181(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n204_), .B(ori_ori_n203_), .C(ori_ori_n41_), .Y(ori_ori_n205_));
  INV        o183(.A(ori_ori_n132_), .Y(ori_ori_n206_));
  OAI210     o184(.A0(ori_ori_n206_), .A1(ori_ori_n205_), .B0(x02), .Y(ori_ori_n207_));
  AOI210     o185(.A0(ori_ori_n207_), .A1(ori_ori_n57_), .B0(ori_ori_n23_), .Y(ori_ori_n208_));
  OAI210     o186(.A0(ori_ori_n201_), .A1(ori_ori_n57_), .B0(ori_ori_n208_), .Y(ori_ori_n209_));
  INV        o187(.A(ori_ori_n132_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n211_));
  OAI210     o189(.A0(ori_ori_n79_), .A1(ori_ori_n36_), .B0(ori_ori_n112_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n102_), .B(x03), .Y(ori_ori_n213_));
  AOI220     o191(.A0(ori_ori_n213_), .A1(ori_ori_n212_), .B0(ori_ori_n76_), .B1(ori_ori_n211_), .Y(ori_ori_n214_));
  NA2        o192(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n215_));
  INV        o193(.A(ori_ori_n148_), .Y(ori_ori_n216_));
  NOi21      o194(.An(x13), .B(x04), .Y(ori_ori_n217_));
  NO3        o195(.A(ori_ori_n217_), .B(ori_ori_n76_), .C(ori_ori_n177_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n218_), .B(x05), .Y(ori_ori_n219_));
  AOI220     o197(.A0(ori_ori_n219_), .A1(ori_ori_n215_), .B0(ori_ori_n216_), .B1(ori_ori_n57_), .Y(ori_ori_n220_));
  OAI210     o198(.A0(ori_ori_n214_), .A1(ori_ori_n210_), .B0(ori_ori_n220_), .Y(ori_ori_n221_));
  INV        o199(.A(ori_ori_n92_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n222_), .B(x12), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n225_), .A1(ori_ori_n169_), .B0(ori_ori_n167_), .Y(ori_ori_n226_));
  AOI210     o204(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n227_));
  NO2        o205(.A(x06), .B(x00), .Y(ori_ori_n228_));
  NO3        o206(.A(ori_ori_n228_), .B(ori_ori_n227_), .C(ori_ori_n41_), .Y(ori_ori_n229_));
  OAI210     o207(.A0(ori_ori_n103_), .A1(ori_ori_n138_), .B0(ori_ori_n72_), .Y(ori_ori_n230_));
  NO2        o208(.A(ori_ori_n230_), .B(ori_ori_n229_), .Y(ori_ori_n231_));
  NA2        o209(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n232_), .B(x03), .Y(ori_ori_n233_));
  OA210      o211(.A0(ori_ori_n233_), .A1(ori_ori_n231_), .B0(ori_ori_n226_), .Y(ori_ori_n234_));
  NA2        o212(.A(x13), .B(ori_ori_n101_), .Y(ori_ori_n235_));
  NA3        o213(.A(ori_ori_n235_), .B(ori_ori_n183_), .C(ori_ori_n93_), .Y(ori_ori_n236_));
  OAI210     o214(.A0(ori_ori_n234_), .A1(ori_ori_n224_), .B0(ori_ori_n236_), .Y(ori_ori_n237_));
  AOI210     o215(.A0(ori_ori_n223_), .A1(ori_ori_n221_), .B0(ori_ori_n237_), .Y(ori_ori_n238_));
  AOI210     o216(.A0(ori_ori_n238_), .A1(ori_ori_n209_), .B0(x07), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n71_), .B(ori_ori_n29_), .Y(ori_ori_n240_));
  NOi31      o218(.An(ori_ori_n128_), .B(ori_ori_n217_), .C(ori_ori_n177_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n241_), .B(ori_ori_n240_), .Y(ori_ori_n242_));
  NO2        o220(.A(x08), .B(x05), .Y(ori_ori_n243_));
  INV        o221(.A(ori_ori_n227_), .Y(ori_ori_n244_));
  OAI210     o222(.A0(ori_ori_n76_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n245_));
  INV        o223(.A(ori_ori_n245_), .Y(ori_ori_n246_));
  NO2        o224(.A(x12), .B(x02), .Y(ori_ori_n247_));
  INV        o225(.A(ori_ori_n247_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n248_), .B(ori_ori_n222_), .Y(ori_ori_n249_));
  OA210      o227(.A0(ori_ori_n246_), .A1(ori_ori_n242_), .B0(ori_ori_n249_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n251_), .B(x01), .Y(ori_ori_n252_));
  NOi21      o230(.An(ori_ori_n84_), .B(ori_ori_n112_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n253_), .B(ori_ori_n252_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n254_), .A1(ori_ori_n123_), .B0(ori_ori_n29_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n102_), .B(x04), .Y(ori_ori_n256_));
  NO2        o234(.A(x02), .B(ori_ori_n111_), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n91_), .B(x12), .C(x03), .Y(ori_ori_n258_));
  OAI210     o236(.A0(ori_ori_n257_), .A1(ori_ori_n255_), .B0(ori_ori_n258_), .Y(ori_ori_n259_));
  AOI210     o237(.A0(ori_ori_n188_), .A1(ori_ori_n182_), .B0(ori_ori_n103_), .Y(ori_ori_n260_));
  NOi21      o238(.An(ori_ori_n240_), .B(ori_ori_n203_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n262_));
  OAI210     o240(.A0(ori_ori_n261_), .A1(ori_ori_n260_), .B0(ori_ori_n262_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n264_));
  NO3        o242(.A(ori_ori_n264_), .B(ori_ori_n204_), .C(ori_ori_n172_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n224_), .B(ori_ori_n28_), .Y(ori_ori_n266_));
  OAI210     o244(.A0(ori_ori_n265_), .A1(ori_ori_n210_), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  NA3        o245(.A(ori_ori_n267_), .B(ori_ori_n263_), .C(ori_ori_n259_), .Y(ori_ori_n268_));
  NO3        o246(.A(ori_ori_n268_), .B(ori_ori_n250_), .C(ori_ori_n239_), .Y(ori_ori_n269_));
  OAI210     o247(.A0(ori_ori_n193_), .A1(ori_ori_n61_), .B0(ori_ori_n269_), .Y(ori02));
  AOI210     o248(.A0(ori_ori_n128_), .A1(ori_ori_n85_), .B0(ori_ori_n121_), .Y(ori_ori_n271_));
  NOi21      o249(.An(ori_ori_n218_), .B(ori_ori_n159_), .Y(ori_ori_n272_));
  NO2        o250(.A(ori_ori_n102_), .B(ori_ori_n35_), .Y(ori_ori_n273_));
  NA3        o251(.A(ori_ori_n273_), .B(ori_ori_n181_), .C(ori_ori_n56_), .Y(ori_ori_n274_));
  OAI210     o252(.A0(ori_ori_n272_), .A1(ori_ori_n32_), .B0(ori_ori_n274_), .Y(ori_ori_n275_));
  OAI210     o253(.A0(ori_ori_n275_), .A1(ori_ori_n271_), .B0(ori_ori_n158_), .Y(ori_ori_n276_));
  INV        o254(.A(ori_ori_n158_), .Y(ori_ori_n277_));
  INV        o255(.A(ori_ori_n204_), .Y(ori_ori_n278_));
  OAI220     o256(.A0(ori_ori_n278_), .A1(ori_ori_n102_), .B0(ori_ori_n85_), .B1(ori_ori_n51_), .Y(ori_ori_n279_));
  AOI220     o257(.A0(ori_ori_n279_), .A1(ori_ori_n277_), .B0(ori_ori_n143_), .B1(ori_ori_n142_), .Y(ori_ori_n280_));
  AOI210     o258(.A0(ori_ori_n280_), .A1(ori_ori_n276_), .B0(ori_ori_n48_), .Y(ori_ori_n281_));
  NO2        o259(.A(x05), .B(x02), .Y(ori_ori_n282_));
  OAI210     o260(.A0(ori_ori_n197_), .A1(ori_ori_n177_), .B0(ori_ori_n282_), .Y(ori_ori_n283_));
  AOI220     o261(.A0(ori_ori_n243_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n284_));
  NOi21      o262(.An(ori_ori_n273_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  AOI210     o263(.A0(ori_ori_n217_), .A1(ori_ori_n79_), .B0(ori_ori_n285_), .Y(ori_ori_n286_));
  AOI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n283_), .B0(ori_ori_n132_), .Y(ori_ori_n287_));
  NAi21      o265(.An(ori_ori_n219_), .B(ori_ori_n214_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n232_), .B(ori_ori_n47_), .Y(ori_ori_n289_));
  NA2        o267(.A(ori_ori_n289_), .B(ori_ori_n288_), .Y(ori_ori_n290_));
  AN2        o268(.A(ori_ori_n213_), .B(ori_ori_n212_), .Y(ori_ori_n291_));
  OAI210     o269(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n292_));
  NA2        o270(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n293_));
  OA210      o271(.A0(ori_ori_n293_), .A1(x08), .B0(ori_ori_n136_), .Y(ori_ori_n294_));
  AOI210     o272(.A0(ori_ori_n294_), .A1(ori_ori_n129_), .B0(ori_ori_n292_), .Y(ori_ori_n295_));
  OAI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n291_), .B0(ori_ori_n96_), .Y(ori_ori_n296_));
  NA3        o274(.A(ori_ori_n96_), .B(ori_ori_n84_), .C(ori_ori_n211_), .Y(ori_ori_n297_));
  NA3        o275(.A(ori_ori_n95_), .B(ori_ori_n83_), .C(ori_ori_n42_), .Y(ori_ori_n298_));
  AOI210     o276(.A0(ori_ori_n298_), .A1(ori_ori_n297_), .B0(x04), .Y(ori_ori_n299_));
  INV        o277(.A(ori_ori_n142_), .Y(ori_ori_n300_));
  OAI220     o278(.A0(ori_ori_n244_), .A1(ori_ori_n104_), .B0(ori_ori_n300_), .B1(ori_ori_n120_), .Y(ori_ori_n301_));
  AOI210     o279(.A0(ori_ori_n301_), .A1(x13), .B0(ori_ori_n299_), .Y(ori_ori_n302_));
  NA3        o280(.A(ori_ori_n302_), .B(ori_ori_n296_), .C(ori_ori_n290_), .Y(ori_ori_n303_));
  NO3        o281(.A(ori_ori_n303_), .B(ori_ori_n287_), .C(ori_ori_n281_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n131_), .B(x03), .Y(ori_ori_n305_));
  INV        o283(.A(ori_ori_n166_), .Y(ori_ori_n306_));
  AOI220     o284(.A0(x08), .A1(ori_ori_n306_), .B0(ori_ori_n189_), .B1(x08), .Y(ori_ori_n307_));
  OAI210     o285(.A0(ori_ori_n307_), .A1(ori_ori_n264_), .B0(ori_ori_n305_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n308_), .B(ori_ori_n105_), .Y(ori_ori_n309_));
  NA2        o287(.A(ori_ori_n157_), .B(ori_ori_n151_), .Y(ori_ori_n310_));
  AN2        o288(.A(ori_ori_n310_), .B(ori_ori_n162_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n121_), .B(ori_ori_n28_), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n311_), .B0(ori_ori_n106_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n256_), .B(ori_ori_n101_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n101_), .B(ori_ori_n41_), .Y(ori_ori_n315_));
  NA3        o293(.A(ori_ori_n315_), .B(ori_ori_n314_), .C(ori_ori_n120_), .Y(ori_ori_n316_));
  NA4        o294(.A(ori_ori_n316_), .B(ori_ori_n313_), .C(ori_ori_n309_), .D(ori_ori_n48_), .Y(ori_ori_n317_));
  INV        o295(.A(ori_ori_n189_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n319_));
  OAI220     o297(.A0(ori_ori_n319_), .A1(ori_ori_n421_), .B0(ori_ori_n318_), .B1(ori_ori_n59_), .Y(ori_ori_n320_));
  NA2        o298(.A(ori_ori_n320_), .B(x02), .Y(ori_ori_n321_));
  INV        o299(.A(ori_ori_n225_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n186_), .B(x04), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n323_), .B(ori_ori_n322_), .Y(ori_ori_n324_));
  NO3        o302(.A(ori_ori_n168_), .B(x13), .C(ori_ori_n31_), .Y(ori_ori_n325_));
  OAI210     o303(.A0(ori_ori_n325_), .A1(ori_ori_n324_), .B0(ori_ori_n96_), .Y(ori_ori_n326_));
  NO3        o304(.A(ori_ori_n186_), .B(ori_ori_n150_), .C(ori_ori_n52_), .Y(ori_ori_n327_));
  OAI210     o305(.A0(ori_ori_n138_), .A1(ori_ori_n36_), .B0(ori_ori_n101_), .Y(ori_ori_n328_));
  OAI210     o306(.A0(ori_ori_n328_), .A1(ori_ori_n178_), .B0(ori_ori_n327_), .Y(ori_ori_n329_));
  NA4        o307(.A(ori_ori_n329_), .B(ori_ori_n326_), .C(ori_ori_n321_), .D(x06), .Y(ori_ori_n330_));
  NA2        o308(.A(x09), .B(x03), .Y(ori_ori_n331_));
  OAI220     o309(.A0(ori_ori_n331_), .A1(ori_ori_n119_), .B0(ori_ori_n196_), .B1(ori_ori_n63_), .Y(ori_ori_n332_));
  OAI220     o310(.A0(ori_ori_n151_), .A1(x09), .B0(x08), .B1(ori_ori_n41_), .Y(ori_ori_n333_));
  NO3        o311(.A(ori_ori_n264_), .B(ori_ori_n118_), .C(x08), .Y(ori_ori_n334_));
  AOI210     o312(.A0(ori_ori_n333_), .A1(ori_ori_n210_), .B0(ori_ori_n334_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n336_));
  NO3        o314(.A(ori_ori_n109_), .B(ori_ori_n119_), .C(ori_ori_n38_), .Y(ori_ori_n337_));
  AOI210     o315(.A0(ori_ori_n327_), .A1(ori_ori_n336_), .B0(ori_ori_n337_), .Y(ori_ori_n338_));
  OAI210     o316(.A0(ori_ori_n335_), .A1(ori_ori_n28_), .B0(ori_ori_n338_), .Y(ori_ori_n339_));
  AO220      o317(.A0(ori_ori_n339_), .A1(x04), .B0(ori_ori_n332_), .B1(x05), .Y(ori_ori_n340_));
  AOI210     o318(.A0(ori_ori_n330_), .A1(ori_ori_n317_), .B0(ori_ori_n340_), .Y(ori_ori_n341_));
  OAI210     o319(.A0(ori_ori_n304_), .A1(x12), .B0(ori_ori_n341_), .Y(ori03));
  OR2        o320(.A(ori_ori_n42_), .B(ori_ori_n211_), .Y(ori_ori_n343_));
  AOI210     o321(.A0(ori_ori_n143_), .A1(ori_ori_n101_), .B0(ori_ori_n343_), .Y(ori_ori_n344_));
  AO210      o322(.A0(ori_ori_n322_), .A1(ori_ori_n86_), .B0(ori_ori_n323_), .Y(ori_ori_n345_));
  NA2        o323(.A(ori_ori_n186_), .B(ori_ori_n142_), .Y(ori_ori_n346_));
  NA3        o324(.A(ori_ori_n346_), .B(ori_ori_n345_), .C(ori_ori_n190_), .Y(ori_ori_n347_));
  OAI210     o325(.A0(ori_ori_n347_), .A1(ori_ori_n344_), .B0(x05), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n343_), .B(x05), .Y(ori_ori_n349_));
  AOI210     o327(.A0(ori_ori_n129_), .A1(ori_ori_n202_), .B0(ori_ori_n349_), .Y(ori_ori_n350_));
  AOI210     o328(.A0(ori_ori_n213_), .A1(ori_ori_n80_), .B0(ori_ori_n114_), .Y(ori_ori_n351_));
  OAI220     o329(.A0(ori_ori_n351_), .A1(ori_ori_n59_), .B0(ori_ori_n293_), .B1(ori_ori_n284_), .Y(ori_ori_n352_));
  OAI210     o330(.A0(ori_ori_n352_), .A1(ori_ori_n350_), .B0(ori_ori_n101_), .Y(ori_ori_n353_));
  AOI210     o331(.A0(ori_ori_n136_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n354_));
  NO2        o332(.A(ori_ori_n159_), .B(ori_ori_n124_), .Y(ori_ori_n355_));
  OAI220     o333(.A0(ori_ori_n355_), .A1(ori_ori_n37_), .B0(ori_ori_n139_), .B1(x13), .Y(ori_ori_n356_));
  OAI210     o334(.A0(ori_ori_n356_), .A1(ori_ori_n354_), .B0(x04), .Y(ori_ori_n357_));
  NO3        o335(.A(ori_ori_n315_), .B(ori_ori_n85_), .C(ori_ori_n59_), .Y(ori_ori_n358_));
  AOI210     o336(.A0(ori_ori_n174_), .A1(ori_ori_n101_), .B0(ori_ori_n136_), .Y(ori_ori_n359_));
  OA210      o337(.A0(ori_ori_n152_), .A1(x12), .B0(ori_ori_n124_), .Y(ori_ori_n360_));
  NO3        o338(.A(ori_ori_n360_), .B(ori_ori_n359_), .C(ori_ori_n358_), .Y(ori_ori_n361_));
  NA4        o339(.A(ori_ori_n361_), .B(ori_ori_n357_), .C(ori_ori_n353_), .D(ori_ori_n348_), .Y(ori04));
  NO2        o340(.A(ori_ori_n89_), .B(ori_ori_n39_), .Y(ori_ori_n363_));
  XO2        o341(.A(ori_ori_n363_), .B(ori_ori_n235_), .Y(ori05));
  NO2        o342(.A(ori_ori_n52_), .B(ori_ori_n199_), .Y(ori_ori_n365_));
  AOI210     o343(.A0(ori_ori_n365_), .A1(ori_ori_n292_), .B0(ori_ori_n25_), .Y(ori_ori_n366_));
  NA3        o344(.A(ori_ori_n132_), .B(ori_ori_n121_), .C(ori_ori_n31_), .Y(ori_ori_n367_));
  INV        o345(.A(ori_ori_n90_), .Y(ori_ori_n368_));
  AOI210     o346(.A0(ori_ori_n368_), .A1(ori_ori_n367_), .B0(ori_ori_n24_), .Y(ori_ori_n369_));
  OAI210     o347(.A0(ori_ori_n369_), .A1(ori_ori_n366_), .B0(ori_ori_n101_), .Y(ori_ori_n370_));
  NA2        o348(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n371_));
  NA2        o349(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n240_), .B(x03), .Y(ori_ori_n373_));
  OAI220     o351(.A0(ori_ori_n373_), .A1(ori_ori_n372_), .B0(ori_ori_n371_), .B1(ori_ori_n81_), .Y(ori_ori_n374_));
  OAI210     o352(.A0(ori_ori_n26_), .A1(ori_ori_n101_), .B0(x07), .Y(ori_ori_n375_));
  AOI210     o353(.A0(ori_ori_n374_), .A1(x06), .B0(ori_ori_n375_), .Y(ori_ori_n376_));
  AOI210     o354(.A0(ori_ori_n81_), .A1(ori_ori_n31_), .B0(ori_ori_n52_), .Y(ori_ori_n377_));
  NO3        o355(.A(ori_ori_n377_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n378_));
  INV        o356(.A(ori_ori_n373_), .Y(ori_ori_n379_));
  OR2        o357(.A(ori_ori_n379_), .B(ori_ori_n224_), .Y(ori_ori_n380_));
  NA2        o358(.A(ori_ori_n228_), .B(ori_ori_n222_), .Y(ori_ori_n381_));
  NA2        o359(.A(ori_ori_n381_), .B(ori_ori_n380_), .Y(ori_ori_n382_));
  OAI210     o360(.A0(ori_ori_n382_), .A1(ori_ori_n378_), .B0(ori_ori_n101_), .Y(ori_ori_n383_));
  NA2        o361(.A(ori_ori_n33_), .B(ori_ori_n101_), .Y(ori_ori_n384_));
  AOI210     o362(.A0(ori_ori_n384_), .A1(ori_ori_n92_), .B0(x07), .Y(ori_ori_n385_));
  AOI220     o363(.A0(ori_ori_n385_), .A1(ori_ori_n383_), .B0(ori_ori_n376_), .B1(ori_ori_n370_), .Y(ori_ori_n386_));
  OR2        o364(.A(ori_ori_n251_), .B(ori_ori_n248_), .Y(ori_ori_n387_));
  NO2        o365(.A(ori_ori_n135_), .B(ori_ori_n28_), .Y(ori_ori_n388_));
  AOI210     o366(.A0(ori_ori_n387_), .A1(ori_ori_n47_), .B0(ori_ori_n388_), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n389_), .B(ori_ori_n102_), .Y(ori_ori_n390_));
  AOI210     o368(.A0(ori_ori_n323_), .A1(ori_ori_n108_), .B0(ori_ori_n247_), .Y(ori_ori_n391_));
  NOi21      o369(.An(ori_ori_n305_), .B(ori_ori_n124_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n392_), .B(ori_ori_n248_), .Y(ori_ori_n393_));
  OAI210     o371(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n394_));
  AOI210     o372(.A0(ori_ori_n235_), .A1(ori_ori_n47_), .B0(ori_ori_n394_), .Y(ori_ori_n395_));
  NO4        o373(.A(ori_ori_n395_), .B(ori_ori_n393_), .C(ori_ori_n391_), .D(x08), .Y(ori_ori_n396_));
  NO2        o374(.A(ori_ori_n121_), .B(ori_ori_n28_), .Y(ori_ori_n397_));
  NO2        o375(.A(ori_ori_n397_), .B(ori_ori_n252_), .Y(ori_ori_n398_));
  OR3        o376(.A(ori_ori_n398_), .B(x12), .C(x03), .Y(ori_ori_n399_));
  NA3        o377(.A(ori_ori_n318_), .B(ori_ori_n115_), .C(x12), .Y(ori_ori_n400_));
  AO210      o378(.A0(ori_ori_n318_), .A1(ori_ori_n115_), .B0(ori_ori_n235_), .Y(ori_ori_n401_));
  NA4        o379(.A(ori_ori_n401_), .B(ori_ori_n400_), .C(ori_ori_n399_), .D(x08), .Y(ori_ori_n402_));
  INV        o380(.A(ori_ori_n402_), .Y(ori_ori_n403_));
  AOI210     o381(.A0(ori_ori_n396_), .A1(ori_ori_n390_), .B0(ori_ori_n403_), .Y(ori_ori_n404_));
  INV        o382(.A(x03), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n135_), .B(ori_ori_n43_), .Y(ori_ori_n406_));
  OAI210     o384(.A0(ori_ori_n406_), .A1(ori_ori_n405_), .B0(ori_ori_n173_), .Y(ori_ori_n407_));
  NA3        o385(.A(ori_ori_n398_), .B(ori_ori_n392_), .C(ori_ori_n314_), .Y(ori_ori_n408_));
  INV        o386(.A(x14), .Y(ori_ori_n409_));
  NO3        o387(.A(ori_ori_n151_), .B(ori_ori_n74_), .C(ori_ori_n57_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n410_), .B(ori_ori_n409_), .Y(ori_ori_n411_));
  NA3        o389(.A(ori_ori_n411_), .B(ori_ori_n408_), .C(ori_ori_n407_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n384_), .B(ori_ori_n61_), .Y(ori_ori_n413_));
  NOi21      o391(.An(ori_ori_n256_), .B(ori_ori_n139_), .Y(ori_ori_n414_));
  NO2        o392(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n415_));
  OAI210     o393(.A0(ori_ori_n415_), .A1(ori_ori_n414_), .B0(ori_ori_n101_), .Y(ori_ori_n416_));
  OAI210     o394(.A0(ori_ori_n413_), .A1(ori_ori_n91_), .B0(ori_ori_n416_), .Y(ori_ori_n417_));
  NO4        o395(.A(ori_ori_n417_), .B(ori_ori_n412_), .C(ori_ori_n404_), .D(ori_ori_n386_), .Y(ori06));
  INV        o396(.A(ori_ori_n40_), .Y(ori_ori_n421_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n61_), .B(mai_mai_n23_), .Y(mai_mai_n71_));
  NA2        m049(.A(x09), .B(x05), .Y(mai_mai_n72_));
  NA2        m050(.A(x10), .B(x06), .Y(mai_mai_n73_));
  NA3        m051(.A(mai_mai_n73_), .B(mai_mai_n72_), .C(mai_mai_n28_), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n61_), .B(mai_mai_n41_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n74_), .A1(mai_mai_n71_), .B0(x03), .Y(mai_mai_n76_));
  NOi31      m054(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n77_));
  NO2        m055(.A(x10), .B(x09), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n450_), .B(mai_mai_n24_), .Y(mai_mai_n79_));
  NO2        m057(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n80_));
  NO2        m058(.A(mai_mai_n80_), .B(mai_mai_n36_), .Y(mai_mai_n81_));
  OAI210     m059(.A0(mai_mai_n80_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n82_));
  AOI210     m060(.A0(mai_mai_n81_), .A1(mai_mai_n48_), .B0(mai_mai_n82_), .Y(mai_mai_n83_));
  NO2        m061(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n84_));
  NO2        m062(.A(x08), .B(x01), .Y(mai_mai_n85_));
  OAI210     m063(.A0(mai_mai_n85_), .A1(mai_mai_n84_), .B0(mai_mai_n35_), .Y(mai_mai_n86_));
  NA2        m064(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n87_));
  NO3        m065(.A(mai_mai_n86_), .B(mai_mai_n83_), .C(mai_mai_n79_), .Y(mai_mai_n88_));
  AN2        m066(.A(mai_mai_n88_), .B(mai_mai_n76_), .Y(mai_mai_n89_));
  INV        m067(.A(mai_mai_n86_), .Y(mai_mai_n90_));
  NO2        m068(.A(x06), .B(x05), .Y(mai_mai_n91_));
  NA2        m069(.A(x11), .B(x00), .Y(mai_mai_n92_));
  NO2        m070(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n93_));
  NOi21      m071(.An(mai_mai_n92_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  NOi21      m072(.An(x01), .B(x10), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n95_), .C(x06), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n97_), .B(mai_mai_n27_), .Y(mai_mai_n98_));
  OAI210     m076(.A0(mai_mai_n452_), .A1(x07), .B0(mai_mai_n98_), .Y(mai_mai_n99_));
  NO3        m077(.A(mai_mai_n99_), .B(mai_mai_n89_), .C(mai_mai_n70_), .Y(mai01));
  INV        m078(.A(x12), .Y(mai_mai_n101_));
  INV        m079(.A(x13), .Y(mai_mai_n102_));
  NA2        m080(.A(x08), .B(x04), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n57_), .Y(mai_mai_n104_));
  NA2        m082(.A(mai_mai_n104_), .B(mai_mai_n91_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n95_), .B(mai_mai_n28_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(mai_mai_n72_), .Y(mai_mai_n107_));
  NO2        m085(.A(x10), .B(x01), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NA2        m088(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n111_));
  NO3        m089(.A(mai_mai_n111_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n112_));
  AOI210     m090(.A0(mai_mai_n112_), .A1(mai_mai_n110_), .B0(mai_mai_n107_), .Y(mai_mai_n113_));
  AOI210     m091(.A0(mai_mai_n113_), .A1(mai_mai_n105_), .B0(mai_mai_n102_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n115_));
  NOi21      m093(.An(mai_mai_n115_), .B(mai_mai_n58_), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n102_), .B(mai_mai_n36_), .Y(mai_mai_n118_));
  NA3        m096(.A(mai_mai_n118_), .B(mai_mai_n117_), .C(x06), .Y(mai_mai_n119_));
  INV        m097(.A(mai_mai_n119_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n85_), .B(x13), .Y(mai_mai_n121_));
  NA2        m099(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n122_), .B(mai_mai_n121_), .Y(mai_mai_n123_));
  NA2        m101(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n124_));
  NO2        m102(.A(mai_mai_n124_), .B(x05), .Y(mai_mai_n125_));
  NO2        m103(.A(mai_mai_n125_), .B(mai_mai_n123_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n127_));
  INV        m105(.A(mai_mai_n116_), .Y(mai_mai_n128_));
  AOI210     m106(.A0(mai_mai_n128_), .A1(mai_mai_n126_), .B0(mai_mai_n73_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n130_));
  NA2        m108(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(mai_mai_n130_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n36_), .B(x04), .Y(mai_mai_n134_));
  NA3        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(x13), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n127_), .B(mai_mai_n36_), .Y(mai_mai_n136_));
  NO2        m114(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n137_));
  NOi41      m115(.An(mai_mai_n135_), .B(mai_mai_n137_), .C(mai_mai_n136_), .D(mai_mai_n132_), .Y(mai_mai_n138_));
  NO3        m116(.A(mai_mai_n138_), .B(x06), .C(x03), .Y(mai_mai_n139_));
  NO4        m117(.A(mai_mai_n139_), .B(mai_mai_n129_), .C(mai_mai_n120_), .D(mai_mai_n114_), .Y(mai_mai_n140_));
  NA2        m118(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n141_));
  OAI210     m119(.A0(mai_mai_n85_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n35_), .B(mai_mai_n47_), .Y(mai_mai_n144_));
  OA210      m122(.A0(x00), .A1(mai_mai_n78_), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n147_));
  AOI210     m125(.A0(mai_mai_n147_), .A1(mai_mai_n49_), .B0(mai_mai_n146_), .Y(mai_mai_n148_));
  OA210      m126(.A0(mai_mai_n148_), .A1(mai_mai_n145_), .B0(mai_mai_n143_), .Y(mai_mai_n149_));
  NO2        m127(.A(x09), .B(x05), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n150_), .B(mai_mai_n47_), .Y(mai_mai_n151_));
  AOI210     m129(.A0(mai_mai_n151_), .A1(mai_mai_n110_), .B0(mai_mai_n49_), .Y(mai_mai_n152_));
  NA2        m130(.A(x09), .B(x00), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n115_), .B(mai_mai_n153_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n77_), .B(mai_mai_n51_), .Y(mai_mai_n155_));
  AOI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n154_), .B0(mai_mai_n147_), .Y(mai_mai_n156_));
  NO3        m134(.A(mai_mai_n156_), .B(mai_mai_n152_), .C(mai_mai_n149_), .Y(mai_mai_n157_));
  NO2        m135(.A(x03), .B(x02), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n86_), .B(mai_mai_n102_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n116_), .B0(mai_mai_n158_), .Y(mai_mai_n160_));
  OA210      m138(.A0(mai_mai_n157_), .A1(x11), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  OAI210     m139(.A0(mai_mai_n140_), .A1(mai_mai_n23_), .B0(mai_mai_n161_), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n110_), .B(mai_mai_n40_), .Y(mai_mai_n163_));
  NAi21      m141(.An(x06), .B(x10), .Y(mai_mai_n164_));
  NOi21      m142(.An(x01), .B(x13), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  BUFFER     m144(.A(mai_mai_n166_), .Y(mai_mai_n167_));
  AOI210     m145(.A0(mai_mai_n167_), .A1(mai_mai_n163_), .B0(mai_mai_n41_), .Y(mai_mai_n168_));
  NO2        m146(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n102_), .B(x01), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n170_), .B(x08), .Y(mai_mai_n171_));
  NO2        m149(.A(mai_mai_n169_), .B(mai_mai_n48_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n173_));
  OAI210     m151(.A0(mai_mai_n172_), .A1(mai_mai_n168_), .B0(mai_mai_n173_), .Y(mai_mai_n174_));
  NA2        m152(.A(x04), .B(x02), .Y(mai_mai_n175_));
  NA2        m153(.A(x10), .B(x05), .Y(mai_mai_n176_));
  INV        m154(.A(x06), .Y(mai_mai_n177_));
  NO2        m155(.A(x09), .B(x01), .Y(mai_mai_n178_));
  NO3        m156(.A(mai_mai_n178_), .B(mai_mai_n108_), .C(mai_mai_n31_), .Y(mai_mai_n179_));
  NA2        m157(.A(mai_mai_n179_), .B(x00), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n115_), .B(x08), .Y(mai_mai_n181_));
  NA3        m159(.A(mai_mai_n165_), .B(mai_mai_n164_), .C(mai_mai_n51_), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n95_), .B(x05), .Y(mai_mai_n183_));
  OAI210     m161(.A0(mai_mai_n183_), .A1(mai_mai_n118_), .B0(mai_mai_n182_), .Y(mai_mai_n184_));
  AOI210     m162(.A0(mai_mai_n181_), .A1(x06), .B0(mai_mai_n184_), .Y(mai_mai_n185_));
  OAI210     m163(.A0(mai_mai_n185_), .A1(x11), .B0(mai_mai_n180_), .Y(mai_mai_n186_));
  NAi21      m164(.An(mai_mai_n175_), .B(mai_mai_n186_), .Y(mai_mai_n187_));
  INV        m165(.A(mai_mai_n25_), .Y(mai_mai_n188_));
  NAi21      m166(.An(x13), .B(x00), .Y(mai_mai_n189_));
  BUFFER     m167(.A(mai_mai_n72_), .Y(mai_mai_n190_));
  NO2        m168(.A(mai_mai_n96_), .B(x06), .Y(mai_mai_n191_));
  NO2        m169(.A(mai_mai_n189_), .B(mai_mai_n36_), .Y(mai_mai_n192_));
  INV        m170(.A(mai_mai_n192_), .Y(mai_mai_n193_));
  OAI220     m171(.A0(mai_mai_n193_), .A1(mai_mai_n177_), .B0(mai_mai_n191_), .B1(mai_mai_n190_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(mai_mai_n188_), .Y(mai_mai_n195_));
  NOi21      m173(.An(x09), .B(x00), .Y(mai_mai_n196_));
  NO3        m174(.A(mai_mai_n84_), .B(mai_mai_n196_), .C(mai_mai_n47_), .Y(mai_mai_n197_));
  NA2        m175(.A(mai_mai_n197_), .B(mai_mai_n131_), .Y(mai_mai_n198_));
  NA2        m176(.A(x06), .B(x05), .Y(mai_mai_n199_));
  OAI210     m177(.A0(mai_mai_n199_), .A1(mai_mai_n35_), .B0(mai_mai_n101_), .Y(mai_mai_n200_));
  AOI210     m178(.A0(x10), .A1(mai_mai_n58_), .B0(mai_mai_n200_), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n201_), .B(mai_mai_n198_), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n102_), .B(x12), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n203_), .Y(mai_mai_n204_));
  NA2        m182(.A(mai_mai_n95_), .B(mai_mai_n51_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n206_), .B(x02), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n207_), .B(mai_mai_n205_), .Y(mai_mai_n208_));
  AOI210     m186(.A0(mai_mai_n204_), .A1(mai_mai_n202_), .B0(mai_mai_n208_), .Y(mai_mai_n209_));
  NA4        m187(.A(mai_mai_n209_), .B(mai_mai_n195_), .C(mai_mai_n187_), .D(mai_mai_n174_), .Y(mai_mai_n210_));
  AOI210     m188(.A0(mai_mai_n162_), .A1(mai_mai_n101_), .B0(mai_mai_n210_), .Y(mai_mai_n211_));
  INV        m189(.A(mai_mai_n74_), .Y(mai_mai_n212_));
  NA2        m190(.A(mai_mai_n212_), .B(mai_mai_n143_), .Y(mai_mai_n213_));
  NA2        m191(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n214_), .B(mai_mai_n142_), .Y(mai_mai_n215_));
  AOI210     m193(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n130_), .B(x06), .Y(mai_mai_n217_));
  AOI210     m195(.A0(mai_mai_n216_), .A1(mai_mai_n215_), .B0(mai_mai_n217_), .Y(mai_mai_n218_));
  AOI210     m196(.A0(mai_mai_n218_), .A1(mai_mai_n213_), .B0(x12), .Y(mai_mai_n219_));
  INV        m197(.A(mai_mai_n77_), .Y(mai_mai_n220_));
  NO2        m198(.A(x05), .B(mai_mai_n51_), .Y(mai_mai_n221_));
  OAI210     m199(.A0(mai_mai_n221_), .A1(mai_mai_n166_), .B0(mai_mai_n57_), .Y(mai_mai_n222_));
  NA2        m200(.A(mai_mai_n222_), .B(mai_mai_n220_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n95_), .B(x06), .Y(mai_mai_n224_));
  AOI210     m202(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n225_));
  NO3        m203(.A(mai_mai_n225_), .B(mai_mai_n224_), .C(mai_mai_n41_), .Y(mai_mai_n226_));
  NA4        m204(.A(mai_mai_n164_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n227_));
  NA2        m205(.A(mai_mai_n227_), .B(mai_mai_n147_), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(x02), .Y(mai_mai_n229_));
  AOI210     m207(.A0(mai_mai_n229_), .A1(mai_mai_n223_), .B0(mai_mai_n23_), .Y(mai_mai_n230_));
  OAI210     m208(.A0(mai_mai_n219_), .A1(mai_mai_n57_), .B0(mai_mai_n230_), .Y(mai_mai_n231_));
  INV        m209(.A(mai_mai_n147_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n233_));
  OAI210     m211(.A0(mai_mai_n80_), .A1(mai_mai_n36_), .B0(mai_mai_n122_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n102_), .B(x03), .Y(mai_mai_n235_));
  AOI220     m213(.A0(mai_mai_n235_), .A1(mai_mai_n234_), .B0(mai_mai_n77_), .B1(mai_mai_n233_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n237_));
  INV        m215(.A(mai_mai_n164_), .Y(mai_mai_n238_));
  NOi21      m216(.An(x13), .B(x04), .Y(mai_mai_n239_));
  NO3        m217(.A(mai_mai_n239_), .B(mai_mai_n77_), .C(mai_mai_n196_), .Y(mai_mai_n240_));
  NO2        m218(.A(mai_mai_n240_), .B(x05), .Y(mai_mai_n241_));
  AOI220     m219(.A0(mai_mai_n241_), .A1(mai_mai_n237_), .B0(mai_mai_n238_), .B1(mai_mai_n57_), .Y(mai_mai_n242_));
  OAI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n232_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  INV        m221(.A(mai_mai_n93_), .Y(mai_mai_n244_));
  NO2        m222(.A(mai_mai_n244_), .B(x12), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n248_));
  NO2        m226(.A(x06), .B(x00), .Y(mai_mai_n249_));
  NO3        m227(.A(mai_mai_n249_), .B(mai_mai_n248_), .C(mai_mai_n41_), .Y(mai_mai_n250_));
  INV        m228(.A(mai_mai_n73_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n253_), .B(x03), .Y(mai_mai_n254_));
  OR2        m232(.A(mai_mai_n254_), .B(mai_mai_n252_), .Y(mai_mai_n255_));
  NA2        m233(.A(x13), .B(mai_mai_n101_), .Y(mai_mai_n256_));
  NA3        m234(.A(mai_mai_n256_), .B(mai_mai_n200_), .C(mai_mai_n94_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n255_), .A1(mai_mai_n246_), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  AOI210     m236(.A0(mai_mai_n245_), .A1(mai_mai_n243_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  AOI210     m237(.A0(mai_mai_n259_), .A1(mai_mai_n231_), .B0(x07), .Y(mai_mai_n260_));
  NA2        m238(.A(mai_mai_n72_), .B(mai_mai_n29_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n239_), .B(mai_mai_n196_), .Y(mai_mai_n262_));
  AOI210     m240(.A0(mai_mai_n262_), .A1(mai_mai_n155_), .B0(mai_mai_n261_), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n102_), .B(x06), .Y(mai_mai_n264_));
  INV        m242(.A(mai_mai_n264_), .Y(mai_mai_n265_));
  NO2        m243(.A(x08), .B(x05), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n266_), .B(mai_mai_n248_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n77_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n268_));
  OAI210     m246(.A0(mai_mai_n267_), .A1(mai_mai_n265_), .B0(mai_mai_n268_), .Y(mai_mai_n269_));
  NO2        m247(.A(x12), .B(x02), .Y(mai_mai_n270_));
  INV        m248(.A(mai_mai_n270_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n271_), .B(mai_mai_n244_), .Y(mai_mai_n272_));
  OA210      m250(.A0(mai_mai_n269_), .A1(mai_mai_n263_), .B0(mai_mai_n272_), .Y(mai_mai_n273_));
  NA2        m251(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n274_), .B(x01), .Y(mai_mai_n275_));
  INV        m253(.A(mai_mai_n275_), .Y(mai_mai_n276_));
  AOI210     m254(.A0(mai_mai_n276_), .A1(mai_mai_n135_), .B0(mai_mai_n29_), .Y(mai_mai_n277_));
  NA2        m255(.A(mai_mai_n264_), .B(mai_mai_n234_), .Y(mai_mai_n278_));
  NA2        m256(.A(mai_mai_n102_), .B(x04), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n279_), .B(mai_mai_n28_), .Y(mai_mai_n280_));
  OAI210     m258(.A0(mai_mai_n280_), .A1(mai_mai_n121_), .B0(mai_mai_n278_), .Y(mai_mai_n281_));
  NO3        m259(.A(mai_mai_n92_), .B(x12), .C(x03), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n281_), .A1(mai_mai_n277_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  NOi21      m261(.An(mai_mai_n261_), .B(mai_mai_n224_), .Y(mai_mai_n284_));
  NO2        m262(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n285_));
  NA2        m263(.A(mai_mai_n284_), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  NO2        m264(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n287_));
  NO3        m265(.A(mai_mai_n287_), .B(mai_mai_n225_), .C(mai_mai_n191_), .Y(mai_mai_n288_));
  NO2        m266(.A(mai_mai_n246_), .B(mai_mai_n28_), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n288_), .A1(mai_mai_n232_), .B0(mai_mai_n289_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n290_), .B(mai_mai_n286_), .C(mai_mai_n283_), .Y(mai_mai_n291_));
  NO3        m269(.A(mai_mai_n291_), .B(mai_mai_n273_), .C(mai_mai_n260_), .Y(mai_mai_n292_));
  OAI210     m270(.A0(mai_mai_n211_), .A1(mai_mai_n61_), .B0(mai_mai_n292_), .Y(mai02));
  AOI210     m271(.A0(mai_mai_n141_), .A1(mai_mai_n86_), .B0(mai_mai_n133_), .Y(mai_mai_n294_));
  NOi21      m272(.An(mai_mai_n240_), .B(mai_mai_n178_), .Y(mai_mai_n295_));
  NO2        m273(.A(mai_mai_n295_), .B(mai_mai_n32_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n296_), .A1(mai_mai_n294_), .B0(mai_mai_n176_), .Y(mai_mai_n297_));
  INV        m275(.A(mai_mai_n176_), .Y(mai_mai_n298_));
  AOI210     m276(.A0(mai_mai_n117_), .A1(mai_mai_n87_), .B0(mai_mai_n225_), .Y(mai_mai_n299_));
  OAI220     m277(.A0(mai_mai_n299_), .A1(mai_mai_n102_), .B0(mai_mai_n86_), .B1(mai_mai_n51_), .Y(mai_mai_n300_));
  AOI220     m278(.A0(mai_mai_n300_), .A1(mai_mai_n298_), .B0(mai_mai_n159_), .B1(mai_mai_n158_), .Y(mai_mai_n301_));
  AOI210     m279(.A0(mai_mai_n301_), .A1(mai_mai_n297_), .B0(mai_mai_n48_), .Y(mai_mai_n302_));
  NO2        m280(.A(x05), .B(x02), .Y(mai_mai_n303_));
  OAI210     m281(.A0(mai_mai_n215_), .A1(mai_mai_n196_), .B0(mai_mai_n303_), .Y(mai_mai_n304_));
  AOI220     m282(.A0(mai_mai_n266_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n305_));
  NA2        m283(.A(mai_mai_n239_), .B(mai_mai_n80_), .Y(mai_mai_n306_));
  AOI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n304_), .B0(mai_mai_n147_), .Y(mai_mai_n307_));
  NAi21      m285(.An(mai_mai_n241_), .B(mai_mai_n236_), .Y(mai_mai_n308_));
  NO2        m286(.A(mai_mai_n253_), .B(mai_mai_n47_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  AN2        m288(.A(mai_mai_n235_), .B(mai_mai_n234_), .Y(mai_mai_n311_));
  OAI210     m289(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n312_));
  NA2        m290(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n313_));
  OA210      m291(.A0(mai_mai_n313_), .A1(x08), .B0(mai_mai_n151_), .Y(mai_mai_n314_));
  AOI210     m292(.A0(mai_mai_n314_), .A1(mai_mai_n142_), .B0(mai_mai_n312_), .Y(mai_mai_n315_));
  OAI210     m293(.A0(mai_mai_n315_), .A1(mai_mai_n311_), .B0(mai_mai_n96_), .Y(mai_mai_n316_));
  NA3        m294(.A(mai_mai_n96_), .B(mai_mai_n85_), .C(mai_mai_n233_), .Y(mai_mai_n317_));
  NA3        m295(.A(mai_mai_n95_), .B(mai_mai_n84_), .C(mai_mai_n42_), .Y(mai_mai_n318_));
  AOI210     m296(.A0(mai_mai_n318_), .A1(mai_mai_n317_), .B0(x04), .Y(mai_mai_n319_));
  INV        m297(.A(mai_mai_n158_), .Y(mai_mai_n320_));
  OAI220     m298(.A0(mai_mai_n267_), .A1(mai_mai_n106_), .B0(mai_mai_n320_), .B1(mai_mai_n132_), .Y(mai_mai_n321_));
  AOI210     m299(.A0(mai_mai_n321_), .A1(x13), .B0(mai_mai_n319_), .Y(mai_mai_n322_));
  NA3        m300(.A(mai_mai_n322_), .B(mai_mai_n316_), .C(mai_mai_n310_), .Y(mai_mai_n323_));
  NO3        m301(.A(mai_mai_n323_), .B(mai_mai_n307_), .C(mai_mai_n302_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n146_), .B(x03), .Y(mai_mai_n325_));
  INV        m303(.A(mai_mai_n189_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n51_), .A1(mai_mai_n35_), .B0(mai_mai_n36_), .Y(mai_mai_n327_));
  AOI220     m305(.A0(mai_mai_n327_), .A1(mai_mai_n326_), .B0(mai_mai_n206_), .B1(x08), .Y(mai_mai_n328_));
  OAI210     m306(.A0(mai_mai_n328_), .A1(mai_mai_n287_), .B0(mai_mai_n325_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(mai_mai_n108_), .Y(mai_mai_n330_));
  NA2        m308(.A(mai_mai_n175_), .B(mai_mai_n170_), .Y(mai_mai_n331_));
  AN2        m309(.A(mai_mai_n331_), .B(mai_mai_n181_), .Y(mai_mai_n332_));
  INV        m310(.A(mai_mai_n56_), .Y(mai_mai_n333_));
  OAI220     m311(.A0(mai_mai_n279_), .A1(mai_mai_n333_), .B0(mai_mai_n133_), .B1(mai_mai_n28_), .Y(mai_mai_n334_));
  OAI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n332_), .B0(mai_mai_n109_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n279_), .B(mai_mai_n101_), .Y(mai_mai_n336_));
  NA2        m314(.A(mai_mai_n101_), .B(mai_mai_n41_), .Y(mai_mai_n337_));
  NA3        m315(.A(mai_mai_n337_), .B(mai_mai_n336_), .C(mai_mai_n132_), .Y(mai_mai_n338_));
  NA4        m316(.A(mai_mai_n338_), .B(mai_mai_n335_), .C(mai_mai_n330_), .D(mai_mai_n48_), .Y(mai_mai_n339_));
  INV        m317(.A(mai_mai_n206_), .Y(mai_mai_n340_));
  NO2        m318(.A(mai_mai_n171_), .B(mai_mai_n40_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n342_));
  OAI220     m320(.A0(mai_mai_n342_), .A1(mai_mai_n341_), .B0(mai_mai_n340_), .B1(mai_mai_n59_), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n343_), .B(x02), .Y(mai_mai_n344_));
  INV        m322(.A(mai_mai_n247_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n203_), .B(x04), .Y(mai_mai_n346_));
  NO3        m324(.A(mai_mai_n203_), .B(mai_mai_n169_), .C(mai_mai_n52_), .Y(mai_mai_n347_));
  OAI210     m325(.A0(mai_mai_n153_), .A1(mai_mai_n36_), .B0(mai_mai_n101_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(mai_mai_n348_), .A1(mai_mai_n197_), .B0(mai_mai_n347_), .Y(mai_mai_n349_));
  NA3        m327(.A(mai_mai_n349_), .B(mai_mai_n344_), .C(x06), .Y(mai_mai_n350_));
  NA2        m328(.A(x09), .B(x03), .Y(mai_mai_n351_));
  OAI220     m329(.A0(mai_mai_n351_), .A1(mai_mai_n131_), .B0(mai_mai_n214_), .B1(mai_mai_n64_), .Y(mai_mai_n352_));
  OAI220     m330(.A0(mai_mai_n170_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n353_));
  NO3        m331(.A(mai_mai_n287_), .B(mai_mai_n130_), .C(x08), .Y(mai_mai_n354_));
  AOI210     m332(.A0(mai_mai_n353_), .A1(mai_mai_n232_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NO2        m333(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n356_));
  NO3        m334(.A(mai_mai_n115_), .B(mai_mai_n131_), .C(mai_mai_n38_), .Y(mai_mai_n357_));
  AOI210     m335(.A0(mai_mai_n347_), .A1(mai_mai_n356_), .B0(mai_mai_n357_), .Y(mai_mai_n358_));
  OAI210     m336(.A0(mai_mai_n355_), .A1(mai_mai_n28_), .B0(mai_mai_n358_), .Y(mai_mai_n359_));
  AO220      m337(.A0(mai_mai_n359_), .A1(x04), .B0(mai_mai_n352_), .B1(x05), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n350_), .A1(mai_mai_n339_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  OAI210     m339(.A0(mai_mai_n324_), .A1(x12), .B0(mai_mai_n361_), .Y(mai03));
  OR2        m340(.A(mai_mai_n42_), .B(mai_mai_n233_), .Y(mai_mai_n363_));
  AOI210     m341(.A0(mai_mai_n159_), .A1(mai_mai_n101_), .B0(mai_mai_n363_), .Y(mai_mai_n364_));
  AO210      m342(.A0(mai_mai_n345_), .A1(mai_mai_n87_), .B0(mai_mai_n346_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n203_), .B(mai_mai_n158_), .Y(mai_mai_n366_));
  NA3        m344(.A(mai_mai_n366_), .B(mai_mai_n365_), .C(mai_mai_n207_), .Y(mai_mai_n367_));
  OAI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n364_), .B0(x05), .Y(mai_mai_n368_));
  NA2        m346(.A(mai_mai_n363_), .B(x05), .Y(mai_mai_n369_));
  AOI210     m347(.A0(mai_mai_n142_), .A1(mai_mai_n220_), .B0(mai_mai_n369_), .Y(mai_mai_n370_));
  AOI210     m348(.A0(mai_mai_n235_), .A1(mai_mai_n81_), .B0(mai_mai_n125_), .Y(mai_mai_n371_));
  OAI220     m349(.A0(mai_mai_n371_), .A1(mai_mai_n59_), .B0(mai_mai_n313_), .B1(mai_mai_n305_), .Y(mai_mai_n372_));
  OAI210     m350(.A0(mai_mai_n372_), .A1(mai_mai_n370_), .B0(mai_mai_n101_), .Y(mai_mai_n373_));
  AOI210     m351(.A0(mai_mai_n151_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n374_));
  NO2        m352(.A(mai_mai_n178_), .B(mai_mai_n137_), .Y(mai_mai_n375_));
  OAI220     m353(.A0(mai_mai_n375_), .A1(mai_mai_n37_), .B0(mai_mai_n154_), .B1(x13), .Y(mai_mai_n376_));
  OAI210     m354(.A0(mai_mai_n376_), .A1(mai_mai_n374_), .B0(x04), .Y(mai_mai_n377_));
  NO3        m355(.A(mai_mai_n337_), .B(mai_mai_n86_), .C(mai_mai_n59_), .Y(mai_mai_n378_));
  AOI210     m356(.A0(mai_mai_n193_), .A1(mai_mai_n101_), .B0(mai_mai_n151_), .Y(mai_mai_n379_));
  OA210      m357(.A0(mai_mai_n171_), .A1(x12), .B0(mai_mai_n137_), .Y(mai_mai_n380_));
  NO3        m358(.A(mai_mai_n380_), .B(mai_mai_n379_), .C(mai_mai_n378_), .Y(mai_mai_n381_));
  NA4        m359(.A(mai_mai_n381_), .B(mai_mai_n377_), .C(mai_mai_n373_), .D(mai_mai_n368_), .Y(mai04));
  NO2        m360(.A(mai_mai_n90_), .B(mai_mai_n39_), .Y(mai_mai_n383_));
  XO2        m361(.A(mai_mai_n383_), .B(mai_mai_n256_), .Y(mai05));
  AOI210     m362(.A0(mai_mai_n72_), .A1(mai_mai_n52_), .B0(mai_mai_n217_), .Y(mai_mai_n385_));
  AOI210     m363(.A0(mai_mai_n385_), .A1(mai_mai_n312_), .B0(mai_mai_n25_), .Y(mai_mai_n386_));
  NO2        m364(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n387_));
  OAI210     m365(.A0(mai_mai_n387_), .A1(mai_mai_n386_), .B0(mai_mai_n101_), .Y(mai_mai_n388_));
  OAI210     m366(.A0(mai_mai_n26_), .A1(mai_mai_n101_), .B0(x07), .Y(mai_mai_n389_));
  INV        m367(.A(mai_mai_n389_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n82_), .B(mai_mai_n31_), .Y(mai_mai_n391_));
  NO3        m369(.A(mai_mai_n391_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n392_));
  NO2        m370(.A(mai_mai_n451_), .B(mai_mai_n264_), .Y(mai_mai_n393_));
  OR2        m371(.A(mai_mai_n393_), .B(mai_mai_n246_), .Y(mai_mai_n394_));
  NA2        m372(.A(mai_mai_n165_), .B(x05), .Y(mai_mai_n395_));
  NA3        m373(.A(mai_mai_n395_), .B(mai_mai_n249_), .C(mai_mai_n244_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n397_));
  OAI210     m375(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n398_));
  OR3        m376(.A(mai_mai_n398_), .B(mai_mai_n397_), .C(mai_mai_n44_), .Y(mai_mai_n399_));
  NA3        m377(.A(mai_mai_n399_), .B(mai_mai_n396_), .C(mai_mai_n394_), .Y(mai_mai_n400_));
  OAI210     m378(.A0(mai_mai_n400_), .A1(mai_mai_n392_), .B0(mai_mai_n101_), .Y(mai_mai_n401_));
  NA2        m379(.A(mai_mai_n33_), .B(mai_mai_n101_), .Y(mai_mai_n402_));
  AOI210     m380(.A0(mai_mai_n402_), .A1(mai_mai_n93_), .B0(x07), .Y(mai_mai_n403_));
  AOI220     m381(.A0(mai_mai_n403_), .A1(mai_mai_n401_), .B0(mai_mai_n390_), .B1(mai_mai_n388_), .Y(mai_mai_n404_));
  NA3        m382(.A(mai_mai_n23_), .B(mai_mai_n61_), .C(mai_mai_n48_), .Y(mai_mai_n405_));
  AOI210     m383(.A0(mai_mai_n397_), .A1(mai_mai_n75_), .B0(mai_mai_n146_), .Y(mai_mai_n406_));
  OR2        m384(.A(mai_mai_n406_), .B(x03), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n356_), .B(mai_mai_n61_), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n408_), .B(x11), .Y(mai_mai_n409_));
  NO3        m387(.A(mai_mai_n409_), .B(mai_mai_n150_), .C(mai_mai_n28_), .Y(mai_mai_n410_));
  AOI210     m388(.A0(mai_mai_n410_), .A1(mai_mai_n407_), .B0(mai_mai_n47_), .Y(mai_mai_n411_));
  NO4        m389(.A(mai_mai_n337_), .B(mai_mai_n32_), .C(x11), .D(x09), .Y(mai_mai_n412_));
  OAI210     m390(.A0(mai_mai_n412_), .A1(mai_mai_n411_), .B0(mai_mai_n102_), .Y(mai_mai_n413_));
  AOI210     m391(.A0(mai_mai_n346_), .A1(mai_mai_n111_), .B0(mai_mai_n270_), .Y(mai_mai_n414_));
  NOi21      m392(.An(mai_mai_n325_), .B(mai_mai_n137_), .Y(mai_mai_n415_));
  NO2        m393(.A(mai_mai_n415_), .B(mai_mai_n271_), .Y(mai_mai_n416_));
  OAI210     m394(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n417_));
  AOI210     m395(.A0(mai_mai_n256_), .A1(mai_mai_n47_), .B0(mai_mai_n417_), .Y(mai_mai_n418_));
  NO4        m396(.A(mai_mai_n418_), .B(mai_mai_n416_), .C(mai_mai_n414_), .D(x08), .Y(mai_mai_n419_));
  NA2        m397(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n420_));
  NO2        m398(.A(mai_mai_n420_), .B(x03), .Y(mai_mai_n421_));
  NO2        m399(.A(x13), .B(x12), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n133_), .B(mai_mai_n28_), .Y(mai_mai_n423_));
  NO2        m401(.A(mai_mai_n423_), .B(mai_mai_n275_), .Y(mai_mai_n424_));
  OR3        m402(.A(mai_mai_n424_), .B(x12), .C(x03), .Y(mai_mai_n425_));
  NA3        m403(.A(mai_mai_n340_), .B(mai_mai_n127_), .C(x12), .Y(mai_mai_n426_));
  AO210      m404(.A0(mai_mai_n340_), .A1(mai_mai_n127_), .B0(mai_mai_n256_), .Y(mai_mai_n427_));
  NA4        m405(.A(mai_mai_n427_), .B(mai_mai_n426_), .C(mai_mai_n425_), .D(x08), .Y(mai_mai_n428_));
  AOI210     m406(.A0(mai_mai_n422_), .A1(mai_mai_n421_), .B0(mai_mai_n428_), .Y(mai_mai_n429_));
  AOI210     m407(.A0(mai_mai_n419_), .A1(mai_mai_n413_), .B0(mai_mai_n429_), .Y(mai_mai_n430_));
  OAI210     m408(.A0(mai_mai_n408_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n431_));
  OAI220     m409(.A0(mai_mai_n176_), .A1(x02), .B0(mai_mai_n150_), .B1(mai_mai_n43_), .Y(mai_mai_n432_));
  OAI210     m410(.A0(mai_mai_n432_), .A1(mai_mai_n431_), .B0(mai_mai_n192_), .Y(mai_mai_n433_));
  NA3        m411(.A(mai_mai_n424_), .B(mai_mai_n415_), .C(mai_mai_n336_), .Y(mai_mai_n434_));
  INV        m412(.A(x14), .Y(mai_mai_n435_));
  NO3        m413(.A(mai_mai_n325_), .B(mai_mai_n106_), .C(x11), .Y(mai_mai_n436_));
  NO3        m414(.A(mai_mai_n170_), .B(mai_mai_n75_), .C(mai_mai_n57_), .Y(mai_mai_n437_));
  NO3        m415(.A(mai_mai_n405_), .B(mai_mai_n337_), .C(mai_mai_n189_), .Y(mai_mai_n438_));
  NO4        m416(.A(mai_mai_n438_), .B(mai_mai_n437_), .C(mai_mai_n436_), .D(mai_mai_n435_), .Y(mai_mai_n439_));
  NA3        m417(.A(mai_mai_n439_), .B(mai_mai_n434_), .C(mai_mai_n433_), .Y(mai_mai_n440_));
  AOI220     m418(.A0(mai_mai_n402_), .A1(mai_mai_n61_), .B0(mai_mai_n423_), .B1(mai_mai_n169_), .Y(mai_mai_n441_));
  NOi21      m419(.An(mai_mai_n279_), .B(mai_mai_n154_), .Y(mai_mai_n442_));
  NA2        m420(.A(mai_mai_n285_), .B(mai_mai_n238_), .Y(mai_mai_n443_));
  OAI210     m421(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n443_), .Y(mai_mai_n444_));
  OAI210     m422(.A0(mai_mai_n444_), .A1(mai_mai_n442_), .B0(mai_mai_n101_), .Y(mai_mai_n445_));
  OAI210     m423(.A0(mai_mai_n441_), .A1(mai_mai_n92_), .B0(mai_mai_n445_), .Y(mai_mai_n446_));
  NO4        m424(.A(mai_mai_n446_), .B(mai_mai_n440_), .C(mai_mai_n430_), .D(mai_mai_n404_), .Y(mai06));
  INV        m425(.A(x07), .Y(mai_mai_n450_));
  INV        m426(.A(x02), .Y(mai_mai_n451_));
  INV        m427(.A(mai_mai_n94_), .Y(mai_mai_n452_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  INV        u027(.A(x09), .Y(men_men_n50_));
  NO2        u028(.A(x10), .B(x02), .Y(men_men_n51_));
  NOi21      u029(.An(x01), .B(x09), .Y(men_men_n52_));
  INV        u030(.A(x00), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n54_), .B(men_men_n52_), .Y(men_men_n55_));
  NA2        u033(.A(x09), .B(men_men_n53_), .Y(men_men_n56_));
  INV        u034(.A(x07), .Y(men_men_n57_));
  AOI220     u035(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n57_), .Y(men_men_n58_));
  INV        u036(.A(men_men_n55_), .Y(men_men_n59_));
  NA2        u037(.A(men_men_n29_), .B(x02), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n60_), .B(men_men_n24_), .Y(men_men_n61_));
  OAI220     u039(.A0(men_men_n61_), .A1(men_men_n59_), .B0(men_men_n58_), .B1(men_men_n56_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n57_), .B(men_men_n48_), .Y(men_men_n63_));
  OAI210     u041(.A0(men_men_n30_), .A1(x11), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u042(.A0(men_men_n64_), .A1(men_men_n55_), .B0(men_men_n62_), .B1(men_men_n31_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n65_), .B(x05), .Y(men_men_n66_));
  NA2        u044(.A(x10), .B(x09), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n57_), .B(men_men_n23_), .Y(men_men_n68_));
  NA2        u046(.A(x09), .B(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x06), .Y(men_men_n70_));
  NA3        u048(.A(men_men_n70_), .B(men_men_n69_), .C(men_men_n28_), .Y(men_men_n71_));
  OAI210     u049(.A0(men_men_n71_), .A1(men_men_n68_), .B0(x03), .Y(men_men_n72_));
  NOi31      u050(.An(x08), .B(x04), .C(x00), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n458_), .B(men_men_n24_), .Y(men_men_n74_));
  NO2        u052(.A(x09), .B(men_men_n41_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n75_), .B(men_men_n36_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n77_));
  AOI210     u055(.A0(men_men_n76_), .A1(men_men_n48_), .B0(men_men_n77_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n36_), .B(x00), .Y(men_men_n79_));
  NO2        u057(.A(x08), .B(x01), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n80_), .A1(men_men_n79_), .B0(men_men_n35_), .Y(men_men_n81_));
  NA2        u059(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n82_));
  NO3        u060(.A(men_men_n81_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n83_));
  AN2        u061(.A(men_men_n83_), .B(men_men_n72_), .Y(men_men_n84_));
  INV        u062(.A(men_men_n81_), .Y(men_men_n85_));
  NO2        u063(.A(x06), .B(x05), .Y(men_men_n86_));
  NA2        u064(.A(x11), .B(x00), .Y(men_men_n87_));
  NO2        u065(.A(x11), .B(men_men_n47_), .Y(men_men_n88_));
  NOi21      u066(.An(men_men_n87_), .B(men_men_n88_), .Y(men_men_n89_));
  AOI210     u067(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n89_), .Y(men_men_n90_));
  NOi21      u068(.An(x01), .B(x10), .Y(men_men_n91_));
  NO2        u069(.A(men_men_n29_), .B(men_men_n53_), .Y(men_men_n92_));
  NO3        u070(.A(men_men_n92_), .B(men_men_n91_), .C(x06), .Y(men_men_n93_));
  NA2        u071(.A(men_men_n93_), .B(men_men_n27_), .Y(men_men_n94_));
  OAI210     u072(.A0(men_men_n90_), .A1(x07), .B0(men_men_n94_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n84_), .C(men_men_n66_), .Y(men01));
  INV        u074(.A(x12), .Y(men_men_n97_));
  INV        u075(.A(x13), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n86_), .B(x01), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n99_), .B(men_men_n67_), .Y(men_men_n100_));
  NA2        u078(.A(x08), .B(x04), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n101_), .B(men_men_n53_), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n102_), .B(men_men_n100_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n91_), .B(men_men_n28_), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n69_), .Y(men_men_n105_));
  NO2        u083(.A(x10), .B(x01), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n29_), .B(x00), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NA2        u086(.A(x04), .B(men_men_n28_), .Y(men_men_n109_));
  NO3        u087(.A(men_men_n109_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n110_));
  AOI210     u088(.A0(men_men_n110_), .A1(men_men_n108_), .B0(men_men_n105_), .Y(men_men_n111_));
  AOI210     u089(.A0(men_men_n111_), .A1(men_men_n103_), .B0(men_men_n98_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n52_), .B(x05), .Y(men_men_n113_));
  NOi21      u091(.An(men_men_n113_), .B(men_men_n54_), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n35_), .B(x02), .Y(men_men_n115_));
  NA3        u093(.A(x13), .B(men_men_n115_), .C(x06), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n116_), .B(men_men_n114_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n80_), .B(x13), .Y(men_men_n118_));
  NA2        u096(.A(x09), .B(men_men_n35_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u098(.A(x13), .B(men_men_n35_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(x05), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(men_men_n120_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n35_), .B(men_men_n53_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n124_), .B(men_men_n98_), .Y(men_men_n125_));
  AOI210     u103(.A0(men_men_n125_), .A1(men_men_n76_), .B0(men_men_n114_), .Y(men_men_n126_));
  AOI210     u104(.A0(men_men_n126_), .A1(men_men_n123_), .B0(men_men_n70_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n128_));
  NA2        u106(.A(x10), .B(men_men_n53_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n129_), .B(men_men_n128_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n50_), .B(x05), .Y(men_men_n131_));
  NO3        u109(.A(men_men_n124_), .B(men_men_n75_), .C(men_men_n36_), .Y(men_men_n132_));
  NO2        u110(.A(men_men_n56_), .B(x05), .Y(men_men_n133_));
  NO3        u111(.A(men_men_n133_), .B(men_men_n132_), .C(men_men_n130_), .Y(men_men_n134_));
  NO3        u112(.A(men_men_n134_), .B(x06), .C(x03), .Y(men_men_n135_));
  NO4        u113(.A(men_men_n135_), .B(men_men_n127_), .C(men_men_n117_), .D(men_men_n112_), .Y(men_men_n136_));
  NA2        u114(.A(x13), .B(men_men_n36_), .Y(men_men_n137_));
  OAI210     u115(.A0(men_men_n80_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n138_), .B(men_men_n137_), .Y(men_men_n139_));
  NO2        u117(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n140_));
  AN2        u118(.A(men_men_n86_), .B(men_men_n140_), .Y(men_men_n141_));
  NO2        u119(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n142_));
  NA2        u120(.A(men_men_n29_), .B(x06), .Y(men_men_n143_));
  AOI210     u121(.A0(men_men_n143_), .A1(men_men_n49_), .B0(men_men_n142_), .Y(men_men_n144_));
  OA210      u122(.A0(men_men_n144_), .A1(men_men_n141_), .B0(men_men_n139_), .Y(men_men_n145_));
  NO2        u123(.A(x09), .B(x05), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n146_), .B(men_men_n47_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n108_), .B(men_men_n49_), .Y(men_men_n148_));
  NA2        u126(.A(x09), .B(x00), .Y(men_men_n149_));
  NA2        u127(.A(men_men_n113_), .B(men_men_n149_), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n73_), .B(men_men_n50_), .Y(men_men_n151_));
  AOI210     u129(.A0(men_men_n151_), .A1(men_men_n150_), .B0(men_men_n143_), .Y(men_men_n152_));
  NO3        u130(.A(men_men_n152_), .B(men_men_n148_), .C(men_men_n145_), .Y(men_men_n153_));
  NO2        u131(.A(x03), .B(x02), .Y(men_men_n154_));
  NA2        u132(.A(men_men_n81_), .B(men_men_n98_), .Y(men_men_n155_));
  OAI210     u133(.A0(men_men_n155_), .A1(men_men_n114_), .B0(men_men_n154_), .Y(men_men_n156_));
  OA210      u134(.A0(men_men_n153_), .A1(x11), .B0(men_men_n156_), .Y(men_men_n157_));
  OAI210     u135(.A0(men_men_n136_), .A1(men_men_n23_), .B0(men_men_n157_), .Y(men_men_n158_));
  NA2        u136(.A(men_men_n108_), .B(men_men_n40_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n160_));
  NAi21      u138(.An(x06), .B(x10), .Y(men_men_n161_));
  NOi21      u139(.An(x01), .B(x13), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  OR2        u141(.A(men_men_n163_), .B(men_men_n160_), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n159_), .B0(men_men_n41_), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n29_), .B(x03), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n98_), .B(x01), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n167_), .B(x08), .Y(men_men_n168_));
  OAI210     u146(.A0(x05), .A1(men_men_n168_), .B0(men_men_n50_), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n169_), .A1(men_men_n166_), .B0(men_men_n48_), .Y(men_men_n170_));
  AOI210     u148(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n170_), .A1(men_men_n165_), .B0(men_men_n171_), .Y(men_men_n172_));
  NA2        u150(.A(x04), .B(x02), .Y(men_men_n173_));
  NA2        u151(.A(x10), .B(x05), .Y(men_men_n174_));
  NA2        u152(.A(x09), .B(x06), .Y(men_men_n175_));
  AOI210     u153(.A0(men_men_n175_), .A1(men_men_n174_), .B0(men_men_n160_), .Y(men_men_n176_));
  NO2        u154(.A(x09), .B(x01), .Y(men_men_n177_));
  NA2        u155(.A(men_men_n176_), .B(x00), .Y(men_men_n178_));
  NO2        u156(.A(men_men_n113_), .B(x08), .Y(men_men_n179_));
  NA3        u157(.A(men_men_n162_), .B(men_men_n161_), .C(men_men_n50_), .Y(men_men_n180_));
  NA2        u158(.A(men_men_n91_), .B(x05), .Y(men_men_n181_));
  NA2        u159(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  AOI210     u160(.A0(men_men_n179_), .A1(x06), .B0(men_men_n182_), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n183_), .A1(x11), .B0(men_men_n178_), .Y(men_men_n184_));
  NAi21      u162(.An(men_men_n173_), .B(men_men_n184_), .Y(men_men_n185_));
  INV        u163(.A(men_men_n25_), .Y(men_men_n186_));
  NAi21      u164(.An(x13), .B(x00), .Y(men_men_n187_));
  AOI210     u165(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n187_), .Y(men_men_n188_));
  AOI220     u166(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n174_), .A1(men_men_n35_), .B0(men_men_n189_), .Y(men_men_n190_));
  AN2        u168(.A(men_men_n190_), .B(men_men_n188_), .Y(men_men_n191_));
  NO2        u169(.A(men_men_n92_), .B(x06), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n187_), .B(men_men_n36_), .Y(men_men_n193_));
  INV        u171(.A(men_men_n193_), .Y(men_men_n194_));
  OAI210     u172(.A0(men_men_n194_), .A1(men_men_n175_), .B0(men_men_n70_), .Y(men_men_n195_));
  OAI210     u173(.A0(men_men_n195_), .A1(men_men_n191_), .B0(men_men_n186_), .Y(men_men_n196_));
  NOi21      u174(.An(x09), .B(x00), .Y(men_men_n197_));
  NO3        u175(.A(men_men_n79_), .B(men_men_n197_), .C(men_men_n47_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n198_), .B(men_men_n129_), .Y(men_men_n199_));
  NA2        u177(.A(x10), .B(x08), .Y(men_men_n200_));
  INV        u178(.A(men_men_n200_), .Y(men_men_n201_));
  NA2        u179(.A(x06), .B(x05), .Y(men_men_n202_));
  OAI210     u180(.A0(men_men_n202_), .A1(men_men_n35_), .B0(men_men_n97_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n201_), .A1(men_men_n54_), .B0(men_men_n203_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n204_), .B(men_men_n199_), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n98_), .B(x12), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n206_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n91_), .B(men_men_n50_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n209_), .B(x02), .Y(men_men_n210_));
  NO2        u188(.A(men_men_n210_), .B(men_men_n208_), .Y(men_men_n211_));
  AOI210     u189(.A0(men_men_n207_), .A1(men_men_n205_), .B0(men_men_n211_), .Y(men_men_n212_));
  NA4        u190(.A(men_men_n212_), .B(men_men_n196_), .C(men_men_n185_), .D(men_men_n172_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n158_), .A1(men_men_n97_), .B0(men_men_n213_), .Y(men_men_n214_));
  INV        u192(.A(men_men_n71_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(men_men_n139_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n138_), .Y(men_men_n218_));
  AOI210     u196(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n128_), .B(x06), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n219_), .A1(men_men_n218_), .B0(men_men_n220_), .Y(men_men_n221_));
  AOI210     u199(.A0(men_men_n221_), .A1(men_men_n216_), .B0(x12), .Y(men_men_n222_));
  INV        u200(.A(men_men_n73_), .Y(men_men_n223_));
  NO2        u201(.A(x05), .B(men_men_n50_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n224_), .A1(men_men_n163_), .B0(men_men_n53_), .Y(men_men_n225_));
  NA2        u203(.A(men_men_n225_), .B(men_men_n223_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n91_), .B(x06), .Y(men_men_n227_));
  AOI210     u205(.A0(men_men_n36_), .A1(x04), .B0(men_men_n50_), .Y(men_men_n228_));
  NO3        u206(.A(men_men_n228_), .B(men_men_n227_), .C(men_men_n41_), .Y(men_men_n229_));
  NA4        u207(.A(men_men_n161_), .B(men_men_n52_), .C(men_men_n36_), .D(x04), .Y(men_men_n230_));
  NA2        u208(.A(men_men_n230_), .B(men_men_n143_), .Y(men_men_n231_));
  OAI210     u209(.A0(men_men_n231_), .A1(men_men_n229_), .B0(x02), .Y(men_men_n232_));
  AOI210     u210(.A0(men_men_n232_), .A1(men_men_n226_), .B0(men_men_n23_), .Y(men_men_n233_));
  OAI210     u211(.A0(men_men_n222_), .A1(men_men_n53_), .B0(men_men_n233_), .Y(men_men_n234_));
  INV        u212(.A(men_men_n143_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n50_), .B(x03), .Y(men_men_n236_));
  OAI210     u214(.A0(men_men_n75_), .A1(men_men_n36_), .B0(men_men_n119_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n98_), .B(x03), .Y(men_men_n238_));
  AOI220     u216(.A0(men_men_n238_), .A1(men_men_n237_), .B0(men_men_n73_), .B1(men_men_n236_), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n32_), .B(x06), .Y(men_men_n240_));
  INV        u218(.A(men_men_n161_), .Y(men_men_n241_));
  NOi21      u219(.An(x13), .B(x04), .Y(men_men_n242_));
  NO3        u220(.A(men_men_n242_), .B(men_men_n73_), .C(men_men_n197_), .Y(men_men_n243_));
  NO2        u221(.A(men_men_n243_), .B(x05), .Y(men_men_n244_));
  AOI220     u222(.A0(men_men_n244_), .A1(men_men_n240_), .B0(men_men_n241_), .B1(men_men_n53_), .Y(men_men_n245_));
  OAI210     u223(.A0(men_men_n239_), .A1(men_men_n235_), .B0(men_men_n245_), .Y(men_men_n246_));
  INV        u224(.A(men_men_n88_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n247_), .B(x12), .Y(men_men_n248_));
  NA2        u226(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n249_));
  NO2        u227(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n250_), .A1(men_men_n190_), .B0(men_men_n188_), .Y(men_men_n251_));
  AOI210     u229(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n252_));
  NA2        u230(.A(men_men_n149_), .B(men_men_n70_), .Y(men_men_n253_));
  INV        u231(.A(men_men_n253_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n255_), .B(x03), .Y(men_men_n256_));
  OA210      u234(.A0(men_men_n256_), .A1(men_men_n254_), .B0(men_men_n251_), .Y(men_men_n257_));
  NA2        u235(.A(x13), .B(men_men_n97_), .Y(men_men_n258_));
  NA3        u236(.A(men_men_n258_), .B(men_men_n203_), .C(men_men_n89_), .Y(men_men_n259_));
  OAI210     u237(.A0(men_men_n257_), .A1(men_men_n249_), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n248_), .A1(men_men_n246_), .B0(men_men_n260_), .Y(men_men_n261_));
  AOI210     u239(.A0(men_men_n261_), .A1(men_men_n234_), .B0(x07), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n69_), .B(men_men_n29_), .Y(men_men_n263_));
  NOi21      u241(.An(men_men_n137_), .B(men_men_n197_), .Y(men_men_n264_));
  AOI210     u242(.A0(men_men_n264_), .A1(men_men_n151_), .B0(men_men_n263_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n98_), .B(x06), .Y(men_men_n266_));
  INV        u244(.A(men_men_n266_), .Y(men_men_n267_));
  NO2        u245(.A(x08), .B(x05), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n268_), .B(men_men_n252_), .Y(men_men_n269_));
  NA2        u247(.A(x13), .B(men_men_n31_), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n269_), .A1(men_men_n267_), .B0(men_men_n270_), .Y(men_men_n271_));
  NO2        u249(.A(x12), .B(x02), .Y(men_men_n272_));
  INV        u250(.A(men_men_n272_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n273_), .B(men_men_n247_), .Y(men_men_n274_));
  OA210      u252(.A0(men_men_n271_), .A1(men_men_n265_), .B0(men_men_n274_), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n276_), .B(x01), .Y(men_men_n277_));
  NOi21      u255(.An(men_men_n80_), .B(men_men_n119_), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n278_), .B(men_men_n277_), .Y(men_men_n279_));
  NO2        u257(.A(men_men_n279_), .B(men_men_n29_), .Y(men_men_n280_));
  NA2        u258(.A(men_men_n266_), .B(men_men_n237_), .Y(men_men_n281_));
  NA2        u259(.A(men_men_n98_), .B(x04), .Y(men_men_n282_));
  NA2        u260(.A(men_men_n282_), .B(men_men_n28_), .Y(men_men_n283_));
  OAI210     u261(.A0(men_men_n283_), .A1(men_men_n118_), .B0(men_men_n281_), .Y(men_men_n284_));
  NO3        u262(.A(men_men_n87_), .B(x12), .C(x03), .Y(men_men_n285_));
  OAI210     u263(.A0(men_men_n284_), .A1(men_men_n280_), .B0(men_men_n285_), .Y(men_men_n286_));
  AOI210     u264(.A0(men_men_n208_), .A1(men_men_n202_), .B0(men_men_n101_), .Y(men_men_n287_));
  NOi21      u265(.An(men_men_n263_), .B(men_men_n227_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n25_), .B(x00), .Y(men_men_n289_));
  OAI210     u267(.A0(men_men_n288_), .A1(men_men_n287_), .B0(men_men_n289_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n54_), .B(x05), .Y(men_men_n291_));
  NO3        u269(.A(men_men_n291_), .B(men_men_n228_), .C(men_men_n192_), .Y(men_men_n292_));
  NO2        u270(.A(men_men_n249_), .B(men_men_n28_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n292_), .A1(men_men_n235_), .B0(men_men_n293_), .Y(men_men_n294_));
  NA3        u272(.A(men_men_n294_), .B(men_men_n290_), .C(men_men_n286_), .Y(men_men_n295_));
  NO3        u273(.A(men_men_n295_), .B(men_men_n275_), .C(men_men_n262_), .Y(men_men_n296_));
  OAI210     u274(.A0(men_men_n214_), .A1(men_men_n57_), .B0(men_men_n296_), .Y(men02));
  AOI210     u275(.A0(men_men_n137_), .A1(men_men_n81_), .B0(men_men_n131_), .Y(men_men_n298_));
  NOi21      u276(.An(men_men_n243_), .B(men_men_n177_), .Y(men_men_n299_));
  NO2        u277(.A(men_men_n98_), .B(men_men_n35_), .Y(men_men_n300_));
  NA3        u278(.A(men_men_n300_), .B(men_men_n201_), .C(men_men_n52_), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n299_), .A1(men_men_n32_), .B0(men_men_n301_), .Y(men_men_n302_));
  OAI210     u280(.A0(men_men_n302_), .A1(men_men_n298_), .B0(men_men_n174_), .Y(men_men_n303_));
  INV        u281(.A(men_men_n174_), .Y(men_men_n304_));
  AOI210     u282(.A0(men_men_n115_), .A1(men_men_n82_), .B0(men_men_n228_), .Y(men_men_n305_));
  OAI220     u283(.A0(men_men_n305_), .A1(men_men_n98_), .B0(men_men_n81_), .B1(men_men_n50_), .Y(men_men_n306_));
  AOI220     u284(.A0(men_men_n306_), .A1(men_men_n304_), .B0(men_men_n155_), .B1(men_men_n154_), .Y(men_men_n307_));
  AOI210     u285(.A0(men_men_n307_), .A1(men_men_n303_), .B0(men_men_n48_), .Y(men_men_n308_));
  NO2        u286(.A(x05), .B(x02), .Y(men_men_n309_));
  OAI210     u287(.A0(men_men_n218_), .A1(men_men_n197_), .B0(men_men_n309_), .Y(men_men_n310_));
  AOI220     u288(.A0(men_men_n268_), .A1(men_men_n54_), .B0(men_men_n52_), .B1(men_men_n36_), .Y(men_men_n311_));
  NOi21      u289(.An(men_men_n300_), .B(men_men_n311_), .Y(men_men_n312_));
  INV        u290(.A(men_men_n312_), .Y(men_men_n313_));
  AOI210     u291(.A0(men_men_n313_), .A1(men_men_n310_), .B0(men_men_n143_), .Y(men_men_n314_));
  NAi21      u292(.An(men_men_n244_), .B(men_men_n239_), .Y(men_men_n315_));
  NO2        u293(.A(men_men_n255_), .B(men_men_n47_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n316_), .B(men_men_n315_), .Y(men_men_n317_));
  AN2        u295(.A(men_men_n238_), .B(men_men_n237_), .Y(men_men_n318_));
  OAI210     u296(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n319_));
  NA2        u297(.A(x13), .B(men_men_n28_), .Y(men_men_n320_));
  AOI210     u298(.A0(men_men_n147_), .A1(men_men_n138_), .B0(men_men_n319_), .Y(men_men_n321_));
  OAI210     u299(.A0(men_men_n321_), .A1(men_men_n318_), .B0(men_men_n92_), .Y(men_men_n322_));
  INV        u300(.A(men_men_n154_), .Y(men_men_n323_));
  OAI220     u301(.A0(men_men_n269_), .A1(men_men_n104_), .B0(men_men_n323_), .B1(men_men_n130_), .Y(men_men_n324_));
  NA2        u302(.A(men_men_n324_), .B(x13), .Y(men_men_n325_));
  NA3        u303(.A(men_men_n325_), .B(men_men_n322_), .C(men_men_n317_), .Y(men_men_n326_));
  NO3        u304(.A(men_men_n326_), .B(men_men_n314_), .C(men_men_n308_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n142_), .B(x03), .Y(men_men_n328_));
  INV        u306(.A(men_men_n187_), .Y(men_men_n329_));
  OAI210     u307(.A0(men_men_n50_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n330_));
  AOI220     u308(.A0(men_men_n330_), .A1(men_men_n329_), .B0(men_men_n209_), .B1(x08), .Y(men_men_n331_));
  OAI210     u309(.A0(men_men_n331_), .A1(men_men_n291_), .B0(men_men_n328_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n332_), .B(men_men_n106_), .Y(men_men_n333_));
  NA2        u311(.A(men_men_n173_), .B(men_men_n167_), .Y(men_men_n334_));
  AN2        u312(.A(men_men_n334_), .B(men_men_n179_), .Y(men_men_n335_));
  INV        u313(.A(men_men_n52_), .Y(men_men_n336_));
  OAI220     u314(.A0(men_men_n282_), .A1(men_men_n336_), .B0(men_men_n131_), .B1(men_men_n28_), .Y(men_men_n337_));
  OAI210     u315(.A0(men_men_n337_), .A1(men_men_n335_), .B0(men_men_n107_), .Y(men_men_n338_));
  NA2        u316(.A(men_men_n282_), .B(men_men_n97_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n97_), .B(men_men_n41_), .Y(men_men_n340_));
  NA3        u318(.A(men_men_n340_), .B(men_men_n339_), .C(men_men_n130_), .Y(men_men_n341_));
  NA4        u319(.A(men_men_n341_), .B(men_men_n338_), .C(men_men_n333_), .D(men_men_n48_), .Y(men_men_n342_));
  INV        u320(.A(men_men_n209_), .Y(men_men_n343_));
  NO2        u321(.A(men_men_n168_), .B(men_men_n40_), .Y(men_men_n344_));
  NA2        u322(.A(men_men_n32_), .B(x05), .Y(men_men_n345_));
  OAI220     u323(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n343_), .B1(men_men_n55_), .Y(men_men_n346_));
  NA2        u324(.A(men_men_n346_), .B(x02), .Y(men_men_n347_));
  INV        u325(.A(men_men_n250_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n206_), .B(x04), .Y(men_men_n349_));
  NO2        u327(.A(men_men_n349_), .B(men_men_n348_), .Y(men_men_n350_));
  NO3        u328(.A(men_men_n189_), .B(x13), .C(men_men_n31_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n351_), .A1(men_men_n350_), .B0(men_men_n92_), .Y(men_men_n352_));
  NO3        u330(.A(men_men_n206_), .B(men_men_n166_), .C(men_men_n51_), .Y(men_men_n353_));
  OAI210     u331(.A0(men_men_n149_), .A1(men_men_n36_), .B0(men_men_n97_), .Y(men_men_n354_));
  OAI210     u332(.A0(men_men_n354_), .A1(men_men_n198_), .B0(men_men_n353_), .Y(men_men_n355_));
  NA4        u333(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n347_), .D(x06), .Y(men_men_n356_));
  NA2        u334(.A(x09), .B(x03), .Y(men_men_n357_));
  OAI220     u335(.A0(men_men_n357_), .A1(men_men_n129_), .B0(men_men_n217_), .B1(men_men_n60_), .Y(men_men_n358_));
  NO3        u336(.A(men_men_n291_), .B(men_men_n128_), .C(x08), .Y(men_men_n359_));
  INV        u337(.A(men_men_n359_), .Y(men_men_n360_));
  NO3        u338(.A(men_men_n113_), .B(men_men_n129_), .C(men_men_n38_), .Y(men_men_n361_));
  INV        u339(.A(men_men_n361_), .Y(men_men_n362_));
  OAI210     u340(.A0(men_men_n360_), .A1(men_men_n28_), .B0(men_men_n362_), .Y(men_men_n363_));
  AO220      u341(.A0(men_men_n363_), .A1(x04), .B0(men_men_n358_), .B1(x05), .Y(men_men_n364_));
  AOI210     u342(.A0(men_men_n356_), .A1(men_men_n342_), .B0(men_men_n364_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n327_), .A1(x12), .B0(men_men_n365_), .Y(men03));
  OR2        u344(.A(men_men_n42_), .B(men_men_n236_), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n155_), .A1(men_men_n97_), .B0(men_men_n367_), .Y(men_men_n368_));
  AO210      u346(.A0(men_men_n348_), .A1(men_men_n82_), .B0(men_men_n349_), .Y(men_men_n369_));
  NA2        u347(.A(men_men_n206_), .B(men_men_n154_), .Y(men_men_n370_));
  NA3        u348(.A(men_men_n370_), .B(men_men_n369_), .C(men_men_n210_), .Y(men_men_n371_));
  OAI210     u349(.A0(men_men_n371_), .A1(men_men_n368_), .B0(x05), .Y(men_men_n372_));
  NA2        u350(.A(men_men_n367_), .B(x05), .Y(men_men_n373_));
  AOI210     u351(.A0(men_men_n138_), .A1(men_men_n223_), .B0(men_men_n373_), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n238_), .A1(men_men_n76_), .B0(men_men_n122_), .Y(men_men_n375_));
  OAI220     u353(.A0(men_men_n375_), .A1(men_men_n55_), .B0(men_men_n320_), .B1(men_men_n311_), .Y(men_men_n376_));
  OAI210     u354(.A0(men_men_n376_), .A1(men_men_n374_), .B0(men_men_n97_), .Y(men_men_n377_));
  AOI210     u355(.A0(men_men_n147_), .A1(men_men_n56_), .B0(men_men_n38_), .Y(men_men_n378_));
  NO2        u356(.A(men_men_n177_), .B(men_men_n133_), .Y(men_men_n379_));
  OAI220     u357(.A0(men_men_n379_), .A1(men_men_n37_), .B0(men_men_n150_), .B1(x13), .Y(men_men_n380_));
  OAI210     u358(.A0(men_men_n380_), .A1(men_men_n378_), .B0(x04), .Y(men_men_n381_));
  NO3        u359(.A(men_men_n340_), .B(men_men_n81_), .C(men_men_n55_), .Y(men_men_n382_));
  AOI210     u360(.A0(men_men_n194_), .A1(men_men_n97_), .B0(men_men_n147_), .Y(men_men_n383_));
  OA210      u361(.A0(men_men_n168_), .A1(x12), .B0(men_men_n133_), .Y(men_men_n384_));
  NO3        u362(.A(men_men_n384_), .B(men_men_n383_), .C(men_men_n382_), .Y(men_men_n385_));
  NA4        u363(.A(men_men_n385_), .B(men_men_n381_), .C(men_men_n377_), .D(men_men_n372_), .Y(men04));
  NO2        u364(.A(men_men_n85_), .B(men_men_n39_), .Y(men_men_n387_));
  XO2        u365(.A(men_men_n387_), .B(men_men_n258_), .Y(men05));
  NO2        u366(.A(men_men_n319_), .B(men_men_n25_), .Y(men_men_n389_));
  NA3        u367(.A(men_men_n143_), .B(men_men_n131_), .C(men_men_n31_), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n241_), .A1(men_men_n53_), .B0(men_men_n86_), .Y(men_men_n391_));
  AOI210     u369(.A0(men_men_n391_), .A1(men_men_n390_), .B0(men_men_n24_), .Y(men_men_n392_));
  OAI210     u370(.A0(men_men_n392_), .A1(men_men_n389_), .B0(men_men_n97_), .Y(men_men_n393_));
  NA2        u371(.A(x11), .B(men_men_n31_), .Y(men_men_n394_));
  NA2        u372(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n395_));
  NA2        u373(.A(men_men_n263_), .B(x03), .Y(men_men_n396_));
  OAI220     u374(.A0(men_men_n396_), .A1(men_men_n395_), .B0(men_men_n394_), .B1(men_men_n77_), .Y(men_men_n397_));
  OAI210     u375(.A0(men_men_n26_), .A1(men_men_n97_), .B0(x07), .Y(men_men_n398_));
  AOI210     u376(.A0(men_men_n397_), .A1(x06), .B0(men_men_n398_), .Y(men_men_n399_));
  AOI220     u377(.A0(men_men_n77_), .A1(men_men_n31_), .B0(men_men_n51_), .B1(men_men_n50_), .Y(men_men_n400_));
  NO3        u378(.A(men_men_n400_), .B(men_men_n23_), .C(x00), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n67_), .B(x02), .Y(men_men_n402_));
  AOI210     u380(.A0(men_men_n402_), .A1(men_men_n396_), .B0(men_men_n266_), .Y(men_men_n403_));
  OR2        u381(.A(men_men_n403_), .B(men_men_n249_), .Y(men_men_n404_));
  NO2        u382(.A(men_men_n23_), .B(x10), .Y(men_men_n405_));
  OAI210     u383(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n406_));
  OR3        u384(.A(men_men_n406_), .B(men_men_n405_), .C(men_men_n44_), .Y(men_men_n407_));
  NA2        u385(.A(men_men_n407_), .B(men_men_n404_), .Y(men_men_n408_));
  OAI210     u386(.A0(men_men_n408_), .A1(men_men_n401_), .B0(men_men_n97_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n33_), .B(men_men_n97_), .Y(men_men_n410_));
  AOI210     u388(.A0(men_men_n410_), .A1(men_men_n88_), .B0(x07), .Y(men_men_n411_));
  AOI220     u389(.A0(men_men_n411_), .A1(men_men_n409_), .B0(men_men_n399_), .B1(men_men_n393_), .Y(men_men_n412_));
  NA3        u390(.A(men_men_n23_), .B(men_men_n57_), .C(men_men_n48_), .Y(men_men_n413_));
  AO210      u391(.A0(men_men_n413_), .A1(men_men_n276_), .B0(men_men_n273_), .Y(men_men_n414_));
  AOI210     u392(.A0(men_men_n405_), .A1(x07), .B0(men_men_n142_), .Y(men_men_n415_));
  OR2        u393(.A(men_men_n415_), .B(x03), .Y(men_men_n416_));
  NO2        u394(.A(x07), .B(x11), .Y(men_men_n417_));
  NO3        u395(.A(men_men_n417_), .B(men_men_n146_), .C(men_men_n28_), .Y(men_men_n418_));
  AOI220     u396(.A0(men_men_n418_), .A1(men_men_n416_), .B0(men_men_n414_), .B1(men_men_n47_), .Y(men_men_n419_));
  NO3        u397(.A(men_men_n340_), .B(men_men_n32_), .C(x11), .Y(men_men_n420_));
  OAI210     u398(.A0(men_men_n420_), .A1(men_men_n419_), .B0(men_men_n98_), .Y(men_men_n421_));
  AOI210     u399(.A0(men_men_n349_), .A1(men_men_n109_), .B0(men_men_n272_), .Y(men_men_n422_));
  NOi21      u400(.An(men_men_n328_), .B(men_men_n133_), .Y(men_men_n423_));
  NO2        u401(.A(men_men_n423_), .B(men_men_n273_), .Y(men_men_n424_));
  OAI210     u402(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n425_));
  AOI210     u403(.A0(men_men_n258_), .A1(men_men_n47_), .B0(men_men_n425_), .Y(men_men_n426_));
  NO4        u404(.A(men_men_n426_), .B(men_men_n424_), .C(men_men_n422_), .D(x08), .Y(men_men_n427_));
  NO2        u405(.A(men_men_n405_), .B(men_men_n31_), .Y(men_men_n428_));
  OAI220     u406(.A0(x05), .A1(men_men_n428_), .B0(men_men_n394_), .B1(men_men_n63_), .Y(men_men_n429_));
  NO2        u407(.A(x13), .B(x12), .Y(men_men_n430_));
  NO2        u408(.A(men_men_n131_), .B(men_men_n28_), .Y(men_men_n431_));
  NO2        u409(.A(men_men_n431_), .B(men_men_n277_), .Y(men_men_n432_));
  OR3        u410(.A(men_men_n432_), .B(x12), .C(x03), .Y(men_men_n433_));
  NA3        u411(.A(men_men_n343_), .B(men_men_n124_), .C(x12), .Y(men_men_n434_));
  AO210      u412(.A0(men_men_n343_), .A1(men_men_n124_), .B0(men_men_n258_), .Y(men_men_n435_));
  NA4        u413(.A(men_men_n435_), .B(men_men_n434_), .C(men_men_n433_), .D(x08), .Y(men_men_n436_));
  AOI210     u414(.A0(men_men_n430_), .A1(men_men_n429_), .B0(men_men_n436_), .Y(men_men_n437_));
  AOI210     u415(.A0(men_men_n427_), .A1(men_men_n421_), .B0(men_men_n437_), .Y(men_men_n438_));
  OAI210     u416(.A0(x07), .A1(men_men_n23_), .B0(x03), .Y(men_men_n439_));
  NO2        u417(.A(men_men_n459_), .B(men_men_n395_), .Y(men_men_n440_));
  OAI210     u418(.A0(men_men_n440_), .A1(men_men_n439_), .B0(men_men_n193_), .Y(men_men_n441_));
  NA3        u419(.A(men_men_n432_), .B(men_men_n423_), .C(men_men_n339_), .Y(men_men_n442_));
  INV        u420(.A(x14), .Y(men_men_n443_));
  NO3        u421(.A(men_men_n328_), .B(men_men_n104_), .C(x11), .Y(men_men_n444_));
  NO3        u422(.A(men_men_n413_), .B(men_men_n340_), .C(men_men_n187_), .Y(men_men_n445_));
  NO3        u423(.A(men_men_n445_), .B(men_men_n444_), .C(men_men_n443_), .Y(men_men_n446_));
  NA3        u424(.A(men_men_n446_), .B(men_men_n442_), .C(men_men_n441_), .Y(men_men_n447_));
  AOI220     u425(.A0(men_men_n410_), .A1(men_men_n57_), .B0(men_men_n431_), .B1(men_men_n166_), .Y(men_men_n448_));
  NOi21      u426(.An(men_men_n282_), .B(men_men_n150_), .Y(men_men_n449_));
  NO3        u427(.A(men_men_n128_), .B(men_men_n24_), .C(x06), .Y(men_men_n450_));
  AOI210     u428(.A0(men_men_n289_), .A1(men_men_n241_), .B0(men_men_n450_), .Y(men_men_n451_));
  OAI210     u429(.A0(men_men_n44_), .A1(x04), .B0(men_men_n451_), .Y(men_men_n452_));
  OAI210     u430(.A0(men_men_n452_), .A1(men_men_n449_), .B0(men_men_n97_), .Y(men_men_n453_));
  OAI210     u431(.A0(men_men_n448_), .A1(men_men_n87_), .B0(men_men_n453_), .Y(men_men_n454_));
  NO4        u432(.A(men_men_n454_), .B(men_men_n447_), .C(men_men_n438_), .D(men_men_n412_), .Y(men06));
  INV        u433(.A(x07), .Y(men_men_n458_));
  INV        u434(.A(x07), .Y(men_men_n459_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule