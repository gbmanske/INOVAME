//Benchmark atmr_intb_466_0.0625

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n319_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n370_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n339_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n362_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  AOI220     o039(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o040(.A(ori_ori_n59_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n64_), .B(ori_ori_n24_), .Y(ori_ori_n65_));
  OAI220     o043(.A0(ori_ori_n65_), .A1(ori_ori_n63_), .B0(ori_ori_n62_), .B1(ori_ori_n60_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n67_));
  OAI210     o045(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n67_), .Y(ori_ori_n68_));
  AOI220     o046(.A0(ori_ori_n68_), .A1(ori_ori_n59_), .B0(ori_ori_n66_), .B1(ori_ori_n31_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(ori_ori_n69_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n61_), .B(ori_ori_n23_), .Y(ori_ori_n71_));
  NA2        o049(.A(x09), .B(x05), .Y(ori_ori_n72_));
  NA2        o050(.A(x10), .B(x06), .Y(ori_ori_n73_));
  NA2        o051(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n74_), .A1(ori_ori_n71_), .B0(x03), .Y(ori_ori_n76_));
  NOi31      o054(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n77_));
  NO2        o055(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n36_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n80_));
  NO2        o058(.A(x08), .B(x01), .Y(ori_ori_n81_));
  OAI210     o059(.A0(ori_ori_n81_), .A1(ori_ori_n80_), .B0(ori_ori_n35_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n82_), .B(x02), .Y(ori_ori_n83_));
  AN2        o061(.A(ori_ori_n83_), .B(ori_ori_n76_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n82_), .Y(ori_ori_n85_));
  NA2        o063(.A(x11), .B(x00), .Y(ori_ori_n86_));
  NO2        o064(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n87_));
  NOi21      o065(.An(ori_ori_n86_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  INV        o066(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  NOi21      o067(.An(x01), .B(x10), .Y(ori_ori_n90_));
  NO2        o068(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n91_));
  NO3        o069(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(x06), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n92_), .B(ori_ori_n27_), .Y(ori_ori_n93_));
  OAI210     o071(.A0(ori_ori_n89_), .A1(x07), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NO3        o072(.A(ori_ori_n94_), .B(ori_ori_n84_), .C(ori_ori_n70_), .Y(ori01));
  INV        o073(.A(x12), .Y(ori_ori_n96_));
  INV        o074(.A(x13), .Y(ori_ori_n97_));
  NA2        o075(.A(x08), .B(x04), .Y(ori_ori_n98_));
  NO2        o076(.A(x10), .B(x01), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n100_), .B(ori_ori_n99_), .Y(ori_ori_n101_));
  NA2        o079(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n103_));
  NA2        o081(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n104_));
  NA2        o082(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n105_), .B(x05), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n108_));
  NA2        o086(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n109_), .B(ori_ori_n108_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n112_));
  NA3        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .C(x13), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n114_));
  NOi31      o092(.An(ori_ori_n113_), .B(ori_ori_n114_), .C(ori_ori_n110_), .Y(ori_ori_n115_));
  NO3        o093(.A(ori_ori_n115_), .B(x06), .C(x03), .Y(ori_ori_n116_));
  INV        o094(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NA2        o095(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n118_));
  OAI210     o096(.A0(ori_ori_n81_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n122_));
  AOI210     o100(.A0(ori_ori_n122_), .A1(ori_ori_n49_), .B0(ori_ori_n121_), .Y(ori_ori_n123_));
  AN2        o101(.A(ori_ori_n123_), .B(ori_ori_n120_), .Y(ori_ori_n124_));
  NO2        o102(.A(x09), .B(x05), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(ori_ori_n47_), .Y(ori_ori_n126_));
  AOI210     o104(.A0(ori_ori_n126_), .A1(ori_ori_n101_), .B0(ori_ori_n49_), .Y(ori_ori_n127_));
  NA2        o105(.A(x09), .B(x00), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n103_), .B(ori_ori_n128_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n127_), .B(ori_ori_n124_), .Y(ori_ori_n130_));
  NO2        o108(.A(x03), .B(x02), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n82_), .B(ori_ori_n97_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n131_), .Y(ori_ori_n133_));
  OA210      o111(.A0(ori_ori_n130_), .A1(x11), .B0(ori_ori_n133_), .Y(ori_ori_n134_));
  OAI210     o112(.A0(ori_ori_n117_), .A1(ori_ori_n23_), .B0(ori_ori_n134_), .Y(ori_ori_n135_));
  NAi21      o113(.An(x06), .B(x10), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n97_), .B(x01), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n138_), .B(x08), .Y(ori_ori_n139_));
  OAI210     o117(.A0(x05), .A1(ori_ori_n139_), .B0(ori_ori_n51_), .Y(ori_ori_n140_));
  AOI210     o118(.A0(ori_ori_n140_), .A1(ori_ori_n137_), .B0(ori_ori_n48_), .Y(ori_ori_n141_));
  AOI210     o119(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n141_), .B(ori_ori_n142_), .Y(ori_ori_n143_));
  NA2        o121(.A(x10), .B(x05), .Y(ori_ori_n144_));
  NO2        o122(.A(x09), .B(x01), .Y(ori_ori_n145_));
  INV        o123(.A(ori_ori_n25_), .Y(ori_ori_n146_));
  NAi21      o124(.An(x13), .B(x00), .Y(ori_ori_n147_));
  AN2        o125(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n91_), .B(x06), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n147_), .B(ori_ori_n36_), .Y(ori_ori_n150_));
  INV        o128(.A(ori_ori_n150_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n149_), .B(ori_ori_n148_), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n152_), .B(ori_ori_n146_), .Y(ori_ori_n153_));
  NOi21      o131(.An(x09), .B(x00), .Y(ori_ori_n154_));
  NO3        o132(.A(ori_ori_n80_), .B(ori_ori_n154_), .C(ori_ori_n47_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n155_), .B(ori_ori_n109_), .Y(ori_ori_n156_));
  NA2        o134(.A(x10), .B(x08), .Y(ori_ori_n157_));
  INV        o135(.A(ori_ori_n157_), .Y(ori_ori_n158_));
  NA2        o136(.A(x06), .B(x05), .Y(ori_ori_n159_));
  OAI210     o137(.A0(ori_ori_n159_), .A1(ori_ori_n35_), .B0(ori_ori_n96_), .Y(ori_ori_n160_));
  AOI210     o138(.A0(ori_ori_n158_), .A1(ori_ori_n58_), .B0(ori_ori_n160_), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n161_), .B(ori_ori_n156_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n97_), .B(x12), .Y(ori_ori_n163_));
  AOI210     o141(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n163_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n90_), .B(ori_ori_n51_), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n166_), .B(x02), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n164_), .B(ori_ori_n162_), .Y(ori_ori_n168_));
  NA3        o146(.A(ori_ori_n168_), .B(ori_ori_n153_), .C(ori_ori_n143_), .Y(ori_ori_n169_));
  AOI210     o147(.A0(ori_ori_n135_), .A1(ori_ori_n96_), .B0(ori_ori_n169_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n28_), .B(ori_ori_n120_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(ori_ori_n119_), .Y(ori_ori_n173_));
  AOI210     o151(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n108_), .B(x06), .Y(ori_ori_n175_));
  AOI210     o153(.A0(ori_ori_n174_), .A1(ori_ori_n173_), .B0(ori_ori_n175_), .Y(ori_ori_n176_));
  AOI210     o154(.A0(ori_ori_n176_), .A1(ori_ori_n171_), .B0(x12), .Y(ori_ori_n177_));
  INV        o155(.A(ori_ori_n77_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n90_), .B(x06), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n180_));
  NO3        o158(.A(ori_ori_n180_), .B(ori_ori_n179_), .C(ori_ori_n41_), .Y(ori_ori_n181_));
  INV        o159(.A(ori_ori_n122_), .Y(ori_ori_n182_));
  OAI210     o160(.A0(ori_ori_n182_), .A1(ori_ori_n181_), .B0(x02), .Y(ori_ori_n183_));
  AOI210     o161(.A0(ori_ori_n183_), .A1(ori_ori_n57_), .B0(ori_ori_n23_), .Y(ori_ori_n184_));
  OAI210     o162(.A0(ori_ori_n177_), .A1(ori_ori_n57_), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  INV        o163(.A(ori_ori_n122_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n187_));
  OAI210     o165(.A0(ori_ori_n78_), .A1(ori_ori_n36_), .B0(ori_ori_n104_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n97_), .B(x03), .Y(ori_ori_n189_));
  AOI220     o167(.A0(ori_ori_n189_), .A1(ori_ori_n188_), .B0(ori_ori_n77_), .B1(ori_ori_n187_), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n191_));
  INV        o169(.A(ori_ori_n136_), .Y(ori_ori_n192_));
  NOi21      o170(.An(x13), .B(x04), .Y(ori_ori_n193_));
  NO3        o171(.A(ori_ori_n193_), .B(ori_ori_n77_), .C(ori_ori_n154_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n194_), .B(x05), .Y(ori_ori_n195_));
  AOI220     o173(.A0(ori_ori_n195_), .A1(ori_ori_n191_), .B0(ori_ori_n192_), .B1(ori_ori_n57_), .Y(ori_ori_n196_));
  OAI210     o174(.A0(ori_ori_n190_), .A1(ori_ori_n186_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  INV        o175(.A(ori_ori_n87_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n198_), .B(x12), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n200_));
  NO2        o178(.A(x06), .B(x00), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n41_), .Y(ori_ori_n202_));
  INV        o180(.A(ori_ori_n73_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n203_), .B(ori_ori_n202_), .Y(ori_ori_n204_));
  NA2        o182(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n205_), .B(x03), .Y(ori_ori_n206_));
  OR2        o184(.A(ori_ori_n206_), .B(ori_ori_n204_), .Y(ori_ori_n207_));
  NA2        o185(.A(x13), .B(ori_ori_n96_), .Y(ori_ori_n208_));
  NA3        o186(.A(ori_ori_n208_), .B(ori_ori_n160_), .C(ori_ori_n88_), .Y(ori_ori_n209_));
  OAI210     o187(.A0(ori_ori_n207_), .A1(ori_ori_n200_), .B0(ori_ori_n209_), .Y(ori_ori_n210_));
  AOI210     o188(.A0(ori_ori_n199_), .A1(ori_ori_n197_), .B0(ori_ori_n210_), .Y(ori_ori_n211_));
  AOI210     o189(.A0(ori_ori_n211_), .A1(ori_ori_n185_), .B0(x07), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n72_), .B(ori_ori_n29_), .Y(ori_ori_n213_));
  NOi31      o191(.An(ori_ori_n118_), .B(ori_ori_n193_), .C(ori_ori_n154_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n214_), .B(ori_ori_n213_), .Y(ori_ori_n215_));
  NO2        o193(.A(x08), .B(x05), .Y(ori_ori_n216_));
  OAI210     o194(.A0(ori_ori_n77_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n217_));
  INV        o195(.A(ori_ori_n217_), .Y(ori_ori_n218_));
  NO2        o196(.A(x12), .B(x02), .Y(ori_ori_n219_));
  INV        o197(.A(ori_ori_n219_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(ori_ori_n198_), .Y(ori_ori_n221_));
  OA210      o199(.A0(ori_ori_n218_), .A1(ori_ori_n215_), .B0(ori_ori_n221_), .Y(ori_ori_n222_));
  NA2        o200(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(x01), .Y(ori_ori_n224_));
  INV        o202(.A(ori_ori_n224_), .Y(ori_ori_n225_));
  AOI210     o203(.A0(ori_ori_n225_), .A1(ori_ori_n113_), .B0(ori_ori_n29_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n97_), .B(x04), .Y(ori_ori_n227_));
  NO3        o205(.A(ori_ori_n86_), .B(x12), .C(x03), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n226_), .B(ori_ori_n228_), .Y(ori_ori_n229_));
  AOI210     o207(.A0(ori_ori_n165_), .A1(ori_ori_n159_), .B0(ori_ori_n98_), .Y(ori_ori_n230_));
  NOi21      o208(.An(ori_ori_n213_), .B(ori_ori_n179_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n232_));
  OAI210     o210(.A0(ori_ori_n231_), .A1(ori_ori_n230_), .B0(ori_ori_n232_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n234_));
  NO3        o212(.A(ori_ori_n234_), .B(ori_ori_n180_), .C(ori_ori_n149_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n200_), .B(ori_ori_n28_), .Y(ori_ori_n236_));
  OAI210     o214(.A0(ori_ori_n235_), .A1(ori_ori_n186_), .B0(ori_ori_n236_), .Y(ori_ori_n237_));
  NA3        o215(.A(ori_ori_n237_), .B(ori_ori_n233_), .C(ori_ori_n229_), .Y(ori_ori_n238_));
  NO3        o216(.A(ori_ori_n238_), .B(ori_ori_n222_), .C(ori_ori_n212_), .Y(ori_ori_n239_));
  OAI210     o217(.A0(ori_ori_n170_), .A1(ori_ori_n61_), .B0(ori_ori_n239_), .Y(ori02));
  AOI210     o218(.A0(ori_ori_n118_), .A1(ori_ori_n82_), .B0(ori_ori_n111_), .Y(ori_ori_n241_));
  NOi21      o219(.An(ori_ori_n194_), .B(ori_ori_n145_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n97_), .B(ori_ori_n35_), .Y(ori_ori_n243_));
  NA3        o221(.A(ori_ori_n243_), .B(ori_ori_n158_), .C(ori_ori_n56_), .Y(ori_ori_n244_));
  OAI210     o222(.A0(ori_ori_n242_), .A1(ori_ori_n32_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  OAI210     o223(.A0(ori_ori_n245_), .A1(ori_ori_n241_), .B0(ori_ori_n144_), .Y(ori_ori_n246_));
  INV        o224(.A(ori_ori_n144_), .Y(ori_ori_n247_));
  NO2        o225(.A(ori_ori_n82_), .B(ori_ori_n51_), .Y(ori_ori_n248_));
  AOI220     o226(.A0(ori_ori_n248_), .A1(ori_ori_n247_), .B0(ori_ori_n132_), .B1(ori_ori_n131_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n249_), .A1(ori_ori_n246_), .B0(ori_ori_n48_), .Y(ori_ori_n250_));
  NO2        o228(.A(x05), .B(x02), .Y(ori_ori_n251_));
  OAI210     o229(.A0(ori_ori_n173_), .A1(ori_ori_n154_), .B0(ori_ori_n251_), .Y(ori_ori_n252_));
  AOI220     o230(.A0(ori_ori_n216_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n253_));
  NOi21      o231(.An(ori_ori_n243_), .B(ori_ori_n253_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n193_), .A1(ori_ori_n78_), .B0(ori_ori_n254_), .Y(ori_ori_n255_));
  AOI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n252_), .B0(ori_ori_n122_), .Y(ori_ori_n256_));
  NAi21      o234(.An(ori_ori_n195_), .B(ori_ori_n190_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n205_), .B(ori_ori_n47_), .Y(ori_ori_n258_));
  NA2        o236(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  AN2        o237(.A(ori_ori_n189_), .B(ori_ori_n188_), .Y(ori_ori_n260_));
  OAI210     o238(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n261_));
  NA2        o239(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n262_));
  BUFFER     o240(.A(ori_ori_n126_), .Y(ori_ori_n263_));
  AOI210     o241(.A0(ori_ori_n263_), .A1(ori_ori_n119_), .B0(ori_ori_n261_), .Y(ori_ori_n264_));
  OAI210     o242(.A0(ori_ori_n264_), .A1(ori_ori_n260_), .B0(ori_ori_n91_), .Y(ori_ori_n265_));
  INV        o243(.A(ori_ori_n131_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n266_), .B(ori_ori_n110_), .Y(ori_ori_n267_));
  NA2        o245(.A(ori_ori_n267_), .B(x13), .Y(ori_ori_n268_));
  NA3        o246(.A(ori_ori_n268_), .B(ori_ori_n265_), .C(ori_ori_n259_), .Y(ori_ori_n269_));
  NO3        o247(.A(ori_ori_n269_), .B(ori_ori_n256_), .C(ori_ori_n250_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n121_), .B(x03), .Y(ori_ori_n271_));
  OAI210     o249(.A0(ori_ori_n35_), .A1(ori_ori_n234_), .B0(ori_ori_n271_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n272_), .B(ori_ori_n99_), .Y(ori_ori_n273_));
  INV        o251(.A(ori_ori_n56_), .Y(ori_ori_n274_));
  OAI220     o252(.A0(ori_ori_n227_), .A1(ori_ori_n274_), .B0(ori_ori_n111_), .B1(ori_ori_n28_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n275_), .B(ori_ori_n100_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n227_), .B(ori_ori_n96_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n96_), .B(ori_ori_n41_), .Y(ori_ori_n278_));
  NA3        o256(.A(ori_ori_n278_), .B(ori_ori_n277_), .C(ori_ori_n110_), .Y(ori_ori_n279_));
  NA4        o257(.A(ori_ori_n279_), .B(ori_ori_n276_), .C(ori_ori_n273_), .D(ori_ori_n48_), .Y(ori_ori_n280_));
  INV        o258(.A(ori_ori_n166_), .Y(ori_ori_n281_));
  OAI220     o259(.A0(ori_ori_n370_), .A1(ori_ori_n31_), .B0(ori_ori_n281_), .B1(ori_ori_n59_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(x02), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n163_), .B(x04), .Y(ori_ori_n284_));
  NO3        o262(.A(ori_ori_n163_), .B(ori_ori_n137_), .C(ori_ori_n52_), .Y(ori_ori_n285_));
  OAI210     o263(.A0(ori_ori_n128_), .A1(ori_ori_n36_), .B0(ori_ori_n96_), .Y(ori_ori_n286_));
  OAI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n155_), .B0(ori_ori_n285_), .Y(ori_ori_n287_));
  NA3        o265(.A(ori_ori_n287_), .B(ori_ori_n283_), .C(x06), .Y(ori_ori_n288_));
  NA2        o266(.A(x09), .B(x03), .Y(ori_ori_n289_));
  OAI220     o267(.A0(ori_ori_n289_), .A1(ori_ori_n109_), .B0(ori_ori_n172_), .B1(ori_ori_n64_), .Y(ori_ori_n290_));
  OAI220     o268(.A0(ori_ori_n138_), .A1(x09), .B0(x08), .B1(ori_ori_n41_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n291_), .B(ori_ori_n186_), .Y(ori_ori_n292_));
  NO2        o270(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n293_));
  NO3        o271(.A(ori_ori_n103_), .B(ori_ori_n109_), .C(ori_ori_n38_), .Y(ori_ori_n294_));
  AOI210     o272(.A0(ori_ori_n285_), .A1(ori_ori_n293_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  OAI210     o273(.A0(ori_ori_n292_), .A1(ori_ori_n28_), .B0(ori_ori_n295_), .Y(ori_ori_n296_));
  AO220      o274(.A0(ori_ori_n296_), .A1(x04), .B0(ori_ori_n290_), .B1(x05), .Y(ori_ori_n297_));
  AOI210     o275(.A0(ori_ori_n288_), .A1(ori_ori_n280_), .B0(ori_ori_n297_), .Y(ori_ori_n298_));
  OAI210     o276(.A0(ori_ori_n270_), .A1(x12), .B0(ori_ori_n298_), .Y(ori03));
  OR2        o277(.A(ori_ori_n42_), .B(ori_ori_n187_), .Y(ori_ori_n300_));
  AOI210     o278(.A0(ori_ori_n132_), .A1(ori_ori_n96_), .B0(ori_ori_n300_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n163_), .B(ori_ori_n131_), .Y(ori_ori_n302_));
  NA2        o280(.A(ori_ori_n302_), .B(ori_ori_n167_), .Y(ori_ori_n303_));
  OAI210     o281(.A0(ori_ori_n303_), .A1(ori_ori_n301_), .B0(x05), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n300_), .B(x05), .Y(ori_ori_n305_));
  AOI210     o283(.A0(ori_ori_n119_), .A1(ori_ori_n178_), .B0(ori_ori_n305_), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n189_), .A1(ori_ori_n79_), .B0(ori_ori_n106_), .Y(ori_ori_n307_));
  OAI220     o285(.A0(ori_ori_n307_), .A1(ori_ori_n59_), .B0(ori_ori_n262_), .B1(ori_ori_n253_), .Y(ori_ori_n308_));
  OAI210     o286(.A0(ori_ori_n308_), .A1(ori_ori_n306_), .B0(ori_ori_n96_), .Y(ori_ori_n309_));
  AOI210     o287(.A0(ori_ori_n126_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n145_), .B(ori_ori_n114_), .Y(ori_ori_n311_));
  OAI220     o289(.A0(ori_ori_n311_), .A1(ori_ori_n37_), .B0(ori_ori_n129_), .B1(x13), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n310_), .B0(x04), .Y(ori_ori_n313_));
  NO3        o291(.A(ori_ori_n278_), .B(ori_ori_n82_), .C(ori_ori_n59_), .Y(ori_ori_n314_));
  AOI210     o292(.A0(ori_ori_n151_), .A1(ori_ori_n96_), .B0(ori_ori_n126_), .Y(ori_ori_n315_));
  OA210      o293(.A0(ori_ori_n139_), .A1(x12), .B0(ori_ori_n114_), .Y(ori_ori_n316_));
  NO3        o294(.A(ori_ori_n316_), .B(ori_ori_n315_), .C(ori_ori_n314_), .Y(ori_ori_n317_));
  NA4        o295(.A(ori_ori_n317_), .B(ori_ori_n313_), .C(ori_ori_n309_), .D(ori_ori_n304_), .Y(ori04));
  NO2        o296(.A(ori_ori_n85_), .B(ori_ori_n39_), .Y(ori_ori_n319_));
  XO2        o297(.A(ori_ori_n319_), .B(ori_ori_n208_), .Y(ori05));
  AOI210     o298(.A0(ori_ori_n72_), .A1(ori_ori_n52_), .B0(ori_ori_n175_), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n321_), .A1(ori_ori_n261_), .B0(ori_ori_n25_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n111_), .B(ori_ori_n31_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n192_), .B(ori_ori_n57_), .Y(ori_ori_n324_));
  AOI210     o302(.A0(ori_ori_n324_), .A1(ori_ori_n323_), .B0(ori_ori_n24_), .Y(ori_ori_n325_));
  OAI210     o303(.A0(ori_ori_n325_), .A1(ori_ori_n322_), .B0(ori_ori_n96_), .Y(ori_ori_n326_));
  OAI210     o304(.A0(ori_ori_n26_), .A1(ori_ori_n96_), .B0(x07), .Y(ori_ori_n327_));
  INV        o305(.A(ori_ori_n327_), .Y(ori_ori_n328_));
  NO2        o306(.A(ori_ori_n31_), .B(ori_ori_n52_), .Y(ori_ori_n329_));
  NO3        o307(.A(ori_ori_n329_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n330_));
  OR2        o308(.A(x03), .B(ori_ori_n200_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n201_), .B(ori_ori_n198_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n332_), .B(ori_ori_n331_), .Y(ori_ori_n333_));
  OAI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n330_), .B0(ori_ori_n96_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n33_), .B(ori_ori_n96_), .Y(ori_ori_n335_));
  AOI210     o313(.A0(ori_ori_n335_), .A1(ori_ori_n87_), .B0(x07), .Y(ori_ori_n336_));
  AOI220     o314(.A0(ori_ori_n336_), .A1(ori_ori_n334_), .B0(ori_ori_n328_), .B1(ori_ori_n326_), .Y(ori_ori_n337_));
  AOI210     o315(.A0(ori_ori_n284_), .A1(ori_ori_n102_), .B0(ori_ori_n219_), .Y(ori_ori_n338_));
  NOi21      o316(.An(ori_ori_n271_), .B(ori_ori_n114_), .Y(ori_ori_n339_));
  NO2        o317(.A(ori_ori_n339_), .B(ori_ori_n220_), .Y(ori_ori_n340_));
  OAI210     o318(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n341_));
  AOI210     o319(.A0(ori_ori_n208_), .A1(ori_ori_n47_), .B0(ori_ori_n341_), .Y(ori_ori_n342_));
  NO4        o320(.A(ori_ori_n342_), .B(ori_ori_n340_), .C(ori_ori_n338_), .D(x08), .Y(ori_ori_n343_));
  NO2        o321(.A(x05), .B(x03), .Y(ori_ori_n344_));
  NO2        o322(.A(x13), .B(x12), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n111_), .B(ori_ori_n28_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n346_), .B(ori_ori_n224_), .Y(ori_ori_n347_));
  OR3        o325(.A(ori_ori_n347_), .B(x12), .C(x03), .Y(ori_ori_n348_));
  NA3        o326(.A(ori_ori_n281_), .B(ori_ori_n107_), .C(x12), .Y(ori_ori_n349_));
  AO210      o327(.A0(ori_ori_n281_), .A1(ori_ori_n107_), .B0(ori_ori_n208_), .Y(ori_ori_n350_));
  NA4        o328(.A(ori_ori_n350_), .B(ori_ori_n349_), .C(ori_ori_n348_), .D(x08), .Y(ori_ori_n351_));
  AOI210     o329(.A0(ori_ori_n345_), .A1(ori_ori_n344_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n343_), .B(ori_ori_n352_), .Y(ori_ori_n353_));
  NO2        o331(.A(ori_ori_n125_), .B(ori_ori_n43_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n354_), .B(ori_ori_n150_), .Y(ori_ori_n355_));
  NA3        o333(.A(ori_ori_n347_), .B(ori_ori_n339_), .C(ori_ori_n277_), .Y(ori_ori_n356_));
  INV        o334(.A(x14), .Y(ori_ori_n357_));
  NO3        o335(.A(ori_ori_n138_), .B(ori_ori_n75_), .C(ori_ori_n57_), .Y(ori_ori_n358_));
  NO2        o336(.A(ori_ori_n358_), .B(ori_ori_n357_), .Y(ori_ori_n359_));
  NA3        o337(.A(ori_ori_n359_), .B(ori_ori_n356_), .C(ori_ori_n355_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n335_), .B(ori_ori_n61_), .Y(ori_ori_n361_));
  NOi21      o339(.An(ori_ori_n227_), .B(ori_ori_n129_), .Y(ori_ori_n362_));
  NA2        o340(.A(ori_ori_n232_), .B(ori_ori_n192_), .Y(ori_ori_n363_));
  OAI210     o341(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  OAI210     o342(.A0(ori_ori_n364_), .A1(ori_ori_n362_), .B0(ori_ori_n96_), .Y(ori_ori_n365_));
  OAI210     o343(.A0(ori_ori_n361_), .A1(ori_ori_n86_), .B0(ori_ori_n365_), .Y(ori_ori_n366_));
  NO4        o344(.A(ori_ori_n366_), .B(ori_ori_n360_), .C(ori_ori_n353_), .D(ori_ori_n337_), .Y(ori06));
  INV        o345(.A(x05), .Y(ori_ori_n370_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NOi21      m029(.An(x01), .B(x09), .Y(mai_mai_n52_));
  INV        m030(.A(x00), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  NO2        m032(.A(mai_mai_n54_), .B(mai_mai_n52_), .Y(mai_mai_n55_));
  NA2        m033(.A(x09), .B(mai_mai_n53_), .Y(mai_mai_n56_));
  INV        m034(.A(x07), .Y(mai_mai_n57_));
  AOI210     m035(.A0(x11), .A1(mai_mai_n48_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  INV        m036(.A(mai_mai_n55_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n60_), .B(mai_mai_n24_), .Y(mai_mai_n61_));
  OAI220     m039(.A0(mai_mai_n61_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .B1(mai_mai_n56_), .Y(mai_mai_n62_));
  NO2        m040(.A(mai_mai_n30_), .B(x11), .Y(mai_mai_n63_));
  AOI220     m041(.A0(mai_mai_n63_), .A1(mai_mai_n55_), .B0(mai_mai_n62_), .B1(mai_mai_n31_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(x05), .Y(mai_mai_n65_));
  NA2        m043(.A(x09), .B(x05), .Y(mai_mai_n66_));
  NA2        m044(.A(x10), .B(x06), .Y(mai_mai_n67_));
  NA2        m045(.A(mai_mai_n67_), .B(mai_mai_n66_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n57_), .B(mai_mai_n41_), .Y(mai_mai_n69_));
  OAI210     m047(.A0(mai_mai_n68_), .A1(x07), .B0(x03), .Y(mai_mai_n70_));
  NOi31      m048(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n71_));
  NO2        m049(.A(mai_mai_n403_), .B(mai_mai_n24_), .Y(mai_mai_n72_));
  NO2        m050(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n36_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n73_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n75_));
  AOI210     m053(.A0(mai_mai_n74_), .A1(mai_mai_n48_), .B0(mai_mai_n75_), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n77_));
  NO2        m055(.A(x08), .B(x01), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n78_), .A1(mai_mai_n77_), .B0(mai_mai_n35_), .Y(mai_mai_n79_));
  NA2        m057(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n79_), .B(mai_mai_n76_), .C(mai_mai_n72_), .Y(mai_mai_n81_));
  AN2        m059(.A(mai_mai_n81_), .B(mai_mai_n70_), .Y(mai_mai_n82_));
  INV        m060(.A(mai_mai_n79_), .Y(mai_mai_n83_));
  NA2        m061(.A(x11), .B(x00), .Y(mai_mai_n84_));
  NO2        m062(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n85_));
  NOi21      m063(.An(mai_mai_n84_), .B(mai_mai_n85_), .Y(mai_mai_n86_));
  INV        m064(.A(mai_mai_n86_), .Y(mai_mai_n87_));
  NOi21      m065(.An(x01), .B(x10), .Y(mai_mai_n88_));
  NO2        m066(.A(mai_mai_n29_), .B(mai_mai_n53_), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(x06), .Y(mai_mai_n90_));
  NA2        m068(.A(mai_mai_n90_), .B(mai_mai_n27_), .Y(mai_mai_n91_));
  OAI210     m069(.A0(mai_mai_n87_), .A1(x07), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NO3        m070(.A(mai_mai_n92_), .B(mai_mai_n82_), .C(mai_mai_n65_), .Y(mai01));
  INV        m071(.A(x12), .Y(mai_mai_n94_));
  INV        m072(.A(x13), .Y(mai_mai_n95_));
  NA2        m073(.A(x08), .B(x04), .Y(mai_mai_n96_));
  NA2        m074(.A(mai_mai_n88_), .B(mai_mai_n28_), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n97_), .B(mai_mai_n66_), .Y(mai_mai_n98_));
  NO2        m076(.A(x10), .B(x01), .Y(mai_mai_n99_));
  NO2        m077(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NA2        m079(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(mai_mai_n36_), .Y(mai_mai_n103_));
  AOI210     m081(.A0(mai_mai_n103_), .A1(mai_mai_n101_), .B0(mai_mai_n98_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n104_), .B(mai_mai_n95_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n52_), .B(x05), .Y(mai_mai_n106_));
  NOi21      m084(.An(mai_mai_n106_), .B(mai_mai_n54_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n108_));
  NA3        m086(.A(x13), .B(mai_mai_n108_), .C(x06), .Y(mai_mai_n109_));
  INV        m087(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n78_), .B(x13), .Y(mai_mai_n111_));
  NA2        m089(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n113_));
  NA2        m091(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n114_), .B(x05), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n113_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n35_), .B(mai_mai_n53_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(mai_mai_n95_), .Y(mai_mai_n118_));
  AOI210     m096(.A0(mai_mai_n118_), .A1(mai_mai_n74_), .B0(mai_mai_n107_), .Y(mai_mai_n119_));
  AOI210     m097(.A0(mai_mai_n119_), .A1(mai_mai_n116_), .B0(mai_mai_n67_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n121_));
  NA2        m099(.A(x10), .B(mai_mai_n53_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n122_), .B(mai_mai_n121_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n124_));
  NO3        m102(.A(mai_mai_n117_), .B(mai_mai_n73_), .C(mai_mai_n36_), .Y(mai_mai_n125_));
  NO2        m103(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n126_));
  NO3        m104(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n123_), .Y(mai_mai_n127_));
  NO3        m105(.A(mai_mai_n127_), .B(x06), .C(x03), .Y(mai_mai_n128_));
  NO4        m106(.A(mai_mai_n128_), .B(mai_mai_n120_), .C(mai_mai_n110_), .D(mai_mai_n105_), .Y(mai_mai_n129_));
  OAI210     m107(.A0(mai_mai_n78_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n132_));
  NO2        m110(.A(x09), .B(x05), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n47_), .Y(mai_mai_n134_));
  NO2        m112(.A(mai_mai_n101_), .B(mai_mai_n49_), .Y(mai_mai_n135_));
  NA2        m113(.A(x09), .B(x00), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n106_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  INV        m115(.A(mai_mai_n71_), .Y(mai_mai_n138_));
  AOI210     m116(.A0(mai_mai_n138_), .A1(mai_mai_n137_), .B0(mai_mai_n132_), .Y(mai_mai_n139_));
  NO2        m117(.A(mai_mai_n139_), .B(mai_mai_n135_), .Y(mai_mai_n140_));
  NO2        m118(.A(x03), .B(x02), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n79_), .B(mai_mai_n95_), .Y(mai_mai_n142_));
  OAI210     m120(.A0(mai_mai_n142_), .A1(mai_mai_n107_), .B0(mai_mai_n141_), .Y(mai_mai_n143_));
  OA210      m121(.A0(mai_mai_n140_), .A1(x11), .B0(mai_mai_n143_), .Y(mai_mai_n144_));
  OAI210     m122(.A0(mai_mai_n129_), .A1(mai_mai_n23_), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n101_), .B(mai_mai_n40_), .Y(mai_mai_n146_));
  NOi21      m124(.An(x01), .B(x13), .Y(mai_mai_n147_));
  AOI210     m125(.A0(mai_mai_n407_), .A1(mai_mai_n146_), .B0(mai_mai_n41_), .Y(mai_mai_n148_));
  NO2        m126(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n95_), .B(x01), .Y(mai_mai_n150_));
  NO2        m128(.A(mai_mai_n150_), .B(x08), .Y(mai_mai_n151_));
  NO2        m129(.A(mai_mai_n149_), .B(mai_mai_n48_), .Y(mai_mai_n152_));
  AOI210     m130(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n153_));
  OAI210     m131(.A0(mai_mai_n152_), .A1(mai_mai_n148_), .B0(mai_mai_n153_), .Y(mai_mai_n154_));
  NA2        m132(.A(x04), .B(x02), .Y(mai_mai_n155_));
  NA2        m133(.A(x10), .B(x05), .Y(mai_mai_n156_));
  NA2        m134(.A(x09), .B(x06), .Y(mai_mai_n157_));
  NO2        m135(.A(x09), .B(x01), .Y(mai_mai_n158_));
  NO3        m136(.A(mai_mai_n158_), .B(mai_mai_n99_), .C(mai_mai_n31_), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n159_), .B(x00), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n106_), .B(x08), .Y(mai_mai_n161_));
  OAI210     m139(.A0(mai_mai_n405_), .A1(x11), .B0(mai_mai_n160_), .Y(mai_mai_n162_));
  NAi21      m140(.An(mai_mai_n155_), .B(mai_mai_n162_), .Y(mai_mai_n163_));
  INV        m141(.A(mai_mai_n25_), .Y(mai_mai_n164_));
  NAi21      m142(.An(x13), .B(x00), .Y(mai_mai_n165_));
  AOI210     m143(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n165_), .Y(mai_mai_n166_));
  AOI220     m144(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n167_));
  OAI210     m145(.A0(mai_mai_n156_), .A1(mai_mai_n35_), .B0(mai_mai_n167_), .Y(mai_mai_n168_));
  AN2        m146(.A(mai_mai_n168_), .B(mai_mai_n166_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n89_), .B(x06), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n165_), .B(mai_mai_n36_), .Y(mai_mai_n171_));
  INV        m149(.A(mai_mai_n171_), .Y(mai_mai_n172_));
  OAI210     m150(.A0(mai_mai_n172_), .A1(mai_mai_n157_), .B0(mai_mai_n67_), .Y(mai_mai_n173_));
  OAI210     m151(.A0(mai_mai_n173_), .A1(mai_mai_n169_), .B0(mai_mai_n164_), .Y(mai_mai_n174_));
  NOi21      m152(.An(x09), .B(x00), .Y(mai_mai_n175_));
  NO3        m153(.A(mai_mai_n77_), .B(mai_mai_n175_), .C(mai_mai_n47_), .Y(mai_mai_n176_));
  INV        m154(.A(mai_mai_n176_), .Y(mai_mai_n177_));
  INV        m155(.A(x12), .Y(mai_mai_n178_));
  NA2        m156(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n95_), .B(x12), .Y(mai_mai_n180_));
  AOI210     m158(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n180_), .Y(mai_mai_n181_));
  INV        m159(.A(mai_mai_n88_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n183_));
  NA2        m161(.A(mai_mai_n183_), .B(x02), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n184_), .B(mai_mai_n182_), .Y(mai_mai_n185_));
  AOI210     m163(.A0(mai_mai_n181_), .A1(mai_mai_n179_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NA4        m164(.A(mai_mai_n186_), .B(mai_mai_n174_), .C(mai_mai_n163_), .D(mai_mai_n154_), .Y(mai_mai_n187_));
  AOI210     m165(.A0(mai_mai_n145_), .A1(mai_mai_n94_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n130_), .Y(mai_mai_n190_));
  AOI210     m168(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n191_));
  NO2        m169(.A(mai_mai_n121_), .B(x06), .Y(mai_mai_n192_));
  AOI210     m170(.A0(mai_mai_n191_), .A1(mai_mai_n190_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n193_), .B(x12), .Y(mai_mai_n194_));
  INV        m172(.A(mai_mai_n71_), .Y(mai_mai_n195_));
  NO2        m173(.A(mai_mai_n88_), .B(x06), .Y(mai_mai_n196_));
  AOI210     m174(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n197_));
  AOI210     m175(.A0(mai_mai_n196_), .A1(mai_mai_n53_), .B0(mai_mai_n23_), .Y(mai_mai_n198_));
  OAI210     m176(.A0(mai_mai_n194_), .A1(mai_mai_n53_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n132_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n201_));
  OAI210     m179(.A0(mai_mai_n73_), .A1(mai_mai_n36_), .B0(mai_mai_n112_), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n95_), .B(x03), .Y(mai_mai_n203_));
  NOi21      m181(.An(x13), .B(x04), .Y(mai_mai_n204_));
  NO3        m182(.A(mai_mai_n204_), .B(mai_mai_n71_), .C(mai_mai_n175_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n205_), .B(x05), .Y(mai_mai_n206_));
  INV        m184(.A(mai_mai_n85_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n207_), .B(x12), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n210_));
  OAI210     m188(.A0(mai_mai_n210_), .A1(mai_mai_n168_), .B0(mai_mai_n166_), .Y(mai_mai_n211_));
  AOI210     m189(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n212_));
  NO2        m190(.A(x06), .B(x00), .Y(mai_mai_n213_));
  NO3        m191(.A(mai_mai_n213_), .B(mai_mai_n212_), .C(mai_mai_n41_), .Y(mai_mai_n214_));
  OAI210     m192(.A0(mai_mai_n96_), .A1(mai_mai_n136_), .B0(mai_mai_n67_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n217_), .B(x03), .Y(mai_mai_n218_));
  OA210      m196(.A0(mai_mai_n218_), .A1(mai_mai_n216_), .B0(mai_mai_n211_), .Y(mai_mai_n219_));
  NA2        m197(.A(x13), .B(mai_mai_n94_), .Y(mai_mai_n220_));
  NA3        m198(.A(mai_mai_n220_), .B(x12), .C(mai_mai_n86_), .Y(mai_mai_n221_));
  OAI210     m199(.A0(mai_mai_n219_), .A1(mai_mai_n209_), .B0(mai_mai_n221_), .Y(mai_mai_n222_));
  AOI210     m200(.A0(mai_mai_n208_), .A1(mai_mai_n206_), .B0(mai_mai_n222_), .Y(mai_mai_n223_));
  AOI210     m201(.A0(mai_mai_n223_), .A1(mai_mai_n199_), .B0(x07), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n66_), .B(mai_mai_n29_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n204_), .B(mai_mai_n175_), .Y(mai_mai_n226_));
  AOI210     m204(.A0(mai_mai_n226_), .A1(mai_mai_n138_), .B0(mai_mai_n225_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n95_), .B(x06), .Y(mai_mai_n228_));
  INV        m206(.A(mai_mai_n228_), .Y(mai_mai_n229_));
  NO2        m207(.A(x08), .B(x05), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n230_), .B(mai_mai_n212_), .Y(mai_mai_n231_));
  NA2        m209(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n232_));
  OAI210     m210(.A0(mai_mai_n231_), .A1(mai_mai_n229_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  NO2        m211(.A(x12), .B(x02), .Y(mai_mai_n234_));
  INV        m212(.A(mai_mai_n234_), .Y(mai_mai_n235_));
  NO2        m213(.A(mai_mai_n235_), .B(mai_mai_n207_), .Y(mai_mai_n236_));
  OA210      m214(.A0(mai_mai_n233_), .A1(mai_mai_n227_), .B0(mai_mai_n236_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n238_), .B(x01), .Y(mai_mai_n239_));
  NOi21      m217(.An(mai_mai_n78_), .B(mai_mai_n112_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n228_), .B(mai_mai_n202_), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n95_), .B(x04), .Y(mai_mai_n242_));
  NA2        m220(.A(mai_mai_n242_), .B(mai_mai_n28_), .Y(mai_mai_n243_));
  OAI210     m221(.A0(mai_mai_n243_), .A1(mai_mai_n111_), .B0(mai_mai_n241_), .Y(mai_mai_n244_));
  NO3        m222(.A(mai_mai_n84_), .B(x12), .C(x03), .Y(mai_mai_n245_));
  OAI210     m223(.A0(mai_mai_n244_), .A1(mai_mai_n240_), .B0(mai_mai_n245_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n54_), .B(x05), .Y(mai_mai_n247_));
  NO3        m225(.A(mai_mai_n247_), .B(mai_mai_n197_), .C(mai_mai_n170_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n209_), .B(mai_mai_n28_), .Y(mai_mai_n249_));
  OAI210     m227(.A0(mai_mai_n248_), .A1(mai_mai_n200_), .B0(mai_mai_n249_), .Y(mai_mai_n250_));
  NA2        m228(.A(mai_mai_n250_), .B(mai_mai_n246_), .Y(mai_mai_n251_));
  NO3        m229(.A(mai_mai_n251_), .B(mai_mai_n237_), .C(mai_mai_n224_), .Y(mai_mai_n252_));
  OAI210     m230(.A0(mai_mai_n188_), .A1(mai_mai_n57_), .B0(mai_mai_n252_), .Y(mai02));
  NOi21      m231(.An(mai_mai_n205_), .B(mai_mai_n158_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n254_), .B(mai_mai_n32_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n255_), .B(mai_mai_n156_), .Y(mai_mai_n256_));
  INV        m234(.A(mai_mai_n156_), .Y(mai_mai_n257_));
  AOI210     m235(.A0(mai_mai_n108_), .A1(mai_mai_n80_), .B0(mai_mai_n197_), .Y(mai_mai_n258_));
  NO2        m236(.A(mai_mai_n258_), .B(mai_mai_n95_), .Y(mai_mai_n259_));
  AOI220     m237(.A0(mai_mai_n259_), .A1(mai_mai_n257_), .B0(mai_mai_n142_), .B1(mai_mai_n141_), .Y(mai_mai_n260_));
  AOI210     m238(.A0(mai_mai_n260_), .A1(mai_mai_n256_), .B0(mai_mai_n48_), .Y(mai_mai_n261_));
  NO2        m239(.A(x05), .B(x02), .Y(mai_mai_n262_));
  OAI210     m240(.A0(mai_mai_n190_), .A1(mai_mai_n175_), .B0(mai_mai_n262_), .Y(mai_mai_n263_));
  AOI220     m241(.A0(mai_mai_n230_), .A1(mai_mai_n54_), .B0(mai_mai_n52_), .B1(mai_mai_n36_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n263_), .B(mai_mai_n132_), .Y(mai_mai_n265_));
  NO2        m243(.A(mai_mai_n217_), .B(mai_mai_n47_), .Y(mai_mai_n266_));
  NA2        m244(.A(mai_mai_n266_), .B(mai_mai_n206_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n268_));
  NA2        m246(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n269_));
  OA210      m247(.A0(mai_mai_n269_), .A1(x08), .B0(mai_mai_n134_), .Y(mai_mai_n270_));
  AOI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n130_), .B0(mai_mai_n268_), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n271_), .B(mai_mai_n89_), .Y(mai_mai_n272_));
  NA3        m250(.A(mai_mai_n89_), .B(mai_mai_n78_), .C(mai_mai_n201_), .Y(mai_mai_n273_));
  NA3        m251(.A(mai_mai_n88_), .B(mai_mai_n77_), .C(mai_mai_n42_), .Y(mai_mai_n274_));
  AOI210     m252(.A0(mai_mai_n274_), .A1(mai_mai_n273_), .B0(x04), .Y(mai_mai_n275_));
  INV        m253(.A(mai_mai_n141_), .Y(mai_mai_n276_));
  OAI220     m254(.A0(mai_mai_n231_), .A1(mai_mai_n97_), .B0(mai_mai_n276_), .B1(mai_mai_n123_), .Y(mai_mai_n277_));
  AOI210     m255(.A0(mai_mai_n277_), .A1(x13), .B0(mai_mai_n275_), .Y(mai_mai_n278_));
  NA3        m256(.A(mai_mai_n278_), .B(mai_mai_n272_), .C(mai_mai_n267_), .Y(mai_mai_n279_));
  NO3        m257(.A(mai_mai_n279_), .B(mai_mai_n265_), .C(mai_mai_n261_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n131_), .B(x03), .Y(mai_mai_n281_));
  INV        m259(.A(mai_mai_n165_), .Y(mai_mai_n282_));
  NA2        m260(.A(mai_mai_n35_), .B(mai_mai_n36_), .Y(mai_mai_n283_));
  AOI220     m261(.A0(mai_mai_n283_), .A1(mai_mai_n282_), .B0(mai_mai_n183_), .B1(x08), .Y(mai_mai_n284_));
  OAI210     m262(.A0(mai_mai_n284_), .A1(mai_mai_n247_), .B0(mai_mai_n281_), .Y(mai_mai_n285_));
  NA2        m263(.A(mai_mai_n285_), .B(mai_mai_n99_), .Y(mai_mai_n286_));
  NA2        m264(.A(mai_mai_n155_), .B(mai_mai_n150_), .Y(mai_mai_n287_));
  AN2        m265(.A(mai_mai_n287_), .B(mai_mai_n161_), .Y(mai_mai_n288_));
  INV        m266(.A(mai_mai_n52_), .Y(mai_mai_n289_));
  OAI220     m267(.A0(mai_mai_n242_), .A1(mai_mai_n289_), .B0(mai_mai_n124_), .B1(mai_mai_n28_), .Y(mai_mai_n290_));
  OAI210     m268(.A0(mai_mai_n290_), .A1(mai_mai_n288_), .B0(mai_mai_n100_), .Y(mai_mai_n291_));
  NA2        m269(.A(mai_mai_n242_), .B(mai_mai_n94_), .Y(mai_mai_n292_));
  NA2        m270(.A(mai_mai_n94_), .B(mai_mai_n41_), .Y(mai_mai_n293_));
  NA3        m271(.A(mai_mai_n293_), .B(mai_mai_n292_), .C(mai_mai_n123_), .Y(mai_mai_n294_));
  NA4        m272(.A(mai_mai_n294_), .B(mai_mai_n291_), .C(mai_mai_n286_), .D(mai_mai_n48_), .Y(mai_mai_n295_));
  INV        m273(.A(mai_mai_n183_), .Y(mai_mai_n296_));
  NO2        m274(.A(mai_mai_n151_), .B(mai_mai_n40_), .Y(mai_mai_n297_));
  NA2        m275(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n298_));
  OAI220     m276(.A0(mai_mai_n298_), .A1(mai_mai_n297_), .B0(mai_mai_n296_), .B1(mai_mai_n55_), .Y(mai_mai_n299_));
  NA2        m277(.A(mai_mai_n299_), .B(x02), .Y(mai_mai_n300_));
  INV        m278(.A(mai_mai_n210_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n180_), .B(x04), .Y(mai_mai_n302_));
  NO2        m280(.A(mai_mai_n302_), .B(mai_mai_n301_), .Y(mai_mai_n303_));
  NO3        m281(.A(mai_mai_n167_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n304_));
  OAI210     m282(.A0(mai_mai_n304_), .A1(mai_mai_n303_), .B0(mai_mai_n89_), .Y(mai_mai_n305_));
  NO3        m283(.A(mai_mai_n180_), .B(mai_mai_n149_), .C(mai_mai_n51_), .Y(mai_mai_n306_));
  OAI210     m284(.A0(x12), .A1(mai_mai_n176_), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  NA4        m285(.A(mai_mai_n307_), .B(mai_mai_n305_), .C(mai_mai_n300_), .D(x06), .Y(mai_mai_n308_));
  NA2        m286(.A(x09), .B(x03), .Y(mai_mai_n309_));
  OAI220     m287(.A0(mai_mai_n309_), .A1(mai_mai_n122_), .B0(mai_mai_n189_), .B1(mai_mai_n60_), .Y(mai_mai_n310_));
  NO3        m288(.A(mai_mai_n247_), .B(mai_mai_n121_), .C(x08), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n311_), .Y(mai_mai_n312_));
  NO2        m290(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n313_));
  NA2        m291(.A(mai_mai_n306_), .B(mai_mai_n313_), .Y(mai_mai_n314_));
  OAI210     m292(.A0(mai_mai_n312_), .A1(mai_mai_n28_), .B0(mai_mai_n314_), .Y(mai_mai_n315_));
  AO220      m293(.A0(mai_mai_n315_), .A1(x04), .B0(mai_mai_n310_), .B1(x05), .Y(mai_mai_n316_));
  AOI210     m294(.A0(mai_mai_n308_), .A1(mai_mai_n295_), .B0(mai_mai_n316_), .Y(mai_mai_n317_));
  OAI210     m295(.A0(mai_mai_n280_), .A1(x12), .B0(mai_mai_n317_), .Y(mai03));
  OR2        m296(.A(mai_mai_n42_), .B(mai_mai_n201_), .Y(mai_mai_n319_));
  AOI210     m297(.A0(mai_mai_n142_), .A1(mai_mai_n94_), .B0(mai_mai_n319_), .Y(mai_mai_n320_));
  AO210      m298(.A0(mai_mai_n301_), .A1(mai_mai_n80_), .B0(mai_mai_n302_), .Y(mai_mai_n321_));
  NA2        m299(.A(mai_mai_n180_), .B(mai_mai_n141_), .Y(mai_mai_n322_));
  NA3        m300(.A(mai_mai_n322_), .B(mai_mai_n321_), .C(mai_mai_n184_), .Y(mai_mai_n323_));
  OAI210     m301(.A0(mai_mai_n323_), .A1(mai_mai_n320_), .B0(x05), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n319_), .B(x05), .Y(mai_mai_n325_));
  AOI210     m303(.A0(mai_mai_n130_), .A1(mai_mai_n195_), .B0(mai_mai_n325_), .Y(mai_mai_n326_));
  AOI210     m304(.A0(mai_mai_n203_), .A1(mai_mai_n74_), .B0(mai_mai_n115_), .Y(mai_mai_n327_));
  OAI220     m305(.A0(mai_mai_n327_), .A1(mai_mai_n55_), .B0(mai_mai_n269_), .B1(mai_mai_n264_), .Y(mai_mai_n328_));
  OAI210     m306(.A0(mai_mai_n328_), .A1(mai_mai_n326_), .B0(mai_mai_n94_), .Y(mai_mai_n329_));
  AOI210     m307(.A0(mai_mai_n134_), .A1(mai_mai_n56_), .B0(mai_mai_n38_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n158_), .B(mai_mai_n126_), .Y(mai_mai_n331_));
  OAI220     m309(.A0(mai_mai_n331_), .A1(mai_mai_n37_), .B0(mai_mai_n137_), .B1(x13), .Y(mai_mai_n332_));
  OAI210     m310(.A0(mai_mai_n332_), .A1(mai_mai_n330_), .B0(x04), .Y(mai_mai_n333_));
  NO3        m311(.A(mai_mai_n293_), .B(mai_mai_n79_), .C(mai_mai_n55_), .Y(mai_mai_n334_));
  AOI210     m312(.A0(mai_mai_n172_), .A1(mai_mai_n94_), .B0(mai_mai_n134_), .Y(mai_mai_n335_));
  OA210      m313(.A0(mai_mai_n151_), .A1(x12), .B0(mai_mai_n126_), .Y(mai_mai_n336_));
  NO3        m314(.A(mai_mai_n336_), .B(mai_mai_n335_), .C(mai_mai_n334_), .Y(mai_mai_n337_));
  NA4        m315(.A(mai_mai_n337_), .B(mai_mai_n333_), .C(mai_mai_n329_), .D(mai_mai_n324_), .Y(mai04));
  NO2        m316(.A(mai_mai_n83_), .B(mai_mai_n39_), .Y(mai_mai_n339_));
  XO2        m317(.A(mai_mai_n339_), .B(mai_mai_n220_), .Y(mai05));
  NO2        m318(.A(mai_mai_n268_), .B(mai_mai_n25_), .Y(mai_mai_n341_));
  NA3        m319(.A(mai_mai_n132_), .B(mai_mai_n124_), .C(mai_mai_n31_), .Y(mai_mai_n342_));
  AOI210     m320(.A0(x06), .A1(mai_mai_n342_), .B0(mai_mai_n24_), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(mai_mai_n94_), .Y(mai_mai_n344_));
  NA2        m322(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n346_));
  NA2        m324(.A(mai_mai_n225_), .B(x03), .Y(mai_mai_n347_));
  OAI220     m325(.A0(mai_mai_n347_), .A1(mai_mai_n346_), .B0(mai_mai_n345_), .B1(mai_mai_n75_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(mai_mai_n26_), .A1(mai_mai_n94_), .B0(x07), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n348_), .A1(x06), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  AOI210     m328(.A0(mai_mai_n404_), .A1(mai_mai_n347_), .B0(mai_mai_n228_), .Y(mai_mai_n351_));
  OR2        m329(.A(mai_mai_n351_), .B(mai_mai_n209_), .Y(mai_mai_n352_));
  NA2        m330(.A(mai_mai_n147_), .B(x05), .Y(mai_mai_n353_));
  NA3        m331(.A(mai_mai_n353_), .B(mai_mai_n213_), .C(mai_mai_n207_), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n355_));
  OAI210     m333(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n356_));
  OR3        m334(.A(mai_mai_n356_), .B(mai_mai_n355_), .C(mai_mai_n44_), .Y(mai_mai_n357_));
  NA3        m335(.A(mai_mai_n357_), .B(mai_mai_n354_), .C(mai_mai_n352_), .Y(mai_mai_n358_));
  NA2        m336(.A(mai_mai_n358_), .B(mai_mai_n94_), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n33_), .B(mai_mai_n94_), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n360_), .A1(mai_mai_n85_), .B0(x07), .Y(mai_mai_n361_));
  AOI220     m339(.A0(mai_mai_n361_), .A1(mai_mai_n359_), .B0(mai_mai_n350_), .B1(mai_mai_n344_), .Y(mai_mai_n362_));
  NA3        m340(.A(mai_mai_n23_), .B(mai_mai_n57_), .C(mai_mai_n48_), .Y(mai_mai_n363_));
  AO210      m341(.A0(mai_mai_n363_), .A1(mai_mai_n238_), .B0(mai_mai_n235_), .Y(mai_mai_n364_));
  NO2        m342(.A(mai_mai_n69_), .B(mai_mai_n131_), .Y(mai_mai_n365_));
  OR2        m343(.A(mai_mai_n365_), .B(x03), .Y(mai_mai_n366_));
  NA2        m344(.A(mai_mai_n313_), .B(mai_mai_n57_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n367_), .B(x11), .Y(mai_mai_n368_));
  NO3        m346(.A(mai_mai_n368_), .B(mai_mai_n133_), .C(mai_mai_n28_), .Y(mai_mai_n369_));
  AOI220     m347(.A0(mai_mai_n369_), .A1(mai_mai_n366_), .B0(mai_mai_n364_), .B1(mai_mai_n47_), .Y(mai_mai_n370_));
  NA2        m348(.A(mai_mai_n370_), .B(mai_mai_n95_), .Y(mai_mai_n371_));
  AOI210     m349(.A0(mai_mai_n302_), .A1(mai_mai_n102_), .B0(mai_mai_n234_), .Y(mai_mai_n372_));
  NOi21      m350(.An(mai_mai_n281_), .B(mai_mai_n126_), .Y(mai_mai_n373_));
  NO2        m351(.A(mai_mai_n373_), .B(mai_mai_n235_), .Y(mai_mai_n374_));
  OAI210     m352(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n375_));
  AOI210     m353(.A0(mai_mai_n220_), .A1(mai_mai_n47_), .B0(mai_mai_n375_), .Y(mai_mai_n376_));
  NO4        m354(.A(mai_mai_n376_), .B(mai_mai_n374_), .C(mai_mai_n372_), .D(x08), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n124_), .B(mai_mai_n28_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(mai_mai_n239_), .Y(mai_mai_n379_));
  OR3        m357(.A(mai_mai_n379_), .B(x12), .C(x03), .Y(mai_mai_n380_));
  NA3        m358(.A(mai_mai_n296_), .B(mai_mai_n117_), .C(x12), .Y(mai_mai_n381_));
  AO210      m359(.A0(mai_mai_n296_), .A1(mai_mai_n117_), .B0(mai_mai_n220_), .Y(mai_mai_n382_));
  NA4        m360(.A(mai_mai_n382_), .B(mai_mai_n381_), .C(mai_mai_n380_), .D(x08), .Y(mai_mai_n383_));
  INV        m361(.A(mai_mai_n383_), .Y(mai_mai_n384_));
  AOI210     m362(.A0(mai_mai_n377_), .A1(mai_mai_n371_), .B0(mai_mai_n384_), .Y(mai_mai_n385_));
  OAI210     m363(.A0(mai_mai_n367_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n386_));
  OAI210     m364(.A0(mai_mai_n406_), .A1(mai_mai_n386_), .B0(mai_mai_n171_), .Y(mai_mai_n387_));
  NA3        m365(.A(mai_mai_n379_), .B(mai_mai_n373_), .C(mai_mai_n292_), .Y(mai_mai_n388_));
  INV        m366(.A(x14), .Y(mai_mai_n389_));
  NO3        m367(.A(mai_mai_n281_), .B(mai_mai_n97_), .C(x11), .Y(mai_mai_n390_));
  NO3        m368(.A(mai_mai_n150_), .B(mai_mai_n69_), .C(mai_mai_n53_), .Y(mai_mai_n391_));
  NO3        m369(.A(mai_mai_n363_), .B(mai_mai_n293_), .C(mai_mai_n165_), .Y(mai_mai_n392_));
  NO4        m370(.A(mai_mai_n392_), .B(mai_mai_n391_), .C(mai_mai_n390_), .D(mai_mai_n389_), .Y(mai_mai_n393_));
  NA3        m371(.A(mai_mai_n393_), .B(mai_mai_n388_), .C(mai_mai_n387_), .Y(mai_mai_n394_));
  AOI220     m372(.A0(mai_mai_n360_), .A1(mai_mai_n57_), .B0(mai_mai_n378_), .B1(mai_mai_n149_), .Y(mai_mai_n395_));
  NOi21      m373(.An(mai_mai_n242_), .B(mai_mai_n137_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n397_));
  OAI210     m375(.A0(mai_mai_n397_), .A1(mai_mai_n396_), .B0(mai_mai_n94_), .Y(mai_mai_n398_));
  OAI210     m376(.A0(mai_mai_n395_), .A1(mai_mai_n84_), .B0(mai_mai_n398_), .Y(mai_mai_n399_));
  NO4        m377(.A(mai_mai_n399_), .B(mai_mai_n394_), .C(mai_mai_n385_), .D(mai_mai_n362_), .Y(mai06));
  INV        m378(.A(x07), .Y(mai_mai_n403_));
  INV        m379(.A(x02), .Y(mai_mai_n404_));
  INV        m380(.A(x01), .Y(mai_mai_n405_));
  INV        m381(.A(mai_mai_n156_), .Y(mai_mai_n406_));
  INV        m382(.A(mai_mai_n147_), .Y(mai_mai_n407_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  INV        u039(.A(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  NO2        u042(.A(men_men_n64_), .B(men_men_n62_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  NA3        u050(.A(men_men_n72_), .B(men_men_n71_), .C(men_men_n28_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n73_), .A1(x11), .B0(x03), .Y(men_men_n74_));
  NOi31      u052(.An(x08), .B(x04), .C(x00), .Y(men_men_n75_));
  NO2        u053(.A(x10), .B(x09), .Y(men_men_n76_));
  NO2        u054(.A(men_men_n429_), .B(men_men_n24_), .Y(men_men_n77_));
  NO2        u055(.A(x09), .B(men_men_n41_), .Y(men_men_n78_));
  OAI210     u056(.A0(men_men_n78_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n48_), .B(men_men_n79_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n36_), .B(x00), .Y(men_men_n81_));
  NO2        u059(.A(x08), .B(x01), .Y(men_men_n82_));
  OAI210     u060(.A0(men_men_n82_), .A1(men_men_n81_), .B0(men_men_n35_), .Y(men_men_n83_));
  NA2        u061(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n84_));
  NO3        u062(.A(men_men_n83_), .B(men_men_n80_), .C(men_men_n77_), .Y(men_men_n85_));
  AN2        u063(.A(men_men_n85_), .B(men_men_n74_), .Y(men_men_n86_));
  INV        u064(.A(men_men_n83_), .Y(men_men_n87_));
  NO2        u065(.A(x06), .B(x05), .Y(men_men_n88_));
  NA2        u066(.A(x11), .B(x00), .Y(men_men_n89_));
  NO2        u067(.A(x11), .B(men_men_n47_), .Y(men_men_n90_));
  NOi21      u068(.An(men_men_n89_), .B(men_men_n90_), .Y(men_men_n91_));
  AOI210     u069(.A0(men_men_n88_), .A1(men_men_n87_), .B0(men_men_n91_), .Y(men_men_n92_));
  NOi21      u070(.An(x01), .B(x10), .Y(men_men_n93_));
  NO2        u071(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n94_));
  NO3        u072(.A(men_men_n94_), .B(men_men_n93_), .C(x06), .Y(men_men_n95_));
  NA2        u073(.A(men_men_n95_), .B(men_men_n27_), .Y(men_men_n96_));
  OAI210     u074(.A0(men_men_n92_), .A1(x07), .B0(men_men_n96_), .Y(men_men_n97_));
  NO3        u075(.A(men_men_n97_), .B(men_men_n86_), .C(men_men_n69_), .Y(men01));
  INV        u076(.A(x12), .Y(men_men_n99_));
  INV        u077(.A(x13), .Y(men_men_n100_));
  NA2        u078(.A(men_men_n431_), .B(men_men_n70_), .Y(men_men_n101_));
  NA2        u079(.A(x08), .B(x04), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n102_), .B(men_men_n57_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n103_), .B(men_men_n101_), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n93_), .B(men_men_n28_), .Y(men_men_n105_));
  NO2        u083(.A(x10), .B(x01), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n29_), .B(x00), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NA2        u086(.A(x04), .B(men_men_n28_), .Y(men_men_n109_));
  NO3        u087(.A(men_men_n109_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n110_));
  NA2        u088(.A(men_men_n110_), .B(men_men_n108_), .Y(men_men_n111_));
  AOI210     u089(.A0(men_men_n111_), .A1(men_men_n104_), .B0(men_men_n100_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n56_), .B(x05), .Y(men_men_n113_));
  NOi21      u091(.An(men_men_n113_), .B(men_men_n58_), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n100_), .B(men_men_n36_), .Y(men_men_n115_));
  NA3        u093(.A(men_men_n115_), .B(x04), .C(x06), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n116_), .B(men_men_n114_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n82_), .B(x13), .Y(men_men_n118_));
  NA2        u096(.A(x13), .B(men_men_n35_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(x05), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n121_));
  NO2        u099(.A(x00), .B(men_men_n72_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n123_));
  NA2        u101(.A(x10), .B(men_men_n57_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n51_), .B(x05), .Y(men_men_n126_));
  NO2        u104(.A(men_men_n60_), .B(x05), .Y(men_men_n127_));
  NO3        u105(.A(x00), .B(x06), .C(x03), .Y(men_men_n128_));
  NO4        u106(.A(men_men_n128_), .B(men_men_n122_), .C(men_men_n117_), .D(men_men_n112_), .Y(men_men_n129_));
  NA2        u107(.A(x13), .B(men_men_n36_), .Y(men_men_n130_));
  OAI210     u108(.A0(men_men_n82_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n131_), .B(men_men_n130_), .Y(men_men_n132_));
  OA210      u110(.A0(x00), .A1(men_men_n76_), .B0(x04), .Y(men_men_n133_));
  NO2        u111(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n134_));
  NA2        u112(.A(men_men_n29_), .B(x06), .Y(men_men_n135_));
  AOI210     u113(.A0(men_men_n135_), .A1(men_men_n49_), .B0(men_men_n134_), .Y(men_men_n136_));
  OA210      u114(.A0(men_men_n136_), .A1(men_men_n133_), .B0(men_men_n132_), .Y(men_men_n137_));
  NO2        u115(.A(x09), .B(x05), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n138_), .B(men_men_n47_), .Y(men_men_n139_));
  AOI210     u117(.A0(men_men_n139_), .A1(men_men_n108_), .B0(men_men_n49_), .Y(men_men_n140_));
  NA2        u118(.A(x09), .B(x00), .Y(men_men_n141_));
  NA2        u119(.A(men_men_n113_), .B(men_men_n141_), .Y(men_men_n142_));
  NA2        u120(.A(men_men_n75_), .B(men_men_n51_), .Y(men_men_n143_));
  AOI210     u121(.A0(men_men_n143_), .A1(men_men_n142_), .B0(men_men_n135_), .Y(men_men_n144_));
  NO3        u122(.A(men_men_n144_), .B(men_men_n140_), .C(men_men_n137_), .Y(men_men_n145_));
  NO2        u123(.A(x03), .B(x02), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n83_), .B(men_men_n100_), .Y(men_men_n147_));
  OAI210     u125(.A0(men_men_n147_), .A1(men_men_n114_), .B0(men_men_n146_), .Y(men_men_n148_));
  OA210      u126(.A0(men_men_n145_), .A1(x11), .B0(men_men_n148_), .Y(men_men_n149_));
  OAI210     u127(.A0(men_men_n129_), .A1(men_men_n23_), .B0(men_men_n149_), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n108_), .B(men_men_n40_), .Y(men_men_n151_));
  NAi21      u129(.An(x06), .B(x10), .Y(men_men_n152_));
  NOi21      u130(.An(x01), .B(x13), .Y(men_men_n153_));
  NA2        u131(.A(men_men_n153_), .B(men_men_n152_), .Y(men_men_n154_));
  OR2        u132(.A(men_men_n154_), .B(x08), .Y(men_men_n155_));
  AOI210     u133(.A0(men_men_n155_), .A1(men_men_n151_), .B0(men_men_n41_), .Y(men_men_n156_));
  NO2        u134(.A(men_men_n29_), .B(x03), .Y(men_men_n157_));
  NA2        u135(.A(men_men_n100_), .B(x01), .Y(men_men_n158_));
  NO2        u136(.A(men_men_n158_), .B(x08), .Y(men_men_n159_));
  OAI210     u137(.A0(x05), .A1(men_men_n159_), .B0(men_men_n51_), .Y(men_men_n160_));
  AOI210     u138(.A0(men_men_n160_), .A1(men_men_n157_), .B0(men_men_n48_), .Y(men_men_n161_));
  AOI210     u139(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n161_), .A1(men_men_n156_), .B0(men_men_n162_), .Y(men_men_n163_));
  NA2        u141(.A(x04), .B(x02), .Y(men_men_n164_));
  NA2        u142(.A(x10), .B(x05), .Y(men_men_n165_));
  NO2        u143(.A(x09), .B(x01), .Y(men_men_n166_));
  NA2        u144(.A(x03), .B(x00), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n113_), .B(x08), .Y(men_men_n168_));
  NA3        u146(.A(men_men_n153_), .B(men_men_n152_), .C(men_men_n51_), .Y(men_men_n169_));
  NA2        u147(.A(men_men_n93_), .B(x05), .Y(men_men_n170_));
  OAI210     u148(.A0(men_men_n170_), .A1(men_men_n115_), .B0(men_men_n169_), .Y(men_men_n171_));
  AOI210     u149(.A0(men_men_n168_), .A1(x06), .B0(men_men_n171_), .Y(men_men_n172_));
  OAI210     u150(.A0(men_men_n172_), .A1(x11), .B0(men_men_n167_), .Y(men_men_n173_));
  NAi21      u151(.An(men_men_n164_), .B(men_men_n173_), .Y(men_men_n174_));
  INV        u152(.A(men_men_n25_), .Y(men_men_n175_));
  NAi21      u153(.An(x13), .B(x00), .Y(men_men_n176_));
  AOI210     u154(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n176_), .Y(men_men_n177_));
  AOI220     u155(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n165_), .A1(men_men_n35_), .B0(men_men_n178_), .Y(men_men_n179_));
  BUFFER     u157(.A(men_men_n177_), .Y(men_men_n180_));
  BUFFER     u158(.A(men_men_n71_), .Y(men_men_n181_));
  NO2        u159(.A(men_men_n176_), .B(men_men_n36_), .Y(men_men_n182_));
  INV        u160(.A(men_men_n182_), .Y(men_men_n183_));
  NO2        u161(.A(men_men_n57_), .B(men_men_n181_), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(men_men_n180_), .B0(men_men_n175_), .Y(men_men_n185_));
  NOi21      u163(.An(x09), .B(x00), .Y(men_men_n186_));
  NO3        u164(.A(men_men_n81_), .B(men_men_n186_), .C(men_men_n47_), .Y(men_men_n187_));
  NA2        u165(.A(men_men_n187_), .B(men_men_n124_), .Y(men_men_n188_));
  NA2        u166(.A(x06), .B(x05), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n35_), .B0(men_men_n99_), .Y(men_men_n190_));
  AOI210     u168(.A0(x10), .A1(men_men_n58_), .B0(men_men_n190_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n191_), .B(men_men_n188_), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n100_), .B(x12), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n193_), .Y(men_men_n194_));
  NA2        u172(.A(men_men_n93_), .B(men_men_n51_), .Y(men_men_n195_));
  NO2        u173(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n196_), .B(x02), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n197_), .B(men_men_n195_), .Y(men_men_n198_));
  AOI210     u176(.A0(men_men_n194_), .A1(men_men_n192_), .B0(men_men_n198_), .Y(men_men_n199_));
  NA4        u177(.A(men_men_n199_), .B(men_men_n185_), .C(men_men_n174_), .D(men_men_n163_), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n150_), .A1(men_men_n99_), .B0(men_men_n200_), .Y(men_men_n201_));
  INV        u179(.A(men_men_n73_), .Y(men_men_n202_));
  NA2        u180(.A(men_men_n202_), .B(men_men_n132_), .Y(men_men_n203_));
  NA2        u181(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n204_));
  INV        u182(.A(men_men_n204_), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n123_), .B(x06), .Y(men_men_n206_));
  INV        u184(.A(men_men_n206_), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n207_), .A1(men_men_n203_), .B0(x12), .Y(men_men_n208_));
  INV        u186(.A(men_men_n75_), .Y(men_men_n209_));
  NO2        u187(.A(x05), .B(men_men_n51_), .Y(men_men_n210_));
  OAI210     u188(.A0(men_men_n210_), .A1(men_men_n154_), .B0(men_men_n57_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n211_), .B(men_men_n209_), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n93_), .B(x06), .Y(men_men_n213_));
  NA4        u191(.A(men_men_n152_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n214_));
  NA2        u192(.A(men_men_n214_), .B(men_men_n135_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(x02), .Y(men_men_n216_));
  AOI210     u194(.A0(men_men_n216_), .A1(men_men_n212_), .B0(men_men_n23_), .Y(men_men_n217_));
  OAI210     u195(.A0(men_men_n208_), .A1(men_men_n57_), .B0(men_men_n217_), .Y(men_men_n218_));
  INV        u196(.A(men_men_n135_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n51_), .B(x03), .Y(men_men_n220_));
  NO2        u198(.A(men_men_n100_), .B(x03), .Y(men_men_n221_));
  AOI210     u199(.A0(men_men_n75_), .A1(men_men_n220_), .B0(men_men_n221_), .Y(men_men_n222_));
  INV        u200(.A(men_men_n152_), .Y(men_men_n223_));
  NOi21      u201(.An(x13), .B(x04), .Y(men_men_n224_));
  NO3        u202(.A(men_men_n224_), .B(men_men_n75_), .C(men_men_n186_), .Y(men_men_n225_));
  NO2        u203(.A(men_men_n225_), .B(x05), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n223_), .B(men_men_n57_), .Y(men_men_n227_));
  OAI210     u205(.A0(men_men_n222_), .A1(men_men_n219_), .B0(men_men_n227_), .Y(men_men_n228_));
  INV        u206(.A(men_men_n90_), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n229_), .B(x12), .Y(men_men_n230_));
  NA2        u208(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n232_));
  OAI210     u210(.A0(men_men_n232_), .A1(men_men_n179_), .B0(men_men_n177_), .Y(men_men_n233_));
  AOI210     u211(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n234_));
  NA2        u212(.A(men_men_n141_), .B(men_men_n72_), .Y(men_men_n235_));
  INV        u213(.A(men_men_n235_), .Y(men_men_n236_));
  NA2        u214(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n237_));
  NA2        u215(.A(men_men_n237_), .B(x03), .Y(men_men_n238_));
  OA210      u216(.A0(men_men_n238_), .A1(men_men_n236_), .B0(men_men_n233_), .Y(men_men_n239_));
  NA2        u217(.A(x13), .B(men_men_n99_), .Y(men_men_n240_));
  NA3        u218(.A(men_men_n240_), .B(men_men_n190_), .C(men_men_n91_), .Y(men_men_n241_));
  OAI210     u219(.A0(men_men_n239_), .A1(men_men_n231_), .B0(men_men_n241_), .Y(men_men_n242_));
  AOI210     u220(.A0(men_men_n230_), .A1(men_men_n228_), .B0(men_men_n242_), .Y(men_men_n243_));
  AOI210     u221(.A0(men_men_n243_), .A1(men_men_n218_), .B0(x07), .Y(men_men_n244_));
  NA2        u222(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n245_));
  AOI210     u223(.A0(men_men_n130_), .A1(men_men_n143_), .B0(men_men_n245_), .Y(men_men_n246_));
  NO2        u224(.A(men_men_n100_), .B(x06), .Y(men_men_n247_));
  INV        u225(.A(men_men_n247_), .Y(men_men_n248_));
  NO2        u226(.A(x08), .B(x05), .Y(men_men_n249_));
  NO2        u227(.A(men_men_n249_), .B(men_men_n234_), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n75_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n251_));
  OAI210     u229(.A0(men_men_n250_), .A1(men_men_n248_), .B0(men_men_n251_), .Y(men_men_n252_));
  NO2        u230(.A(x12), .B(x02), .Y(men_men_n253_));
  INV        u231(.A(men_men_n253_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n254_), .B(men_men_n229_), .Y(men_men_n255_));
  OA210      u233(.A0(men_men_n252_), .A1(men_men_n246_), .B0(men_men_n255_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n257_));
  NO2        u235(.A(men_men_n257_), .B(x01), .Y(men_men_n258_));
  BUFFER     u236(.A(men_men_n82_), .Y(men_men_n259_));
  NO2        u237(.A(men_men_n259_), .B(men_men_n258_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n260_), .A1(men_men_n432_), .B0(men_men_n29_), .Y(men_men_n261_));
  INV        u239(.A(men_men_n247_), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n100_), .B(x04), .Y(men_men_n263_));
  OAI210     u241(.A0(x02), .A1(men_men_n118_), .B0(men_men_n262_), .Y(men_men_n264_));
  NO3        u242(.A(men_men_n89_), .B(x12), .C(x03), .Y(men_men_n265_));
  OAI210     u243(.A0(men_men_n264_), .A1(men_men_n261_), .B0(men_men_n265_), .Y(men_men_n266_));
  AOI210     u244(.A0(men_men_n195_), .A1(men_men_n189_), .B0(men_men_n102_), .Y(men_men_n267_));
  NOi21      u245(.An(men_men_n245_), .B(men_men_n213_), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n25_), .B(x00), .Y(men_men_n269_));
  OAI210     u247(.A0(men_men_n268_), .A1(men_men_n267_), .B0(men_men_n269_), .Y(men_men_n270_));
  NO2        u248(.A(men_men_n58_), .B(x05), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n231_), .B(men_men_n28_), .Y(men_men_n272_));
  NA2        u250(.A(men_men_n219_), .B(men_men_n272_), .Y(men_men_n273_));
  NA3        u251(.A(men_men_n273_), .B(men_men_n270_), .C(men_men_n266_), .Y(men_men_n274_));
  NO3        u252(.A(men_men_n274_), .B(men_men_n256_), .C(men_men_n244_), .Y(men_men_n275_));
  OAI210     u253(.A0(men_men_n201_), .A1(men_men_n61_), .B0(men_men_n275_), .Y(men02));
  AOI210     u254(.A0(men_men_n130_), .A1(men_men_n83_), .B0(men_men_n126_), .Y(men_men_n277_));
  NOi21      u255(.An(men_men_n225_), .B(men_men_n166_), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n100_), .B(men_men_n35_), .Y(men_men_n279_));
  NA3        u257(.A(men_men_n279_), .B(x10), .C(men_men_n56_), .Y(men_men_n280_));
  OAI210     u258(.A0(men_men_n278_), .A1(men_men_n32_), .B0(men_men_n280_), .Y(men_men_n281_));
  OAI210     u259(.A0(men_men_n281_), .A1(men_men_n277_), .B0(men_men_n165_), .Y(men_men_n282_));
  INV        u260(.A(men_men_n165_), .Y(men_men_n283_));
  OAI210     u261(.A0(men_men_n83_), .A1(men_men_n51_), .B0(men_men_n100_), .Y(men_men_n284_));
  AOI220     u262(.A0(men_men_n284_), .A1(men_men_n283_), .B0(men_men_n147_), .B1(men_men_n146_), .Y(men_men_n285_));
  AOI210     u263(.A0(men_men_n285_), .A1(men_men_n282_), .B0(men_men_n48_), .Y(men_men_n286_));
  NO2        u264(.A(x05), .B(x02), .Y(men_men_n287_));
  OAI210     u265(.A0(men_men_n205_), .A1(men_men_n186_), .B0(men_men_n287_), .Y(men_men_n288_));
  AOI220     u266(.A0(men_men_n249_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n289_));
  NOi21      u267(.An(men_men_n279_), .B(men_men_n289_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n224_), .A1(men_men_n78_), .B0(men_men_n290_), .Y(men_men_n291_));
  AOI210     u269(.A0(men_men_n291_), .A1(men_men_n288_), .B0(men_men_n135_), .Y(men_men_n292_));
  NAi21      u270(.An(men_men_n226_), .B(men_men_n222_), .Y(men_men_n293_));
  NO2        u271(.A(men_men_n237_), .B(men_men_n47_), .Y(men_men_n294_));
  NA2        u272(.A(men_men_n294_), .B(men_men_n293_), .Y(men_men_n295_));
  OAI210     u273(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n296_));
  NA2        u274(.A(x13), .B(men_men_n28_), .Y(men_men_n297_));
  AOI210     u275(.A0(men_men_n297_), .A1(men_men_n131_), .B0(men_men_n296_), .Y(men_men_n298_));
  OAI210     u276(.A0(men_men_n298_), .A1(men_men_n221_), .B0(men_men_n94_), .Y(men_men_n299_));
  NA3        u277(.A(men_men_n94_), .B(men_men_n82_), .C(men_men_n220_), .Y(men_men_n300_));
  NA3        u278(.A(men_men_n93_), .B(men_men_n81_), .C(men_men_n42_), .Y(men_men_n301_));
  AOI210     u279(.A0(men_men_n301_), .A1(men_men_n300_), .B0(x04), .Y(men_men_n302_));
  NO2        u280(.A(men_men_n250_), .B(men_men_n105_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n303_), .A1(x13), .B0(men_men_n302_), .Y(men_men_n304_));
  NA3        u282(.A(men_men_n304_), .B(men_men_n299_), .C(men_men_n295_), .Y(men_men_n305_));
  NO3        u283(.A(men_men_n305_), .B(men_men_n292_), .C(men_men_n286_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n134_), .B(x03), .Y(men_men_n307_));
  OAI210     u285(.A0(men_men_n176_), .A1(men_men_n271_), .B0(men_men_n307_), .Y(men_men_n308_));
  NA2        u286(.A(men_men_n308_), .B(men_men_n106_), .Y(men_men_n309_));
  NA2        u287(.A(men_men_n164_), .B(men_men_n158_), .Y(men_men_n310_));
  AN2        u288(.A(men_men_n310_), .B(men_men_n168_), .Y(men_men_n311_));
  NO2        u289(.A(men_men_n126_), .B(men_men_n28_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n312_), .A1(men_men_n311_), .B0(men_men_n107_), .Y(men_men_n313_));
  NA2        u291(.A(men_men_n263_), .B(men_men_n99_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n99_), .B(men_men_n41_), .Y(men_men_n315_));
  NA3        u293(.A(men_men_n315_), .B(men_men_n314_), .C(men_men_n125_), .Y(men_men_n316_));
  NA4        u294(.A(men_men_n316_), .B(men_men_n313_), .C(men_men_n309_), .D(men_men_n48_), .Y(men_men_n317_));
  INV        u295(.A(men_men_n196_), .Y(men_men_n318_));
  NO2        u296(.A(men_men_n159_), .B(men_men_n40_), .Y(men_men_n319_));
  NA2        u297(.A(men_men_n32_), .B(x05), .Y(men_men_n320_));
  NO2        u298(.A(men_men_n320_), .B(men_men_n319_), .Y(men_men_n321_));
  NA2        u299(.A(men_men_n321_), .B(x02), .Y(men_men_n322_));
  INV        u300(.A(men_men_n232_), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n193_), .B(x04), .Y(men_men_n324_));
  NO2        u302(.A(men_men_n324_), .B(men_men_n323_), .Y(men_men_n325_));
  NO3        u303(.A(men_men_n178_), .B(x13), .C(men_men_n31_), .Y(men_men_n326_));
  OAI210     u304(.A0(men_men_n326_), .A1(men_men_n325_), .B0(men_men_n94_), .Y(men_men_n327_));
  NO3        u305(.A(men_men_n193_), .B(men_men_n157_), .C(men_men_n52_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n141_), .A1(men_men_n36_), .B0(men_men_n99_), .Y(men_men_n329_));
  OAI210     u307(.A0(men_men_n329_), .A1(men_men_n187_), .B0(men_men_n328_), .Y(men_men_n330_));
  NA4        u308(.A(men_men_n330_), .B(men_men_n327_), .C(men_men_n322_), .D(x06), .Y(men_men_n331_));
  NA2        u309(.A(x09), .B(x03), .Y(men_men_n332_));
  OAI220     u310(.A0(men_men_n332_), .A1(men_men_n124_), .B0(men_men_n204_), .B1(men_men_n63_), .Y(men_men_n333_));
  NO3        u311(.A(men_men_n271_), .B(men_men_n123_), .C(x08), .Y(men_men_n334_));
  AOI210     u312(.A0(x01), .A1(men_men_n219_), .B0(men_men_n334_), .Y(men_men_n335_));
  NO3        u313(.A(men_men_n113_), .B(men_men_n124_), .C(men_men_n38_), .Y(men_men_n336_));
  INV        u314(.A(men_men_n336_), .Y(men_men_n337_));
  OAI210     u315(.A0(men_men_n335_), .A1(men_men_n28_), .B0(men_men_n337_), .Y(men_men_n338_));
  AO220      u316(.A0(men_men_n338_), .A1(x04), .B0(men_men_n333_), .B1(x05), .Y(men_men_n339_));
  AOI210     u317(.A0(men_men_n331_), .A1(men_men_n317_), .B0(men_men_n339_), .Y(men_men_n340_));
  OAI210     u318(.A0(men_men_n306_), .A1(x12), .B0(men_men_n340_), .Y(men03));
  OR2        u319(.A(men_men_n42_), .B(men_men_n220_), .Y(men_men_n342_));
  AOI210     u320(.A0(men_men_n147_), .A1(men_men_n99_), .B0(men_men_n342_), .Y(men_men_n343_));
  AO210      u321(.A0(men_men_n323_), .A1(men_men_n84_), .B0(men_men_n324_), .Y(men_men_n344_));
  NA2        u322(.A(men_men_n193_), .B(men_men_n146_), .Y(men_men_n345_));
  NA3        u323(.A(men_men_n345_), .B(men_men_n344_), .C(men_men_n197_), .Y(men_men_n346_));
  OAI210     u324(.A0(men_men_n346_), .A1(men_men_n343_), .B0(x05), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n342_), .B(x05), .Y(men_men_n348_));
  AOI210     u326(.A0(men_men_n131_), .A1(men_men_n209_), .B0(men_men_n348_), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n221_), .A1(x08), .B0(men_men_n120_), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n350_), .A1(men_men_n59_), .B0(men_men_n297_), .B1(men_men_n289_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n351_), .A1(men_men_n349_), .B0(men_men_n99_), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n139_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n353_));
  NO2        u331(.A(men_men_n166_), .B(men_men_n127_), .Y(men_men_n354_));
  OAI220     u332(.A0(men_men_n354_), .A1(men_men_n37_), .B0(men_men_n142_), .B1(x13), .Y(men_men_n355_));
  OAI210     u333(.A0(men_men_n355_), .A1(men_men_n353_), .B0(x04), .Y(men_men_n356_));
  NO3        u334(.A(men_men_n315_), .B(men_men_n83_), .C(men_men_n59_), .Y(men_men_n357_));
  AOI210     u335(.A0(men_men_n183_), .A1(men_men_n99_), .B0(men_men_n139_), .Y(men_men_n358_));
  OA210      u336(.A0(men_men_n159_), .A1(x12), .B0(men_men_n127_), .Y(men_men_n359_));
  NO3        u337(.A(men_men_n359_), .B(men_men_n358_), .C(men_men_n357_), .Y(men_men_n360_));
  NA4        u338(.A(men_men_n360_), .B(men_men_n356_), .C(men_men_n352_), .D(men_men_n347_), .Y(men04));
  NO2        u339(.A(men_men_n87_), .B(men_men_n39_), .Y(men_men_n362_));
  XO2        u340(.A(men_men_n362_), .B(men_men_n240_), .Y(men05));
  NO2        u341(.A(x10), .B(men_men_n25_), .Y(men_men_n364_));
  NO2        u342(.A(men_men_n430_), .B(men_men_n24_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n364_), .B0(men_men_n99_), .Y(men_men_n366_));
  NA2        u344(.A(x11), .B(men_men_n31_), .Y(men_men_n367_));
  NA2        u345(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n368_));
  NA2        u346(.A(men_men_n245_), .B(x03), .Y(men_men_n369_));
  OAI220     u347(.A0(men_men_n369_), .A1(men_men_n368_), .B0(men_men_n367_), .B1(men_men_n79_), .Y(men_men_n370_));
  OAI210     u348(.A0(men_men_n26_), .A1(men_men_n99_), .B0(x07), .Y(men_men_n371_));
  AOI210     u349(.A0(men_men_n370_), .A1(x06), .B0(men_men_n371_), .Y(men_men_n372_));
  AOI220     u350(.A0(men_men_n79_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n373_));
  NO3        u351(.A(men_men_n373_), .B(men_men_n23_), .C(x00), .Y(men_men_n374_));
  NA2        u352(.A(men_men_n70_), .B(x02), .Y(men_men_n375_));
  AOI210     u353(.A0(men_men_n375_), .A1(men_men_n369_), .B0(men_men_n247_), .Y(men_men_n376_));
  OR2        u354(.A(men_men_n376_), .B(men_men_n231_), .Y(men_men_n377_));
  NO2        u355(.A(men_men_n23_), .B(x10), .Y(men_men_n378_));
  OAI210     u356(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n379_));
  OR3        u357(.A(men_men_n379_), .B(men_men_n378_), .C(men_men_n44_), .Y(men_men_n380_));
  NA2        u358(.A(men_men_n380_), .B(men_men_n377_), .Y(men_men_n381_));
  OAI210     u359(.A0(men_men_n381_), .A1(men_men_n374_), .B0(men_men_n99_), .Y(men_men_n382_));
  NA2        u360(.A(men_men_n33_), .B(men_men_n99_), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n383_), .A1(men_men_n90_), .B0(x07), .Y(men_men_n384_));
  AOI220     u362(.A0(men_men_n384_), .A1(men_men_n382_), .B0(men_men_n372_), .B1(men_men_n366_), .Y(men_men_n385_));
  BUFFER     u363(.A(men_men_n254_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n378_), .A1(x07), .B0(men_men_n134_), .Y(men_men_n387_));
  OR2        u365(.A(men_men_n387_), .B(x03), .Y(men_men_n388_));
  NO2        u366(.A(x07), .B(x11), .Y(men_men_n389_));
  NO3        u367(.A(men_men_n389_), .B(men_men_n138_), .C(men_men_n28_), .Y(men_men_n390_));
  AOI220     u368(.A0(men_men_n390_), .A1(men_men_n388_), .B0(men_men_n386_), .B1(men_men_n47_), .Y(men_men_n391_));
  NO3        u369(.A(men_men_n315_), .B(men_men_n32_), .C(x11), .Y(men_men_n392_));
  OAI210     u370(.A0(men_men_n392_), .A1(men_men_n391_), .B0(men_men_n100_), .Y(men_men_n393_));
  AOI210     u371(.A0(men_men_n324_), .A1(men_men_n109_), .B0(men_men_n253_), .Y(men_men_n394_));
  NOi21      u372(.An(men_men_n307_), .B(men_men_n127_), .Y(men_men_n395_));
  OAI210     u373(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n396_));
  AOI210     u374(.A0(men_men_n240_), .A1(men_men_n47_), .B0(men_men_n396_), .Y(men_men_n397_));
  NO3        u375(.A(men_men_n397_), .B(men_men_n394_), .C(x08), .Y(men_men_n398_));
  NA2        u376(.A(x09), .B(men_men_n41_), .Y(men_men_n399_));
  OAI210     u377(.A0(men_men_n367_), .A1(men_men_n66_), .B0(men_men_n399_), .Y(men_men_n400_));
  NO2        u378(.A(x13), .B(x12), .Y(men_men_n401_));
  NO2        u379(.A(men_men_n126_), .B(men_men_n28_), .Y(men_men_n402_));
  NO2        u380(.A(men_men_n402_), .B(men_men_n258_), .Y(men_men_n403_));
  NA3        u381(.A(men_men_n318_), .B(men_men_n121_), .C(x12), .Y(men_men_n404_));
  AO210      u382(.A0(men_men_n318_), .A1(men_men_n121_), .B0(men_men_n240_), .Y(men_men_n405_));
  NA3        u383(.A(men_men_n405_), .B(men_men_n404_), .C(x08), .Y(men_men_n406_));
  AOI210     u384(.A0(men_men_n401_), .A1(men_men_n400_), .B0(men_men_n406_), .Y(men_men_n407_));
  AOI210     u385(.A0(men_men_n398_), .A1(men_men_n393_), .B0(men_men_n407_), .Y(men_men_n408_));
  OAI210     u386(.A0(x07), .A1(men_men_n23_), .B0(x03), .Y(men_men_n409_));
  INV        u387(.A(x07), .Y(men_men_n410_));
  NO2        u388(.A(men_men_n410_), .B(men_men_n368_), .Y(men_men_n411_));
  OAI210     u389(.A0(men_men_n411_), .A1(men_men_n409_), .B0(men_men_n182_), .Y(men_men_n412_));
  NA3        u390(.A(men_men_n403_), .B(men_men_n395_), .C(men_men_n314_), .Y(men_men_n413_));
  INV        u391(.A(x14), .Y(men_men_n414_));
  NO3        u392(.A(men_men_n307_), .B(men_men_n105_), .C(x11), .Y(men_men_n415_));
  NO3        u393(.A(x06), .B(men_men_n315_), .C(men_men_n176_), .Y(men_men_n416_));
  NO3        u394(.A(men_men_n416_), .B(men_men_n415_), .C(men_men_n414_), .Y(men_men_n417_));
  NA3        u395(.A(men_men_n417_), .B(men_men_n413_), .C(men_men_n412_), .Y(men_men_n418_));
  AOI220     u396(.A0(men_men_n383_), .A1(men_men_n61_), .B0(men_men_n402_), .B1(men_men_n157_), .Y(men_men_n419_));
  NOi21      u397(.An(men_men_n263_), .B(men_men_n142_), .Y(men_men_n420_));
  NO3        u398(.A(men_men_n123_), .B(men_men_n24_), .C(x06), .Y(men_men_n421_));
  AOI210     u399(.A0(men_men_n269_), .A1(men_men_n223_), .B0(men_men_n421_), .Y(men_men_n422_));
  OAI210     u400(.A0(men_men_n44_), .A1(x04), .B0(men_men_n422_), .Y(men_men_n423_));
  OAI210     u401(.A0(men_men_n423_), .A1(men_men_n420_), .B0(men_men_n99_), .Y(men_men_n424_));
  OAI210     u402(.A0(men_men_n419_), .A1(men_men_n89_), .B0(men_men_n424_), .Y(men_men_n425_));
  NO4        u403(.A(men_men_n425_), .B(men_men_n418_), .C(men_men_n408_), .D(men_men_n385_), .Y(men06));
  INV        u404(.A(x07), .Y(men_men_n429_));
  INV        u405(.A(men_men_n88_), .Y(men_men_n430_));
  INV        u406(.A(x01), .Y(men_men_n431_));
  INV        u407(.A(x13), .Y(men_men_n432_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule