//Benchmark atmr_intb_466_0.0625

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n302_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n343_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n350_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n412_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n383_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n459_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  INV        o035(.A(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(ori_ori_n24_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n60_), .B(ori_ori_n58_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n62_));
  OAI210     o040(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o041(.A0(ori_ori_n63_), .A1(ori_ori_n55_), .B0(ori_ori_n61_), .B1(ori_ori_n31_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(x05), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n57_), .B(ori_ori_n23_), .Y(ori_ori_n66_));
  NA2        o044(.A(x09), .B(x05), .Y(ori_ori_n67_));
  NA2        o045(.A(x10), .B(x06), .Y(ori_ori_n68_));
  NA3        o046(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(ori_ori_n28_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n57_), .B(ori_ori_n41_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n69_), .A1(ori_ori_n66_), .B0(x03), .Y(ori_ori_n71_));
  NOi31      o049(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n72_));
  INV        o050(.A(x07), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n74_));
  NO2        o052(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n36_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n75_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n77_));
  AOI210     o055(.A0(ori_ori_n76_), .A1(ori_ori_n48_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n79_));
  NO2        o057(.A(x08), .B(x01), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n80_), .A1(ori_ori_n79_), .B0(ori_ori_n35_), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n82_));
  NO3        o060(.A(ori_ori_n81_), .B(ori_ori_n78_), .C(ori_ori_n74_), .Y(ori_ori_n83_));
  AN2        o061(.A(ori_ori_n83_), .B(ori_ori_n71_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n81_), .Y(ori_ori_n85_));
  NA2        o063(.A(x11), .B(x00), .Y(ori_ori_n86_));
  NO2        o064(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n87_));
  NOi21      o065(.An(ori_ori_n86_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  INV        o066(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  NOi21      o067(.An(x01), .B(x10), .Y(ori_ori_n90_));
  NO2        o068(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n91_));
  NO3        o069(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(x06), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n92_), .B(ori_ori_n27_), .Y(ori_ori_n93_));
  OAI210     o071(.A0(ori_ori_n89_), .A1(x07), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NO3        o072(.A(ori_ori_n94_), .B(ori_ori_n84_), .C(ori_ori_n65_), .Y(ori01));
  INV        o073(.A(x12), .Y(ori_ori_n96_));
  INV        o074(.A(x13), .Y(ori_ori_n97_));
  NO2        o075(.A(x10), .B(x01), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  NA2        o078(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n102_));
  NOi21      o080(.An(ori_ori_n102_), .B(ori_ori_n54_), .Y(ori_ori_n103_));
  NA2        o081(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(x05), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n106_));
  INV        o084(.A(ori_ori_n103_), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n107_), .B(ori_ori_n68_), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n109_));
  NA2        o087(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n110_), .B(ori_ori_n109_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n113_));
  INV        o091(.A(ori_ori_n111_), .Y(ori_ori_n114_));
  NO3        o092(.A(ori_ori_n114_), .B(x06), .C(x03), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n115_), .B(ori_ori_n108_), .Y(ori_ori_n116_));
  OAI210     o094(.A0(ori_ori_n80_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n119_));
  NO2        o097(.A(x09), .B(x05), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n47_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n100_), .B(ori_ori_n49_), .Y(ori_ori_n122_));
  NA2        o100(.A(x09), .B(x00), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n102_), .B(ori_ori_n123_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n124_), .B(ori_ori_n119_), .Y(ori_ori_n125_));
  NO2        o103(.A(ori_ori_n125_), .B(ori_ori_n122_), .Y(ori_ori_n126_));
  NO2        o104(.A(x03), .B(x02), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n81_), .B(ori_ori_n97_), .Y(ori_ori_n128_));
  OAI210     o106(.A0(ori_ori_n128_), .A1(ori_ori_n103_), .B0(ori_ori_n127_), .Y(ori_ori_n129_));
  OA210      o107(.A0(ori_ori_n126_), .A1(x11), .B0(ori_ori_n129_), .Y(ori_ori_n130_));
  OAI210     o108(.A0(ori_ori_n116_), .A1(ori_ori_n23_), .B0(ori_ori_n130_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n100_), .B(ori_ori_n40_), .Y(ori_ori_n132_));
  NAi21      o110(.An(x06), .B(x10), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n132_), .B(ori_ori_n41_), .Y(ori_ori_n134_));
  NO2        o112(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n97_), .B(x01), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n136_), .B(x08), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n135_), .B(ori_ori_n48_), .Y(ori_ori_n138_));
  AOI210     o116(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n139_));
  OAI210     o117(.A0(ori_ori_n138_), .A1(ori_ori_n134_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NA2        o118(.A(x04), .B(x02), .Y(ori_ori_n141_));
  NA2        o119(.A(x10), .B(x05), .Y(ori_ori_n142_));
  NO2        o120(.A(x09), .B(x01), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n102_), .B(x08), .Y(ori_ori_n144_));
  NAi21      o122(.An(x13), .B(x00), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n91_), .B(x06), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n145_), .B(ori_ori_n36_), .Y(ori_ori_n147_));
  INV        o125(.A(ori_ori_n147_), .Y(ori_ori_n148_));
  NOi21      o126(.An(x09), .B(x00), .Y(ori_ori_n149_));
  NO3        o127(.A(ori_ori_n79_), .B(ori_ori_n149_), .C(ori_ori_n47_), .Y(ori_ori_n150_));
  NA2        o128(.A(ori_ori_n150_), .B(ori_ori_n110_), .Y(ori_ori_n151_));
  NA2        o129(.A(x06), .B(x05), .Y(ori_ori_n152_));
  OAI210     o130(.A0(ori_ori_n152_), .A1(ori_ori_n35_), .B0(ori_ori_n96_), .Y(ori_ori_n153_));
  AOI210     o131(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n153_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n154_), .B(ori_ori_n151_), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n97_), .B(x12), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n158_));
  NA2        o136(.A(ori_ori_n158_), .B(x02), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n157_), .B(ori_ori_n155_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n140_), .Y(ori_ori_n161_));
  AOI210     o139(.A0(ori_ori_n131_), .A1(ori_ori_n96_), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n163_), .B(ori_ori_n117_), .Y(ori_ori_n164_));
  AOI210     o142(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n109_), .B(x06), .Y(ori_ori_n166_));
  AOI210     o144(.A0(ori_ori_n165_), .A1(ori_ori_n164_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n167_), .B(x12), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n72_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n90_), .B(x06), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n170_), .B(ori_ori_n41_), .Y(ori_ori_n171_));
  INV        o149(.A(ori_ori_n119_), .Y(ori_ori_n172_));
  OAI210     o150(.A0(ori_ori_n172_), .A1(ori_ori_n171_), .B0(x02), .Y(ori_ori_n173_));
  AOI210     o151(.A0(ori_ori_n173_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n174_));
  OAI210     o152(.A0(ori_ori_n168_), .A1(ori_ori_n53_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  INV        o153(.A(ori_ori_n119_), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n177_));
  NO2        o155(.A(ori_ori_n97_), .B(x03), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n179_));
  INV        o157(.A(ori_ori_n133_), .Y(ori_ori_n180_));
  NOi21      o158(.An(x13), .B(x04), .Y(ori_ori_n181_));
  NO3        o159(.A(ori_ori_n181_), .B(ori_ori_n72_), .C(ori_ori_n149_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n182_), .B(x05), .Y(ori_ori_n183_));
  AOI220     o161(.A0(ori_ori_n183_), .A1(ori_ori_n179_), .B0(ori_ori_n180_), .B1(ori_ori_n53_), .Y(ori_ori_n184_));
  INV        o162(.A(ori_ori_n184_), .Y(ori_ori_n185_));
  INV        o163(.A(ori_ori_n87_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n186_), .B(x12), .Y(ori_ori_n187_));
  NA2        o165(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n189_));
  NO2        o167(.A(x06), .B(x00), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n191_));
  INV        o169(.A(x03), .Y(ori_ori_n192_));
  OR2        o170(.A(ori_ori_n192_), .B(ori_ori_n68_), .Y(ori_ori_n193_));
  NA2        o171(.A(x13), .B(ori_ori_n96_), .Y(ori_ori_n194_));
  NA3        o172(.A(ori_ori_n194_), .B(ori_ori_n153_), .C(ori_ori_n88_), .Y(ori_ori_n195_));
  OAI210     o173(.A0(ori_ori_n193_), .A1(ori_ori_n188_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  AOI210     o174(.A0(ori_ori_n187_), .A1(ori_ori_n185_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  AOI210     o175(.A0(ori_ori_n197_), .A1(ori_ori_n175_), .B0(x07), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n67_), .B(ori_ori_n29_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n181_), .B(ori_ori_n149_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n200_), .B(ori_ori_n199_), .Y(ori_ori_n201_));
  NO2        o179(.A(x08), .B(x05), .Y(ori_ori_n202_));
  NA2        o180(.A(x13), .B(ori_ori_n31_), .Y(ori_ori_n203_));
  INV        o181(.A(ori_ori_n203_), .Y(ori_ori_n204_));
  NO2        o182(.A(x12), .B(x02), .Y(ori_ori_n205_));
  INV        o183(.A(ori_ori_n205_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(ori_ori_n186_), .Y(ori_ori_n207_));
  OA210      o185(.A0(ori_ori_n204_), .A1(ori_ori_n201_), .B0(ori_ori_n207_), .Y(ori_ori_n208_));
  NA2        o186(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n209_), .B(x01), .Y(ori_ori_n210_));
  NA2        o188(.A(ori_ori_n97_), .B(x04), .Y(ori_ori_n211_));
  NA2        o189(.A(ori_ori_n211_), .B(ori_ori_n28_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n212_), .B(ori_ori_n343_), .Y(ori_ori_n213_));
  NO3        o191(.A(ori_ori_n86_), .B(x12), .C(x03), .Y(ori_ori_n214_));
  NA2        o192(.A(ori_ori_n213_), .B(ori_ori_n214_), .Y(ori_ori_n215_));
  NOi21      o193(.An(ori_ori_n199_), .B(ori_ori_n170_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n216_), .B(ori_ori_n217_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n219_), .B(ori_ori_n146_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n188_), .B(ori_ori_n28_), .Y(ori_ori_n221_));
  OAI210     o199(.A0(ori_ori_n220_), .A1(ori_ori_n176_), .B0(ori_ori_n221_), .Y(ori_ori_n222_));
  NA3        o200(.A(ori_ori_n222_), .B(ori_ori_n218_), .C(ori_ori_n215_), .Y(ori_ori_n223_));
  NO3        o201(.A(ori_ori_n223_), .B(ori_ori_n208_), .C(ori_ori_n198_), .Y(ori_ori_n224_));
  OAI210     o202(.A0(ori_ori_n162_), .A1(ori_ori_n57_), .B0(ori_ori_n224_), .Y(ori02));
  NOi21      o203(.An(ori_ori_n182_), .B(ori_ori_n143_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(ori_ori_n32_), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n227_), .B(ori_ori_n142_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n229_));
  AOI210     o207(.A0(ori_ori_n229_), .A1(ori_ori_n228_), .B0(ori_ori_n48_), .Y(ori_ori_n230_));
  NO2        o208(.A(x05), .B(x02), .Y(ori_ori_n231_));
  OAI210     o209(.A0(ori_ori_n164_), .A1(ori_ori_n149_), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  AOI220     o210(.A0(ori_ori_n202_), .A1(ori_ori_n54_), .B0(ori_ori_n52_), .B1(ori_ori_n36_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n232_), .B(ori_ori_n119_), .Y(ori_ori_n234_));
  NO2        o212(.A(ori_ori_n191_), .B(ori_ori_n47_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n235_), .B(ori_ori_n183_), .Y(ori_ori_n236_));
  OAI210     o214(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n237_));
  NA2        o215(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n238_));
  BUFFER     o216(.A(ori_ori_n121_), .Y(ori_ori_n239_));
  AOI210     o217(.A0(ori_ori_n239_), .A1(ori_ori_n117_), .B0(ori_ori_n237_), .Y(ori_ori_n240_));
  NA2        o218(.A(ori_ori_n240_), .B(ori_ori_n91_), .Y(ori_ori_n241_));
  INV        o219(.A(ori_ori_n127_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n242_), .B(ori_ori_n111_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n243_), .B(x13), .Y(ori_ori_n244_));
  NA3        o222(.A(ori_ori_n244_), .B(ori_ori_n241_), .C(ori_ori_n236_), .Y(ori_ori_n245_));
  NO3        o223(.A(ori_ori_n245_), .B(ori_ori_n234_), .C(ori_ori_n230_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n118_), .B(x03), .Y(ori_ori_n247_));
  INV        o225(.A(ori_ori_n145_), .Y(ori_ori_n248_));
  AOI220     o226(.A0(x08), .A1(ori_ori_n248_), .B0(ori_ori_n158_), .B1(x08), .Y(ori_ori_n249_));
  OAI210     o227(.A0(ori_ori_n249_), .A1(ori_ori_n219_), .B0(ori_ori_n247_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n250_), .B(ori_ori_n98_), .Y(ori_ori_n251_));
  NA2        o229(.A(ori_ori_n141_), .B(ori_ori_n136_), .Y(ori_ori_n252_));
  AN2        o230(.A(ori_ori_n252_), .B(ori_ori_n144_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n112_), .B(ori_ori_n28_), .Y(ori_ori_n254_));
  OAI210     o232(.A0(ori_ori_n254_), .A1(ori_ori_n253_), .B0(ori_ori_n99_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n211_), .B(ori_ori_n96_), .Y(ori_ori_n256_));
  NA2        o234(.A(ori_ori_n96_), .B(ori_ori_n41_), .Y(ori_ori_n257_));
  NA3        o235(.A(ori_ori_n257_), .B(ori_ori_n256_), .C(ori_ori_n111_), .Y(ori_ori_n258_));
  NA4        o236(.A(ori_ori_n258_), .B(ori_ori_n255_), .C(ori_ori_n251_), .D(ori_ori_n48_), .Y(ori_ori_n259_));
  INV        o237(.A(ori_ori_n158_), .Y(ori_ori_n260_));
  INV        o238(.A(ori_ori_n40_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n262_));
  OAI220     o240(.A0(ori_ori_n262_), .A1(ori_ori_n261_), .B0(ori_ori_n260_), .B1(ori_ori_n55_), .Y(ori_ori_n263_));
  NA2        o241(.A(ori_ori_n263_), .B(x02), .Y(ori_ori_n264_));
  INV        o242(.A(ori_ori_n189_), .Y(ori_ori_n265_));
  NA2        o243(.A(ori_ori_n156_), .B(x04), .Y(ori_ori_n266_));
  NO3        o244(.A(ori_ori_n156_), .B(ori_ori_n135_), .C(ori_ori_n51_), .Y(ori_ori_n267_));
  OAI210     o245(.A0(ori_ori_n123_), .A1(ori_ori_n36_), .B0(ori_ori_n96_), .Y(ori_ori_n268_));
  OAI210     o246(.A0(ori_ori_n268_), .A1(ori_ori_n150_), .B0(ori_ori_n267_), .Y(ori_ori_n269_));
  NA3        o247(.A(ori_ori_n269_), .B(ori_ori_n264_), .C(x06), .Y(ori_ori_n270_));
  NA2        o248(.A(x09), .B(x03), .Y(ori_ori_n271_));
  OAI220     o249(.A0(ori_ori_n271_), .A1(ori_ori_n110_), .B0(ori_ori_n163_), .B1(ori_ori_n59_), .Y(ori_ori_n272_));
  NO3        o250(.A(ori_ori_n219_), .B(ori_ori_n109_), .C(x08), .Y(ori_ori_n273_));
  INV        o251(.A(ori_ori_n273_), .Y(ori_ori_n274_));
  NO2        o252(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n275_));
  NO3        o253(.A(ori_ori_n102_), .B(ori_ori_n110_), .C(ori_ori_n38_), .Y(ori_ori_n276_));
  AOI210     o254(.A0(ori_ori_n267_), .A1(ori_ori_n275_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  OAI210     o255(.A0(ori_ori_n274_), .A1(ori_ori_n28_), .B0(ori_ori_n277_), .Y(ori_ori_n278_));
  AO220      o256(.A0(ori_ori_n278_), .A1(x04), .B0(ori_ori_n272_), .B1(x05), .Y(ori_ori_n279_));
  AOI210     o257(.A0(ori_ori_n270_), .A1(ori_ori_n259_), .B0(ori_ori_n279_), .Y(ori_ori_n280_));
  OAI210     o258(.A0(ori_ori_n246_), .A1(x12), .B0(ori_ori_n280_), .Y(ori03));
  OR2        o259(.A(ori_ori_n42_), .B(ori_ori_n177_), .Y(ori_ori_n282_));
  AOI210     o260(.A0(ori_ori_n128_), .A1(ori_ori_n96_), .B0(ori_ori_n282_), .Y(ori_ori_n283_));
  AO210      o261(.A0(ori_ori_n265_), .A1(ori_ori_n82_), .B0(ori_ori_n266_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n156_), .B(ori_ori_n127_), .Y(ori_ori_n285_));
  NA3        o263(.A(ori_ori_n285_), .B(ori_ori_n284_), .C(ori_ori_n159_), .Y(ori_ori_n286_));
  OAI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n283_), .B0(x05), .Y(ori_ori_n287_));
  NA2        o265(.A(ori_ori_n282_), .B(x05), .Y(ori_ori_n288_));
  AOI210     o266(.A0(ori_ori_n117_), .A1(ori_ori_n169_), .B0(ori_ori_n288_), .Y(ori_ori_n289_));
  AOI210     o267(.A0(ori_ori_n178_), .A1(ori_ori_n76_), .B0(ori_ori_n105_), .Y(ori_ori_n290_));
  OAI220     o268(.A0(ori_ori_n290_), .A1(ori_ori_n55_), .B0(ori_ori_n238_), .B1(ori_ori_n233_), .Y(ori_ori_n291_));
  OAI210     o269(.A0(ori_ori_n291_), .A1(ori_ori_n289_), .B0(ori_ori_n96_), .Y(ori_ori_n292_));
  AOI210     o270(.A0(ori_ori_n121_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n143_), .B(ori_ori_n113_), .Y(ori_ori_n294_));
  OAI220     o272(.A0(ori_ori_n294_), .A1(ori_ori_n37_), .B0(ori_ori_n124_), .B1(x13), .Y(ori_ori_n295_));
  OAI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n293_), .B0(x04), .Y(ori_ori_n296_));
  NO3        o274(.A(ori_ori_n257_), .B(ori_ori_n81_), .C(ori_ori_n55_), .Y(ori_ori_n297_));
  AOI210     o275(.A0(ori_ori_n148_), .A1(ori_ori_n96_), .B0(ori_ori_n121_), .Y(ori_ori_n298_));
  OA210      o276(.A0(ori_ori_n137_), .A1(x12), .B0(ori_ori_n113_), .Y(ori_ori_n299_));
  NO3        o277(.A(ori_ori_n299_), .B(ori_ori_n298_), .C(ori_ori_n297_), .Y(ori_ori_n300_));
  NA4        o278(.A(ori_ori_n300_), .B(ori_ori_n296_), .C(ori_ori_n292_), .D(ori_ori_n287_), .Y(ori04));
  NO2        o279(.A(ori_ori_n85_), .B(ori_ori_n39_), .Y(ori_ori_n302_));
  XO2        o280(.A(ori_ori_n302_), .B(ori_ori_n194_), .Y(ori05));
  OAI210     o281(.A0(ori_ori_n26_), .A1(ori_ori_n96_), .B0(x07), .Y(ori_ori_n304_));
  INV        o282(.A(ori_ori_n304_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n190_), .B(ori_ori_n186_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n306_), .B(ori_ori_n188_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n307_), .B(ori_ori_n96_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n33_), .B(ori_ori_n96_), .Y(ori_ori_n309_));
  AOI210     o287(.A0(ori_ori_n309_), .A1(ori_ori_n87_), .B0(x07), .Y(ori_ori_n310_));
  AOI210     o288(.A0(ori_ori_n310_), .A1(ori_ori_n308_), .B0(ori_ori_n305_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n47_), .B(x02), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n312_), .B(ori_ori_n97_), .Y(ori_ori_n313_));
  AOI210     o291(.A0(ori_ori_n266_), .A1(ori_ori_n101_), .B0(ori_ori_n205_), .Y(ori_ori_n314_));
  NOi21      o292(.An(ori_ori_n247_), .B(ori_ori_n113_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n315_), .B(ori_ori_n206_), .Y(ori_ori_n316_));
  OAI210     o294(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n317_));
  AOI210     o295(.A0(ori_ori_n194_), .A1(ori_ori_n47_), .B0(ori_ori_n317_), .Y(ori_ori_n318_));
  NO4        o296(.A(ori_ori_n318_), .B(ori_ori_n316_), .C(ori_ori_n314_), .D(x08), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n112_), .B(ori_ori_n28_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n320_), .B(ori_ori_n210_), .Y(ori_ori_n321_));
  OR3        o299(.A(ori_ori_n321_), .B(x12), .C(x03), .Y(ori_ori_n322_));
  NA3        o300(.A(ori_ori_n260_), .B(ori_ori_n106_), .C(x12), .Y(ori_ori_n323_));
  AO210      o301(.A0(ori_ori_n260_), .A1(ori_ori_n106_), .B0(ori_ori_n194_), .Y(ori_ori_n324_));
  NA4        o302(.A(ori_ori_n324_), .B(ori_ori_n323_), .C(ori_ori_n322_), .D(x08), .Y(ori_ori_n325_));
  INV        o303(.A(ori_ori_n325_), .Y(ori_ori_n326_));
  AOI210     o304(.A0(ori_ori_n319_), .A1(ori_ori_n313_), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  INV        o305(.A(x03), .Y(ori_ori_n328_));
  NA2        o306(.A(ori_ori_n328_), .B(ori_ori_n147_), .Y(ori_ori_n329_));
  NA3        o307(.A(ori_ori_n321_), .B(ori_ori_n315_), .C(ori_ori_n256_), .Y(ori_ori_n330_));
  INV        o308(.A(x14), .Y(ori_ori_n331_));
  NO3        o309(.A(ori_ori_n136_), .B(ori_ori_n70_), .C(ori_ori_n53_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n332_), .B(ori_ori_n331_), .Y(ori_ori_n333_));
  NA3        o311(.A(ori_ori_n333_), .B(ori_ori_n330_), .C(ori_ori_n329_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n309_), .B(ori_ori_n57_), .Y(ori_ori_n335_));
  INV        o313(.A(ori_ori_n124_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n337_));
  OAI210     o315(.A0(ori_ori_n337_), .A1(ori_ori_n336_), .B0(ori_ori_n96_), .Y(ori_ori_n338_));
  OAI210     o316(.A0(ori_ori_n335_), .A1(ori_ori_n86_), .B0(ori_ori_n338_), .Y(ori_ori_n339_));
  NO4        o317(.A(ori_ori_n339_), .B(ori_ori_n334_), .C(ori_ori_n327_), .D(ori_ori_n311_), .Y(ori06));
  INV        o318(.A(x13), .Y(ori_ori_n343_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA3        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n28_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n61_), .B(mai_mai_n41_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n73_), .A1(x11), .B0(x03), .Y(mai_mai_n75_));
  NOi31      m053(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n76_));
  INV        m054(.A(mai_mai_n24_), .Y(mai_mai_n77_));
  NO2        m055(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n78_), .B(mai_mai_n36_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n78_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n80_));
  AOI210     m058(.A0(mai_mai_n79_), .A1(mai_mai_n48_), .B0(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m059(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n82_));
  NO2        m060(.A(x08), .B(x01), .Y(mai_mai_n83_));
  OAI210     m061(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n35_), .Y(mai_mai_n84_));
  NA2        m062(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n84_), .B(mai_mai_n81_), .C(mai_mai_n77_), .Y(mai_mai_n86_));
  AN2        m064(.A(mai_mai_n86_), .B(mai_mai_n75_), .Y(mai_mai_n87_));
  INV        m065(.A(mai_mai_n84_), .Y(mai_mai_n88_));
  NO2        m066(.A(x06), .B(x05), .Y(mai_mai_n89_));
  NA2        m067(.A(x11), .B(x00), .Y(mai_mai_n90_));
  NO2        m068(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n91_));
  NOi21      m069(.An(mai_mai_n90_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  AOI210     m070(.A0(mai_mai_n89_), .A1(mai_mai_n88_), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  NOi21      m071(.An(x01), .B(x10), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n95_));
  NO3        m073(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(x06), .Y(mai_mai_n96_));
  NA2        m074(.A(mai_mai_n96_), .B(mai_mai_n27_), .Y(mai_mai_n97_));
  OAI210     m075(.A0(mai_mai_n93_), .A1(x07), .B0(mai_mai_n97_), .Y(mai_mai_n98_));
  NO3        m076(.A(mai_mai_n98_), .B(mai_mai_n87_), .C(mai_mai_n70_), .Y(mai01));
  INV        m077(.A(x12), .Y(mai_mai_n100_));
  INV        m078(.A(x13), .Y(mai_mai_n101_));
  NA2        m079(.A(x08), .B(x04), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n94_), .B(mai_mai_n28_), .Y(mai_mai_n103_));
  NO2        m081(.A(x10), .B(x01), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n105_), .B(mai_mai_n104_), .Y(mai_mai_n106_));
  NA2        m084(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n107_));
  NO3        m085(.A(mai_mai_n107_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n101_), .B(mai_mai_n36_), .Y(mai_mai_n110_));
  NA3        m088(.A(mai_mai_n110_), .B(x04), .C(x06), .Y(mai_mai_n111_));
  INV        m089(.A(mai_mai_n111_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n83_), .B(x13), .Y(mai_mai_n113_));
  NA2        m091(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n114_), .B(x05), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n116_));
  AOI210     m094(.A0(x00), .A1(mai_mai_n113_), .B0(mai_mai_n72_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n118_));
  NA2        m096(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n122_));
  NOi41      m100(.An(mai_mai_n412_), .B(mai_mai_n122_), .C(mai_mai_n57_), .D(mai_mai_n120_), .Y(mai_mai_n123_));
  NO3        m101(.A(mai_mai_n123_), .B(x06), .C(x03), .Y(mai_mai_n124_));
  NO4        m102(.A(mai_mai_n124_), .B(mai_mai_n117_), .C(mai_mai_n112_), .D(mai_mai_n108_), .Y(mai_mai_n125_));
  NA2        m103(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n126_));
  OAI210     m104(.A0(mai_mai_n83_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n130_));
  AOI210     m108(.A0(mai_mai_n130_), .A1(mai_mai_n49_), .B0(mai_mai_n129_), .Y(mai_mai_n131_));
  AN2        m109(.A(mai_mai_n131_), .B(mai_mai_n128_), .Y(mai_mai_n132_));
  NO2        m110(.A(x09), .B(x05), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n47_), .Y(mai_mai_n134_));
  AOI210     m112(.A0(mai_mai_n134_), .A1(mai_mai_n106_), .B0(mai_mai_n49_), .Y(mai_mai_n135_));
  NA2        m113(.A(x09), .B(x00), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n109_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n76_), .B(mai_mai_n51_), .Y(mai_mai_n138_));
  AOI210     m116(.A0(mai_mai_n138_), .A1(mai_mai_n137_), .B0(mai_mai_n130_), .Y(mai_mai_n139_));
  NO3        m117(.A(mai_mai_n139_), .B(mai_mai_n135_), .C(mai_mai_n132_), .Y(mai_mai_n140_));
  NO2        m118(.A(x03), .B(x02), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n84_), .B(mai_mai_n101_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  OA210      m121(.A0(mai_mai_n140_), .A1(x11), .B0(mai_mai_n143_), .Y(mai_mai_n144_));
  OAI210     m122(.A0(mai_mai_n125_), .A1(mai_mai_n23_), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n106_), .B(mai_mai_n40_), .Y(mai_mai_n146_));
  NAi21      m124(.An(x06), .B(x10), .Y(mai_mai_n147_));
  NOi21      m125(.An(x01), .B(x13), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n147_), .Y(mai_mai_n149_));
  AOI210     m127(.A0(mai_mai_n149_), .A1(mai_mai_n146_), .B0(mai_mai_n41_), .Y(mai_mai_n150_));
  NO2        m128(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n101_), .B(x01), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n152_), .B(x08), .Y(mai_mai_n153_));
  OAI210     m131(.A0(x05), .A1(mai_mai_n153_), .B0(mai_mai_n51_), .Y(mai_mai_n154_));
  AOI210     m132(.A0(mai_mai_n154_), .A1(mai_mai_n151_), .B0(mai_mai_n48_), .Y(mai_mai_n155_));
  AOI210     m133(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n156_));
  OAI210     m134(.A0(mai_mai_n155_), .A1(mai_mai_n150_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NA2        m135(.A(x04), .B(x02), .Y(mai_mai_n158_));
  NA2        m136(.A(x10), .B(x05), .Y(mai_mai_n159_));
  NO2        m137(.A(x09), .B(x01), .Y(mai_mai_n160_));
  INV        m138(.A(x08), .Y(mai_mai_n161_));
  NA3        m139(.A(mai_mai_n148_), .B(mai_mai_n147_), .C(mai_mai_n51_), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n94_), .B(x05), .Y(mai_mai_n163_));
  OAI210     m141(.A0(mai_mai_n163_), .A1(mai_mai_n110_), .B0(mai_mai_n162_), .Y(mai_mai_n164_));
  AOI210     m142(.A0(mai_mai_n161_), .A1(x06), .B0(mai_mai_n164_), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n165_), .B(x11), .Y(mai_mai_n166_));
  NAi21      m144(.An(mai_mai_n158_), .B(mai_mai_n166_), .Y(mai_mai_n167_));
  INV        m145(.A(mai_mai_n25_), .Y(mai_mai_n168_));
  NAi21      m146(.An(x13), .B(x00), .Y(mai_mai_n169_));
  AOI210     m147(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n169_), .Y(mai_mai_n170_));
  AOI220     m148(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n171_));
  OAI210     m149(.A0(mai_mai_n159_), .A1(mai_mai_n35_), .B0(mai_mai_n171_), .Y(mai_mai_n172_));
  AN2        m150(.A(mai_mai_n172_), .B(mai_mai_n170_), .Y(mai_mai_n173_));
  AN2        m151(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n174_));
  NO2        m152(.A(mai_mai_n169_), .B(mai_mai_n36_), .Y(mai_mai_n175_));
  INV        m153(.A(mai_mai_n175_), .Y(mai_mai_n176_));
  OAI210     m154(.A0(mai_mai_n57_), .A1(mai_mai_n174_), .B0(mai_mai_n176_), .Y(mai_mai_n177_));
  OAI210     m155(.A0(mai_mai_n177_), .A1(mai_mai_n173_), .B0(mai_mai_n168_), .Y(mai_mai_n178_));
  NOi21      m156(.An(x09), .B(x00), .Y(mai_mai_n179_));
  NO3        m157(.A(mai_mai_n82_), .B(mai_mai_n179_), .C(mai_mai_n47_), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n180_), .B(mai_mai_n119_), .Y(mai_mai_n181_));
  NA2        m159(.A(x06), .B(x05), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n100_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n101_), .B(x12), .Y(mai_mai_n184_));
  AOI210     m162(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n184_), .Y(mai_mai_n185_));
  NA2        m163(.A(mai_mai_n94_), .B(mai_mai_n51_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n187_));
  NA2        m165(.A(mai_mai_n187_), .B(x02), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n188_), .B(mai_mai_n186_), .Y(mai_mai_n189_));
  AOI210     m167(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(mai_mai_n189_), .Y(mai_mai_n190_));
  NA4        m168(.A(mai_mai_n190_), .B(mai_mai_n178_), .C(mai_mai_n167_), .D(mai_mai_n157_), .Y(mai_mai_n191_));
  AOI210     m169(.A0(mai_mai_n145_), .A1(mai_mai_n100_), .B0(mai_mai_n191_), .Y(mai_mai_n192_));
  INV        m170(.A(mai_mai_n73_), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n193_), .B(mai_mai_n128_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n195_), .B(mai_mai_n127_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n118_), .B(x06), .Y(mai_mai_n197_));
  INV        m175(.A(mai_mai_n197_), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n198_), .A1(mai_mai_n194_), .B0(x12), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n76_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n149_), .B(mai_mai_n57_), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n201_), .B(mai_mai_n200_), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n94_), .B(x06), .Y(mai_mai_n203_));
  NA4        m181(.A(mai_mai_n147_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n204_));
  NA2        m182(.A(mai_mai_n204_), .B(mai_mai_n130_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n205_), .B(x02), .Y(mai_mai_n206_));
  AOI210     m184(.A0(mai_mai_n206_), .A1(mai_mai_n202_), .B0(mai_mai_n23_), .Y(mai_mai_n207_));
  OAI210     m185(.A0(mai_mai_n199_), .A1(mai_mai_n57_), .B0(mai_mai_n207_), .Y(mai_mai_n208_));
  INV        m186(.A(mai_mai_n130_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n101_), .B(x03), .Y(mai_mai_n211_));
  AOI210     m189(.A0(mai_mai_n76_), .A1(mai_mai_n210_), .B0(mai_mai_n211_), .Y(mai_mai_n212_));
  INV        m190(.A(mai_mai_n147_), .Y(mai_mai_n213_));
  NOi21      m191(.An(x13), .B(x04), .Y(mai_mai_n214_));
  NO3        m192(.A(mai_mai_n214_), .B(mai_mai_n76_), .C(mai_mai_n179_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n215_), .B(x05), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n213_), .B(mai_mai_n57_), .Y(mai_mai_n217_));
  OAI210     m195(.A0(mai_mai_n212_), .A1(mai_mai_n209_), .B0(mai_mai_n217_), .Y(mai_mai_n218_));
  INV        m196(.A(mai_mai_n91_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n219_), .B(x12), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n222_));
  OAI210     m200(.A0(mai_mai_n222_), .A1(mai_mai_n172_), .B0(mai_mai_n170_), .Y(mai_mai_n223_));
  AOI210     m201(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n224_));
  OAI210     m202(.A0(mai_mai_n102_), .A1(mai_mai_n136_), .B0(mai_mai_n72_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n225_), .B(x05), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n227_));
  NA2        m205(.A(mai_mai_n227_), .B(x03), .Y(mai_mai_n228_));
  OA210      m206(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n223_), .Y(mai_mai_n229_));
  NA2        m207(.A(x13), .B(mai_mai_n100_), .Y(mai_mai_n230_));
  NA3        m208(.A(mai_mai_n230_), .B(x12), .C(mai_mai_n92_), .Y(mai_mai_n231_));
  OAI210     m209(.A0(mai_mai_n229_), .A1(mai_mai_n221_), .B0(mai_mai_n231_), .Y(mai_mai_n232_));
  AOI210     m210(.A0(mai_mai_n220_), .A1(mai_mai_n218_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  AOI210     m211(.A0(mai_mai_n233_), .A1(mai_mai_n208_), .B0(x07), .Y(mai_mai_n234_));
  NA2        m212(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n235_));
  AOI210     m213(.A0(mai_mai_n126_), .A1(mai_mai_n138_), .B0(mai_mai_n235_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n101_), .B(x06), .Y(mai_mai_n237_));
  INV        m215(.A(mai_mai_n237_), .Y(mai_mai_n238_));
  NO2        m216(.A(x08), .B(x05), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n239_), .B(mai_mai_n224_), .Y(mai_mai_n240_));
  OAI210     m218(.A0(mai_mai_n76_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n241_));
  OAI210     m219(.A0(mai_mai_n240_), .A1(mai_mai_n238_), .B0(mai_mai_n241_), .Y(mai_mai_n242_));
  NO2        m220(.A(x12), .B(x02), .Y(mai_mai_n243_));
  INV        m221(.A(mai_mai_n243_), .Y(mai_mai_n244_));
  NO2        m222(.A(mai_mai_n244_), .B(mai_mai_n219_), .Y(mai_mai_n245_));
  OA210      m223(.A0(mai_mai_n242_), .A1(mai_mai_n236_), .B0(mai_mai_n245_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n247_));
  NO2        m225(.A(mai_mai_n247_), .B(x01), .Y(mai_mai_n248_));
  BUFFER     m226(.A(mai_mai_n83_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n249_), .B(mai_mai_n248_), .Y(mai_mai_n250_));
  AOI210     m228(.A0(mai_mai_n250_), .A1(mai_mai_n412_), .B0(mai_mai_n29_), .Y(mai_mai_n251_));
  INV        m229(.A(mai_mai_n237_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n101_), .B(x04), .Y(mai_mai_n253_));
  OAI210     m231(.A0(x02), .A1(mai_mai_n113_), .B0(mai_mai_n252_), .Y(mai_mai_n254_));
  NO3        m232(.A(mai_mai_n90_), .B(x12), .C(x03), .Y(mai_mai_n255_));
  OAI210     m233(.A0(mai_mai_n254_), .A1(mai_mai_n251_), .B0(mai_mai_n255_), .Y(mai_mai_n256_));
  AOI210     m234(.A0(mai_mai_n186_), .A1(mai_mai_n182_), .B0(mai_mai_n102_), .Y(mai_mai_n257_));
  NOi21      m235(.An(mai_mai_n235_), .B(mai_mai_n203_), .Y(mai_mai_n258_));
  NO2        m236(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n259_));
  OAI210     m237(.A0(mai_mai_n258_), .A1(mai_mai_n257_), .B0(mai_mai_n259_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n221_), .B(mai_mai_n28_), .Y(mai_mai_n261_));
  NA2        m239(.A(mai_mai_n209_), .B(mai_mai_n261_), .Y(mai_mai_n262_));
  NA3        m240(.A(mai_mai_n262_), .B(mai_mai_n260_), .C(mai_mai_n256_), .Y(mai_mai_n263_));
  NO3        m241(.A(mai_mai_n263_), .B(mai_mai_n246_), .C(mai_mai_n234_), .Y(mai_mai_n264_));
  OAI210     m242(.A0(mai_mai_n192_), .A1(mai_mai_n61_), .B0(mai_mai_n264_), .Y(mai02));
  AOI210     m243(.A0(mai_mai_n126_), .A1(mai_mai_n84_), .B0(mai_mai_n121_), .Y(mai_mai_n266_));
  NOi21      m244(.An(mai_mai_n215_), .B(mai_mai_n160_), .Y(mai_mai_n267_));
  NO2        m245(.A(mai_mai_n101_), .B(mai_mai_n35_), .Y(mai_mai_n268_));
  NA3        m246(.A(mai_mai_n268_), .B(x08), .C(mai_mai_n56_), .Y(mai_mai_n269_));
  OAI210     m247(.A0(mai_mai_n267_), .A1(mai_mai_n32_), .B0(mai_mai_n269_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n266_), .B0(mai_mai_n159_), .Y(mai_mai_n271_));
  INV        m249(.A(mai_mai_n159_), .Y(mai_mai_n272_));
  AOI210     m250(.A0(x04), .A1(mai_mai_n85_), .B0(x09), .Y(mai_mai_n273_));
  OAI220     m251(.A0(mai_mai_n273_), .A1(mai_mai_n101_), .B0(mai_mai_n84_), .B1(mai_mai_n51_), .Y(mai_mai_n274_));
  AOI220     m252(.A0(mai_mai_n274_), .A1(mai_mai_n272_), .B0(mai_mai_n142_), .B1(mai_mai_n141_), .Y(mai_mai_n275_));
  AOI210     m253(.A0(mai_mai_n275_), .A1(mai_mai_n271_), .B0(mai_mai_n48_), .Y(mai_mai_n276_));
  NO2        m254(.A(x05), .B(x02), .Y(mai_mai_n277_));
  OAI210     m255(.A0(mai_mai_n196_), .A1(mai_mai_n179_), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  AOI220     m256(.A0(mai_mai_n239_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n279_));
  NOi21      m257(.An(mai_mai_n268_), .B(mai_mai_n279_), .Y(mai_mai_n280_));
  AOI210     m258(.A0(mai_mai_n214_), .A1(mai_mai_n78_), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  AOI210     m259(.A0(mai_mai_n281_), .A1(mai_mai_n278_), .B0(mai_mai_n130_), .Y(mai_mai_n282_));
  NAi21      m260(.An(mai_mai_n216_), .B(mai_mai_n212_), .Y(mai_mai_n283_));
  NO2        m261(.A(mai_mai_n227_), .B(mai_mai_n47_), .Y(mai_mai_n284_));
  NA2        m262(.A(mai_mai_n284_), .B(mai_mai_n283_), .Y(mai_mai_n285_));
  OAI210     m263(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n286_));
  NA2        m264(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n287_));
  OA210      m265(.A0(mai_mai_n287_), .A1(x08), .B0(mai_mai_n134_), .Y(mai_mai_n288_));
  AOI210     m266(.A0(mai_mai_n288_), .A1(mai_mai_n127_), .B0(mai_mai_n286_), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n289_), .A1(mai_mai_n211_), .B0(mai_mai_n95_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n95_), .B(mai_mai_n83_), .C(mai_mai_n210_), .Y(mai_mai_n291_));
  NA3        m269(.A(mai_mai_n94_), .B(mai_mai_n82_), .C(mai_mai_n42_), .Y(mai_mai_n292_));
  AOI210     m270(.A0(mai_mai_n292_), .A1(mai_mai_n291_), .B0(x04), .Y(mai_mai_n293_));
  NO2        m271(.A(mai_mai_n240_), .B(mai_mai_n103_), .Y(mai_mai_n294_));
  AOI210     m272(.A0(mai_mai_n294_), .A1(x13), .B0(mai_mai_n293_), .Y(mai_mai_n295_));
  NA3        m273(.A(mai_mai_n295_), .B(mai_mai_n290_), .C(mai_mai_n285_), .Y(mai_mai_n296_));
  NO3        m274(.A(mai_mai_n296_), .B(mai_mai_n282_), .C(mai_mai_n276_), .Y(mai_mai_n297_));
  NA2        m275(.A(mai_mai_n129_), .B(x03), .Y(mai_mai_n298_));
  OAI210     m276(.A0(mai_mai_n169_), .A1(mai_mai_n51_), .B0(mai_mai_n298_), .Y(mai_mai_n299_));
  NA2        m277(.A(mai_mai_n299_), .B(mai_mai_n104_), .Y(mai_mai_n300_));
  INV        m278(.A(mai_mai_n56_), .Y(mai_mai_n301_));
  OAI220     m279(.A0(mai_mai_n253_), .A1(mai_mai_n301_), .B0(mai_mai_n121_), .B1(mai_mai_n28_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n302_), .B(mai_mai_n105_), .Y(mai_mai_n303_));
  NA2        m281(.A(mai_mai_n253_), .B(mai_mai_n100_), .Y(mai_mai_n304_));
  NA2        m282(.A(mai_mai_n100_), .B(mai_mai_n41_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n305_), .B(mai_mai_n304_), .C(mai_mai_n120_), .Y(mai_mai_n306_));
  NA4        m284(.A(mai_mai_n306_), .B(mai_mai_n303_), .C(mai_mai_n300_), .D(mai_mai_n48_), .Y(mai_mai_n307_));
  INV        m285(.A(mai_mai_n187_), .Y(mai_mai_n308_));
  NO2        m286(.A(mai_mai_n153_), .B(mai_mai_n40_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n310_));
  OAI220     m288(.A0(mai_mai_n310_), .A1(mai_mai_n309_), .B0(mai_mai_n308_), .B1(mai_mai_n59_), .Y(mai_mai_n311_));
  NA2        m289(.A(mai_mai_n311_), .B(x02), .Y(mai_mai_n312_));
  INV        m290(.A(mai_mai_n222_), .Y(mai_mai_n313_));
  NA2        m291(.A(mai_mai_n184_), .B(x04), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n314_), .B(mai_mai_n313_), .Y(mai_mai_n315_));
  NO3        m293(.A(mai_mai_n171_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n316_));
  OAI210     m294(.A0(mai_mai_n316_), .A1(mai_mai_n315_), .B0(mai_mai_n95_), .Y(mai_mai_n317_));
  NO3        m295(.A(mai_mai_n184_), .B(mai_mai_n151_), .C(mai_mai_n52_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(x12), .A1(mai_mai_n180_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  NA4        m297(.A(mai_mai_n319_), .B(mai_mai_n317_), .C(mai_mai_n312_), .D(x06), .Y(mai_mai_n320_));
  NA2        m298(.A(x09), .B(x03), .Y(mai_mai_n321_));
  OAI220     m299(.A0(mai_mai_n321_), .A1(mai_mai_n119_), .B0(mai_mai_n195_), .B1(mai_mai_n64_), .Y(mai_mai_n322_));
  OAI220     m300(.A0(mai_mai_n152_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n323_), .B(mai_mai_n209_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n324_), .B(mai_mai_n28_), .Y(mai_mai_n326_));
  AO220      m304(.A0(mai_mai_n326_), .A1(x04), .B0(mai_mai_n322_), .B1(x05), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n320_), .A1(mai_mai_n307_), .B0(mai_mai_n327_), .Y(mai_mai_n328_));
  OAI210     m306(.A0(mai_mai_n297_), .A1(x12), .B0(mai_mai_n328_), .Y(mai03));
  OR2        m307(.A(mai_mai_n42_), .B(mai_mai_n210_), .Y(mai_mai_n330_));
  AOI210     m308(.A0(mai_mai_n142_), .A1(mai_mai_n100_), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  AO210      m309(.A0(mai_mai_n313_), .A1(mai_mai_n85_), .B0(mai_mai_n314_), .Y(mai_mai_n332_));
  NA2        m310(.A(mai_mai_n184_), .B(mai_mai_n141_), .Y(mai_mai_n333_));
  NA3        m311(.A(mai_mai_n333_), .B(mai_mai_n332_), .C(mai_mai_n188_), .Y(mai_mai_n334_));
  OAI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n331_), .B0(x05), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n330_), .B(x05), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n127_), .A1(mai_mai_n200_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  AOI210     m315(.A0(mai_mai_n211_), .A1(mai_mai_n79_), .B0(mai_mai_n115_), .Y(mai_mai_n338_));
  OAI220     m316(.A0(mai_mai_n338_), .A1(mai_mai_n59_), .B0(mai_mai_n287_), .B1(mai_mai_n279_), .Y(mai_mai_n339_));
  OAI210     m317(.A0(mai_mai_n339_), .A1(mai_mai_n337_), .B0(mai_mai_n100_), .Y(mai_mai_n340_));
  AOI210     m318(.A0(mai_mai_n134_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n341_));
  NO2        m319(.A(mai_mai_n160_), .B(mai_mai_n122_), .Y(mai_mai_n342_));
  OAI220     m320(.A0(mai_mai_n342_), .A1(mai_mai_n37_), .B0(mai_mai_n137_), .B1(x13), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(x04), .Y(mai_mai_n344_));
  NO3        m322(.A(mai_mai_n305_), .B(mai_mai_n84_), .C(mai_mai_n59_), .Y(mai_mai_n345_));
  AOI210     m323(.A0(mai_mai_n176_), .A1(mai_mai_n100_), .B0(mai_mai_n134_), .Y(mai_mai_n346_));
  OA210      m324(.A0(mai_mai_n153_), .A1(x12), .B0(mai_mai_n122_), .Y(mai_mai_n347_));
  NO3        m325(.A(mai_mai_n347_), .B(mai_mai_n346_), .C(mai_mai_n345_), .Y(mai_mai_n348_));
  NA4        m326(.A(mai_mai_n348_), .B(mai_mai_n344_), .C(mai_mai_n340_), .D(mai_mai_n335_), .Y(mai04));
  NO2        m327(.A(mai_mai_n88_), .B(mai_mai_n39_), .Y(mai_mai_n350_));
  XO2        m328(.A(mai_mai_n350_), .B(mai_mai_n230_), .Y(mai05));
  AOI210     m329(.A0(mai_mai_n71_), .A1(mai_mai_n52_), .B0(mai_mai_n197_), .Y(mai_mai_n352_));
  AOI210     m330(.A0(mai_mai_n352_), .A1(mai_mai_n286_), .B0(mai_mai_n25_), .Y(mai_mai_n353_));
  NA3        m331(.A(mai_mai_n130_), .B(mai_mai_n121_), .C(mai_mai_n31_), .Y(mai_mai_n354_));
  AOI210     m332(.A0(x06), .A1(mai_mai_n354_), .B0(mai_mai_n24_), .Y(mai_mai_n355_));
  OAI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n353_), .B0(mai_mai_n100_), .Y(mai_mai_n356_));
  NA2        m334(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n357_));
  NA2        m335(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n358_));
  NA2        m336(.A(mai_mai_n235_), .B(x03), .Y(mai_mai_n359_));
  OAI220     m337(.A0(mai_mai_n359_), .A1(mai_mai_n358_), .B0(mai_mai_n357_), .B1(mai_mai_n80_), .Y(mai_mai_n360_));
  OAI210     m338(.A0(mai_mai_n26_), .A1(mai_mai_n100_), .B0(x07), .Y(mai_mai_n361_));
  AOI210     m339(.A0(mai_mai_n360_), .A1(x06), .B0(mai_mai_n361_), .Y(mai_mai_n362_));
  AOI220     m340(.A0(mai_mai_n80_), .A1(mai_mai_n31_), .B0(mai_mai_n52_), .B1(mai_mai_n51_), .Y(mai_mai_n363_));
  NO3        m341(.A(mai_mai_n363_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n364_));
  NO2        m342(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n365_));
  OAI210     m343(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n366_));
  OR3        m344(.A(mai_mai_n366_), .B(mai_mai_n365_), .C(mai_mai_n44_), .Y(mai_mai_n367_));
  INV        m345(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  OAI210     m346(.A0(mai_mai_n368_), .A1(mai_mai_n364_), .B0(mai_mai_n100_), .Y(mai_mai_n369_));
  NA2        m347(.A(mai_mai_n33_), .B(mai_mai_n100_), .Y(mai_mai_n370_));
  AOI210     m348(.A0(mai_mai_n370_), .A1(mai_mai_n91_), .B0(x07), .Y(mai_mai_n371_));
  AOI220     m349(.A0(mai_mai_n371_), .A1(mai_mai_n369_), .B0(mai_mai_n362_), .B1(mai_mai_n356_), .Y(mai_mai_n372_));
  AOI210     m350(.A0(mai_mai_n365_), .A1(mai_mai_n74_), .B0(mai_mai_n129_), .Y(mai_mai_n373_));
  OR2        m351(.A(mai_mai_n373_), .B(x03), .Y(mai_mai_n374_));
  NA2        m352(.A(mai_mai_n325_), .B(mai_mai_n61_), .Y(mai_mai_n375_));
  NO2        m353(.A(mai_mai_n375_), .B(x11), .Y(mai_mai_n376_));
  NO3        m354(.A(mai_mai_n376_), .B(mai_mai_n133_), .C(mai_mai_n28_), .Y(mai_mai_n377_));
  AOI210     m355(.A0(mai_mai_n377_), .A1(mai_mai_n374_), .B0(mai_mai_n47_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n378_), .B(mai_mai_n101_), .Y(mai_mai_n379_));
  AOI210     m357(.A0(mai_mai_n314_), .A1(mai_mai_n107_), .B0(mai_mai_n243_), .Y(mai_mai_n380_));
  NOi21      m358(.An(mai_mai_n298_), .B(mai_mai_n122_), .Y(mai_mai_n381_));
  NO2        m359(.A(mai_mai_n381_), .B(mai_mai_n244_), .Y(mai_mai_n382_));
  OAI210     m360(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n383_));
  AOI210     m361(.A0(mai_mai_n230_), .A1(mai_mai_n47_), .B0(mai_mai_n383_), .Y(mai_mai_n384_));
  NO4        m362(.A(mai_mai_n384_), .B(mai_mai_n382_), .C(mai_mai_n380_), .D(x08), .Y(mai_mai_n385_));
  NO2        m363(.A(mai_mai_n121_), .B(mai_mai_n28_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n386_), .B(mai_mai_n248_), .Y(mai_mai_n387_));
  NA3        m365(.A(mai_mai_n308_), .B(mai_mai_n116_), .C(x12), .Y(mai_mai_n388_));
  AO210      m366(.A0(mai_mai_n308_), .A1(mai_mai_n116_), .B0(mai_mai_n230_), .Y(mai_mai_n389_));
  NA3        m367(.A(mai_mai_n389_), .B(mai_mai_n388_), .C(x08), .Y(mai_mai_n390_));
  INV        m368(.A(mai_mai_n390_), .Y(mai_mai_n391_));
  AOI210     m369(.A0(mai_mai_n385_), .A1(mai_mai_n379_), .B0(mai_mai_n391_), .Y(mai_mai_n392_));
  OAI210     m370(.A0(mai_mai_n375_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n393_));
  NA2        m371(.A(mai_mai_n272_), .B(x07), .Y(mai_mai_n394_));
  OAI220     m372(.A0(mai_mai_n394_), .A1(mai_mai_n358_), .B0(mai_mai_n133_), .B1(mai_mai_n43_), .Y(mai_mai_n395_));
  OAI210     m373(.A0(mai_mai_n395_), .A1(mai_mai_n393_), .B0(mai_mai_n175_), .Y(mai_mai_n396_));
  NA3        m374(.A(mai_mai_n387_), .B(mai_mai_n381_), .C(mai_mai_n304_), .Y(mai_mai_n397_));
  INV        m375(.A(x14), .Y(mai_mai_n398_));
  NO3        m376(.A(mai_mai_n298_), .B(mai_mai_n103_), .C(x11), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n399_), .B(mai_mai_n398_), .Y(mai_mai_n400_));
  NA3        m378(.A(mai_mai_n400_), .B(mai_mai_n397_), .C(mai_mai_n396_), .Y(mai_mai_n401_));
  AOI220     m379(.A0(mai_mai_n370_), .A1(mai_mai_n61_), .B0(mai_mai_n386_), .B1(mai_mai_n151_), .Y(mai_mai_n402_));
  NOi21      m380(.An(mai_mai_n253_), .B(mai_mai_n137_), .Y(mai_mai_n403_));
  NO3        m381(.A(mai_mai_n118_), .B(mai_mai_n24_), .C(x06), .Y(mai_mai_n404_));
  AOI210     m382(.A0(mai_mai_n259_), .A1(mai_mai_n213_), .B0(mai_mai_n404_), .Y(mai_mai_n405_));
  OAI210     m383(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n405_), .Y(mai_mai_n406_));
  OAI210     m384(.A0(mai_mai_n406_), .A1(mai_mai_n403_), .B0(mai_mai_n100_), .Y(mai_mai_n407_));
  OAI210     m385(.A0(mai_mai_n402_), .A1(mai_mai_n90_), .B0(mai_mai_n407_), .Y(mai_mai_n408_));
  NO4        m386(.A(mai_mai_n408_), .B(mai_mai_n401_), .C(mai_mai_n392_), .D(mai_mai_n372_), .Y(mai06));
  INV        m387(.A(x13), .Y(mai_mai_n412_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI220     u039(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n61_), .Y(men_men_n62_));
  INV        u040(.A(men_men_n59_), .Y(men_men_n63_));
  OAI220     u041(.A0(x02), .A1(men_men_n63_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n64_));
  NA2        u042(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n65_));
  OAI210     u043(.A0(men_men_n30_), .A1(x11), .B0(men_men_n65_), .Y(men_men_n66_));
  AOI220     u044(.A0(men_men_n66_), .A1(men_men_n59_), .B0(men_men_n64_), .B1(men_men_n31_), .Y(men_men_n67_));
  AOI210     u045(.A0(men_men_n67_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n68_));
  NA2        u046(.A(x10), .B(x09), .Y(men_men_n69_));
  NA2        u047(.A(x09), .B(x05), .Y(men_men_n70_));
  NA2        u048(.A(x10), .B(x06), .Y(men_men_n71_));
  NO2        u049(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n72_));
  OAI210     u050(.A0(x02), .A1(x07), .B0(x03), .Y(men_men_n73_));
  NOi31      u051(.An(x08), .B(x04), .C(x00), .Y(men_men_n74_));
  NO2        u052(.A(x10), .B(x09), .Y(men_men_n75_));
  AOI210     u053(.A0(men_men_n459_), .A1(men_men_n74_), .B0(men_men_n24_), .Y(men_men_n76_));
  NO2        u054(.A(x09), .B(men_men_n41_), .Y(men_men_n77_));
  NO2        u055(.A(men_men_n77_), .B(men_men_n36_), .Y(men_men_n78_));
  OAI210     u056(.A0(men_men_n77_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n79_));
  AOI210     u057(.A0(men_men_n78_), .A1(men_men_n48_), .B0(men_men_n79_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n36_), .B(x00), .Y(men_men_n81_));
  NO2        u059(.A(x08), .B(x01), .Y(men_men_n82_));
  OAI210     u060(.A0(men_men_n82_), .A1(men_men_n81_), .B0(men_men_n35_), .Y(men_men_n83_));
  NO3        u061(.A(men_men_n83_), .B(men_men_n80_), .C(men_men_n76_), .Y(men_men_n84_));
  AN2        u062(.A(men_men_n84_), .B(men_men_n73_), .Y(men_men_n85_));
  INV        u063(.A(men_men_n83_), .Y(men_men_n86_));
  NO2        u064(.A(x06), .B(x05), .Y(men_men_n87_));
  NA2        u065(.A(x11), .B(x00), .Y(men_men_n88_));
  NO2        u066(.A(x11), .B(men_men_n47_), .Y(men_men_n89_));
  NOi21      u067(.An(men_men_n88_), .B(men_men_n89_), .Y(men_men_n90_));
  AOI210     u068(.A0(men_men_n87_), .A1(men_men_n86_), .B0(men_men_n90_), .Y(men_men_n91_));
  NOi21      u069(.An(x01), .B(x10), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n93_));
  NO3        u071(.A(men_men_n93_), .B(men_men_n92_), .C(x06), .Y(men_men_n94_));
  NA2        u072(.A(men_men_n94_), .B(men_men_n27_), .Y(men_men_n95_));
  OAI210     u073(.A0(men_men_n91_), .A1(x07), .B0(men_men_n95_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n85_), .C(men_men_n68_), .Y(men01));
  INV        u075(.A(x12), .Y(men_men_n98_));
  INV        u076(.A(x13), .Y(men_men_n99_));
  NA2        u077(.A(x08), .B(x04), .Y(men_men_n100_));
  NO2        u078(.A(men_men_n100_), .B(men_men_n57_), .Y(men_men_n101_));
  NA2        u079(.A(men_men_n101_), .B(men_men_n87_), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n92_), .B(men_men_n28_), .Y(men_men_n103_));
  NO2        u081(.A(x10), .B(x01), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n29_), .B(x00), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n105_), .B(men_men_n104_), .Y(men_men_n106_));
  NA2        u084(.A(x04), .B(men_men_n28_), .Y(men_men_n107_));
  NO3        u085(.A(men_men_n107_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n108_));
  NA2        u086(.A(men_men_n108_), .B(men_men_n106_), .Y(men_men_n109_));
  AOI210     u087(.A0(men_men_n109_), .A1(men_men_n102_), .B0(men_men_n99_), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n56_), .B(x05), .Y(men_men_n111_));
  NOi21      u089(.An(men_men_n111_), .B(men_men_n58_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n35_), .B(x02), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n99_), .B(men_men_n36_), .Y(men_men_n114_));
  NA3        u092(.A(men_men_n114_), .B(men_men_n113_), .C(x06), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n115_), .B(men_men_n112_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n82_), .B(x13), .Y(men_men_n117_));
  NA2        u095(.A(x09), .B(men_men_n35_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NA2        u097(.A(x13), .B(men_men_n35_), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(x05), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(men_men_n119_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n123_), .B(men_men_n99_), .Y(men_men_n124_));
  AOI210     u102(.A0(men_men_n124_), .A1(men_men_n78_), .B0(men_men_n112_), .Y(men_men_n125_));
  AOI210     u103(.A0(men_men_n125_), .A1(men_men_n122_), .B0(men_men_n71_), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n127_));
  NA2        u105(.A(x10), .B(men_men_n57_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n51_), .B(x05), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n36_), .B(x04), .Y(men_men_n131_));
  NA3        u109(.A(men_men_n131_), .B(men_men_n130_), .C(x13), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n123_), .B(men_men_n77_), .C(men_men_n36_), .Y(men_men_n133_));
  NO2        u111(.A(men_men_n60_), .B(x05), .Y(men_men_n134_));
  NOi41      u112(.An(men_men_n132_), .B(men_men_n134_), .C(men_men_n133_), .D(men_men_n129_), .Y(men_men_n135_));
  NO3        u113(.A(men_men_n135_), .B(x06), .C(x03), .Y(men_men_n136_));
  NO4        u114(.A(men_men_n136_), .B(men_men_n126_), .C(men_men_n116_), .D(men_men_n110_), .Y(men_men_n137_));
  NA2        u115(.A(x13), .B(men_men_n36_), .Y(men_men_n138_));
  OAI210     u116(.A0(men_men_n82_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  OA210      u118(.A0(men_men_n87_), .A1(men_men_n75_), .B0(x04), .Y(men_men_n141_));
  NO2        u119(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n142_));
  NA2        u120(.A(men_men_n29_), .B(x06), .Y(men_men_n143_));
  AOI210     u121(.A0(men_men_n143_), .A1(men_men_n49_), .B0(men_men_n142_), .Y(men_men_n144_));
  OA210      u122(.A0(men_men_n144_), .A1(men_men_n141_), .B0(men_men_n140_), .Y(men_men_n145_));
  NO2        u123(.A(x09), .B(x05), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n146_), .B(men_men_n47_), .Y(men_men_n147_));
  AOI210     u125(.A0(men_men_n147_), .A1(men_men_n106_), .B0(men_men_n49_), .Y(men_men_n148_));
  NA2        u126(.A(x09), .B(x00), .Y(men_men_n149_));
  NA2        u127(.A(men_men_n111_), .B(men_men_n149_), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n74_), .B(men_men_n51_), .Y(men_men_n151_));
  AOI210     u129(.A0(men_men_n151_), .A1(men_men_n150_), .B0(men_men_n143_), .Y(men_men_n152_));
  NO3        u130(.A(men_men_n152_), .B(men_men_n148_), .C(men_men_n145_), .Y(men_men_n153_));
  NO2        u131(.A(x03), .B(x02), .Y(men_men_n154_));
  NA2        u132(.A(men_men_n83_), .B(men_men_n99_), .Y(men_men_n155_));
  OAI210     u133(.A0(men_men_n155_), .A1(men_men_n112_), .B0(men_men_n154_), .Y(men_men_n156_));
  OA210      u134(.A0(men_men_n153_), .A1(x11), .B0(men_men_n156_), .Y(men_men_n157_));
  OAI210     u135(.A0(men_men_n137_), .A1(men_men_n23_), .B0(men_men_n157_), .Y(men_men_n158_));
  NA2        u136(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n159_));
  NAi21      u137(.An(x06), .B(x10), .Y(men_men_n160_));
  NOi21      u138(.An(x01), .B(x13), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  OR2        u140(.A(men_men_n162_), .B(men_men_n159_), .Y(men_men_n163_));
  NO2        u141(.A(men_men_n163_), .B(men_men_n41_), .Y(men_men_n164_));
  NO2        u142(.A(men_men_n29_), .B(x03), .Y(men_men_n165_));
  NA2        u143(.A(men_men_n99_), .B(x01), .Y(men_men_n166_));
  NO2        u144(.A(men_men_n166_), .B(x08), .Y(men_men_n167_));
  OAI210     u145(.A0(x05), .A1(men_men_n167_), .B0(men_men_n51_), .Y(men_men_n168_));
  AOI210     u146(.A0(men_men_n168_), .A1(men_men_n165_), .B0(men_men_n48_), .Y(men_men_n169_));
  AOI210     u147(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n170_));
  OAI210     u148(.A0(men_men_n169_), .A1(men_men_n164_), .B0(men_men_n170_), .Y(men_men_n171_));
  NA2        u149(.A(x04), .B(x02), .Y(men_men_n172_));
  NA2        u150(.A(x10), .B(x05), .Y(men_men_n173_));
  NA2        u151(.A(x09), .B(x06), .Y(men_men_n174_));
  AOI210     u152(.A0(men_men_n174_), .A1(men_men_n173_), .B0(men_men_n159_), .Y(men_men_n175_));
  NO2        u153(.A(x09), .B(x01), .Y(men_men_n176_));
  NO3        u154(.A(men_men_n176_), .B(men_men_n104_), .C(men_men_n31_), .Y(men_men_n177_));
  OAI210     u155(.A0(men_men_n177_), .A1(men_men_n175_), .B0(x00), .Y(men_men_n178_));
  NO2        u156(.A(men_men_n111_), .B(x08), .Y(men_men_n179_));
  NA3        u157(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n51_), .Y(men_men_n180_));
  NA2        u158(.A(men_men_n92_), .B(x05), .Y(men_men_n181_));
  OAI210     u159(.A0(men_men_n181_), .A1(men_men_n114_), .B0(men_men_n180_), .Y(men_men_n182_));
  AOI210     u160(.A0(men_men_n179_), .A1(x06), .B0(men_men_n182_), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n183_), .A1(x11), .B0(men_men_n178_), .Y(men_men_n184_));
  NAi21      u162(.An(men_men_n172_), .B(men_men_n184_), .Y(men_men_n185_));
  INV        u163(.A(men_men_n25_), .Y(men_men_n186_));
  NAi21      u164(.An(x13), .B(x00), .Y(men_men_n187_));
  AOI210     u165(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n187_), .Y(men_men_n188_));
  AOI220     u166(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n173_), .A1(men_men_n35_), .B0(men_men_n189_), .Y(men_men_n190_));
  AN2        u168(.A(men_men_n190_), .B(men_men_n188_), .Y(men_men_n191_));
  AN2        u169(.A(men_men_n71_), .B(men_men_n70_), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n93_), .B(x06), .Y(men_men_n193_));
  NO2        u171(.A(men_men_n187_), .B(men_men_n36_), .Y(men_men_n194_));
  INV        u172(.A(men_men_n194_), .Y(men_men_n195_));
  OAI220     u173(.A0(men_men_n195_), .A1(men_men_n174_), .B0(men_men_n193_), .B1(men_men_n192_), .Y(men_men_n196_));
  OAI210     u174(.A0(men_men_n196_), .A1(men_men_n191_), .B0(men_men_n186_), .Y(men_men_n197_));
  NOi21      u175(.An(x09), .B(x00), .Y(men_men_n198_));
  NO3        u176(.A(men_men_n81_), .B(men_men_n198_), .C(men_men_n47_), .Y(men_men_n199_));
  NA2        u177(.A(men_men_n199_), .B(men_men_n128_), .Y(men_men_n200_));
  NA2        u178(.A(x10), .B(x08), .Y(men_men_n201_));
  INV        u179(.A(men_men_n201_), .Y(men_men_n202_));
  NA2        u180(.A(x06), .B(x05), .Y(men_men_n203_));
  OAI210     u181(.A0(men_men_n203_), .A1(men_men_n35_), .B0(men_men_n98_), .Y(men_men_n204_));
  AOI210     u182(.A0(men_men_n202_), .A1(men_men_n58_), .B0(men_men_n204_), .Y(men_men_n205_));
  NA2        u183(.A(men_men_n205_), .B(men_men_n200_), .Y(men_men_n206_));
  NO2        u184(.A(men_men_n99_), .B(x12), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n207_), .Y(men_men_n208_));
  NA2        u186(.A(men_men_n92_), .B(men_men_n51_), .Y(men_men_n209_));
  NO2        u187(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n210_));
  NA2        u188(.A(men_men_n210_), .B(x02), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n211_), .B(men_men_n209_), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n208_), .A1(men_men_n206_), .B0(men_men_n212_), .Y(men_men_n213_));
  NA4        u191(.A(men_men_n213_), .B(men_men_n197_), .C(men_men_n185_), .D(men_men_n171_), .Y(men_men_n214_));
  AOI210     u192(.A0(men_men_n158_), .A1(men_men_n98_), .B0(men_men_n214_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n28_), .B(men_men_n140_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n139_), .Y(men_men_n218_));
  AOI210     u196(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n127_), .B(x06), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n219_), .A1(men_men_n218_), .B0(men_men_n220_), .Y(men_men_n221_));
  AOI210     u199(.A0(men_men_n221_), .A1(men_men_n216_), .B0(x12), .Y(men_men_n222_));
  INV        u200(.A(men_men_n74_), .Y(men_men_n223_));
  AOI210     u201(.A0(men_men_n201_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n224_), .A1(men_men_n162_), .B0(men_men_n57_), .Y(men_men_n225_));
  NA2        u203(.A(men_men_n225_), .B(men_men_n223_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n92_), .B(x06), .Y(men_men_n227_));
  AOI210     u205(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n228_));
  NO3        u206(.A(men_men_n228_), .B(men_men_n227_), .C(men_men_n41_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n56_), .A1(men_men_n229_), .B0(x02), .Y(men_men_n230_));
  AOI210     u208(.A0(men_men_n230_), .A1(men_men_n226_), .B0(men_men_n23_), .Y(men_men_n231_));
  OAI210     u209(.A0(men_men_n222_), .A1(men_men_n57_), .B0(men_men_n231_), .Y(men_men_n232_));
  INV        u210(.A(men_men_n143_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n51_), .B(x03), .Y(men_men_n234_));
  OAI210     u212(.A0(men_men_n77_), .A1(men_men_n36_), .B0(men_men_n118_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n99_), .B(x03), .Y(men_men_n236_));
  AOI220     u214(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n74_), .B1(men_men_n234_), .Y(men_men_n237_));
  NA2        u215(.A(men_men_n32_), .B(x06), .Y(men_men_n238_));
  INV        u216(.A(men_men_n160_), .Y(men_men_n239_));
  NOi21      u217(.An(x13), .B(x04), .Y(men_men_n240_));
  NO3        u218(.A(men_men_n240_), .B(men_men_n74_), .C(men_men_n198_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n241_), .B(x05), .Y(men_men_n242_));
  AOI220     u220(.A0(men_men_n242_), .A1(men_men_n238_), .B0(men_men_n239_), .B1(men_men_n57_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n237_), .A1(men_men_n233_), .B0(men_men_n243_), .Y(men_men_n244_));
  INV        u222(.A(men_men_n89_), .Y(men_men_n245_));
  NO2        u223(.A(men_men_n245_), .B(x12), .Y(men_men_n246_));
  NA2        u224(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n248_));
  OAI210     u226(.A0(men_men_n248_), .A1(men_men_n190_), .B0(men_men_n188_), .Y(men_men_n249_));
  AOI210     u227(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n250_));
  NO2        u228(.A(x06), .B(x00), .Y(men_men_n251_));
  NO3        u229(.A(men_men_n251_), .B(men_men_n250_), .C(men_men_n41_), .Y(men_men_n252_));
  OAI210     u230(.A0(men_men_n100_), .A1(men_men_n149_), .B0(men_men_n71_), .Y(men_men_n253_));
  NO2        u231(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n255_), .B(x03), .Y(men_men_n256_));
  OA210      u234(.A0(men_men_n256_), .A1(men_men_n254_), .B0(men_men_n249_), .Y(men_men_n257_));
  NA2        u235(.A(x13), .B(men_men_n98_), .Y(men_men_n258_));
  NA3        u236(.A(men_men_n258_), .B(men_men_n204_), .C(men_men_n90_), .Y(men_men_n259_));
  OAI210     u237(.A0(men_men_n257_), .A1(men_men_n247_), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n246_), .A1(men_men_n244_), .B0(men_men_n260_), .Y(men_men_n261_));
  AOI210     u239(.A0(men_men_n261_), .A1(men_men_n232_), .B0(x07), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n70_), .B(men_men_n29_), .Y(men_men_n263_));
  NOi31      u241(.An(men_men_n138_), .B(men_men_n240_), .C(men_men_n198_), .Y(men_men_n264_));
  AOI210     u242(.A0(men_men_n264_), .A1(men_men_n151_), .B0(men_men_n263_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n99_), .B(x06), .Y(men_men_n266_));
  INV        u244(.A(men_men_n266_), .Y(men_men_n267_));
  NO2        u245(.A(x08), .B(x05), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n268_), .B(men_men_n250_), .Y(men_men_n269_));
  OAI210     u247(.A0(men_men_n74_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n269_), .A1(men_men_n267_), .B0(men_men_n270_), .Y(men_men_n271_));
  NO2        u249(.A(x12), .B(x02), .Y(men_men_n272_));
  INV        u250(.A(men_men_n272_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n273_), .B(men_men_n245_), .Y(men_men_n274_));
  OA210      u252(.A0(men_men_n271_), .A1(men_men_n265_), .B0(men_men_n274_), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n276_), .B(x01), .Y(men_men_n277_));
  NOi21      u255(.An(men_men_n82_), .B(men_men_n118_), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n278_), .B(men_men_n277_), .Y(men_men_n279_));
  AOI210     u257(.A0(men_men_n279_), .A1(men_men_n132_), .B0(men_men_n29_), .Y(men_men_n280_));
  NA2        u258(.A(men_men_n266_), .B(men_men_n235_), .Y(men_men_n281_));
  NA2        u259(.A(men_men_n99_), .B(x04), .Y(men_men_n282_));
  NA2        u260(.A(men_men_n282_), .B(men_men_n28_), .Y(men_men_n283_));
  OAI210     u261(.A0(men_men_n283_), .A1(men_men_n117_), .B0(men_men_n281_), .Y(men_men_n284_));
  NO3        u262(.A(men_men_n88_), .B(x12), .C(x03), .Y(men_men_n285_));
  OAI210     u263(.A0(men_men_n284_), .A1(men_men_n280_), .B0(men_men_n285_), .Y(men_men_n286_));
  AOI210     u264(.A0(men_men_n209_), .A1(men_men_n203_), .B0(men_men_n100_), .Y(men_men_n287_));
  NOi21      u265(.An(men_men_n263_), .B(men_men_n227_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n25_), .B(x00), .Y(men_men_n289_));
  OAI210     u267(.A0(men_men_n288_), .A1(men_men_n287_), .B0(men_men_n289_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n58_), .B(x05), .Y(men_men_n291_));
  NO3        u269(.A(men_men_n291_), .B(men_men_n228_), .C(men_men_n193_), .Y(men_men_n292_));
  NO2        u270(.A(men_men_n247_), .B(men_men_n28_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n292_), .A1(men_men_n233_), .B0(men_men_n293_), .Y(men_men_n294_));
  NA3        u272(.A(men_men_n294_), .B(men_men_n290_), .C(men_men_n286_), .Y(men_men_n295_));
  NO3        u273(.A(men_men_n295_), .B(men_men_n275_), .C(men_men_n262_), .Y(men_men_n296_));
  OAI210     u274(.A0(men_men_n215_), .A1(men_men_n61_), .B0(men_men_n296_), .Y(men02));
  AOI210     u275(.A0(men_men_n138_), .A1(men_men_n83_), .B0(men_men_n130_), .Y(men_men_n298_));
  NO2        u276(.A(men_men_n99_), .B(men_men_n35_), .Y(men_men_n299_));
  NA3        u277(.A(men_men_n299_), .B(men_men_n202_), .C(men_men_n56_), .Y(men_men_n300_));
  OAI210     u278(.A0(men_men_n241_), .A1(men_men_n32_), .B0(men_men_n300_), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n301_), .A1(men_men_n298_), .B0(men_men_n173_), .Y(men_men_n302_));
  INV        u280(.A(men_men_n173_), .Y(men_men_n303_));
  NO2        u281(.A(men_men_n113_), .B(men_men_n228_), .Y(men_men_n304_));
  OAI220     u282(.A0(men_men_n304_), .A1(men_men_n99_), .B0(men_men_n83_), .B1(men_men_n51_), .Y(men_men_n305_));
  AOI220     u283(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n155_), .B1(men_men_n154_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n306_), .A1(men_men_n302_), .B0(men_men_n48_), .Y(men_men_n307_));
  NO2        u285(.A(x05), .B(x02), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n218_), .A1(men_men_n198_), .B0(men_men_n308_), .Y(men_men_n309_));
  AOI220     u287(.A0(men_men_n268_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n310_));
  NOi21      u288(.An(men_men_n299_), .B(men_men_n310_), .Y(men_men_n311_));
  AOI210     u289(.A0(men_men_n240_), .A1(men_men_n77_), .B0(men_men_n311_), .Y(men_men_n312_));
  AOI210     u290(.A0(men_men_n312_), .A1(men_men_n309_), .B0(men_men_n143_), .Y(men_men_n313_));
  NAi21      u291(.An(men_men_n242_), .B(men_men_n237_), .Y(men_men_n314_));
  NO2        u292(.A(men_men_n255_), .B(men_men_n47_), .Y(men_men_n315_));
  NA2        u293(.A(men_men_n315_), .B(men_men_n314_), .Y(men_men_n316_));
  AN2        u294(.A(men_men_n236_), .B(men_men_n235_), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n318_));
  NA2        u296(.A(x13), .B(men_men_n28_), .Y(men_men_n319_));
  AOI210     u297(.A0(men_men_n319_), .A1(men_men_n139_), .B0(men_men_n318_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n320_), .A1(men_men_n317_), .B0(men_men_n93_), .Y(men_men_n321_));
  NA3        u299(.A(men_men_n93_), .B(men_men_n82_), .C(men_men_n234_), .Y(men_men_n322_));
  NA3        u300(.A(men_men_n92_), .B(men_men_n81_), .C(men_men_n42_), .Y(men_men_n323_));
  AOI210     u301(.A0(men_men_n323_), .A1(men_men_n322_), .B0(x04), .Y(men_men_n324_));
  NO2        u302(.A(men_men_n269_), .B(men_men_n103_), .Y(men_men_n325_));
  AOI210     u303(.A0(men_men_n325_), .A1(x13), .B0(men_men_n324_), .Y(men_men_n326_));
  NA3        u304(.A(men_men_n326_), .B(men_men_n321_), .C(men_men_n316_), .Y(men_men_n327_));
  NO3        u305(.A(men_men_n327_), .B(men_men_n313_), .C(men_men_n307_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n142_), .B(x03), .Y(men_men_n329_));
  INV        u307(.A(men_men_n187_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n331_));
  AOI220     u309(.A0(men_men_n331_), .A1(men_men_n330_), .B0(men_men_n210_), .B1(x08), .Y(men_men_n332_));
  OAI210     u310(.A0(men_men_n332_), .A1(men_men_n291_), .B0(men_men_n329_), .Y(men_men_n333_));
  NA2        u311(.A(men_men_n333_), .B(men_men_n104_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n56_), .A1(men_men_n179_), .B0(men_men_n105_), .Y(men_men_n335_));
  NA2        u313(.A(men_men_n282_), .B(men_men_n98_), .Y(men_men_n336_));
  NA2        u314(.A(men_men_n98_), .B(men_men_n41_), .Y(men_men_n337_));
  NA3        u315(.A(men_men_n337_), .B(men_men_n336_), .C(men_men_n129_), .Y(men_men_n338_));
  NA4        u316(.A(men_men_n338_), .B(men_men_n335_), .C(men_men_n334_), .D(men_men_n48_), .Y(men_men_n339_));
  INV        u317(.A(men_men_n210_), .Y(men_men_n340_));
  NO2        u318(.A(men_men_n167_), .B(men_men_n40_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n32_), .B(x05), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  NA2        u321(.A(men_men_n343_), .B(x02), .Y(men_men_n344_));
  INV        u322(.A(men_men_n248_), .Y(men_men_n345_));
  NA2        u323(.A(men_men_n207_), .B(x04), .Y(men_men_n346_));
  NO2        u324(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  NO3        u325(.A(men_men_n189_), .B(x13), .C(men_men_n31_), .Y(men_men_n348_));
  OAI210     u326(.A0(men_men_n348_), .A1(men_men_n347_), .B0(men_men_n93_), .Y(men_men_n349_));
  NO3        u327(.A(men_men_n207_), .B(men_men_n165_), .C(men_men_n52_), .Y(men_men_n350_));
  OAI210     u328(.A0(men_men_n149_), .A1(men_men_n36_), .B0(men_men_n98_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n351_), .A1(men_men_n199_), .B0(men_men_n350_), .Y(men_men_n352_));
  NA4        u330(.A(men_men_n352_), .B(men_men_n349_), .C(men_men_n344_), .D(x06), .Y(men_men_n353_));
  OAI220     u331(.A0(men_men_n166_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n354_));
  NO3        u332(.A(men_men_n291_), .B(men_men_n127_), .C(x08), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n354_), .A1(men_men_n233_), .B0(men_men_n355_), .Y(men_men_n356_));
  NO2        u334(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n357_));
  NO3        u335(.A(men_men_n111_), .B(men_men_n128_), .C(men_men_n38_), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n350_), .A1(men_men_n357_), .B0(men_men_n358_), .Y(men_men_n359_));
  OAI210     u337(.A0(men_men_n356_), .A1(men_men_n28_), .B0(men_men_n359_), .Y(men_men_n360_));
  AN2        u338(.A(men_men_n360_), .B(x04), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n353_), .A1(men_men_n339_), .B0(men_men_n361_), .Y(men_men_n362_));
  OAI210     u340(.A0(men_men_n328_), .A1(x12), .B0(men_men_n362_), .Y(men03));
  OR2        u341(.A(men_men_n42_), .B(men_men_n234_), .Y(men_men_n364_));
  AOI210     u342(.A0(men_men_n155_), .A1(men_men_n98_), .B0(men_men_n364_), .Y(men_men_n365_));
  NA2        u343(.A(men_men_n207_), .B(men_men_n154_), .Y(men_men_n366_));
  NA2        u344(.A(men_men_n366_), .B(men_men_n211_), .Y(men_men_n367_));
  OAI210     u345(.A0(men_men_n367_), .A1(men_men_n365_), .B0(x05), .Y(men_men_n368_));
  NA2        u346(.A(men_men_n364_), .B(x05), .Y(men_men_n369_));
  AOI210     u347(.A0(men_men_n139_), .A1(men_men_n223_), .B0(men_men_n369_), .Y(men_men_n370_));
  AOI210     u348(.A0(men_men_n236_), .A1(men_men_n78_), .B0(men_men_n121_), .Y(men_men_n371_));
  OAI220     u349(.A0(men_men_n371_), .A1(men_men_n59_), .B0(men_men_n319_), .B1(men_men_n310_), .Y(men_men_n372_));
  OAI210     u350(.A0(men_men_n372_), .A1(men_men_n370_), .B0(men_men_n98_), .Y(men_men_n373_));
  AOI210     u351(.A0(men_men_n147_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n374_));
  NO2        u352(.A(men_men_n176_), .B(men_men_n134_), .Y(men_men_n375_));
  OAI220     u353(.A0(men_men_n375_), .A1(men_men_n37_), .B0(men_men_n150_), .B1(x13), .Y(men_men_n376_));
  OAI210     u354(.A0(men_men_n376_), .A1(men_men_n374_), .B0(x04), .Y(men_men_n377_));
  NO3        u355(.A(men_men_n337_), .B(men_men_n83_), .C(men_men_n59_), .Y(men_men_n378_));
  AOI210     u356(.A0(men_men_n195_), .A1(men_men_n98_), .B0(men_men_n147_), .Y(men_men_n379_));
  OA210      u357(.A0(men_men_n167_), .A1(x12), .B0(men_men_n134_), .Y(men_men_n380_));
  NO3        u358(.A(men_men_n380_), .B(men_men_n379_), .C(men_men_n378_), .Y(men_men_n381_));
  NA4        u359(.A(men_men_n381_), .B(men_men_n377_), .C(men_men_n373_), .D(men_men_n368_), .Y(men04));
  NO2        u360(.A(men_men_n86_), .B(men_men_n39_), .Y(men_men_n383_));
  XO2        u361(.A(men_men_n383_), .B(men_men_n258_), .Y(men05));
  AOI210     u362(.A0(men_men_n70_), .A1(men_men_n52_), .B0(men_men_n220_), .Y(men_men_n385_));
  AOI210     u363(.A0(men_men_n385_), .A1(men_men_n318_), .B0(men_men_n25_), .Y(men_men_n386_));
  NAi41      u364(.An(men_men_n75_), .B(men_men_n143_), .C(men_men_n130_), .D(men_men_n31_), .Y(men_men_n387_));
  AOI210     u365(.A0(men_men_n239_), .A1(men_men_n57_), .B0(men_men_n87_), .Y(men_men_n388_));
  AOI210     u366(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n24_), .Y(men_men_n389_));
  OAI210     u367(.A0(men_men_n389_), .A1(men_men_n386_), .B0(men_men_n98_), .Y(men_men_n390_));
  NA2        u368(.A(x11), .B(men_men_n31_), .Y(men_men_n391_));
  NA2        u369(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n392_));
  NA2        u370(.A(men_men_n263_), .B(x03), .Y(men_men_n393_));
  OAI220     u371(.A0(men_men_n393_), .A1(men_men_n392_), .B0(men_men_n391_), .B1(men_men_n79_), .Y(men_men_n394_));
  OAI210     u372(.A0(men_men_n26_), .A1(men_men_n98_), .B0(x07), .Y(men_men_n395_));
  AOI210     u373(.A0(men_men_n394_), .A1(x06), .B0(men_men_n395_), .Y(men_men_n396_));
  AOI220     u374(.A0(men_men_n79_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n397_));
  NO3        u375(.A(men_men_n397_), .B(men_men_n23_), .C(x00), .Y(men_men_n398_));
  NA2        u376(.A(men_men_n69_), .B(x02), .Y(men_men_n399_));
  AOI210     u377(.A0(men_men_n399_), .A1(men_men_n393_), .B0(men_men_n266_), .Y(men_men_n400_));
  OR2        u378(.A(men_men_n400_), .B(men_men_n247_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n161_), .B(x05), .Y(men_men_n402_));
  NA3        u380(.A(men_men_n402_), .B(men_men_n251_), .C(men_men_n245_), .Y(men_men_n403_));
  NO2        u381(.A(men_men_n23_), .B(x10), .Y(men_men_n404_));
  OAI210     u382(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n405_));
  OR3        u383(.A(men_men_n405_), .B(men_men_n404_), .C(men_men_n44_), .Y(men_men_n406_));
  NA3        u384(.A(men_men_n406_), .B(men_men_n403_), .C(men_men_n401_), .Y(men_men_n407_));
  OAI210     u385(.A0(men_men_n407_), .A1(men_men_n398_), .B0(men_men_n98_), .Y(men_men_n408_));
  NA2        u386(.A(men_men_n33_), .B(men_men_n98_), .Y(men_men_n409_));
  AOI210     u387(.A0(men_men_n409_), .A1(men_men_n89_), .B0(x07), .Y(men_men_n410_));
  AOI220     u388(.A0(men_men_n410_), .A1(men_men_n408_), .B0(men_men_n396_), .B1(men_men_n390_), .Y(men_men_n411_));
  NA3        u389(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n412_));
  AO210      u390(.A0(men_men_n412_), .A1(men_men_n276_), .B0(men_men_n273_), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n404_), .A1(men_men_n72_), .B0(men_men_n142_), .Y(men_men_n414_));
  OR2        u392(.A(men_men_n414_), .B(x03), .Y(men_men_n415_));
  NA2        u393(.A(men_men_n357_), .B(men_men_n61_), .Y(men_men_n416_));
  NO3        u394(.A(men_men_n357_), .B(men_men_n146_), .C(men_men_n28_), .Y(men_men_n417_));
  AOI220     u395(.A0(men_men_n417_), .A1(men_men_n415_), .B0(men_men_n413_), .B1(men_men_n47_), .Y(men_men_n418_));
  NO4        u396(.A(men_men_n337_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n419_));
  OAI210     u397(.A0(men_men_n419_), .A1(men_men_n418_), .B0(men_men_n99_), .Y(men_men_n420_));
  AOI210     u398(.A0(men_men_n346_), .A1(men_men_n107_), .B0(men_men_n272_), .Y(men_men_n421_));
  NOi21      u399(.An(men_men_n329_), .B(men_men_n134_), .Y(men_men_n422_));
  OAI210     u400(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n423_));
  AOI210     u401(.A0(men_men_n258_), .A1(men_men_n47_), .B0(men_men_n423_), .Y(men_men_n424_));
  NO3        u402(.A(men_men_n424_), .B(men_men_n421_), .C(x08), .Y(men_men_n425_));
  AOI210     u403(.A0(men_men_n404_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n426_));
  NA2        u404(.A(x09), .B(men_men_n41_), .Y(men_men_n427_));
  OAI210     u405(.A0(men_men_n427_), .A1(men_men_n426_), .B0(men_men_n391_), .Y(men_men_n428_));
  NO2        u406(.A(x13), .B(x12), .Y(men_men_n429_));
  NO2        u407(.A(men_men_n130_), .B(men_men_n28_), .Y(men_men_n430_));
  NO2        u408(.A(men_men_n430_), .B(men_men_n277_), .Y(men_men_n431_));
  OR3        u409(.A(men_men_n431_), .B(x12), .C(x03), .Y(men_men_n432_));
  NA3        u410(.A(men_men_n340_), .B(men_men_n123_), .C(x12), .Y(men_men_n433_));
  AO210      u411(.A0(men_men_n340_), .A1(men_men_n123_), .B0(men_men_n258_), .Y(men_men_n434_));
  NA4        u412(.A(men_men_n434_), .B(men_men_n433_), .C(men_men_n432_), .D(x08), .Y(men_men_n435_));
  AOI210     u413(.A0(men_men_n429_), .A1(men_men_n428_), .B0(men_men_n435_), .Y(men_men_n436_));
  AOI210     u414(.A0(men_men_n425_), .A1(men_men_n420_), .B0(men_men_n436_), .Y(men_men_n437_));
  OAI210     u415(.A0(men_men_n416_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n438_));
  NA2        u416(.A(men_men_n303_), .B(x07), .Y(men_men_n439_));
  OAI220     u417(.A0(men_men_n439_), .A1(men_men_n392_), .B0(men_men_n146_), .B1(men_men_n43_), .Y(men_men_n440_));
  OAI210     u418(.A0(men_men_n440_), .A1(men_men_n438_), .B0(men_men_n194_), .Y(men_men_n441_));
  NA3        u419(.A(men_men_n431_), .B(men_men_n422_), .C(men_men_n336_), .Y(men_men_n442_));
  INV        u420(.A(x14), .Y(men_men_n443_));
  NO3        u421(.A(men_men_n329_), .B(men_men_n103_), .C(x11), .Y(men_men_n444_));
  NO3        u422(.A(men_men_n166_), .B(men_men_n72_), .C(men_men_n57_), .Y(men_men_n445_));
  NO3        u423(.A(men_men_n412_), .B(men_men_n337_), .C(men_men_n187_), .Y(men_men_n446_));
  NO4        u424(.A(men_men_n446_), .B(men_men_n445_), .C(men_men_n444_), .D(men_men_n443_), .Y(men_men_n447_));
  NA3        u425(.A(men_men_n447_), .B(men_men_n442_), .C(men_men_n441_), .Y(men_men_n448_));
  AOI220     u426(.A0(men_men_n409_), .A1(men_men_n61_), .B0(men_men_n430_), .B1(men_men_n165_), .Y(men_men_n449_));
  NOi21      u427(.An(men_men_n282_), .B(men_men_n150_), .Y(men_men_n450_));
  NO3        u428(.A(men_men_n127_), .B(men_men_n24_), .C(x06), .Y(men_men_n451_));
  AOI210     u429(.A0(men_men_n289_), .A1(men_men_n239_), .B0(men_men_n451_), .Y(men_men_n452_));
  OAI210     u430(.A0(men_men_n44_), .A1(x04), .B0(men_men_n452_), .Y(men_men_n453_));
  OAI210     u431(.A0(men_men_n453_), .A1(men_men_n450_), .B0(men_men_n98_), .Y(men_men_n454_));
  OAI210     u432(.A0(men_men_n449_), .A1(men_men_n88_), .B0(men_men_n454_), .Y(men_men_n455_));
  NO4        u433(.A(men_men_n455_), .B(men_men_n448_), .C(men_men_n437_), .D(men_men_n411_), .Y(men06));
  INV        u434(.A(x07), .Y(men_men_n459_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule