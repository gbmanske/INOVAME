module sum(a,b,scanin,scan_en,c,scanout);
input a,b,scanin,scan_en;
output c,scanout;

assign c = a+b;
endmodule
