//Benchmark atmr_9sym_175_0.125

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n104_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n136_, ori00, mai00, men00;
  INV        o00(.A(i_3_), .Y(ori_ori_n11_));
  INV        o01(.A(i_6_), .Y(ori_ori_n12_));
  INV        o02(.A(i_5_), .Y(ori_ori_n13_));
  INV        o03(.A(i_0_), .Y(ori_ori_n14_));
  INV        o04(.A(i_4_), .Y(ori_ori_n15_));
  NA2        o05(.A(i_0_), .B(ori_ori_n15_), .Y(ori_ori_n16_));
  INV        o06(.A(i_7_), .Y(ori_ori_n17_));
  AOI210     o07(.A0(i_1_), .A1(i_2_), .B0(i_5_), .Y(ori_ori_n18_));
  NO2        o08(.A(ori_ori_n18_), .B(ori_ori_n16_), .Y(ori_ori_n19_));
  NA2        o09(.A(ori_ori_n19_), .B(ori_ori_n11_), .Y(ori_ori_n20_));
  NA2        o10(.A(ori_ori_n14_), .B(i_5_), .Y(ori_ori_n21_));
  NO2        o11(.A(i_2_), .B(i_4_), .Y(ori_ori_n22_));
  NA3        o12(.A(ori_ori_n22_), .B(i_6_), .C(i_8_), .Y(ori_ori_n23_));
  AOI210     o13(.A0(ori_ori_n21_), .A1(i_5_), .B0(ori_ori_n23_), .Y(ori_ori_n24_));
  INV        o14(.A(i_2_), .Y(ori_ori_n25_));
  NOi21      o15(.An(i_6_), .B(i_8_), .Y(ori_ori_n26_));
  NOi21      o16(.An(i_7_), .B(i_1_), .Y(ori_ori_n27_));
  NOi21      o17(.An(i_5_), .B(i_6_), .Y(ori_ori_n28_));
  NA2        o18(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n29_));
  NO3        o19(.A(ori_ori_n29_), .B(ori_ori_n25_), .C(i_4_), .Y(ori_ori_n30_));
  NOi21      o20(.An(i_0_), .B(i_4_), .Y(ori_ori_n31_));
  INV        o21(.A(i_1_), .Y(ori_ori_n32_));
  NOi21      o22(.An(i_3_), .B(i_0_), .Y(ori_ori_n33_));
  NO2        o23(.A(ori_ori_n30_), .B(ori_ori_n24_), .Y(ori_ori_n34_));
  NOi21      o24(.An(i_4_), .B(i_0_), .Y(ori_ori_n35_));
  INV        o25(.A(i_8_), .Y(ori_ori_n36_));
  INV        o26(.A(ori_ori_n31_), .Y(ori_ori_n37_));
  NO3        o27(.A(ori_ori_n37_), .B(i_5_), .C(ori_ori_n36_), .Y(ori_ori_n38_));
  INV        o28(.A(ori_ori_n38_), .Y(ori_ori_n39_));
  NOi21      o29(.An(i_2_), .B(i_1_), .Y(ori_ori_n40_));
  NOi21      o30(.An(i_4_), .B(i_3_), .Y(ori_ori_n41_));
  NOi21      o31(.An(i_1_), .B(i_4_), .Y(ori_ori_n42_));
  AN2        o32(.A(i_8_), .B(i_7_), .Y(ori_ori_n43_));
  NOi21      o33(.An(i_8_), .B(i_7_), .Y(ori_ori_n44_));
  NA2        o34(.A(ori_ori_n42_), .B(ori_ori_n28_), .Y(ori_ori_n45_));
  NA4        o35(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .D(ori_ori_n20_), .Y(ori_ori_n46_));
  NOi21      o36(.An(i_1_), .B(i_2_), .Y(ori_ori_n47_));
  NA3        o37(.A(ori_ori_n44_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n48_));
  NA2        o38(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n49_));
  NA2        o39(.A(ori_ori_n49_), .B(ori_ori_n48_), .Y(ori_ori_n50_));
  NA2        o40(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n51_));
  INV        o41(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  INV        o42(.A(i_6_), .Y(ori_ori_n53_));
  NOi21      o43(.An(i_7_), .B(i_8_), .Y(ori_ori_n54_));
  NO2        o44(.A(i_8_), .B(ori_ori_n11_), .Y(ori_ori_n55_));
  NA2        o45(.A(ori_ori_n55_), .B(ori_ori_n47_), .Y(ori_ori_n56_));
  NA2        o46(.A(ori_ori_n33_), .B(ori_ori_n32_), .Y(ori_ori_n57_));
  NA3        o47(.A(ori_ori_n15_), .B(i_5_), .C(i_7_), .Y(ori_ori_n58_));
  NO2        o48(.A(ori_ori_n58_), .B(ori_ori_n57_), .Y(ori_ori_n59_));
  INV        o49(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NA3        o50(.A(ori_ori_n44_), .B(ori_ori_n25_), .C(i_3_), .Y(ori_ori_n61_));
  NA2        o51(.A(ori_ori_n32_), .B(i_6_), .Y(ori_ori_n62_));
  INV        o52(.A(i_1_), .Y(ori_ori_n63_));
  INV        o53(.A(i_0_), .Y(ori_ori_n64_));
  NOi31      o54(.An(ori_ori_n35_), .B(ori_ori_n104_), .C(i_2_), .Y(ori_ori_n65_));
  NOi21      o55(.An(i_3_), .B(i_1_), .Y(ori_ori_n66_));
  NA2        o56(.A(ori_ori_n66_), .B(i_4_), .Y(ori_ori_n67_));
  NO2        o57(.A(i_8_), .B(ori_ori_n67_), .Y(ori_ori_n68_));
  NOi31      o58(.An(ori_ori_n33_), .B(i_5_), .C(ori_ori_n25_), .Y(ori_ori_n69_));
  NO3        o59(.A(ori_ori_n69_), .B(ori_ori_n68_), .C(ori_ori_n65_), .Y(ori_ori_n70_));
  NA3        o60(.A(ori_ori_n70_), .B(ori_ori_n60_), .C(ori_ori_n56_), .Y(ori_ori_n71_));
  NA2        o61(.A(ori_ori_n26_), .B(ori_ori_n31_), .Y(ori_ori_n72_));
  INV        o62(.A(ori_ori_n41_), .Y(ori_ori_n73_));
  AOI210     o63(.A0(ori_ori_n73_), .A1(ori_ori_n48_), .B0(ori_ori_n21_), .Y(ori_ori_n74_));
  NA3        o64(.A(ori_ori_n43_), .B(ori_ori_n63_), .C(ori_ori_n12_), .Y(ori_ori_n75_));
  NAi31      o65(.An(ori_ori_n64_), .B(ori_ori_n54_), .C(ori_ori_n63_), .Y(ori_ori_n76_));
  NA3        o66(.A(ori_ori_n44_), .B(ori_ori_n40_), .C(i_6_), .Y(ori_ori_n77_));
  NA3        o67(.A(ori_ori_n77_), .B(ori_ori_n76_), .C(ori_ori_n75_), .Y(ori_ori_n78_));
  NOi21      o68(.An(i_0_), .B(i_2_), .Y(ori_ori_n79_));
  NA2        o69(.A(ori_ori_n79_), .B(ori_ori_n27_), .Y(ori_ori_n80_));
  INV        o70(.A(ori_ori_n80_), .Y(ori_ori_n81_));
  NO3        o71(.A(ori_ori_n81_), .B(ori_ori_n78_), .C(ori_ori_n74_), .Y(ori_ori_n82_));
  INV        o72(.A(ori_ori_n54_), .Y(ori_ori_n83_));
  NO2        o73(.A(ori_ori_n83_), .B(ori_ori_n62_), .Y(ori_ori_n84_));
  NO3        o74(.A(i_2_), .B(ori_ori_n15_), .C(ori_ori_n13_), .Y(ori_ori_n85_));
  NA2        o75(.A(i_2_), .B(i_4_), .Y(ori_ori_n86_));
  AOI210     o76(.A0(ori_ori_n64_), .A1(ori_ori_n53_), .B0(ori_ori_n86_), .Y(ori_ori_n87_));
  NO2        o77(.A(i_8_), .B(i_7_), .Y(ori_ori_n88_));
  OA210      o78(.A0(ori_ori_n87_), .A1(ori_ori_n85_), .B0(ori_ori_n88_), .Y(ori_ori_n89_));
  NA3        o79(.A(ori_ori_n66_), .B(i_0_), .C(ori_ori_n17_), .Y(ori_ori_n90_));
  INV        o80(.A(ori_ori_n90_), .Y(ori_ori_n91_));
  NO3        o81(.A(ori_ori_n91_), .B(ori_ori_n89_), .C(ori_ori_n84_), .Y(ori_ori_n92_));
  NA2        o82(.A(ori_ori_n54_), .B(ori_ori_n12_), .Y(ori_ori_n93_));
  NA2        o83(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n94_));
  INV        o84(.A(ori_ori_n35_), .Y(ori_ori_n95_));
  AOI210     o85(.A0(ori_ori_n95_), .A1(ori_ori_n94_), .B0(ori_ori_n93_), .Y(ori_ori_n96_));
  NA2        o86(.A(ori_ori_n79_), .B(ori_ori_n44_), .Y(ori_ori_n97_));
  NA2        o87(.A(ori_ori_n61_), .B(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o88(.A(ori_ori_n98_), .B(ori_ori_n96_), .Y(ori_ori_n99_));
  NA4        o89(.A(ori_ori_n99_), .B(ori_ori_n92_), .C(ori_ori_n82_), .D(ori_ori_n72_), .Y(ori_ori_n100_));
  OR4        o90(.A(ori_ori_n100_), .B(ori_ori_n71_), .C(ori_ori_n52_), .D(ori_ori_n46_), .Y(ori00));
  INV        o91(.A(i_7_), .Y(ori_ori_n104_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  NA3        m006(.A(mai_mai_n16_), .B(mai_mai_n15_), .C(i_2_), .Y(mai_mai_n17_));
  NO2        m007(.A(mai_mai_n17_), .B(i_6_), .Y(mai_mai_n18_));
  INV        m008(.A(i_4_), .Y(mai_mai_n19_));
  NA2        m009(.A(i_0_), .B(mai_mai_n19_), .Y(mai_mai_n20_));
  INV        m010(.A(i_7_), .Y(mai_mai_n21_));
  NA3        m011(.A(i_6_), .B(i_5_), .C(mai_mai_n21_), .Y(mai_mai_n22_));
  NOi21      m012(.An(i_8_), .B(i_6_), .Y(mai_mai_n23_));
  NA2        m013(.A(mai_mai_n23_), .B(i_5_), .Y(mai_mai_n24_));
  AOI210     m014(.A0(mai_mai_n24_), .A1(mai_mai_n22_), .B0(mai_mai_n20_), .Y(mai_mai_n25_));
  AOI210     m015(.A0(mai_mai_n25_), .A1(mai_mai_n11_), .B0(mai_mai_n18_), .Y(mai_mai_n26_));
  NA2        m016(.A(i_0_), .B(mai_mai_n13_), .Y(mai_mai_n27_));
  NA2        m017(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n28_));
  NO2        m018(.A(i_2_), .B(i_4_), .Y(mai_mai_n29_));
  NA3        m019(.A(mai_mai_n29_), .B(i_6_), .C(i_8_), .Y(mai_mai_n30_));
  AOI210     m020(.A0(mai_mai_n28_), .A1(mai_mai_n27_), .B0(mai_mai_n30_), .Y(mai_mai_n31_));
  INV        m021(.A(i_2_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_5_), .B(i_0_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_6_), .B(i_8_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_0_), .B(i_4_), .Y(mai_mai_n35_));
  XO2        m025(.A(i_1_), .B(i_3_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_5_), .Y(mai_mai_n37_));
  AN3        m027(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(mai_mai_n35_), .Y(mai_mai_n38_));
  INV        m028(.A(i_1_), .Y(mai_mai_n39_));
  NOi21      m029(.An(i_3_), .B(i_0_), .Y(mai_mai_n40_));
  NA2        m030(.A(mai_mai_n40_), .B(mai_mai_n39_), .Y(mai_mai_n41_));
  NA3        m031(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n42_));
  AOI210     m032(.A0(mai_mai_n42_), .A1(mai_mai_n22_), .B0(mai_mai_n41_), .Y(mai_mai_n43_));
  NO3        m033(.A(mai_mai_n43_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n44_));
  NOi21      m034(.An(i_4_), .B(i_0_), .Y(mai_mai_n45_));
  INV        m035(.A(mai_mai_n14_), .Y(mai_mai_n46_));
  NA2        m036(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n47_));
  NOi21      m037(.An(i_2_), .B(i_8_), .Y(mai_mai_n48_));
  NO3        m038(.A(mai_mai_n48_), .B(mai_mai_n45_), .C(mai_mai_n35_), .Y(mai_mai_n49_));
  NO3        m039(.A(mai_mai_n49_), .B(mai_mai_n47_), .C(mai_mai_n46_), .Y(mai_mai_n50_));
  INV        m040(.A(mai_mai_n50_), .Y(mai_mai_n51_));
  NOi31      m041(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_4_), .B(i_3_), .Y(mai_mai_n53_));
  NOi21      m043(.An(i_1_), .B(i_4_), .Y(mai_mai_n54_));
  AN2        m044(.A(i_8_), .B(i_7_), .Y(mai_mai_n55_));
  INV        m045(.A(mai_mai_n55_), .Y(mai_mai_n56_));
  NOi21      m046(.An(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NO2        m047(.A(mai_mai_n56_), .B(mai_mai_n47_), .Y(mai_mai_n58_));
  NA2        m048(.A(mai_mai_n58_), .B(mai_mai_n32_), .Y(mai_mai_n59_));
  NA4        m049(.A(mai_mai_n59_), .B(mai_mai_n51_), .C(mai_mai_n44_), .D(mai_mai_n26_), .Y(mai_mai_n60_));
  NA2        m050(.A(i_8_), .B(mai_mai_n21_), .Y(mai_mai_n61_));
  AOI220     m051(.A0(mai_mai_n40_), .A1(i_1_), .B0(mai_mai_n36_), .B1(i_2_), .Y(mai_mai_n62_));
  NOi21      m052(.An(i_1_), .B(i_2_), .Y(mai_mai_n63_));
  NO2        m053(.A(mai_mai_n62_), .B(mai_mai_n61_), .Y(mai_mai_n64_));
  NA2        m054(.A(mai_mai_n64_), .B(mai_mai_n13_), .Y(mai_mai_n65_));
  NA3        m055(.A(mai_mai_n16_), .B(i_2_), .C(i_6_), .Y(mai_mai_n66_));
  INV        m056(.A(mai_mai_n66_), .Y(mai_mai_n67_));
  NO2        m057(.A(i_0_), .B(i_4_), .Y(mai_mai_n68_));
  AOI220     m058(.A0(mai_mai_n68_), .A1(mai_mai_n67_), .B0(mai_mai_n57_), .B1(mai_mai_n53_), .Y(mai_mai_n69_));
  NA2        m059(.A(mai_mai_n69_), .B(mai_mai_n65_), .Y(mai_mai_n70_));
  NAi21      m060(.An(i_3_), .B(i_6_), .Y(mai_mai_n71_));
  NO2        m061(.A(mai_mai_n71_), .B(i_0_), .Y(mai_mai_n72_));
  NOi21      m062(.An(i_7_), .B(i_8_), .Y(mai_mai_n73_));
  NOi21      m063(.An(i_6_), .B(i_5_), .Y(mai_mai_n74_));
  OAI210     m064(.A0(mai_mai_n74_), .A1(mai_mai_n72_), .B0(mai_mai_n63_), .Y(mai_mai_n75_));
  NA3        m065(.A(mai_mai_n23_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n76_));
  INV        m066(.A(mai_mai_n76_), .Y(mai_mai_n77_));
  AOI220     m067(.A0(mai_mai_n40_), .A1(mai_mai_n39_), .B0(mai_mai_n16_), .B1(mai_mai_n32_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n19_), .B(i_5_), .C(i_7_), .Y(mai_mai_n79_));
  NO2        m069(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NO2        m070(.A(mai_mai_n80_), .B(mai_mai_n77_), .Y(mai_mai_n81_));
  NA3        m071(.A(mai_mai_n57_), .B(mai_mai_n32_), .C(i_3_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n39_), .B(i_6_), .Y(mai_mai_n83_));
  AOI210     m073(.A0(mai_mai_n83_), .A1(mai_mai_n20_), .B0(mai_mai_n82_), .Y(mai_mai_n84_));
  NAi21      m074(.An(i_6_), .B(i_0_), .Y(mai_mai_n85_));
  NA3        m075(.A(mai_mai_n54_), .B(i_5_), .C(mai_mai_n21_), .Y(mai_mai_n86_));
  NOi21      m076(.An(i_4_), .B(i_6_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_5_), .B(i_3_), .Y(mai_mai_n88_));
  NO2        m078(.A(mai_mai_n86_), .B(mai_mai_n85_), .Y(mai_mai_n89_));
  NO2        m079(.A(mai_mai_n89_), .B(mai_mai_n84_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n57_), .B(mai_mai_n12_), .Y(mai_mai_n91_));
  NA2        m081(.A(mai_mai_n34_), .B(mai_mai_n13_), .Y(mai_mai_n92_));
  NOi21      m082(.An(i_3_), .B(i_1_), .Y(mai_mai_n93_));
  NA2        m083(.A(mai_mai_n93_), .B(i_4_), .Y(mai_mai_n94_));
  AOI210     m084(.A0(mai_mai_n92_), .A1(mai_mai_n91_), .B0(mai_mai_n94_), .Y(mai_mai_n95_));
  INV        m085(.A(mai_mai_n95_), .Y(mai_mai_n96_));
  NA4        m086(.A(mai_mai_n96_), .B(mai_mai_n90_), .C(mai_mai_n81_), .D(mai_mai_n75_), .Y(mai_mai_n97_));
  NA2        m087(.A(mai_mai_n48_), .B(mai_mai_n14_), .Y(mai_mai_n98_));
  NOi21      m088(.An(i_0_), .B(i_2_), .Y(mai_mai_n99_));
  NA2        m089(.A(mai_mai_n99_), .B(mai_mai_n87_), .Y(mai_mai_n100_));
  NA3        m090(.A(mai_mai_n45_), .B(mai_mai_n37_), .C(mai_mai_n16_), .Y(mai_mai_n101_));
  NA3        m091(.A(mai_mai_n99_), .B(mai_mai_n53_), .C(mai_mai_n34_), .Y(mai_mai_n102_));
  NA3        m092(.A(mai_mai_n102_), .B(mai_mai_n101_), .C(mai_mai_n100_), .Y(mai_mai_n103_));
  NA3        m093(.A(mai_mai_n52_), .B(i_6_), .C(i_7_), .Y(mai_mai_n104_));
  NA3        m094(.A(mai_mai_n54_), .B(mai_mai_n40_), .C(i_5_), .Y(mai_mai_n105_));
  NA2        m095(.A(mai_mai_n105_), .B(mai_mai_n104_), .Y(mai_mai_n106_));
  NO2        m096(.A(mai_mai_n106_), .B(mai_mai_n103_), .Y(mai_mai_n107_));
  NOi21      m097(.An(i_5_), .B(i_2_), .Y(mai_mai_n108_));
  AOI220     m098(.A0(mai_mai_n108_), .A1(mai_mai_n73_), .B0(mai_mai_n55_), .B1(mai_mai_n29_), .Y(mai_mai_n109_));
  AOI210     m099(.A0(mai_mai_n109_), .A1(mai_mai_n98_), .B0(mai_mai_n83_), .Y(mai_mai_n110_));
  NO4        m100(.A(i_2_), .B(mai_mai_n19_), .C(mai_mai_n11_), .D(mai_mai_n13_), .Y(mai_mai_n111_));
  NA2        m101(.A(i_2_), .B(i_4_), .Y(mai_mai_n112_));
  AOI210     m102(.A0(mai_mai_n85_), .A1(mai_mai_n71_), .B0(mai_mai_n112_), .Y(mai_mai_n113_));
  NO2        m103(.A(i_8_), .B(i_7_), .Y(mai_mai_n114_));
  OA210      m104(.A0(mai_mai_n113_), .A1(mai_mai_n111_), .B0(mai_mai_n114_), .Y(mai_mai_n115_));
  NA3        m105(.A(mai_mai_n93_), .B(i_0_), .C(i_5_), .Y(mai_mai_n116_));
  NO2        m106(.A(mai_mai_n116_), .B(i_4_), .Y(mai_mai_n117_));
  NO3        m107(.A(mai_mai_n117_), .B(mai_mai_n115_), .C(mai_mai_n110_), .Y(mai_mai_n118_));
  NA2        m108(.A(mai_mai_n73_), .B(mai_mai_n12_), .Y(mai_mai_n119_));
  INV        m109(.A(i_2_), .Y(mai_mai_n120_));
  NA2        m110(.A(mai_mai_n45_), .B(i_3_), .Y(mai_mai_n121_));
  AOI210     m111(.A0(mai_mai_n121_), .A1(mai_mai_n120_), .B0(mai_mai_n119_), .Y(mai_mai_n122_));
  NO2        m112(.A(mai_mai_n82_), .B(mai_mai_n28_), .Y(mai_mai_n123_));
  NA3        m113(.A(mai_mai_n88_), .B(mai_mai_n55_), .C(mai_mai_n39_), .Y(mai_mai_n124_));
  NA2        m114(.A(mai_mai_n48_), .B(mai_mai_n33_), .Y(mai_mai_n125_));
  NA2        m115(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n126_));
  NO3        m116(.A(mai_mai_n126_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n127_));
  NA3        m117(.A(mai_mai_n127_), .B(mai_mai_n118_), .C(mai_mai_n107_), .Y(mai_mai_n128_));
  OR4        m118(.A(mai_mai_n128_), .B(mai_mai_n97_), .C(mai_mai_n70_), .D(mai_mai_n60_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  INV        u005(.A(i_0_), .Y(men_men_n16_));
  NOi21      u006(.An(i_1_), .B(i_3_), .Y(men_men_n17_));
  INV        u007(.A(i_4_), .Y(men_men_n18_));
  NA2        u008(.A(i_0_), .B(men_men_n18_), .Y(men_men_n19_));
  INV        u009(.A(i_7_), .Y(men_men_n20_));
  NA3        u010(.A(i_6_), .B(i_5_), .C(men_men_n20_), .Y(men_men_n21_));
  NOi21      u011(.An(i_8_), .B(i_6_), .Y(men_men_n22_));
  NOi21      u012(.An(i_1_), .B(i_8_), .Y(men_men_n23_));
  AOI220     u013(.A0(men_men_n23_), .A1(i_2_), .B0(men_men_n22_), .B1(i_5_), .Y(men_men_n24_));
  AOI210     u014(.A0(men_men_n24_), .A1(men_men_n21_), .B0(men_men_n19_), .Y(men_men_n25_));
  NA2        u015(.A(men_men_n25_), .B(men_men_n11_), .Y(men_men_n26_));
  NA2        u016(.A(men_men_n16_), .B(i_5_), .Y(men_men_n27_));
  INV        u017(.A(i_2_), .Y(men_men_n28_));
  NOi21      u018(.An(i_5_), .B(i_0_), .Y(men_men_n29_));
  NOi21      u019(.An(i_6_), .B(i_8_), .Y(men_men_n30_));
  NOi21      u020(.An(i_7_), .B(i_1_), .Y(men_men_n31_));
  NOi21      u021(.An(i_5_), .B(i_6_), .Y(men_men_n32_));
  AOI220     u022(.A0(men_men_n32_), .A1(men_men_n31_), .B0(men_men_n30_), .B1(men_men_n29_), .Y(men_men_n33_));
  NO3        u023(.A(men_men_n33_), .B(men_men_n28_), .C(i_4_), .Y(men_men_n34_));
  NOi21      u024(.An(i_0_), .B(i_4_), .Y(men_men_n35_));
  XO2        u025(.A(i_1_), .B(i_3_), .Y(men_men_n36_));
  NOi21      u026(.An(i_7_), .B(i_5_), .Y(men_men_n37_));
  AN3        u027(.A(men_men_n37_), .B(men_men_n36_), .C(men_men_n35_), .Y(men_men_n38_));
  INV        u028(.A(i_1_), .Y(men_men_n39_));
  NO2        u029(.A(men_men_n38_), .B(men_men_n34_), .Y(men_men_n40_));
  NA2        u030(.A(i_1_), .B(men_men_n11_), .Y(men_men_n41_));
  NOi21      u031(.An(i_4_), .B(i_0_), .Y(men_men_n42_));
  NA2        u032(.A(i_1_), .B(men_men_n14_), .Y(men_men_n43_));
  NOi21      u033(.An(i_2_), .B(i_8_), .Y(men_men_n44_));
  NOi31      u034(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n45_));
  NA2        u035(.A(men_men_n45_), .B(i_0_), .Y(men_men_n46_));
  NOi21      u036(.An(i_4_), .B(i_3_), .Y(men_men_n47_));
  NOi21      u037(.An(i_1_), .B(i_4_), .Y(men_men_n48_));
  OAI210     u038(.A0(men_men_n48_), .A1(men_men_n47_), .B0(men_men_n44_), .Y(men_men_n49_));
  NA2        u039(.A(men_men_n49_), .B(men_men_n46_), .Y(men_men_n50_));
  NA2        u040(.A(i_8_), .B(men_men_n12_), .Y(men_men_n51_));
  NOi21      u041(.An(i_8_), .B(i_7_), .Y(men_men_n52_));
  NA3        u042(.A(men_men_n52_), .B(men_men_n47_), .C(i_6_), .Y(men_men_n53_));
  OAI210     u043(.A0(men_men_n51_), .A1(men_men_n43_), .B0(men_men_n53_), .Y(men_men_n54_));
  AOI220     u044(.A0(men_men_n54_), .A1(men_men_n28_), .B0(men_men_n50_), .B1(men_men_n32_), .Y(men_men_n55_));
  NA3        u045(.A(men_men_n55_), .B(men_men_n40_), .C(men_men_n26_), .Y(men_men_n56_));
  NA2        u046(.A(i_8_), .B(i_7_), .Y(men_men_n57_));
  NO3        u047(.A(men_men_n57_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n58_));
  NA2        u048(.A(i_8_), .B(men_men_n20_), .Y(men_men_n59_));
  NOi21      u049(.An(i_1_), .B(i_2_), .Y(men_men_n60_));
  NO2        u050(.A(men_men_n136_), .B(men_men_n59_), .Y(men_men_n61_));
  OAI210     u051(.A0(men_men_n61_), .A1(men_men_n58_), .B0(men_men_n14_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n23_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n63_));
  INV        u053(.A(men_men_n63_), .Y(men_men_n64_));
  NOi32      u054(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(i_3_), .Y(men_men_n66_));
  NA3        u056(.A(men_men_n17_), .B(i_2_), .C(i_6_), .Y(men_men_n67_));
  NA2        u057(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n68_));
  NO2        u058(.A(i_0_), .B(i_4_), .Y(men_men_n69_));
  AOI210     u059(.A0(men_men_n69_), .A1(men_men_n68_), .B0(men_men_n64_), .Y(men_men_n70_));
  NA2        u060(.A(men_men_n70_), .B(men_men_n62_), .Y(men_men_n71_));
  NA2        u061(.A(men_men_n30_), .B(men_men_n29_), .Y(men_men_n72_));
  NOi21      u062(.An(i_7_), .B(i_8_), .Y(men_men_n73_));
  NOi31      u063(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n74_));
  AOI210     u064(.A0(men_men_n73_), .A1(men_men_n12_), .B0(men_men_n74_), .Y(men_men_n75_));
  OAI210     u065(.A0(men_men_n75_), .A1(men_men_n11_), .B0(men_men_n72_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n76_), .B(men_men_n60_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n22_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n78_));
  AOI210     u068(.A0(men_men_n19_), .A1(men_men_n41_), .B0(men_men_n78_), .Y(men_men_n79_));
  NA3        u069(.A(men_men_n18_), .B(i_5_), .C(i_7_), .Y(men_men_n80_));
  OAI210     u070(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n81_));
  NA3        u071(.A(men_men_n57_), .B(men_men_n17_), .C(men_men_n16_), .Y(men_men_n82_));
  OAI220     u072(.A0(men_men_n82_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(i_2_), .Y(men_men_n83_));
  NO2        u073(.A(men_men_n83_), .B(men_men_n79_), .Y(men_men_n84_));
  NA3        u074(.A(men_men_n52_), .B(men_men_n28_), .C(i_3_), .Y(men_men_n85_));
  NO2        u075(.A(men_men_n19_), .B(men_men_n85_), .Y(men_men_n86_));
  NOi21      u076(.An(i_2_), .B(i_1_), .Y(men_men_n87_));
  AN2        u077(.A(men_men_n87_), .B(men_men_n42_), .Y(men_men_n88_));
  NOi21      u078(.An(i_4_), .B(i_6_), .Y(men_men_n89_));
  NOi21      u079(.An(i_5_), .B(i_3_), .Y(men_men_n90_));
  NA3        u080(.A(men_men_n90_), .B(men_men_n60_), .C(men_men_n89_), .Y(men_men_n91_));
  INV        u081(.A(men_men_n91_), .Y(men_men_n92_));
  NA2        u082(.A(men_men_n60_), .B(men_men_n30_), .Y(men_men_n93_));
  NOi21      u083(.An(men_men_n37_), .B(men_men_n93_), .Y(men_men_n94_));
  NO4        u084(.A(men_men_n94_), .B(men_men_n92_), .C(men_men_n88_), .D(men_men_n86_), .Y(men_men_n95_));
  NOi21      u085(.An(i_6_), .B(i_1_), .Y(men_men_n96_));
  AOI220     u086(.A0(men_men_n96_), .A1(i_7_), .B0(men_men_n22_), .B1(i_5_), .Y(men_men_n97_));
  NOi31      u087(.An(men_men_n42_), .B(men_men_n97_), .C(i_2_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n73_), .B(men_men_n14_), .Y(men_men_n99_));
  NOi21      u089(.An(i_3_), .B(men_men_n99_), .Y(men_men_n100_));
  NO2        u090(.A(men_men_n100_), .B(men_men_n98_), .Y(men_men_n101_));
  NA4        u091(.A(men_men_n101_), .B(men_men_n95_), .C(men_men_n84_), .D(men_men_n77_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n44_), .B(men_men_n15_), .Y(men_men_n103_));
  NOi31      u093(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n104_), .B(i_7_), .Y(men_men_n105_));
  NA2        u095(.A(men_men_n105_), .B(men_men_n103_), .Y(men_men_n106_));
  NA2        u096(.A(men_men_n106_), .B(men_men_n35_), .Y(men_men_n107_));
  NA2        u097(.A(men_men_n47_), .B(men_men_n31_), .Y(men_men_n108_));
  NO2        u098(.A(men_men_n108_), .B(men_men_n27_), .Y(men_men_n109_));
  NA3        u099(.A(men_men_n42_), .B(men_men_n37_), .C(men_men_n17_), .Y(men_men_n110_));
  NOi32      u100(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n111_), .B(men_men_n104_), .Y(men_men_n112_));
  NA3        u102(.A(i_0_), .B(men_men_n47_), .C(men_men_n30_), .Y(men_men_n113_));
  NA3        u103(.A(men_men_n113_), .B(men_men_n112_), .C(men_men_n110_), .Y(men_men_n114_));
  NA3        u104(.A(men_men_n45_), .B(i_6_), .C(men_men_n14_), .Y(men_men_n115_));
  NA4        u105(.A(men_men_n48_), .B(men_men_n32_), .C(men_men_n16_), .D(i_8_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NO3        u107(.A(men_men_n117_), .B(men_men_n114_), .C(men_men_n109_), .Y(men_men_n118_));
  NO3        u108(.A(i_2_), .B(men_men_n11_), .C(men_men_n14_), .Y(men_men_n119_));
  NA2        u109(.A(i_2_), .B(i_4_), .Y(men_men_n120_));
  AOI210     u110(.A0(i_6_), .A1(i_3_), .B0(men_men_n120_), .Y(men_men_n121_));
  NO2        u111(.A(i_8_), .B(i_7_), .Y(men_men_n122_));
  OA210      u112(.A0(men_men_n121_), .A1(men_men_n119_), .B0(men_men_n122_), .Y(men_men_n123_));
  INV        u113(.A(men_men_n123_), .Y(men_men_n124_));
  NA4        u114(.A(men_men_n90_), .B(i_8_), .C(men_men_n39_), .D(men_men_n18_), .Y(men_men_n125_));
  NA3        u115(.A(men_men_n74_), .B(i_3_), .C(i_0_), .Y(men_men_n126_));
  NA2        u116(.A(men_men_n29_), .B(men_men_n15_), .Y(men_men_n127_));
  NOi31      u117(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n128_));
  OAI210     u118(.A0(men_men_n111_), .A1(men_men_n65_), .B0(men_men_n128_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n129_), .B(men_men_n127_), .C(men_men_n126_), .D(men_men_n125_), .Y(men_men_n130_));
  INV        u120(.A(men_men_n130_), .Y(men_men_n131_));
  NA4        u121(.A(men_men_n131_), .B(men_men_n124_), .C(men_men_n118_), .D(men_men_n107_), .Y(men_men_n132_));
  OR4        u122(.A(men_men_n132_), .B(men_men_n102_), .C(men_men_n71_), .D(men_men_n56_), .Y(men00));
  INV        u123(.A(i_1_), .Y(men_men_n136_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule