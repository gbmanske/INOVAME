// Benchmark "top" written by ABC on Fri Jun 21 17:49:28 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n139_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n961_, new_new_n962_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  NO2        g036(.A(new_new_n58_), .B(new_new_n57_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA3        g041(.A(new_new_n63_), .B(new_new_n61_), .C(new_new_n31_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_10_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(i_6_), .Y(new_new_n66_));
  NAi31      g044(.An(new_new_n66_), .B(new_new_n64_), .C(new_new_n60_), .Y(new_new_n67_));
  NA2        g045(.A(new_new_n50_), .B(i_2_), .Y(new_new_n68_));
  AOI210     g046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n69_));
  NA2        g047(.A(i_1_), .B(i_6_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n25_), .Y(new_new_n71_));
  INV        g049(.A(i_0_), .Y(new_new_n72_));
  NAi21      g050(.An(i_5_), .B(i_10_), .Y(new_new_n73_));
  NA2        g051(.A(i_5_), .B(i_9_), .Y(new_new_n74_));
  AOI210     g052(.A0(new_new_n74_), .A1(new_new_n73_), .B0(new_new_n72_), .Y(new_new_n75_));
  NO2        g053(.A(new_new_n75_), .B(new_new_n71_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n76_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n77_), .A1(new_new_n67_), .B0(i_0_), .Y(new_new_n78_));
  NA2        g056(.A(i_12_), .B(i_5_), .Y(new_new_n79_));
  NA2        g057(.A(i_2_), .B(i_8_), .Y(new_new_n80_));
  NO2        g058(.A(new_new_n80_), .B(new_new_n57_), .Y(new_new_n81_));
  NO2        g059(.A(i_3_), .B(i_9_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_7_), .Y(new_new_n83_));
  NO2        g061(.A(new_new_n82_), .B(new_new_n62_), .Y(new_new_n84_));
  INV        g062(.A(i_6_), .Y(new_new_n85_));
  NO2        g063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  INV        g064(.A(new_new_n86_), .Y(new_new_n87_));
  OAI210     g065(.A0(new_new_n84_), .A1(new_new_n81_), .B0(new_new_n87_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n62_), .Y(new_new_n91_));
  NA2        g069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g070(.A(new_new_n92_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n79_), .Y(new_new_n95_));
  AN3        g073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g077(.A0(new_new_n99_), .A1(new_new_n61_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g078(.A(i_7_), .Y(new_new_n101_));
  NA2        g079(.A(new_new_n46_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n103_), .B(new_new_n85_), .Y(new_new_n104_));
  NA2        g082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  NO3        g086(.A(new_new_n108_), .B(new_new_n89_), .C(new_new_n53_), .Y(new_new_n109_));
  AN2        g087(.A(i_2_), .B(i_10_), .Y(new_new_n110_));
  NO2        g088(.A(new_new_n110_), .B(i_7_), .Y(new_new_n111_));
  OR2        g089(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n112_));
  NO2        g090(.A(i_8_), .B(new_new_n101_), .Y(new_new_n113_));
  NO3        g091(.A(new_new_n113_), .B(new_new_n112_), .C(new_new_n111_), .Y(new_new_n114_));
  NA2        g092(.A(i_12_), .B(i_7_), .Y(new_new_n115_));
  NO2        g093(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(i_0_), .Y(new_new_n117_));
  NA2        g095(.A(i_11_), .B(i_12_), .Y(new_new_n118_));
  OAI210     g096(.A0(new_new_n117_), .A1(new_new_n115_), .B0(new_new_n118_), .Y(new_new_n119_));
  NO2        g097(.A(new_new_n119_), .B(new_new_n114_), .Y(new_new_n120_));
  NAi41      g098(.An(new_new_n109_), .B(new_new_n120_), .C(new_new_n107_), .D(new_new_n100_), .Y(new_new_n121_));
  NOi21      g099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g104(.A(new_new_n126_), .B(new_new_n46_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n128_));
  NAi21      g106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n129_), .B(new_new_n61_), .Y(new_new_n130_));
  NOi31      g108(.An(new_new_n130_), .B(new_new_n128_), .C(new_new_n127_), .Y(new_new_n131_));
  NO2        g109(.A(i_1_), .B(new_new_n85_), .Y(new_new_n132_));
  NO2        g110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  AO210      g112(.A0(new_new_n134_), .A1(new_new_n47_), .B0(new_new_n132_), .Y(new_new_n135_));
  OAI220     g113(.A0(new_new_n135_), .A1(new_new_n108_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n136_));
  NO3        g114(.A(new_new_n136_), .B(new_new_n121_), .C(new_new_n95_), .Y(new_new_n137_));
  NA3        g115(.A(new_new_n137_), .B(new_new_n78_), .C(new_new_n56_), .Y(ori2));
  NO2        g116(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n139_));
  NA2        g117(.A(i_6_), .B(new_new_n25_), .Y(new_new_n140_));
  NA2        g118(.A(new_new_n140_), .B(new_new_n139_), .Y(new_new_n141_));
  NA4        g119(.A(new_new_n141_), .B(new_new_n76_), .C(new_new_n68_), .D(new_new_n30_), .Y(ori0));
  AN2        g120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  AN2        g129(.A(new_new_n145_), .B(new_new_n82_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n72_), .B(new_new_n46_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g136(.A(new_new_n158_), .B(new_new_n79_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g142(.A(new_new_n72_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  NO2        g146(.A(new_new_n168_), .B(new_new_n144_), .Y(new_new_n169_));
  NOi21      g147(.An(i_4_), .B(i_9_), .Y(new_new_n170_));
  NOi21      g148(.An(i_11_), .B(i_13_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n171_), .B(new_new_n170_), .Y(new_new_n172_));
  NO2        g150(.A(i_4_), .B(i_5_), .Y(new_new_n173_));
  NAi21      g151(.An(i_12_), .B(i_11_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n72_), .B(new_new_n62_), .Y(new_new_n175_));
  NA2        g153(.A(new_new_n175_), .B(new_new_n46_), .Y(new_new_n176_));
  NAi31      g154(.An(i_4_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n177_));
  NA2        g155(.A(i_3_), .B(i_5_), .Y(new_new_n178_));
  OR2        g156(.A(new_new_n178_), .B(new_new_n172_), .Y(new_new_n179_));
  AOI210     g157(.A0(new_new_n179_), .A1(new_new_n177_), .B0(new_new_n176_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n72_), .B(i_5_), .Y(new_new_n181_));
  NO2        g159(.A(i_13_), .B(i_10_), .Y(new_new_n182_));
  NA3        g160(.A(new_new_n182_), .B(new_new_n181_), .C(new_new_n44_), .Y(new_new_n183_));
  NO2        g161(.A(i_2_), .B(i_1_), .Y(new_new_n184_));
  NA2        g162(.A(new_new_n184_), .B(i_3_), .Y(new_new_n185_));
  NAi21      g163(.An(i_4_), .B(i_12_), .Y(new_new_n186_));
  INV        g164(.A(new_new_n180_), .Y(new_new_n187_));
  INV        g165(.A(i_8_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n188_), .B(i_7_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n189_), .B(i_6_), .Y(new_new_n190_));
  NO3        g168(.A(i_3_), .B(new_new_n85_), .C(new_new_n48_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(new_new_n113_), .Y(new_new_n192_));
  NO3        g170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n194_));
  NO3        g172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n195_));
  OAI210     g173(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n195_), .Y(new_new_n196_));
  AOI210     g174(.A0(new_new_n196_), .A1(new_new_n194_), .B0(new_new_n192_), .Y(new_new_n197_));
  NO2        g175(.A(i_3_), .B(i_8_), .Y(new_new_n198_));
  NO3        g176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(new_new_n198_), .C(new_new_n40_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n103_), .B(new_new_n57_), .Y(new_new_n201_));
  INV        g179(.A(new_new_n201_), .Y(new_new_n202_));
  NO2        g180(.A(i_13_), .B(i_9_), .Y(new_new_n203_));
  NAi21      g181(.An(i_12_), .B(i_3_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n44_), .B(i_5_), .Y(new_new_n205_));
  NO3        g183(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n202_), .B(new_new_n200_), .Y(new_new_n207_));
  AOI210     g185(.A0(new_new_n207_), .A1(i_7_), .B0(new_new_n197_), .Y(new_new_n208_));
  OAI220     g186(.A0(new_new_n208_), .A1(i_4_), .B0(new_new_n190_), .B1(new_new_n187_), .Y(new_new_n209_));
  NAi21      g187(.An(i_12_), .B(i_7_), .Y(new_new_n210_));
  NA3        g188(.A(i_13_), .B(new_new_n188_), .C(i_10_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(new_new_n210_), .Y(new_new_n212_));
  NA2        g190(.A(i_0_), .B(i_5_), .Y(new_new_n213_));
  NA2        g191(.A(new_new_n213_), .B(new_new_n104_), .Y(new_new_n214_));
  OAI220     g192(.A0(new_new_n214_), .A1(new_new_n185_), .B0(new_new_n176_), .B1(new_new_n134_), .Y(new_new_n215_));
  NAi31      g193(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n36_), .B(i_13_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n218_));
  INV        g196(.A(i_13_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n219_), .Y(new_new_n220_));
  NA2        g198(.A(new_new_n215_), .B(new_new_n212_), .Y(new_new_n221_));
  NO2        g199(.A(i_12_), .B(new_new_n37_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n178_), .B(i_4_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  OR2        g202(.A(i_8_), .B(i_7_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n225_), .B(new_new_n85_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n53_), .B(i_1_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n228_));
  INV        g206(.A(i_12_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n44_), .B(new_new_n229_), .Y(new_new_n230_));
  NO3        g208(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n231_));
  NA2        g209(.A(i_2_), .B(i_1_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n228_), .B(new_new_n224_), .Y(new_new_n233_));
  NO3        g211(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n234_));
  NAi21      g212(.An(i_4_), .B(i_3_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n235_), .B(new_new_n74_), .Y(new_new_n236_));
  NO2        g214(.A(i_0_), .B(i_6_), .Y(new_new_n237_));
  NOi41      g215(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n232_), .B(new_new_n178_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n233_), .Y(new_new_n240_));
  NO2        g218(.A(i_11_), .B(new_new_n219_), .Y(new_new_n241_));
  NOi21      g219(.An(i_1_), .B(i_6_), .Y(new_new_n242_));
  NAi21      g220(.An(i_3_), .B(i_7_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n229_), .B(i_9_), .Y(new_new_n244_));
  NO2        g222(.A(i_12_), .B(i_3_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n72_), .B(i_5_), .Y(new_new_n246_));
  NA2        g224(.A(i_3_), .B(i_9_), .Y(new_new_n247_));
  NAi21      g225(.An(i_7_), .B(i_10_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n248_), .B(new_new_n247_), .Y(new_new_n249_));
  NA3        g227(.A(new_new_n249_), .B(new_new_n246_), .C(new_new_n63_), .Y(new_new_n250_));
  INV        g228(.A(new_new_n250_), .Y(new_new_n251_));
  INV        g229(.A(new_new_n144_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n229_), .B(i_13_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n253_), .B(new_new_n74_), .Y(new_new_n254_));
  AOI220     g232(.A0(new_new_n254_), .A1(new_new_n252_), .B0(new_new_n251_), .B1(new_new_n241_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n225_), .B(new_new_n37_), .Y(new_new_n256_));
  NA2        g234(.A(i_12_), .B(i_6_), .Y(new_new_n257_));
  OR2        g235(.A(i_13_), .B(i_9_), .Y(new_new_n258_));
  NO3        g236(.A(new_new_n258_), .B(new_new_n257_), .C(new_new_n48_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n235_), .B(i_2_), .Y(new_new_n260_));
  NA3        g238(.A(new_new_n260_), .B(new_new_n259_), .C(new_new_n44_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n241_), .B(i_9_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n246_), .B(new_new_n63_), .Y(new_new_n263_));
  OAI210     g241(.A0(new_new_n263_), .A1(new_new_n262_), .B0(new_new_n261_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n155_), .B(new_new_n62_), .Y(new_new_n265_));
  NO3        g243(.A(i_11_), .B(new_new_n219_), .C(new_new_n25_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n243_), .B(i_8_), .Y(new_new_n267_));
  NO2        g245(.A(i_6_), .B(new_new_n48_), .Y(new_new_n268_));
  NA3        g246(.A(new_new_n268_), .B(new_new_n267_), .C(new_new_n266_), .Y(new_new_n269_));
  NO3        g247(.A(new_new_n26_), .B(new_new_n85_), .C(i_5_), .Y(new_new_n270_));
  NA3        g248(.A(new_new_n270_), .B(new_new_n256_), .C(new_new_n220_), .Y(new_new_n271_));
  AOI210     g249(.A0(new_new_n271_), .A1(new_new_n269_), .B0(new_new_n265_), .Y(new_new_n272_));
  AOI210     g250(.A0(new_new_n264_), .A1(new_new_n256_), .B0(new_new_n272_), .Y(new_new_n273_));
  NA4        g251(.A(new_new_n273_), .B(new_new_n255_), .C(new_new_n240_), .D(new_new_n221_), .Y(new_new_n274_));
  NO3        g252(.A(i_12_), .B(new_new_n219_), .C(new_new_n37_), .Y(new_new_n275_));
  INV        g253(.A(new_new_n275_), .Y(new_new_n276_));
  NA2        g254(.A(i_8_), .B(new_new_n101_), .Y(new_new_n277_));
  NO3        g255(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n278_));
  AOI220     g256(.A0(new_new_n278_), .A1(new_new_n191_), .B0(new_new_n164_), .B1(new_new_n227_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(new_new_n277_), .Y(new_new_n280_));
  NO3        g258(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n232_), .B(i_0_), .Y(new_new_n282_));
  AOI220     g260(.A0(new_new_n282_), .A1(new_new_n189_), .B0(new_new_n281_), .B1(new_new_n143_), .Y(new_new_n283_));
  NA2        g261(.A(new_new_n268_), .B(new_new_n26_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(new_new_n283_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n58_), .B(i_6_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n166_), .B(new_new_n144_), .Y(new_new_n287_));
  NO3        g265(.A(new_new_n287_), .B(new_new_n285_), .C(new_new_n280_), .Y(new_new_n288_));
  NO2        g266(.A(i_3_), .B(i_10_), .Y(new_new_n289_));
  NA3        g267(.A(new_new_n289_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n290_));
  NO2        g268(.A(i_2_), .B(new_new_n101_), .Y(new_new_n291_));
  NA2        g269(.A(i_1_), .B(new_new_n36_), .Y(new_new_n292_));
  AN2        g270(.A(i_3_), .B(i_10_), .Y(new_new_n293_));
  NO2        g271(.A(i_5_), .B(new_new_n37_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n288_), .B(new_new_n276_), .Y(new_new_n296_));
  NO4        g274(.A(new_new_n296_), .B(new_new_n274_), .C(new_new_n209_), .D(new_new_n169_), .Y(new_new_n297_));
  NO3        g275(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n298_));
  NO3        g276(.A(i_6_), .B(new_new_n188_), .C(i_7_), .Y(new_new_n299_));
  NA2        g277(.A(new_new_n299_), .B(new_new_n193_), .Y(new_new_n300_));
  INV        g278(.A(new_new_n300_), .Y(new_new_n301_));
  NO2        g279(.A(i_2_), .B(i_3_), .Y(new_new_n302_));
  OR2        g280(.A(i_0_), .B(i_5_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n213_), .B(new_new_n303_), .Y(new_new_n304_));
  NA4        g282(.A(new_new_n304_), .B(new_new_n226_), .C(new_new_n302_), .D(i_1_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n282_), .B(new_new_n164_), .C(new_new_n113_), .Y(new_new_n306_));
  NAi21      g284(.An(i_8_), .B(i_7_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n158_), .B(new_new_n46_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n306_), .B(new_new_n305_), .Y(new_new_n309_));
  OAI210     g287(.A0(new_new_n309_), .A1(new_new_n301_), .B0(i_4_), .Y(new_new_n310_));
  NO2        g288(.A(i_12_), .B(i_10_), .Y(new_new_n311_));
  NOi21      g289(.An(i_5_), .B(i_0_), .Y(new_new_n312_));
  NO2        g290(.A(i_2_), .B(new_new_n101_), .Y(new_new_n313_));
  NO4        g291(.A(new_new_n313_), .B(new_new_n292_), .C(new_new_n312_), .D(new_new_n129_), .Y(new_new_n314_));
  NA4        g292(.A(new_new_n83_), .B(new_new_n36_), .C(new_new_n85_), .D(i_8_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n314_), .B(new_new_n311_), .Y(new_new_n316_));
  NO2        g294(.A(i_6_), .B(i_8_), .Y(new_new_n317_));
  NOi21      g295(.An(i_0_), .B(i_2_), .Y(new_new_n318_));
  AN2        g296(.A(new_new_n318_), .B(new_new_n317_), .Y(new_new_n319_));
  NO2        g297(.A(i_1_), .B(i_7_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n316_), .B(new_new_n310_), .Y(new_new_n321_));
  NO3        g299(.A(new_new_n225_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n322_));
  NO3        g300(.A(new_new_n307_), .B(i_2_), .C(i_1_), .Y(new_new_n323_));
  OAI210     g301(.A0(new_new_n323_), .A1(new_new_n322_), .B0(i_6_), .Y(new_new_n324_));
  NA3        g302(.A(new_new_n242_), .B(new_new_n291_), .C(new_new_n188_), .Y(new_new_n325_));
  AOI210     g303(.A0(new_new_n325_), .A1(new_new_n324_), .B0(new_new_n304_), .Y(new_new_n326_));
  NOi21      g304(.An(new_new_n154_), .B(new_new_n104_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(new_new_n125_), .Y(new_new_n328_));
  OAI210     g306(.A0(new_new_n328_), .A1(new_new_n326_), .B0(i_3_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n188_), .B(i_9_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n330_), .B(new_new_n201_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n331_), .B(new_new_n46_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n332_), .B(new_new_n285_), .Y(new_new_n333_));
  AOI210     g311(.A0(new_new_n333_), .A1(new_new_n329_), .B0(new_new_n163_), .Y(new_new_n334_));
  AOI210     g312(.A0(new_new_n321_), .A1(new_new_n298_), .B0(new_new_n334_), .Y(new_new_n335_));
  NOi32      g313(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n336_));
  INV        g314(.A(new_new_n336_), .Y(new_new_n337_));
  NAi21      g315(.An(i_0_), .B(i_6_), .Y(new_new_n338_));
  NAi21      g316(.An(i_1_), .B(i_5_), .Y(new_new_n339_));
  NA2        g317(.A(new_new_n339_), .B(new_new_n338_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n340_), .B(new_new_n25_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(new_new_n160_), .Y(new_new_n342_));
  NAi41      g320(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n343_));
  OAI220     g321(.A0(new_new_n343_), .A1(new_new_n339_), .B0(new_new_n216_), .B1(new_new_n160_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n343_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n345_));
  NOi32      g323(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n346_));
  NAi21      g324(.An(i_6_), .B(i_1_), .Y(new_new_n347_));
  NA3        g325(.A(new_new_n347_), .B(new_new_n346_), .C(new_new_n46_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(i_0_), .Y(new_new_n349_));
  OR3        g327(.A(new_new_n349_), .B(new_new_n345_), .C(new_new_n344_), .Y(new_new_n350_));
  NO2        g328(.A(i_1_), .B(new_new_n101_), .Y(new_new_n351_));
  NAi21      g329(.An(i_3_), .B(i_4_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n352_), .B(i_9_), .Y(new_new_n353_));
  AN2        g331(.A(i_6_), .B(i_7_), .Y(new_new_n354_));
  OAI210     g332(.A0(new_new_n354_), .A1(new_new_n351_), .B0(new_new_n353_), .Y(new_new_n355_));
  NA2        g333(.A(i_2_), .B(i_7_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n352_), .B(i_10_), .Y(new_new_n357_));
  NA3        g335(.A(new_new_n357_), .B(new_new_n356_), .C(new_new_n237_), .Y(new_new_n358_));
  AOI210     g336(.A0(new_new_n358_), .A1(new_new_n355_), .B0(new_new_n181_), .Y(new_new_n359_));
  AOI210     g337(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n360_));
  OAI210     g338(.A0(new_new_n360_), .A1(new_new_n184_), .B0(new_new_n357_), .Y(new_new_n361_));
  AOI220     g339(.A0(new_new_n357_), .A1(new_new_n320_), .B0(new_new_n231_), .B1(new_new_n184_), .Y(new_new_n362_));
  AOI210     g340(.A0(new_new_n362_), .A1(new_new_n361_), .B0(i_5_), .Y(new_new_n363_));
  NO4        g341(.A(new_new_n363_), .B(new_new_n359_), .C(new_new_n350_), .D(new_new_n342_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n364_), .B(new_new_n337_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n366_));
  AN2        g344(.A(i_12_), .B(i_5_), .Y(new_new_n367_));
  NO2        g345(.A(i_4_), .B(new_new_n26_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n368_), .B(new_new_n367_), .Y(new_new_n369_));
  NO2        g347(.A(i_11_), .B(i_6_), .Y(new_new_n370_));
  NA3        g348(.A(new_new_n370_), .B(new_new_n308_), .C(new_new_n219_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n371_), .B(new_new_n369_), .Y(new_new_n372_));
  NO2        g350(.A(new_new_n235_), .B(i_5_), .Y(new_new_n373_));
  NO2        g351(.A(i_5_), .B(i_10_), .Y(new_new_n374_));
  AOI220     g352(.A0(new_new_n374_), .A1(new_new_n260_), .B0(new_new_n373_), .B1(new_new_n193_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n145_), .B(new_new_n45_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n377_));
  OAI210     g355(.A0(new_new_n377_), .A1(new_new_n372_), .B0(new_new_n366_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n151_), .B(new_new_n85_), .Y(new_new_n380_));
  OAI210     g358(.A0(new_new_n380_), .A1(new_new_n372_), .B0(new_new_n379_), .Y(new_new_n381_));
  NO3        g359(.A(new_new_n85_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n382_));
  NA3        g360(.A(new_new_n289_), .B(new_new_n74_), .C(new_new_n54_), .Y(new_new_n383_));
  NO2        g361(.A(i_11_), .B(i_12_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n384_), .B(new_new_n36_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n383_), .B(new_new_n385_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n374_), .B(new_new_n229_), .Y(new_new_n387_));
  NAi21      g365(.An(i_13_), .B(i_0_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n388_), .B(new_new_n232_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n386_), .B(new_new_n389_), .Y(new_new_n390_));
  NA3        g368(.A(new_new_n390_), .B(new_new_n381_), .C(new_new_n378_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n44_), .B(new_new_n219_), .Y(new_new_n392_));
  NO2        g370(.A(i_0_), .B(i_11_), .Y(new_new_n393_));
  AN2        g371(.A(i_1_), .B(i_6_), .Y(new_new_n394_));
  NOi21      g372(.An(i_2_), .B(i_12_), .Y(new_new_n395_));
  NAi21      g373(.An(i_9_), .B(i_4_), .Y(new_new_n396_));
  OR2        g374(.A(i_13_), .B(i_10_), .Y(new_new_n397_));
  NO3        g375(.A(new_new_n397_), .B(new_new_n118_), .C(new_new_n396_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n172_), .B(new_new_n124_), .Y(new_new_n399_));
  OR2        g377(.A(new_new_n211_), .B(new_new_n210_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n275_), .B(new_new_n401_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n268_), .B(new_new_n206_), .Y(new_new_n403_));
  OAI220     g381(.A0(new_new_n403_), .A1(new_new_n400_), .B0(new_new_n402_), .B1(new_new_n327_), .Y(new_new_n404_));
  INV        g382(.A(new_new_n404_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(new_new_n26_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n306_), .B(new_new_n305_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n178_), .B(new_new_n85_), .Y(new_new_n408_));
  AOI220     g386(.A0(new_new_n408_), .A1(i_1_), .B0(new_new_n270_), .B1(new_new_n206_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n277_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n410_), .B(new_new_n407_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n191_), .B(new_new_n96_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n308_), .B(new_new_n164_), .Y(new_new_n413_));
  AOI210     g391(.A0(new_new_n413_), .A1(new_new_n412_), .B0(new_new_n307_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n188_), .B(i_10_), .Y(new_new_n415_));
  NA3        g393(.A(new_new_n246_), .B(new_new_n63_), .C(i_2_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n286_), .B(new_new_n227_), .Y(new_new_n417_));
  OAI220     g395(.A0(new_new_n417_), .A1(new_new_n178_), .B0(new_new_n416_), .B1(new_new_n415_), .Y(new_new_n418_));
  NO2        g396(.A(i_3_), .B(new_new_n48_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n418_), .B(new_new_n414_), .Y(new_new_n420_));
  AOI210     g398(.A0(new_new_n420_), .A1(new_new_n411_), .B0(new_new_n262_), .Y(new_new_n421_));
  NO4        g399(.A(new_new_n421_), .B(new_new_n406_), .C(new_new_n391_), .D(new_new_n365_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n72_), .B(i_13_), .Y(new_new_n423_));
  NO2        g401(.A(i_10_), .B(i_9_), .Y(new_new_n424_));
  NAi21      g402(.An(i_12_), .B(i_8_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(i_3_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n46_), .B(i_4_), .Y(new_new_n427_));
  NA2        g405(.A(new_new_n427_), .B(new_new_n104_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n428_), .B(new_new_n200_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n257_), .B(new_new_n97_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n431_), .B(new_new_n430_), .Y(new_new_n432_));
  NA2        g410(.A(i_8_), .B(i_9_), .Y(new_new_n433_));
  AOI210     g411(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n434_));
  OR2        g412(.A(new_new_n434_), .B(new_new_n433_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n275_), .B(new_new_n201_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n435_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n241_), .B(new_new_n294_), .Y(new_new_n438_));
  NO3        g416(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n439_));
  INV        g417(.A(new_new_n439_), .Y(new_new_n440_));
  NA3        g418(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n441_));
  NA4        g419(.A(new_new_n146_), .B(new_new_n116_), .C(new_new_n79_), .D(new_new_n23_), .Y(new_new_n442_));
  OAI220     g420(.A0(new_new_n442_), .A1(new_new_n441_), .B0(new_new_n440_), .B1(new_new_n438_), .Y(new_new_n443_));
  NO3        g421(.A(new_new_n443_), .B(new_new_n437_), .C(new_new_n429_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n96_), .B(i_13_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n408_), .B(new_new_n366_), .Y(new_new_n446_));
  NO2        g424(.A(i_2_), .B(i_13_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n446_), .B(new_new_n445_), .Y(new_new_n448_));
  NO3        g426(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n449_));
  NO2        g427(.A(i_6_), .B(i_7_), .Y(new_new_n450_));
  NO2        g428(.A(i_11_), .B(i_1_), .Y(new_new_n451_));
  OR2        g429(.A(i_11_), .B(i_8_), .Y(new_new_n452_));
  NOi21      g430(.An(i_2_), .B(i_7_), .Y(new_new_n453_));
  NO2        g431(.A(i_3_), .B(new_new_n188_), .Y(new_new_n454_));
  NO2        g432(.A(i_6_), .B(i_10_), .Y(new_new_n455_));
  NA4        g433(.A(new_new_n455_), .B(new_new_n298_), .C(new_new_n454_), .D(new_new_n229_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n456_), .B(new_new_n156_), .Y(new_new_n457_));
  NA3        g435(.A(new_new_n238_), .B(new_new_n171_), .C(new_new_n133_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n158_), .B(i_3_), .Y(new_new_n460_));
  NAi31      g438(.An(new_new_n459_), .B(new_new_n460_), .C(new_new_n220_), .Y(new_new_n461_));
  NA3        g439(.A(new_new_n379_), .B(new_new_n175_), .C(new_new_n150_), .Y(new_new_n462_));
  NA3        g440(.A(new_new_n462_), .B(new_new_n461_), .C(new_new_n458_), .Y(new_new_n463_));
  NO3        g441(.A(new_new_n463_), .B(new_new_n457_), .C(new_new_n448_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n430_), .B(new_new_n367_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n439_), .B(new_new_n374_), .Y(new_new_n466_));
  NAi21      g444(.An(new_new_n211_), .B(new_new_n384_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n26_), .B(i_5_), .Y(new_new_n468_));
  NO2        g446(.A(i_0_), .B(new_new_n85_), .Y(new_new_n469_));
  NA3        g447(.A(new_new_n469_), .B(new_new_n468_), .C(new_new_n143_), .Y(new_new_n470_));
  OR3        g448(.A(new_new_n292_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n471_), .B(new_new_n470_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n27_), .B(i_10_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n298_), .B(new_new_n231_), .Y(new_new_n474_));
  OAI220     g452(.A0(new_new_n474_), .A1(new_new_n416_), .B0(new_new_n473_), .B1(new_new_n445_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n475_), .B(new_new_n472_), .Y(new_new_n476_));
  NA3        g454(.A(new_new_n476_), .B(new_new_n464_), .C(new_new_n444_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n123_), .B(new_new_n112_), .Y(new_new_n478_));
  AN2        g456(.A(new_new_n478_), .B(new_new_n430_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(new_new_n295_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n367_), .B(new_new_n219_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n336_), .B(new_new_n72_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n354_), .B(new_new_n346_), .Y(new_new_n483_));
  OR2        g461(.A(new_new_n481_), .B(new_new_n483_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n36_), .B(i_8_), .Y(new_new_n485_));
  AOI210     g463(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n398_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(new_new_n484_), .Y(new_new_n487_));
  INV        g465(.A(new_new_n487_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n246_), .B(new_new_n63_), .Y(new_new_n489_));
  OAI210     g467(.A0(i_8_), .A1(new_new_n489_), .B0(new_new_n135_), .Y(new_new_n490_));
  AOI210     g468(.A0(new_new_n189_), .A1(i_9_), .B0(new_new_n256_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n491_), .B(new_new_n194_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n178_), .B(new_new_n85_), .Y(new_new_n493_));
  AOI220     g471(.A0(new_new_n493_), .A1(new_new_n492_), .B0(new_new_n490_), .B1(new_new_n399_), .Y(new_new_n494_));
  NA3        g472(.A(new_new_n494_), .B(new_new_n488_), .C(new_new_n480_), .Y(new_new_n495_));
  NO2        g473(.A(i_12_), .B(new_new_n188_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n496_), .B(new_new_n219_), .Y(new_new_n497_));
  NO2        g475(.A(i_8_), .B(i_7_), .Y(new_new_n498_));
  OAI210     g476(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n499_), .B(new_new_n218_), .Y(new_new_n500_));
  AOI220     g478(.A0(new_new_n308_), .A1(new_new_n40_), .B0(new_new_n227_), .B1(new_new_n203_), .Y(new_new_n501_));
  OAI220     g479(.A0(new_new_n501_), .A1(new_new_n178_), .B0(new_new_n500_), .B1(new_new_n235_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n44_), .B(i_10_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(i_6_), .Y(new_new_n504_));
  NA3        g482(.A(new_new_n504_), .B(new_new_n502_), .C(new_new_n498_), .Y(new_new_n505_));
  AOI220     g483(.A0(new_new_n408_), .A1(new_new_n308_), .B0(new_new_n239_), .B1(new_new_n237_), .Y(new_new_n506_));
  OAI220     g484(.A0(new_new_n506_), .A1(new_new_n253_), .B0(new_new_n445_), .B1(new_new_n134_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n507_), .B(new_new_n256_), .Y(new_new_n508_));
  NOi31      g486(.An(new_new_n282_), .B(new_new_n290_), .C(i_4_), .Y(new_new_n509_));
  NA3        g487(.A(new_new_n293_), .B(new_new_n173_), .C(new_new_n96_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n217_), .B(new_new_n44_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n158_), .B(i_5_), .Y(new_new_n512_));
  NA3        g490(.A(new_new_n512_), .B(new_new_n392_), .C(new_new_n302_), .Y(new_new_n513_));
  OAI210     g491(.A0(new_new_n513_), .A1(new_new_n511_), .B0(new_new_n510_), .Y(new_new_n514_));
  OAI210     g492(.A0(new_new_n514_), .A1(new_new_n509_), .B0(new_new_n439_), .Y(new_new_n515_));
  NA3        g493(.A(new_new_n515_), .B(new_new_n508_), .C(new_new_n505_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n286_), .B(new_new_n278_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n517_), .B(new_new_n172_), .Y(new_new_n518_));
  AOI210     g496(.A0(new_new_n347_), .A1(new_new_n46_), .B0(new_new_n351_), .Y(new_new_n519_));
  NA2        g497(.A(i_0_), .B(new_new_n48_), .Y(new_new_n520_));
  NA3        g498(.A(new_new_n496_), .B(new_new_n266_), .C(new_new_n520_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n519_), .B(new_new_n521_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n522_), .B(new_new_n518_), .Y(new_new_n523_));
  NO3        g501(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n225_), .B(new_new_n36_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n397_), .B(i_1_), .Y(new_new_n526_));
  NOi31      g504(.An(new_new_n526_), .B(new_new_n431_), .C(new_new_n72_), .Y(new_new_n527_));
  NOi21      g505(.An(i_10_), .B(i_6_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n530_));
  NA2        g508(.A(new_new_n299_), .B(new_new_n165_), .Y(new_new_n531_));
  AOI220     g509(.A0(new_new_n531_), .A1(new_new_n417_), .B0(new_new_n179_), .B1(new_new_n177_), .Y(new_new_n532_));
  NO2        g510(.A(new_new_n193_), .B(new_new_n37_), .Y(new_new_n533_));
  NOi31      g511(.An(new_new_n147_), .B(new_new_n533_), .C(new_new_n315_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n534_), .B(new_new_n532_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n482_), .B(new_new_n362_), .Y(new_new_n536_));
  INV        g514(.A(new_new_n302_), .Y(new_new_n537_));
  NO2        g515(.A(i_12_), .B(new_new_n85_), .Y(new_new_n538_));
  NA3        g516(.A(new_new_n538_), .B(new_new_n266_), .C(new_new_n520_), .Y(new_new_n539_));
  NA3        g517(.A(new_new_n370_), .B(new_new_n275_), .C(new_new_n213_), .Y(new_new_n540_));
  AOI210     g518(.A0(new_new_n540_), .A1(new_new_n539_), .B0(new_new_n537_), .Y(new_new_n541_));
  NO3        g519(.A(i_4_), .B(new_new_n324_), .C(new_new_n290_), .Y(new_new_n542_));
  OR2        g520(.A(i_2_), .B(i_5_), .Y(new_new_n543_));
  OR2        g521(.A(new_new_n543_), .B(new_new_n394_), .Y(new_new_n544_));
  AOI210     g522(.A0(new_new_n356_), .A1(new_new_n237_), .B0(new_new_n193_), .Y(new_new_n545_));
  AOI210     g523(.A0(new_new_n545_), .A1(new_new_n544_), .B0(new_new_n467_), .Y(new_new_n546_));
  NO4        g524(.A(new_new_n546_), .B(new_new_n542_), .C(new_new_n541_), .D(new_new_n536_), .Y(new_new_n547_));
  NA3        g525(.A(new_new_n547_), .B(new_new_n535_), .C(new_new_n523_), .Y(new_new_n548_));
  NO4        g526(.A(new_new_n548_), .B(new_new_n516_), .C(new_new_n495_), .D(new_new_n477_), .Y(new_new_n549_));
  NA4        g527(.A(new_new_n549_), .B(new_new_n422_), .C(new_new_n335_), .D(new_new_n297_), .Y(ori7));
  NO2        g528(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n552_));
  NA2        g530(.A(new_new_n368_), .B(new_new_n552_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n455_), .B(new_new_n83_), .Y(new_new_n554_));
  NA2        g532(.A(i_11_), .B(new_new_n188_), .Y(new_new_n555_));
  NA2        g533(.A(new_new_n145_), .B(new_new_n555_), .Y(new_new_n556_));
  OAI210     g534(.A0(new_new_n556_), .A1(new_new_n554_), .B0(new_new_n553_), .Y(new_new_n557_));
  NA3        g535(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n229_), .B(i_4_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n559_), .B(i_8_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n105_), .B(new_new_n558_), .Y(new_new_n561_));
  NA2        g539(.A(i_2_), .B(new_new_n85_), .Y(new_new_n562_));
  OAI210     g540(.A0(new_new_n86_), .A1(new_new_n198_), .B0(new_new_n199_), .Y(new_new_n563_));
  NO2        g541(.A(i_7_), .B(new_new_n37_), .Y(new_new_n564_));
  NA2        g542(.A(i_4_), .B(i_8_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n565_), .A1(new_new_n293_), .B0(new_new_n564_), .Y(new_new_n566_));
  OAI220     g544(.A0(new_new_n566_), .A1(new_new_n562_), .B0(new_new_n563_), .B1(i_13_), .Y(new_new_n567_));
  NO4        g545(.A(new_new_n567_), .B(new_new_n561_), .C(new_new_n557_), .D(new_new_n551_), .Y(new_new_n568_));
  AOI210     g546(.A0(new_new_n129_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n569_), .A1(new_new_n229_), .B0(new_new_n162_), .Y(new_new_n570_));
  OR2        g548(.A(i_6_), .B(i_10_), .Y(new_new_n571_));
  OR3        g549(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n572_));
  INV        g550(.A(new_new_n195_), .Y(new_new_n573_));
  OR2        g551(.A(new_new_n570_), .B(new_new_n258_), .Y(new_new_n574_));
  AOI210     g552(.A0(new_new_n574_), .A1(new_new_n568_), .B0(new_new_n62_), .Y(new_new_n575_));
  NOi21      g553(.An(i_11_), .B(i_7_), .Y(new_new_n576_));
  AO210      g554(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n577_), .B(new_new_n576_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n578_), .B(new_new_n203_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n579_), .B(new_new_n62_), .Y(new_new_n580_));
  OR2        g558(.A(new_new_n362_), .B(new_new_n41_), .Y(new_new_n581_));
  NO3        g559(.A(new_new_n248_), .B(new_new_n204_), .C(new_new_n555_), .Y(new_new_n582_));
  OAI210     g560(.A0(new_new_n582_), .A1(new_new_n220_), .B0(new_new_n62_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n395_), .B(new_new_n31_), .Y(new_new_n584_));
  OR2        g562(.A(new_new_n204_), .B(new_new_n108_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n585_), .B(new_new_n584_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n62_), .B(i_9_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n587_), .B(i_4_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(new_new_n586_), .Y(new_new_n589_));
  NO2        g567(.A(i_1_), .B(i_12_), .Y(new_new_n590_));
  NA3        g568(.A(new_new_n590_), .B(new_new_n110_), .C(new_new_n24_), .Y(new_new_n591_));
  BUFFER     g569(.A(new_new_n591_), .Y(new_new_n592_));
  NA4        g570(.A(new_new_n592_), .B(new_new_n589_), .C(new_new_n583_), .D(new_new_n581_), .Y(new_new_n593_));
  OAI210     g571(.A0(new_new_n593_), .A1(new_new_n580_), .B0(i_6_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n229_), .B(new_new_n85_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n595_), .B(i_11_), .Y(new_new_n596_));
  INV        g574(.A(new_new_n432_), .Y(new_new_n597_));
  NA2        g575(.A(new_new_n229_), .B(i_6_), .Y(new_new_n598_));
  NO3        g576(.A(new_new_n571_), .B(new_new_n225_), .C(new_new_n23_), .Y(new_new_n599_));
  AOI210     g577(.A0(i_1_), .A1(new_new_n249_), .B0(new_new_n599_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n600_), .B(new_new_n44_), .Y(new_new_n601_));
  NA3        g579(.A(new_new_n498_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n602_));
  INV        g580(.A(i_2_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n139_), .B(i_9_), .Y(new_new_n604_));
  NO2        g582(.A(new_new_n46_), .B(i_1_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n604_), .B(new_new_n603_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n587_), .B(new_new_n302_), .C(i_6_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n607_), .B(new_new_n23_), .Y(new_new_n608_));
  AOI210     g586(.A0(new_new_n451_), .A1(new_new_n401_), .B0(new_new_n234_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n609_), .B(new_new_n562_), .Y(new_new_n610_));
  NAi21      g588(.An(new_new_n602_), .B(new_new_n91_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n605_), .B(new_new_n257_), .Y(new_new_n612_));
  NO2        g590(.A(i_11_), .B(new_new_n37_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n24_), .Y(new_new_n614_));
  OAI210     g592(.A0(new_new_n614_), .A1(new_new_n612_), .B0(new_new_n611_), .Y(new_new_n615_));
  OR4        g593(.A(new_new_n615_), .B(new_new_n610_), .C(new_new_n608_), .D(new_new_n606_), .Y(new_new_n616_));
  NO3        g594(.A(new_new_n616_), .B(new_new_n601_), .C(new_new_n597_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n229_), .B(new_new_n101_), .Y(new_new_n618_));
  NO2        g596(.A(new_new_n618_), .B(new_new_n576_), .Y(new_new_n619_));
  NA2        g597(.A(new_new_n619_), .B(i_1_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n620_), .B(new_new_n572_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n396_), .B(new_new_n85_), .Y(new_new_n622_));
  NA2        g600(.A(new_new_n621_), .B(new_new_n46_), .Y(new_new_n623_));
  NA2        g601(.A(i_3_), .B(new_new_n188_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n225_), .B(new_new_n44_), .Y(new_new_n625_));
  NO3        g603(.A(new_new_n625_), .B(new_new_n295_), .C(new_new_n230_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n118_), .B(new_new_n37_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n627_), .B(i_6_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n85_), .B(i_9_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n62_), .Y(new_new_n630_));
  NO2        g608(.A(new_new_n630_), .B(new_new_n590_), .Y(new_new_n631_));
  NO4        g609(.A(new_new_n631_), .B(new_new_n628_), .C(new_new_n626_), .D(i_4_), .Y(new_new_n632_));
  NA2        g610(.A(i_1_), .B(i_3_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n433_), .B(new_new_n92_), .Y(new_new_n634_));
  AOI210     g612(.A0(new_new_n625_), .A1(new_new_n528_), .B0(new_new_n634_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n635_), .B(new_new_n633_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n636_), .B(new_new_n632_), .Y(new_new_n637_));
  NA4        g615(.A(new_new_n637_), .B(new_new_n623_), .C(new_new_n617_), .D(new_new_n594_), .Y(new_new_n638_));
  NO3        g616(.A(new_new_n452_), .B(i_3_), .C(i_7_), .Y(new_new_n639_));
  NA2        g617(.A(new_new_n354_), .B(new_new_n353_), .Y(new_new_n640_));
  NA3        g618(.A(new_new_n455_), .B(new_new_n485_), .C(new_new_n46_), .Y(new_new_n641_));
  NA3        g619(.A(new_new_n162_), .B(new_new_n83_), .C(new_new_n85_), .Y(new_new_n642_));
  NA3        g620(.A(new_new_n642_), .B(new_new_n641_), .C(new_new_n640_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n643_), .B(i_1_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n257_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n352_), .B(i_2_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  OAI210     g625(.A0(new_new_n607_), .A1(new_new_n425_), .B0(new_new_n647_), .Y(new_new_n648_));
  INV        g626(.A(new_new_n648_), .Y(new_new_n649_));
  AOI210     g627(.A0(new_new_n649_), .A1(new_new_n644_), .B0(i_13_), .Y(new_new_n650_));
  OR2        g628(.A(i_11_), .B(i_7_), .Y(new_new_n651_));
  NA3        g629(.A(new_new_n651_), .B(new_new_n106_), .C(new_new_n139_), .Y(new_new_n652_));
  AOI220     g630(.A0(new_new_n447_), .A1(new_new_n162_), .B0(new_new_n427_), .B1(new_new_n139_), .Y(new_new_n653_));
  OAI210     g631(.A0(new_new_n653_), .A1(new_new_n44_), .B0(new_new_n652_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n54_), .B(i_12_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n453_), .B(new_new_n24_), .Y(new_new_n656_));
  AOI220     g634(.A0(new_new_n656_), .A1(new_new_n622_), .B0(new_new_n238_), .B1(new_new_n132_), .Y(new_new_n657_));
  OAI220     g635(.A0(new_new_n657_), .A1(new_new_n41_), .B0(new_new_n961_), .B1(new_new_n92_), .Y(new_new_n658_));
  AOI210     g636(.A0(new_new_n654_), .A1(new_new_n317_), .B0(new_new_n658_), .Y(new_new_n659_));
  INV        g637(.A(new_new_n115_), .Y(new_new_n660_));
  AOI220     g638(.A0(new_new_n660_), .A1(new_new_n71_), .B0(new_new_n370_), .B1(new_new_n605_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n661_), .B(new_new_n235_), .Y(new_new_n662_));
  AOI210     g640(.A0(new_new_n425_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n663_));
  NOi31      g641(.An(new_new_n663_), .B(new_new_n554_), .C(new_new_n44_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n128_), .B(i_13_), .Y(new_new_n665_));
  NO2        g643(.A(new_new_n665_), .B(new_new_n645_), .Y(new_new_n666_));
  NO3        g644(.A(new_new_n70_), .B(new_new_n32_), .C(new_new_n101_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n26_), .B(new_new_n188_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n668_), .B(i_7_), .Y(new_new_n669_));
  NO3        g647(.A(new_new_n453_), .B(new_new_n229_), .C(new_new_n85_), .Y(new_new_n670_));
  AOI210     g648(.A0(new_new_n670_), .A1(new_new_n669_), .B0(new_new_n667_), .Y(new_new_n671_));
  AOI220     g649(.A0(new_new_n370_), .A1(new_new_n605_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n672_));
  OAI220     g650(.A0(new_new_n672_), .A1(new_new_n560_), .B0(new_new_n671_), .B1(new_new_n573_), .Y(new_new_n673_));
  NO4        g651(.A(new_new_n673_), .B(new_new_n666_), .C(new_new_n664_), .D(new_new_n662_), .Y(new_new_n674_));
  OR2        g652(.A(i_11_), .B(i_6_), .Y(new_new_n675_));
  NA3        g653(.A(new_new_n559_), .B(new_new_n668_), .C(i_7_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n676_), .B(new_new_n675_), .Y(new_new_n677_));
  NA3        g655(.A(new_new_n395_), .B(new_new_n564_), .C(new_new_n97_), .Y(new_new_n678_));
  NA2        g656(.A(new_new_n596_), .B(i_13_), .Y(new_new_n679_));
  NAi21      g657(.An(i_11_), .B(i_12_), .Y(new_new_n680_));
  NOi41      g658(.An(new_new_n111_), .B(new_new_n680_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n681_));
  NO3        g659(.A(new_new_n453_), .B(new_new_n538_), .C(new_new_n565_), .Y(new_new_n682_));
  AOI220     g660(.A0(new_new_n682_), .A1(new_new_n298_), .B0(new_new_n681_), .B1(new_new_n46_), .Y(new_new_n683_));
  NA3        g661(.A(new_new_n683_), .B(new_new_n679_), .C(new_new_n678_), .Y(new_new_n684_));
  OAI210     g662(.A0(new_new_n684_), .A1(new_new_n677_), .B0(new_new_n62_), .Y(new_new_n685_));
  NO2        g663(.A(i_2_), .B(i_12_), .Y(new_new_n686_));
  NA2        g664(.A(new_new_n351_), .B(new_new_n686_), .Y(new_new_n687_));
  NO2        g665(.A(new_new_n129_), .B(i_2_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n688_), .B(new_new_n590_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n689_), .B(new_new_n687_), .Y(new_new_n690_));
  NA3        g668(.A(new_new_n690_), .B(new_new_n45_), .C(new_new_n219_), .Y(new_new_n691_));
  NA4        g669(.A(new_new_n691_), .B(new_new_n685_), .C(new_new_n674_), .D(new_new_n659_), .Y(new_new_n692_));
  OR4        g670(.A(new_new_n692_), .B(new_new_n650_), .C(new_new_n638_), .D(new_new_n575_), .Y(ori5));
  NA2        g671(.A(new_new_n619_), .B(new_new_n260_), .Y(new_new_n694_));
  AN2        g672(.A(new_new_n24_), .B(i_10_), .Y(new_new_n695_));
  NA3        g673(.A(new_new_n695_), .B(new_new_n686_), .C(new_new_n108_), .Y(new_new_n696_));
  NO2        g674(.A(new_new_n560_), .B(i_11_), .Y(new_new_n697_));
  NA2        g675(.A(new_new_n86_), .B(new_new_n697_), .Y(new_new_n698_));
  NA3        g676(.A(new_new_n698_), .B(new_new_n696_), .C(new_new_n694_), .Y(new_new_n699_));
  NO3        g677(.A(i_11_), .B(new_new_n229_), .C(i_13_), .Y(new_new_n700_));
  NO2        g678(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n701_));
  NA2        g679(.A(i_12_), .B(i_8_), .Y(new_new_n702_));
  OAI210     g680(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n702_), .Y(new_new_n703_));
  INV        g681(.A(new_new_n424_), .Y(new_new_n704_));
  AOI220     g682(.A0(new_new_n302_), .A1(new_new_n530_), .B0(new_new_n703_), .B1(new_new_n701_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n705_), .Y(new_new_n706_));
  NO2        g684(.A(new_new_n706_), .B(new_new_n699_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n171_), .Y(new_new_n708_));
  INV        g686(.A(new_new_n238_), .Y(new_new_n709_));
  OAI210     g687(.A0(new_new_n646_), .A1(new_new_n426_), .B0(new_new_n111_), .Y(new_new_n710_));
  AOI210     g688(.A0(new_new_n710_), .A1(new_new_n709_), .B0(new_new_n708_), .Y(new_new_n711_));
  NO2        g689(.A(new_new_n433_), .B(new_new_n26_), .Y(new_new_n712_));
  NO2        g690(.A(new_new_n712_), .B(new_new_n401_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n713_), .B(i_2_), .Y(new_new_n714_));
  INV        g692(.A(new_new_n714_), .Y(new_new_n715_));
  AOI210     g693(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n397_), .Y(new_new_n716_));
  AOI210     g694(.A0(new_new_n716_), .A1(new_new_n715_), .B0(new_new_n711_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n186_), .B(new_new_n126_), .Y(new_new_n718_));
  OAI210     g696(.A0(new_new_n718_), .A1(new_new_n701_), .B0(i_2_), .Y(new_new_n719_));
  INV        g697(.A(new_new_n172_), .Y(new_new_n720_));
  NO3        g698(.A(new_new_n577_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n721_));
  AOI210     g699(.A0(new_new_n720_), .A1(new_new_n86_), .B0(new_new_n721_), .Y(new_new_n722_));
  AOI210     g700(.A0(new_new_n722_), .A1(new_new_n719_), .B0(new_new_n188_), .Y(new_new_n723_));
  OA210      g701(.A0(new_new_n578_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n195_), .B(new_new_n198_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n152_), .B(new_new_n555_), .Y(new_new_n726_));
  AOI210     g704(.A0(new_new_n726_), .A1(new_new_n725_), .B0(new_new_n356_), .Y(new_new_n727_));
  AOI210     g705(.A0(new_new_n204_), .A1(new_new_n149_), .B0(new_new_n485_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n728_), .B(new_new_n401_), .Y(new_new_n729_));
  NO2        g707(.A(new_new_n102_), .B(new_new_n44_), .Y(new_new_n730_));
  INV        g708(.A(new_new_n291_), .Y(new_new_n731_));
  NA4        g709(.A(new_new_n731_), .B(new_new_n293_), .C(new_new_n125_), .D(new_new_n42_), .Y(new_new_n732_));
  OAI210     g710(.A0(new_new_n732_), .A1(new_new_n730_), .B0(new_new_n729_), .Y(new_new_n733_));
  NO4        g711(.A(new_new_n733_), .B(new_new_n727_), .C(new_new_n724_), .D(new_new_n723_), .Y(new_new_n734_));
  NA2        g712(.A(new_new_n530_), .B(new_new_n28_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n700_), .B(new_new_n267_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n736_), .B(new_new_n735_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n61_), .B(i_12_), .Y(new_new_n738_));
  NO2        g716(.A(new_new_n738_), .B(new_new_n127_), .Y(new_new_n739_));
  NO2        g717(.A(new_new_n739_), .B(new_new_n555_), .Y(new_new_n740_));
  AOI220     g718(.A0(new_new_n740_), .A1(new_new_n36_), .B0(new_new_n737_), .B1(new_new_n46_), .Y(new_new_n741_));
  NA4        g719(.A(new_new_n741_), .B(new_new_n734_), .C(new_new_n717_), .D(new_new_n707_), .Y(ori6));
  NO3        g720(.A(i_9_), .B(new_new_n294_), .C(i_1_), .Y(new_new_n743_));
  NO2        g721(.A(new_new_n181_), .B(new_new_n140_), .Y(new_new_n744_));
  OAI210     g722(.A0(new_new_n744_), .A1(new_new_n743_), .B0(new_new_n688_), .Y(new_new_n745_));
  NO2        g723(.A(new_new_n216_), .B(new_new_n459_), .Y(new_new_n746_));
  NO2        g724(.A(i_11_), .B(i_9_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n312_), .Y(new_new_n748_));
  AO210      g726(.A0(new_new_n748_), .A1(new_new_n745_), .B0(i_12_), .Y(new_new_n749_));
  NA2        g727(.A(new_new_n538_), .B(new_new_n62_), .Y(new_new_n750_));
  INV        g728(.A(new_new_n750_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n192_), .Y(new_new_n752_));
  AOI220     g730(.A0(new_new_n752_), .A1(new_new_n747_), .B0(new_new_n751_), .B1(new_new_n72_), .Y(new_new_n753_));
  INV        g731(.A(new_new_n311_), .Y(new_new_n754_));
  NA2        g732(.A(new_new_n74_), .B(new_new_n132_), .Y(new_new_n755_));
  INV        g733(.A(new_new_n125_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n756_), .B(new_new_n46_), .Y(new_new_n757_));
  AOI210     g735(.A0(new_new_n757_), .A1(new_new_n755_), .B0(new_new_n754_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n242_), .B(i_9_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n759_), .B(new_new_n738_), .Y(new_new_n760_));
  AOI210     g738(.A0(new_new_n760_), .A1(new_new_n483_), .B0(new_new_n181_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n32_), .B(i_11_), .Y(new_new_n762_));
  NAi32      g740(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n763_));
  NO2        g741(.A(new_new_n675_), .B(new_new_n763_), .Y(new_new_n764_));
  OAI210     g742(.A0(new_new_n639_), .A1(new_new_n525_), .B0(new_new_n524_), .Y(new_new_n765_));
  NAi21      g743(.An(new_new_n764_), .B(new_new_n765_), .Y(new_new_n766_));
  OR3        g744(.A(new_new_n766_), .B(new_new_n761_), .C(new_new_n758_), .Y(new_new_n767_));
  NO2        g745(.A(new_new_n651_), .B(i_2_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n769_));
  NO2        g747(.A(new_new_n769_), .B(new_new_n394_), .Y(new_new_n770_));
  NA2        g748(.A(new_new_n770_), .B(new_new_n768_), .Y(new_new_n771_));
  AO220      g749(.A0(new_new_n340_), .A1(new_new_n330_), .B0(new_new_n382_), .B1(new_new_n555_), .Y(new_new_n772_));
  NA3        g750(.A(new_new_n772_), .B(new_new_n245_), .C(i_7_), .Y(new_new_n773_));
  OR2        g751(.A(new_new_n578_), .B(new_new_n426_), .Y(new_new_n774_));
  NA3        g752(.A(new_new_n774_), .B(new_new_n148_), .C(new_new_n68_), .Y(new_new_n775_));
  AO210      g753(.A0(new_new_n466_), .A1(new_new_n704_), .B0(new_new_n36_), .Y(new_new_n776_));
  NA4        g754(.A(new_new_n776_), .B(new_new_n775_), .C(new_new_n773_), .D(new_new_n771_), .Y(new_new_n777_));
  NO2        g755(.A(new_new_n595_), .B(i_11_), .Y(new_new_n778_));
  AOI220     g756(.A0(new_new_n778_), .A1(new_new_n524_), .B0(new_new_n746_), .B1(new_new_n669_), .Y(new_new_n779_));
  NA3        g757(.A(new_new_n356_), .B(new_new_n231_), .C(new_new_n148_), .Y(new_new_n780_));
  NA2        g758(.A(new_new_n382_), .B(new_new_n69_), .Y(new_new_n781_));
  NA4        g759(.A(new_new_n781_), .B(new_new_n780_), .C(new_new_n779_), .D(new_new_n563_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n426_), .B(new_new_n424_), .Y(new_new_n783_));
  NO2        g761(.A(new_new_n571_), .B(new_new_n102_), .Y(new_new_n784_));
  OAI210     g762(.A0(new_new_n784_), .A1(new_new_n112_), .B0(new_new_n393_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n237_), .B(new_new_n46_), .Y(new_new_n786_));
  INV        g764(.A(new_new_n544_), .Y(new_new_n787_));
  NA3        g765(.A(new_new_n787_), .B(new_new_n311_), .C(i_7_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n788_), .B(new_new_n785_), .C(new_new_n783_), .Y(new_new_n789_));
  NO4        g767(.A(new_new_n789_), .B(new_new_n782_), .C(new_new_n777_), .D(new_new_n767_), .Y(new_new_n790_));
  NA4        g768(.A(new_new_n790_), .B(new_new_n753_), .C(new_new_n749_), .D(new_new_n364_), .Y(ori3));
  NA2        g769(.A(i_12_), .B(i_10_), .Y(new_new_n792_));
  NO2        g770(.A(i_11_), .B(new_new_n229_), .Y(new_new_n793_));
  NA2        g771(.A(new_new_n780_), .B(new_new_n563_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n794_), .B(new_new_n40_), .Y(new_new_n795_));
  NOi21      g773(.An(new_new_n96_), .B(new_new_n713_), .Y(new_new_n796_));
  NO3        g774(.A(new_new_n585_), .B(new_new_n433_), .C(new_new_n132_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n395_), .B(new_new_n45_), .Y(new_new_n798_));
  AN2        g776(.A(new_new_n431_), .B(new_new_n55_), .Y(new_new_n799_));
  NO3        g777(.A(new_new_n799_), .B(new_new_n797_), .C(new_new_n796_), .Y(new_new_n800_));
  AOI210     g778(.A0(new_new_n800_), .A1(new_new_n795_), .B0(new_new_n48_), .Y(new_new_n801_));
  NO4        g779(.A(new_new_n360_), .B(new_new_n367_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n181_), .B(new_new_n528_), .Y(new_new_n803_));
  NOi21      g781(.An(new_new_n803_), .B(new_new_n802_), .Y(new_new_n804_));
  NA2        g782(.A(new_new_n663_), .B(new_new_n629_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n318_), .B(new_new_n419_), .Y(new_new_n806_));
  OAI220     g784(.A0(new_new_n806_), .A1(new_new_n805_), .B0(new_new_n804_), .B1(new_new_n62_), .Y(new_new_n807_));
  NOi21      g785(.An(i_5_), .B(i_9_), .Y(new_new_n808_));
  NA2        g786(.A(new_new_n808_), .B(new_new_n423_), .Y(new_new_n809_));
  BUFFER     g787(.A(new_new_n257_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n810_), .B(new_new_n451_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n811_), .B(new_new_n809_), .Y(new_new_n812_));
  NO3        g790(.A(new_new_n812_), .B(new_new_n807_), .C(new_new_n801_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n181_), .B(new_new_n24_), .Y(new_new_n814_));
  NO2        g792(.A(new_new_n627_), .B(new_new_n552_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n815_), .B(new_new_n814_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n298_), .B(new_new_n130_), .Y(new_new_n817_));
  NAi21      g795(.An(new_new_n163_), .B(new_new_n419_), .Y(new_new_n818_));
  OAI220     g796(.A0(new_new_n818_), .A1(new_new_n786_), .B0(new_new_n817_), .B1(new_new_n387_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(new_new_n816_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n529_), .B(i_0_), .Y(new_new_n821_));
  NO3        g799(.A(new_new_n821_), .B(new_new_n369_), .C(new_new_n86_), .Y(new_new_n822_));
  NO4        g800(.A(new_new_n543_), .B(new_new_n210_), .C(new_new_n397_), .D(new_new_n394_), .Y(new_new_n823_));
  AOI210     g801(.A0(new_new_n823_), .A1(i_11_), .B0(new_new_n822_), .Y(new_new_n824_));
  INV        g802(.A(new_new_n450_), .Y(new_new_n825_));
  AN2        g803(.A(new_new_n96_), .B(new_new_n236_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n700_), .B(new_new_n312_), .Y(new_new_n827_));
  AOI210     g805(.A0(new_new_n455_), .A1(new_new_n86_), .B0(new_new_n57_), .Y(new_new_n828_));
  OAI220     g806(.A0(new_new_n828_), .A1(new_new_n827_), .B0(new_new_n614_), .B1(new_new_n500_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n244_), .B(new_new_n154_), .Y(new_new_n830_));
  NA2        g808(.A(i_0_), .B(i_10_), .Y(new_new_n831_));
  INV        g809(.A(new_new_n503_), .Y(new_new_n832_));
  NO4        g810(.A(new_new_n115_), .B(new_new_n57_), .C(new_new_n624_), .D(i_5_), .Y(new_new_n833_));
  AO220      g811(.A0(new_new_n833_), .A1(new_new_n832_), .B0(new_new_n830_), .B1(i_6_), .Y(new_new_n834_));
  NO3        g812(.A(new_new_n834_), .B(new_new_n829_), .C(new_new_n826_), .Y(new_new_n835_));
  NA3        g813(.A(new_new_n835_), .B(new_new_n824_), .C(new_new_n820_), .Y(new_new_n836_));
  NA2        g814(.A(i_11_), .B(i_9_), .Y(new_new_n837_));
  NA2        g815(.A(new_new_n379_), .B(new_new_n175_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n161_), .Y(new_new_n839_));
  NO2        g817(.A(new_new_n837_), .B(new_new_n72_), .Y(new_new_n840_));
  NO2        g818(.A(new_new_n174_), .B(i_0_), .Y(new_new_n841_));
  INV        g819(.A(new_new_n841_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n450_), .B(new_new_n223_), .Y(new_new_n843_));
  NO2        g821(.A(new_new_n843_), .B(new_new_n842_), .Y(new_new_n844_));
  NO2        g822(.A(new_new_n844_), .B(new_new_n839_), .Y(new_new_n845_));
  NA2        g823(.A(new_new_n613_), .B(new_new_n122_), .Y(new_new_n846_));
  NO2        g824(.A(i_6_), .B(new_new_n846_), .Y(new_new_n847_));
  AOI210     g825(.A0(new_new_n425_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n848_));
  NA2        g826(.A(new_new_n171_), .B(new_new_n103_), .Y(new_new_n849_));
  NOi32      g827(.An(new_new_n848_), .Bn(new_new_n184_), .C(new_new_n849_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n564_), .B(new_new_n312_), .Y(new_new_n851_));
  NO2        g829(.A(new_new_n851_), .B(new_new_n798_), .Y(new_new_n852_));
  NO3        g830(.A(new_new_n852_), .B(new_new_n850_), .C(new_new_n847_), .Y(new_new_n853_));
  INV        g831(.A(new_new_n303_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n853_), .B(new_new_n845_), .Y(new_new_n855_));
  NO2        g833(.A(new_new_n792_), .B(new_new_n302_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n856_), .B(new_new_n840_), .Y(new_new_n857_));
  NA3        g835(.A(new_new_n449_), .B(new_new_n395_), .C(new_new_n45_), .Y(new_new_n858_));
  OAI210     g836(.A0(new_new_n818_), .A1(new_new_n825_), .B0(new_new_n858_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n840_), .B(new_new_n293_), .Y(new_new_n860_));
  NA2        g838(.A(new_new_n183_), .B(new_new_n860_), .Y(new_new_n861_));
  AOI220     g839(.A0(new_new_n861_), .A1(new_new_n450_), .B0(new_new_n859_), .B1(new_new_n72_), .Y(new_new_n862_));
  NA3        g840(.A(new_new_n769_), .B(new_new_n366_), .C(new_new_n595_), .Y(new_new_n863_));
  NA2        g841(.A(new_new_n92_), .B(new_new_n44_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n74_), .B(new_new_n702_), .Y(new_new_n865_));
  AOI220     g843(.A0(new_new_n865_), .A1(new_new_n864_), .B0(new_new_n173_), .B1(new_new_n552_), .Y(new_new_n866_));
  AOI210     g844(.A0(new_new_n866_), .A1(new_new_n863_), .B0(new_new_n47_), .Y(new_new_n867_));
  NO3        g845(.A(new_new_n543_), .B(new_new_n338_), .C(new_new_n24_), .Y(new_new_n868_));
  AOI210     g846(.A0(new_new_n656_), .A1(new_new_n512_), .B0(new_new_n868_), .Y(new_new_n869_));
  NAi21      g847(.An(i_9_), .B(i_5_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n869_), .B(new_new_n172_), .Y(new_new_n871_));
  NO3        g849(.A(new_new_n871_), .B(new_new_n867_), .C(new_new_n487_), .Y(new_new_n872_));
  NA3        g850(.A(new_new_n872_), .B(new_new_n862_), .C(new_new_n857_), .Y(new_new_n873_));
  NO3        g851(.A(new_new_n873_), .B(new_new_n855_), .C(new_new_n836_), .Y(new_new_n874_));
  NO2        g852(.A(i_0_), .B(new_new_n680_), .Y(new_new_n875_));
  NA2        g853(.A(new_new_n72_), .B(new_new_n44_), .Y(new_new_n876_));
  AOI210     g854(.A0(new_new_n750_), .A1(new_new_n640_), .B0(new_new_n849_), .Y(new_new_n877_));
  INV        g855(.A(new_new_n877_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n765_), .B(new_new_n388_), .Y(new_new_n879_));
  NA2        g857(.A(new_new_n793_), .B(i_9_), .Y(new_new_n880_));
  NO2        g858(.A(new_new_n470_), .B(new_new_n880_), .Y(new_new_n881_));
  NA2        g859(.A(new_new_n237_), .B(new_new_n222_), .Y(new_new_n882_));
  AOI210     g860(.A0(new_new_n882_), .A1(new_new_n821_), .B0(new_new_n154_), .Y(new_new_n883_));
  NO3        g861(.A(new_new_n883_), .B(new_new_n881_), .C(new_new_n879_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n884_), .B(new_new_n878_), .Y(new_new_n885_));
  NO3        g863(.A(new_new_n831_), .B(new_new_n808_), .C(new_new_n186_), .Y(new_new_n886_));
  AOI220     g864(.A0(new_new_n886_), .A1(i_11_), .B0(new_new_n527_), .B1(new_new_n74_), .Y(new_new_n887_));
  NO3        g865(.A(new_new_n205_), .B(new_new_n367_), .C(i_0_), .Y(new_new_n888_));
  OAI210     g866(.A0(new_new_n888_), .A1(new_new_n75_), .B0(i_13_), .Y(new_new_n889_));
  INV        g867(.A(new_new_n213_), .Y(new_new_n890_));
  OAI220     g868(.A0(new_new_n497_), .A1(new_new_n140_), .B0(new_new_n598_), .B1(new_new_n573_), .Y(new_new_n891_));
  NA3        g869(.A(new_new_n891_), .B(i_7_), .C(new_new_n890_), .Y(new_new_n892_));
  NA3        g870(.A(new_new_n892_), .B(new_new_n889_), .C(new_new_n887_), .Y(new_new_n893_));
  NO2        g871(.A(new_new_n235_), .B(new_new_n92_), .Y(new_new_n894_));
  AOI210     g872(.A0(new_new_n894_), .A1(new_new_n875_), .B0(new_new_n109_), .Y(new_new_n895_));
  OR2        g873(.A(new_new_n895_), .B(i_5_), .Y(new_new_n896_));
  INV        g874(.A(new_new_n510_), .Y(new_new_n897_));
  NO3        g875(.A(new_new_n798_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n465_), .B(new_new_n458_), .Y(new_new_n899_));
  NO3        g877(.A(new_new_n899_), .B(new_new_n898_), .C(new_new_n897_), .Y(new_new_n900_));
  NA3        g878(.A(new_new_n374_), .B(new_new_n171_), .C(new_new_n170_), .Y(new_new_n901_));
  INV        g879(.A(new_new_n901_), .Y(new_new_n902_));
  NA3        g880(.A(new_new_n374_), .B(new_new_n319_), .C(new_new_n217_), .Y(new_new_n903_));
  INV        g881(.A(new_new_n903_), .Y(new_new_n904_));
  NOi31      g882(.An(new_new_n373_), .B(new_new_n876_), .C(new_new_n232_), .Y(new_new_n905_));
  NO3        g883(.A(new_new_n837_), .B(new_new_n213_), .C(new_new_n186_), .Y(new_new_n906_));
  NO4        g884(.A(new_new_n906_), .B(new_new_n905_), .C(new_new_n904_), .D(new_new_n902_), .Y(new_new_n907_));
  NA3        g885(.A(new_new_n907_), .B(new_new_n900_), .C(new_new_n896_), .Y(new_new_n908_));
  NO2        g886(.A(new_new_n85_), .B(i_5_), .Y(new_new_n909_));
  NA3        g887(.A(new_new_n793_), .B(new_new_n110_), .C(new_new_n125_), .Y(new_new_n910_));
  INV        g888(.A(new_new_n910_), .Y(new_new_n911_));
  NA2        g889(.A(new_new_n911_), .B(new_new_n909_), .Y(new_new_n912_));
  NAi21      g890(.An(new_new_n234_), .B(new_new_n235_), .Y(new_new_n913_));
  NO4        g891(.A(new_new_n232_), .B(new_new_n205_), .C(i_0_), .D(i_12_), .Y(new_new_n914_));
  NA2        g892(.A(new_new_n914_), .B(new_new_n913_), .Y(new_new_n915_));
  AN2        g893(.A(new_new_n831_), .B(new_new_n154_), .Y(new_new_n916_));
  NO4        g894(.A(new_new_n916_), .B(i_12_), .C(new_new_n602_), .D(new_new_n132_), .Y(new_new_n917_));
  NA2        g895(.A(new_new_n917_), .B(new_new_n213_), .Y(new_new_n918_));
  NA3        g896(.A(new_new_n98_), .B(new_new_n528_), .C(i_11_), .Y(new_new_n919_));
  NO2        g897(.A(new_new_n919_), .B(new_new_n156_), .Y(new_new_n920_));
  INV        g898(.A(new_new_n920_), .Y(new_new_n921_));
  NA4        g899(.A(new_new_n921_), .B(new_new_n918_), .C(new_new_n915_), .D(new_new_n912_), .Y(new_new_n922_));
  NO4        g900(.A(new_new_n922_), .B(new_new_n908_), .C(new_new_n893_), .D(new_new_n885_), .Y(new_new_n923_));
  OAI210     g901(.A0(new_new_n768_), .A1(new_new_n762_), .B0(new_new_n37_), .Y(new_new_n924_));
  NA3        g902(.A(new_new_n848_), .B(new_new_n351_), .C(i_5_), .Y(new_new_n925_));
  NA3        g903(.A(new_new_n925_), .B(new_new_n924_), .C(new_new_n570_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n926_), .B(new_new_n203_), .Y(new_new_n927_));
  AN2        g905(.A(new_new_n651_), .B(new_new_n352_), .Y(new_new_n928_));
  NA2        g906(.A(new_new_n182_), .B(new_new_n184_), .Y(new_new_n929_));
  AO210      g907(.A0(new_new_n928_), .A1(new_new_n33_), .B0(new_new_n929_), .Y(new_new_n930_));
  INV        g908(.A(new_new_n930_), .Y(new_new_n931_));
  INV        g909(.A(new_new_n823_), .Y(new_new_n932_));
  OAI210     g910(.A0(new_new_n919_), .A1(new_new_n149_), .B0(new_new_n932_), .Y(new_new_n933_));
  AOI210     g911(.A0(new_new_n931_), .A1(new_new_n48_), .B0(new_new_n933_), .Y(new_new_n934_));
  AOI210     g912(.A0(new_new_n934_), .A1(new_new_n927_), .B0(new_new_n72_), .Y(new_new_n935_));
  INV        g913(.A(new_new_n363_), .Y(new_new_n936_));
  NO2        g914(.A(new_new_n936_), .B(new_new_n708_), .Y(new_new_n937_));
  OAI210     g915(.A0(new_new_n79_), .A1(new_new_n54_), .B0(new_new_n108_), .Y(new_new_n938_));
  NA2        g916(.A(new_new_n938_), .B(new_new_n75_), .Y(new_new_n939_));
  NO2        g917(.A(new_new_n939_), .B(new_new_n633_), .Y(new_new_n940_));
  INV        g918(.A(new_new_n940_), .Y(new_new_n941_));
  OAI210     g919(.A0(new_new_n259_), .A1(new_new_n159_), .B0(new_new_n86_), .Y(new_new_n942_));
  NA3        g920(.A(new_new_n712_), .B(new_new_n282_), .C(new_new_n79_), .Y(new_new_n943_));
  AOI210     g921(.A0(new_new_n943_), .A1(new_new_n942_), .B0(i_11_), .Y(new_new_n944_));
  OAI210     g922(.A0(new_new_n962_), .A1(new_new_n848_), .B0(new_new_n203_), .Y(new_new_n945_));
  NA2        g923(.A(new_new_n165_), .B(i_5_), .Y(new_new_n946_));
  NO2        g924(.A(new_new_n945_), .B(new_new_n946_), .Y(new_new_n947_));
  NO3        g925(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n948_));
  OAI210     g926(.A0(new_new_n854_), .A1(new_new_n294_), .B0(new_new_n948_), .Y(new_new_n949_));
  NO2        g927(.A(new_new_n949_), .B(new_new_n680_), .Y(new_new_n950_));
  NO4        g928(.A(new_new_n870_), .B(new_new_n452_), .C(new_new_n243_), .D(new_new_n242_), .Y(new_new_n951_));
  INV        g929(.A(new_new_n951_), .Y(new_new_n952_));
  INV        g930(.A(new_new_n344_), .Y(new_new_n953_));
  AOI210     g931(.A0(new_new_n953_), .A1(new_new_n952_), .B0(new_new_n41_), .Y(new_new_n954_));
  NO4        g932(.A(new_new_n954_), .B(new_new_n950_), .C(new_new_n947_), .D(new_new_n944_), .Y(new_new_n955_));
  OAI210     g933(.A0(new_new_n941_), .A1(i_4_), .B0(new_new_n955_), .Y(new_new_n956_));
  NO3        g934(.A(new_new_n956_), .B(new_new_n937_), .C(new_new_n935_), .Y(new_new_n957_));
  NA4        g935(.A(new_new_n957_), .B(new_new_n923_), .C(new_new_n874_), .D(new_new_n813_), .Y(ori4));
  INV        g936(.A(new_new_n655_), .Y(new_new_n961_));
  INV        g937(.A(i_12_), .Y(new_new_n962_));
endmodule


