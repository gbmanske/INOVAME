//Benchmark atmr_misex3_1774_0.0313

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1375_, ori_ori_n1379_, ori_ori_n1380_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1499_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1511_, men_men_n1512_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(g), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(g), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(g), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO2        o0025(.A(ori_ori_n53_), .B(ori_ori_n39_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NA2        o0031(.A(g), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NAi21      o0032(.An(i), .B(h), .Y(ori_ori_n61_));
  NAi31      o0033(.An(i), .B(l), .C(j), .Y(ori_ori_n62_));
  OAI220     o0034(.A0(ori_ori_n62_), .A1(ori_ori_n49_), .B0(ori_ori_n61_), .B1(ori_ori_n44_), .Y(ori_ori_n63_));
  NAi31      o0035(.An(ori_ori_n60_), .B(ori_ori_n63_), .C(ori_ori_n58_), .Y(ori_ori_n64_));
  NAi41      o0036(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n65_));
  NA2        o0037(.A(g), .B(f), .Y(ori_ori_n66_));
  NO2        o0038(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NAi21      o0039(.An(i), .B(j), .Y(ori_ori_n68_));
  NAi32      o0040(.An(n), .Bn(k), .C(m), .Y(ori_ori_n69_));
  NAi31      o0041(.An(l), .B(m), .C(k), .Y(ori_ori_n70_));
  NAi41      o0042(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n71_));
  INV        o0043(.A(m), .Y(ori_ori_n72_));
  NOi21      o0044(.An(k), .B(l), .Y(ori_ori_n73_));
  NA2        o0045(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  AN4        o0046(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n75_));
  NOi31      o0047(.An(h), .B(g), .C(f), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  NAi32      o0049(.An(m), .Bn(k), .C(j), .Y(ori_ori_n78_));
  NOi32      o0050(.An(h), .Bn(g), .C(f), .Y(ori_ori_n79_));
  NA2        o0051(.A(ori_ori_n79_), .B(ori_ori_n75_), .Y(ori_ori_n80_));
  OR2        o0052(.A(ori_ori_n80_), .B(ori_ori_n78_), .Y(ori_ori_n81_));
  NA2        o0053(.A(ori_ori_n81_), .B(ori_ori_n64_), .Y(ori_ori_n82_));
  INV        o0054(.A(n), .Y(ori_ori_n83_));
  NOi32      o0055(.An(e), .Bn(b), .C(d), .Y(ori_ori_n84_));
  NA2        o0056(.A(ori_ori_n84_), .B(ori_ori_n83_), .Y(ori_ori_n85_));
  INV        o0057(.A(j), .Y(ori_ori_n86_));
  AN3        o0058(.A(m), .B(k), .C(i), .Y(ori_ori_n87_));
  NA3        o0059(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(g), .Y(ori_ori_n88_));
  NO2        o0060(.A(ori_ori_n88_), .B(f), .Y(ori_ori_n89_));
  NAi32      o0061(.An(g), .Bn(f), .C(h), .Y(ori_ori_n90_));
  NAi31      o0062(.An(j), .B(m), .C(l), .Y(ori_ori_n91_));
  NO2        o0063(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n92_));
  NA2        o0064(.A(m), .B(l), .Y(ori_ori_n93_));
  NAi31      o0065(.An(k), .B(j), .C(g), .Y(ori_ori_n94_));
  NO3        o0066(.A(ori_ori_n94_), .B(ori_ori_n93_), .C(f), .Y(ori_ori_n95_));
  AN2        o0067(.A(j), .B(g), .Y(ori_ori_n96_));
  NOi32      o0068(.An(m), .Bn(l), .C(i), .Y(ori_ori_n97_));
  NOi21      o0069(.An(g), .B(i), .Y(ori_ori_n98_));
  NOi32      o0070(.An(m), .Bn(j), .C(k), .Y(ori_ori_n99_));
  AOI220     o0071(.A0(ori_ori_n99_), .A1(ori_ori_n98_), .B0(ori_ori_n97_), .B1(ori_ori_n96_), .Y(ori_ori_n100_));
  NO2        o0072(.A(ori_ori_n100_), .B(f), .Y(ori_ori_n101_));
  NO3        o0073(.A(ori_ori_n101_), .B(ori_ori_n92_), .C(ori_ori_n89_), .Y(ori_ori_n102_));
  NAi41      o0074(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n103_));
  AN2        o0075(.A(e), .B(b), .Y(ori_ori_n104_));
  NOi31      o0076(.An(c), .B(h), .C(f), .Y(ori_ori_n105_));
  NA2        o0077(.A(ori_ori_n105_), .B(ori_ori_n104_), .Y(ori_ori_n106_));
  NO2        o0078(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n107_));
  NOi21      o0079(.An(g), .B(f), .Y(ori_ori_n108_));
  NOi21      o0080(.An(i), .B(h), .Y(ori_ori_n109_));
  NA3        o0081(.A(ori_ori_n109_), .B(ori_ori_n108_), .C(ori_ori_n36_), .Y(ori_ori_n110_));
  INV        o0082(.A(a), .Y(ori_ori_n111_));
  NA2        o0083(.A(ori_ori_n104_), .B(ori_ori_n111_), .Y(ori_ori_n112_));
  INV        o0084(.A(l), .Y(ori_ori_n113_));
  NOi21      o0085(.An(m), .B(n), .Y(ori_ori_n114_));
  AN2        o0086(.A(k), .B(h), .Y(ori_ori_n115_));
  NO2        o0087(.A(ori_ori_n110_), .B(ori_ori_n85_), .Y(ori_ori_n116_));
  INV        o0088(.A(b), .Y(ori_ori_n117_));
  NA2        o0089(.A(l), .B(j), .Y(ori_ori_n118_));
  AN2        o0090(.A(k), .B(i), .Y(ori_ori_n119_));
  NA2        o0091(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NA2        o0092(.A(g), .B(e), .Y(ori_ori_n121_));
  NOi32      o0093(.An(c), .Bn(a), .C(d), .Y(ori_ori_n122_));
  NA2        o0094(.A(ori_ori_n122_), .B(ori_ori_n114_), .Y(ori_ori_n123_));
  NO2        o0095(.A(ori_ori_n116_), .B(ori_ori_n107_), .Y(ori_ori_n124_));
  OAI210     o0096(.A0(ori_ori_n102_), .A1(ori_ori_n85_), .B0(ori_ori_n124_), .Y(ori_ori_n125_));
  NOi31      o0097(.An(k), .B(m), .C(j), .Y(ori_ori_n126_));
  NA3        o0098(.A(ori_ori_n126_), .B(ori_ori_n76_), .C(ori_ori_n75_), .Y(ori_ori_n127_));
  NOi31      o0099(.An(k), .B(m), .C(i), .Y(ori_ori_n128_));
  NA3        o0100(.A(ori_ori_n128_), .B(ori_ori_n79_), .C(ori_ori_n75_), .Y(ori_ori_n129_));
  NA2        o0101(.A(ori_ori_n129_), .B(ori_ori_n127_), .Y(ori_ori_n130_));
  NOi32      o0102(.An(f), .Bn(b), .C(e), .Y(ori_ori_n131_));
  NAi21      o0103(.An(g), .B(h), .Y(ori_ori_n132_));
  NAi21      o0104(.An(m), .B(n), .Y(ori_ori_n133_));
  NAi21      o0105(.An(j), .B(k), .Y(ori_ori_n134_));
  NO3        o0106(.A(ori_ori_n134_), .B(ori_ori_n133_), .C(ori_ori_n132_), .Y(ori_ori_n135_));
  NAi41      o0107(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n136_));
  NAi31      o0108(.An(j), .B(k), .C(h), .Y(ori_ori_n137_));
  NO3        o0109(.A(ori_ori_n137_), .B(ori_ori_n136_), .C(ori_ori_n133_), .Y(ori_ori_n138_));
  AOI210     o0110(.A0(ori_ori_n135_), .A1(ori_ori_n131_), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  NO2        o0111(.A(k), .B(j), .Y(ori_ori_n140_));
  NO2        o0112(.A(ori_ori_n140_), .B(ori_ori_n133_), .Y(ori_ori_n141_));
  AN2        o0113(.A(k), .B(j), .Y(ori_ori_n142_));
  NAi21      o0114(.An(c), .B(b), .Y(ori_ori_n143_));
  NA2        o0115(.A(f), .B(d), .Y(ori_ori_n144_));
  NO4        o0116(.A(ori_ori_n144_), .B(ori_ori_n143_), .C(ori_ori_n142_), .D(ori_ori_n132_), .Y(ori_ori_n145_));
  NA2        o0117(.A(h), .B(c), .Y(ori_ori_n146_));
  NAi31      o0118(.An(f), .B(e), .C(b), .Y(ori_ori_n147_));
  NA2        o0119(.A(ori_ori_n145_), .B(ori_ori_n141_), .Y(ori_ori_n148_));
  NA2        o0120(.A(d), .B(b), .Y(ori_ori_n149_));
  NAi21      o0121(.An(e), .B(f), .Y(ori_ori_n150_));
  NO2        o0122(.A(ori_ori_n150_), .B(ori_ori_n149_), .Y(ori_ori_n151_));
  NA2        o0123(.A(b), .B(a), .Y(ori_ori_n152_));
  NAi21      o0124(.An(e), .B(g), .Y(ori_ori_n153_));
  NAi21      o0125(.An(c), .B(d), .Y(ori_ori_n154_));
  NAi31      o0126(.An(l), .B(k), .C(h), .Y(ori_ori_n155_));
  NO2        o0127(.A(ori_ori_n133_), .B(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o0128(.A(ori_ori_n156_), .B(ori_ori_n151_), .Y(ori_ori_n157_));
  NAi41      o0129(.An(ori_ori_n130_), .B(ori_ori_n157_), .C(ori_ori_n148_), .D(ori_ori_n139_), .Y(ori_ori_n158_));
  NAi31      o0130(.An(e), .B(f), .C(b), .Y(ori_ori_n159_));
  NOi21      o0131(.An(g), .B(d), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NOi21      o0133(.An(h), .B(i), .Y(ori_ori_n162_));
  NOi21      o0134(.An(k), .B(m), .Y(ori_ori_n163_));
  NA3        o0135(.A(ori_ori_n163_), .B(ori_ori_n162_), .C(n), .Y(ori_ori_n164_));
  NOi21      o0136(.An(ori_ori_n161_), .B(ori_ori_n164_), .Y(ori_ori_n165_));
  NOi21      o0137(.An(h), .B(g), .Y(ori_ori_n166_));
  NO2        o0138(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n167_));
  NAi31      o0139(.An(l), .B(j), .C(h), .Y(ori_ori_n168_));
  NO2        o0140(.A(ori_ori_n168_), .B(ori_ori_n49_), .Y(ori_ori_n169_));
  NA2        o0141(.A(ori_ori_n169_), .B(ori_ori_n67_), .Y(ori_ori_n170_));
  NOi32      o0142(.An(n), .Bn(k), .C(m), .Y(ori_ori_n171_));
  NA2        o0143(.A(l), .B(i), .Y(ori_ori_n172_));
  INV        o0144(.A(ori_ori_n170_), .Y(ori_ori_n173_));
  NAi31      o0145(.An(d), .B(f), .C(c), .Y(ori_ori_n174_));
  NAi31      o0146(.An(e), .B(f), .C(c), .Y(ori_ori_n175_));
  NA2        o0147(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  NA2        o0148(.A(j), .B(h), .Y(ori_ori_n177_));
  OR3        o0149(.A(n), .B(m), .C(k), .Y(ori_ori_n178_));
  NO2        o0150(.A(ori_ori_n178_), .B(ori_ori_n177_), .Y(ori_ori_n179_));
  NAi32      o0151(.An(m), .Bn(k), .C(n), .Y(ori_ori_n180_));
  NO2        o0152(.A(ori_ori_n180_), .B(ori_ori_n177_), .Y(ori_ori_n181_));
  AOI220     o0153(.A0(ori_ori_n181_), .A1(ori_ori_n161_), .B0(ori_ori_n179_), .B1(ori_ori_n176_), .Y(ori_ori_n182_));
  NO2        o0154(.A(n), .B(m), .Y(ori_ori_n183_));
  NA2        o0155(.A(ori_ori_n183_), .B(ori_ori_n50_), .Y(ori_ori_n184_));
  NAi21      o0156(.An(f), .B(e), .Y(ori_ori_n185_));
  NA2        o0157(.A(d), .B(c), .Y(ori_ori_n186_));
  NO2        o0158(.A(ori_ori_n186_), .B(ori_ori_n185_), .Y(ori_ori_n187_));
  NOi21      o0159(.An(ori_ori_n187_), .B(ori_ori_n184_), .Y(ori_ori_n188_));
  NAi31      o0160(.An(m), .B(n), .C(b), .Y(ori_ori_n189_));
  NA2        o0161(.A(k), .B(i), .Y(ori_ori_n190_));
  NAi21      o0162(.An(h), .B(f), .Y(ori_ori_n191_));
  NO2        o0163(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n192_));
  NO2        o0164(.A(ori_ori_n189_), .B(ori_ori_n154_), .Y(ori_ori_n193_));
  NA2        o0165(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NOi32      o0166(.An(f), .Bn(c), .C(d), .Y(ori_ori_n195_));
  NOi32      o0167(.An(f), .Bn(c), .C(e), .Y(ori_ori_n196_));
  NO2        o0168(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  NO3        o0169(.A(n), .B(m), .C(j), .Y(ori_ori_n198_));
  NA2        o0170(.A(ori_ori_n198_), .B(ori_ori_n115_), .Y(ori_ori_n199_));
  AO210      o0171(.A0(ori_ori_n199_), .A1(ori_ori_n184_), .B0(ori_ori_n197_), .Y(ori_ori_n200_));
  NAi41      o0172(.An(ori_ori_n188_), .B(ori_ori_n200_), .C(ori_ori_n194_), .D(ori_ori_n182_), .Y(ori_ori_n201_));
  OR4        o0173(.A(ori_ori_n201_), .B(ori_ori_n173_), .C(ori_ori_n165_), .D(ori_ori_n158_), .Y(ori_ori_n202_));
  NO4        o0174(.A(ori_ori_n202_), .B(ori_ori_n125_), .C(ori_ori_n82_), .D(ori_ori_n55_), .Y(ori_ori_n203_));
  NA3        o0175(.A(m), .B(ori_ori_n113_), .C(j), .Y(ori_ori_n204_));
  NAi31      o0176(.An(n), .B(h), .C(g), .Y(ori_ori_n205_));
  NO2        o0177(.A(ori_ori_n205_), .B(ori_ori_n204_), .Y(ori_ori_n206_));
  NOi32      o0178(.An(m), .Bn(k), .C(l), .Y(ori_ori_n207_));
  NA3        o0179(.A(ori_ori_n207_), .B(ori_ori_n86_), .C(g), .Y(ori_ori_n208_));
  NO2        o0180(.A(ori_ori_n208_), .B(n), .Y(ori_ori_n209_));
  NOi21      o0181(.An(k), .B(j), .Y(ori_ori_n210_));
  NA4        o0182(.A(ori_ori_n210_), .B(ori_ori_n114_), .C(i), .D(g), .Y(ori_ori_n211_));
  AN2        o0183(.A(i), .B(g), .Y(ori_ori_n212_));
  NA3        o0184(.A(ori_ori_n73_), .B(ori_ori_n212_), .C(ori_ori_n114_), .Y(ori_ori_n213_));
  NA2        o0185(.A(ori_ori_n213_), .B(ori_ori_n211_), .Y(ori_ori_n214_));
  NO3        o0186(.A(ori_ori_n214_), .B(ori_ori_n209_), .C(ori_ori_n206_), .Y(ori_ori_n215_));
  NAi41      o0187(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n216_));
  INV        o0188(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  INV        o0189(.A(f), .Y(ori_ori_n218_));
  INV        o0190(.A(g), .Y(ori_ori_n219_));
  NOi31      o0191(.An(i), .B(j), .C(h), .Y(ori_ori_n220_));
  NOi21      o0192(.An(l), .B(m), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NO3        o0194(.A(ori_ori_n222_), .B(ori_ori_n219_), .C(ori_ori_n218_), .Y(ori_ori_n223_));
  NA2        o0195(.A(ori_ori_n223_), .B(ori_ori_n217_), .Y(ori_ori_n224_));
  OAI210     o0196(.A0(ori_ori_n215_), .A1(ori_ori_n32_), .B0(ori_ori_n224_), .Y(ori_ori_n225_));
  NOi21      o0197(.An(n), .B(m), .Y(ori_ori_n226_));
  NOi32      o0198(.An(l), .Bn(i), .C(j), .Y(ori_ori_n227_));
  NA2        o0199(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  OA220      o0200(.A0(ori_ori_n228_), .A1(ori_ori_n106_), .B0(ori_ori_n78_), .B1(ori_ori_n77_), .Y(ori_ori_n229_));
  NAi21      o0201(.An(j), .B(h), .Y(ori_ori_n230_));
  XN2        o0202(.A(i), .B(h), .Y(ori_ori_n231_));
  NA2        o0203(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NOi31      o0204(.An(k), .B(n), .C(m), .Y(ori_ori_n233_));
  NOi31      o0205(.An(ori_ori_n233_), .B(ori_ori_n186_), .C(ori_ori_n185_), .Y(ori_ori_n234_));
  NA2        o0206(.A(ori_ori_n234_), .B(ori_ori_n232_), .Y(ori_ori_n235_));
  NAi31      o0207(.An(f), .B(e), .C(c), .Y(ori_ori_n236_));
  NO4        o0208(.A(ori_ori_n236_), .B(ori_ori_n178_), .C(ori_ori_n177_), .D(ori_ori_n59_), .Y(ori_ori_n237_));
  NA4        o0209(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n238_));
  NAi32      o0210(.An(m), .Bn(i), .C(k), .Y(ori_ori_n239_));
  NO3        o0211(.A(ori_ori_n239_), .B(ori_ori_n90_), .C(ori_ori_n238_), .Y(ori_ori_n240_));
  INV        o0212(.A(k), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n240_), .B(ori_ori_n237_), .Y(ori_ori_n242_));
  NAi21      o0214(.An(n), .B(a), .Y(ori_ori_n243_));
  NO2        o0215(.A(ori_ori_n243_), .B(ori_ori_n149_), .Y(ori_ori_n244_));
  NAi41      o0216(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(e), .Y(ori_ori_n246_));
  NA2        o0218(.A(ori_ori_n246_), .B(ori_ori_n244_), .Y(ori_ori_n247_));
  AN4        o0219(.A(ori_ori_n247_), .B(ori_ori_n242_), .C(ori_ori_n235_), .D(ori_ori_n229_), .Y(ori_ori_n248_));
  OR2        o0220(.A(h), .B(g), .Y(ori_ori_n249_));
  NO2        o0221(.A(ori_ori_n249_), .B(ori_ori_n103_), .Y(ori_ori_n250_));
  NA2        o0222(.A(ori_ori_n250_), .B(ori_ori_n131_), .Y(ori_ori_n251_));
  NAi41      o0223(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n252_));
  NO2        o0224(.A(ori_ori_n252_), .B(ori_ori_n218_), .Y(ori_ori_n253_));
  NA2        o0225(.A(ori_ori_n163_), .B(ori_ori_n109_), .Y(ori_ori_n254_));
  NAi21      o0226(.An(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n255_));
  NO2        o0227(.A(n), .B(a), .Y(ori_ori_n256_));
  NAi31      o0228(.An(ori_ori_n245_), .B(ori_ori_n256_), .C(ori_ori_n104_), .Y(ori_ori_n257_));
  AN2        o0229(.A(ori_ori_n257_), .B(ori_ori_n255_), .Y(ori_ori_n258_));
  NAi21      o0230(.An(h), .B(i), .Y(ori_ori_n259_));
  NA2        o0231(.A(ori_ori_n183_), .B(k), .Y(ori_ori_n260_));
  NO2        o0232(.A(ori_ori_n260_), .B(ori_ori_n259_), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n261_), .B(ori_ori_n195_), .Y(ori_ori_n262_));
  NA3        o0234(.A(ori_ori_n262_), .B(ori_ori_n258_), .C(ori_ori_n251_), .Y(ori_ori_n263_));
  NOi21      o0235(.An(g), .B(e), .Y(ori_ori_n264_));
  NO2        o0236(.A(ori_ori_n71_), .B(ori_ori_n72_), .Y(ori_ori_n265_));
  NA2        o0237(.A(ori_ori_n265_), .B(ori_ori_n264_), .Y(ori_ori_n266_));
  NOi32      o0238(.An(l), .Bn(j), .C(i), .Y(ori_ori_n267_));
  AOI210     o0239(.A0(ori_ori_n73_), .A1(ori_ori_n86_), .B0(ori_ori_n267_), .Y(ori_ori_n268_));
  NO2        o0240(.A(ori_ori_n259_), .B(ori_ori_n44_), .Y(ori_ori_n269_));
  NAi21      o0241(.An(f), .B(g), .Y(ori_ori_n270_));
  NO2        o0242(.A(ori_ori_n270_), .B(ori_ori_n65_), .Y(ori_ori_n271_));
  NA2        o0243(.A(ori_ori_n269_), .B(ori_ori_n67_), .Y(ori_ori_n272_));
  OAI210     o0244(.A0(ori_ori_n268_), .A1(ori_ori_n266_), .B0(ori_ori_n272_), .Y(ori_ori_n273_));
  NO2        o0245(.A(ori_ori_n134_), .B(ori_ori_n49_), .Y(ori_ori_n274_));
  NOi41      o0246(.An(ori_ori_n248_), .B(ori_ori_n273_), .C(ori_ori_n263_), .D(ori_ori_n225_), .Y(ori_ori_n275_));
  NO4        o0247(.A(ori_ori_n206_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n276_));
  NO2        o0248(.A(ori_ori_n276_), .B(ori_ori_n112_), .Y(ori_ori_n277_));
  NA3        o0249(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n278_));
  NAi21      o0250(.An(h), .B(g), .Y(ori_ori_n279_));
  OR4        o0251(.A(ori_ori_n279_), .B(ori_ori_n278_), .C(ori_ori_n228_), .D(e), .Y(ori_ori_n280_));
  NAi31      o0252(.An(g), .B(k), .C(h), .Y(ori_ori_n281_));
  NAi31      o0253(.An(e), .B(d), .C(a), .Y(ori_ori_n282_));
  INV        o0254(.A(ori_ori_n280_), .Y(ori_ori_n283_));
  NA4        o0255(.A(ori_ori_n163_), .B(ori_ori_n79_), .C(ori_ori_n75_), .D(ori_ori_n118_), .Y(ori_ori_n284_));
  NA3        o0256(.A(ori_ori_n163_), .B(ori_ori_n162_), .C(ori_ori_n83_), .Y(ori_ori_n285_));
  NO2        o0257(.A(ori_ori_n285_), .B(ori_ori_n197_), .Y(ori_ori_n286_));
  NOi21      o0258(.An(ori_ori_n284_), .B(ori_ori_n286_), .Y(ori_ori_n287_));
  NA3        o0259(.A(e), .B(c), .C(b), .Y(ori_ori_n288_));
  NO2        o0260(.A(ori_ori_n60_), .B(ori_ori_n288_), .Y(ori_ori_n289_));
  NAi32      o0261(.An(k), .Bn(i), .C(j), .Y(ori_ori_n290_));
  NAi31      o0262(.An(h), .B(l), .C(i), .Y(ori_ori_n291_));
  NA3        o0263(.A(ori_ori_n291_), .B(ori_ori_n290_), .C(ori_ori_n168_), .Y(ori_ori_n292_));
  NOi21      o0264(.An(ori_ori_n292_), .B(ori_ori_n49_), .Y(ori_ori_n293_));
  OAI210     o0265(.A0(ori_ori_n271_), .A1(ori_ori_n289_), .B0(ori_ori_n293_), .Y(ori_ori_n294_));
  NAi21      o0266(.An(l), .B(k), .Y(ori_ori_n295_));
  NO2        o0267(.A(ori_ori_n295_), .B(ori_ori_n49_), .Y(ori_ori_n296_));
  NOi21      o0268(.An(l), .B(j), .Y(ori_ori_n297_));
  NA2        o0269(.A(ori_ori_n166_), .B(ori_ori_n297_), .Y(ori_ori_n298_));
  NAi32      o0270(.An(j), .Bn(h), .C(i), .Y(ori_ori_n299_));
  NAi21      o0271(.An(m), .B(l), .Y(ori_ori_n300_));
  NO3        o0272(.A(ori_ori_n300_), .B(ori_ori_n299_), .C(ori_ori_n83_), .Y(ori_ori_n301_));
  NA2        o0273(.A(h), .B(g), .Y(ori_ori_n302_));
  NA2        o0274(.A(ori_ori_n171_), .B(ori_ori_n45_), .Y(ori_ori_n303_));
  NO2        o0275(.A(ori_ori_n303_), .B(ori_ori_n302_), .Y(ori_ori_n304_));
  NA2        o0276(.A(ori_ori_n304_), .B(ori_ori_n167_), .Y(ori_ori_n305_));
  NA3        o0277(.A(ori_ori_n305_), .B(ori_ori_n294_), .C(ori_ori_n287_), .Y(ori_ori_n306_));
  NO2        o0278(.A(ori_ori_n147_), .B(d), .Y(ori_ori_n307_));
  NA2        o0279(.A(ori_ori_n307_), .B(ori_ori_n53_), .Y(ori_ori_n308_));
  NO2        o0280(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n309_));
  NAi32      o0281(.An(n), .Bn(m), .C(l), .Y(ori_ori_n310_));
  NO2        o0282(.A(ori_ori_n310_), .B(ori_ori_n299_), .Y(ori_ori_n311_));
  NA2        o0283(.A(ori_ori_n311_), .B(ori_ori_n187_), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n123_), .B(ori_ori_n117_), .Y(ori_ori_n313_));
  NAi31      o0285(.An(k), .B(l), .C(j), .Y(ori_ori_n314_));
  OAI210     o0286(.A0(ori_ori_n295_), .A1(j), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  NOi21      o0287(.An(ori_ori_n315_), .B(ori_ori_n121_), .Y(ori_ori_n316_));
  NA2        o0288(.A(ori_ori_n316_), .B(ori_ori_n313_), .Y(ori_ori_n317_));
  NA3        o0289(.A(ori_ori_n317_), .B(ori_ori_n312_), .C(ori_ori_n308_), .Y(ori_ori_n318_));
  NO4        o0290(.A(ori_ori_n318_), .B(ori_ori_n306_), .C(ori_ori_n283_), .D(ori_ori_n277_), .Y(ori_ori_n319_));
  NA2        o0291(.A(ori_ori_n261_), .B(ori_ori_n196_), .Y(ori_ori_n320_));
  NAi21      o0292(.An(m), .B(k), .Y(ori_ori_n321_));
  NO2        o0293(.A(ori_ori_n231_), .B(ori_ori_n321_), .Y(ori_ori_n322_));
  NAi41      o0294(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n323_));
  NO2        o0295(.A(ori_ori_n323_), .B(ori_ori_n153_), .Y(ori_ori_n324_));
  NA2        o0296(.A(ori_ori_n324_), .B(ori_ori_n322_), .Y(ori_ori_n325_));
  NA2        o0297(.A(e), .B(c), .Y(ori_ori_n326_));
  NO3        o0298(.A(ori_ori_n326_), .B(n), .C(d), .Y(ori_ori_n327_));
  NOi21      o0299(.An(f), .B(h), .Y(ori_ori_n328_));
  NAi31      o0300(.An(d), .B(e), .C(b), .Y(ori_ori_n329_));
  NA2        o0301(.A(ori_ori_n325_), .B(ori_ori_n320_), .Y(ori_ori_n330_));
  NA2        o0302(.A(ori_ori_n256_), .B(ori_ori_n104_), .Y(ori_ori_n331_));
  OR2        o0303(.A(ori_ori_n331_), .B(ori_ori_n208_), .Y(ori_ori_n332_));
  NOi31      o0304(.An(l), .B(n), .C(m), .Y(ori_ori_n333_));
  NA2        o0305(.A(ori_ori_n333_), .B(ori_ori_n220_), .Y(ori_ori_n334_));
  NO2        o0306(.A(ori_ori_n334_), .B(ori_ori_n197_), .Y(ori_ori_n335_));
  NAi21      o0307(.An(ori_ori_n335_), .B(ori_ori_n332_), .Y(ori_ori_n336_));
  NAi32      o0308(.An(m), .Bn(j), .C(k), .Y(ori_ori_n337_));
  NAi41      o0309(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n338_));
  NOi31      o0310(.An(j), .B(m), .C(k), .Y(ori_ori_n339_));
  NO2        o0311(.A(ori_ori_n126_), .B(ori_ori_n339_), .Y(ori_ori_n340_));
  AN3        o0312(.A(h), .B(g), .C(f), .Y(ori_ori_n341_));
  NOi32      o0313(.An(m), .Bn(j), .C(l), .Y(ori_ori_n342_));
  NO2        o0314(.A(ori_ori_n342_), .B(ori_ori_n97_), .Y(ori_ori_n343_));
  NO2        o0315(.A(ori_ori_n300_), .B(ori_ori_n299_), .Y(ori_ori_n344_));
  NA2        o0316(.A(ori_ori_n253_), .B(ori_ori_n344_), .Y(ori_ori_n345_));
  NA2        o0317(.A(ori_ori_n239_), .B(ori_ori_n78_), .Y(ori_ori_n346_));
  NA3        o0318(.A(ori_ori_n346_), .B(ori_ori_n341_), .C(ori_ori_n217_), .Y(ori_ori_n347_));
  NA2        o0319(.A(ori_ori_n347_), .B(ori_ori_n345_), .Y(ori_ori_n348_));
  NA3        o0320(.A(h), .B(g), .C(f), .Y(ori_ori_n349_));
  NO2        o0321(.A(ori_ori_n349_), .B(ori_ori_n74_), .Y(ori_ori_n350_));
  NA2        o0322(.A(ori_ori_n338_), .B(ori_ori_n216_), .Y(ori_ori_n351_));
  NA2        o0323(.A(ori_ori_n166_), .B(e), .Y(ori_ori_n352_));
  NO2        o0324(.A(ori_ori_n352_), .B(ori_ori_n41_), .Y(ori_ori_n353_));
  AOI220     o0325(.A0(ori_ori_n353_), .A1(ori_ori_n313_), .B0(ori_ori_n351_), .B1(ori_ori_n350_), .Y(ori_ori_n354_));
  NOi32      o0326(.An(j), .Bn(g), .C(i), .Y(ori_ori_n355_));
  NA3        o0327(.A(ori_ori_n355_), .B(ori_ori_n295_), .C(ori_ori_n114_), .Y(ori_ori_n356_));
  AO210      o0328(.A0(ori_ori_n112_), .A1(ori_ori_n32_), .B0(ori_ori_n356_), .Y(ori_ori_n357_));
  NOi32      o0329(.An(e), .Bn(b), .C(a), .Y(ori_ori_n358_));
  AN2        o0330(.A(l), .B(j), .Y(ori_ori_n359_));
  NA3        o0331(.A(ori_ori_n213_), .B(ori_ori_n211_), .C(ori_ori_n35_), .Y(ori_ori_n360_));
  NA2        o0332(.A(ori_ori_n360_), .B(ori_ori_n358_), .Y(ori_ori_n361_));
  NO2        o0333(.A(ori_ori_n329_), .B(n), .Y(ori_ori_n362_));
  NA2        o0334(.A(ori_ori_n212_), .B(k), .Y(ori_ori_n363_));
  NA3        o0335(.A(m), .B(ori_ori_n113_), .C(ori_ori_n218_), .Y(ori_ori_n364_));
  NA4        o0336(.A(ori_ori_n207_), .B(ori_ori_n86_), .C(g), .D(ori_ori_n218_), .Y(ori_ori_n365_));
  OAI210     o0337(.A0(ori_ori_n364_), .A1(ori_ori_n363_), .B0(ori_ori_n365_), .Y(ori_ori_n366_));
  NAi41      o0338(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n367_));
  NA2        o0339(.A(ori_ori_n51_), .B(ori_ori_n114_), .Y(ori_ori_n368_));
  NO2        o0340(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n369_));
  AOI220     o0341(.A0(ori_ori_n369_), .A1(b), .B0(ori_ori_n366_), .B1(ori_ori_n362_), .Y(ori_ori_n370_));
  NA4        o0342(.A(ori_ori_n370_), .B(ori_ori_n361_), .C(ori_ori_n357_), .D(ori_ori_n354_), .Y(ori_ori_n371_));
  NO4        o0343(.A(ori_ori_n371_), .B(ori_ori_n348_), .C(ori_ori_n336_), .D(ori_ori_n330_), .Y(ori_ori_n372_));
  NA4        o0344(.A(ori_ori_n372_), .B(ori_ori_n319_), .C(ori_ori_n275_), .D(ori_ori_n203_), .Y(ori10));
  NA3        o0345(.A(m), .B(k), .C(i), .Y(ori_ori_n374_));
  NOi21      o0346(.An(e), .B(f), .Y(ori_ori_n375_));
  NO4        o0347(.A(ori_ori_n154_), .B(ori_ori_n375_), .C(n), .D(ori_ori_n111_), .Y(ori_ori_n376_));
  NAi31      o0348(.An(b), .B(f), .C(c), .Y(ori_ori_n377_));
  INV        o0349(.A(ori_ori_n377_), .Y(ori_ori_n378_));
  NOi32      o0350(.An(k), .Bn(h), .C(j), .Y(ori_ori_n379_));
  NA2        o0351(.A(ori_ori_n379_), .B(ori_ori_n226_), .Y(ori_ori_n380_));
  NA2        o0352(.A(ori_ori_n164_), .B(ori_ori_n380_), .Y(ori_ori_n381_));
  NA2        o0353(.A(ori_ori_n381_), .B(ori_ori_n378_), .Y(ori_ori_n382_));
  AN2        o0354(.A(j), .B(h), .Y(ori_ori_n383_));
  NO3        o0355(.A(n), .B(m), .C(k), .Y(ori_ori_n384_));
  NA2        o0356(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n385_));
  NO3        o0357(.A(ori_ori_n385_), .B(ori_ori_n154_), .C(ori_ori_n218_), .Y(ori_ori_n386_));
  OR2        o0358(.A(m), .B(k), .Y(ori_ori_n387_));
  NO2        o0359(.A(ori_ori_n177_), .B(ori_ori_n387_), .Y(ori_ori_n388_));
  NA4        o0360(.A(n), .B(f), .C(c), .D(ori_ori_n117_), .Y(ori_ori_n389_));
  NOi21      o0361(.An(ori_ori_n388_), .B(ori_ori_n389_), .Y(ori_ori_n390_));
  NOi32      o0362(.An(d), .Bn(a), .C(c), .Y(ori_ori_n391_));
  NA2        o0363(.A(ori_ori_n391_), .B(ori_ori_n185_), .Y(ori_ori_n392_));
  NAi21      o0364(.An(i), .B(g), .Y(ori_ori_n393_));
  NAi31      o0365(.An(k), .B(m), .C(j), .Y(ori_ori_n394_));
  NO3        o0366(.A(ori_ori_n394_), .B(ori_ori_n393_), .C(n), .Y(ori_ori_n395_));
  NOi21      o0367(.An(ori_ori_n395_), .B(ori_ori_n392_), .Y(ori_ori_n396_));
  NO3        o0368(.A(ori_ori_n396_), .B(ori_ori_n390_), .C(ori_ori_n386_), .Y(ori_ori_n397_));
  NO2        o0369(.A(ori_ori_n389_), .B(ori_ori_n300_), .Y(ori_ori_n398_));
  NOi32      o0370(.An(f), .Bn(d), .C(c), .Y(ori_ori_n399_));
  AOI220     o0371(.A0(ori_ori_n399_), .A1(ori_ori_n311_), .B0(ori_ori_n398_), .B1(ori_ori_n220_), .Y(ori_ori_n400_));
  NA3        o0372(.A(ori_ori_n400_), .B(ori_ori_n397_), .C(ori_ori_n382_), .Y(ori_ori_n401_));
  NO2        o0373(.A(ori_ori_n59_), .B(ori_ori_n117_), .Y(ori_ori_n402_));
  NA2        o0374(.A(ori_ori_n256_), .B(ori_ori_n402_), .Y(ori_ori_n403_));
  INV        o0375(.A(e), .Y(ori_ori_n404_));
  NA2        o0376(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n405_));
  OAI220     o0377(.A0(ori_ori_n405_), .A1(ori_ori_n204_), .B0(ori_ori_n208_), .B1(ori_ori_n404_), .Y(ori_ori_n406_));
  AN2        o0378(.A(g), .B(e), .Y(ori_ori_n407_));
  NA3        o0379(.A(ori_ori_n407_), .B(ori_ori_n207_), .C(i), .Y(ori_ori_n408_));
  OAI210     o0380(.A0(ori_ori_n88_), .A1(ori_ori_n404_), .B0(ori_ori_n408_), .Y(ori_ori_n409_));
  NO2        o0381(.A(ori_ori_n100_), .B(ori_ori_n404_), .Y(ori_ori_n410_));
  NO3        o0382(.A(ori_ori_n410_), .B(ori_ori_n409_), .C(ori_ori_n406_), .Y(ori_ori_n411_));
  NOi32      o0383(.An(h), .Bn(e), .C(g), .Y(ori_ori_n412_));
  NA3        o0384(.A(ori_ori_n412_), .B(ori_ori_n297_), .C(m), .Y(ori_ori_n413_));
  NOi21      o0385(.An(g), .B(h), .Y(ori_ori_n414_));
  AN3        o0386(.A(m), .B(l), .C(i), .Y(ori_ori_n415_));
  NA3        o0387(.A(ori_ori_n415_), .B(ori_ori_n414_), .C(e), .Y(ori_ori_n416_));
  AN3        o0388(.A(h), .B(g), .C(e), .Y(ori_ori_n417_));
  NA2        o0389(.A(ori_ori_n417_), .B(ori_ori_n97_), .Y(ori_ori_n418_));
  AN3        o0390(.A(ori_ori_n418_), .B(ori_ori_n416_), .C(ori_ori_n413_), .Y(ori_ori_n419_));
  AOI210     o0391(.A0(ori_ori_n419_), .A1(ori_ori_n411_), .B0(ori_ori_n403_), .Y(ori_ori_n420_));
  NA3        o0392(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(e), .Y(ori_ori_n421_));
  NO2        o0393(.A(ori_ori_n421_), .B(ori_ori_n403_), .Y(ori_ori_n422_));
  NA3        o0394(.A(ori_ori_n391_), .B(ori_ori_n185_), .C(ori_ori_n83_), .Y(ori_ori_n423_));
  NAi31      o0395(.An(b), .B(c), .C(a), .Y(ori_ori_n424_));
  NO2        o0396(.A(ori_ori_n424_), .B(n), .Y(ori_ori_n425_));
  NA2        o0397(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n426_));
  NO2        o0398(.A(ori_ori_n426_), .B(ori_ori_n150_), .Y(ori_ori_n427_));
  NA2        o0399(.A(ori_ori_n427_), .B(ori_ori_n425_), .Y(ori_ori_n428_));
  INV        o0400(.A(ori_ori_n428_), .Y(ori_ori_n429_));
  NO4        o0401(.A(ori_ori_n429_), .B(ori_ori_n422_), .C(ori_ori_n420_), .D(ori_ori_n401_), .Y(ori_ori_n430_));
  NA2        o0402(.A(i), .B(g), .Y(ori_ori_n431_));
  NOi21      o0403(.An(d), .B(c), .Y(ori_ori_n432_));
  NA3        o0404(.A(i), .B(g), .C(f), .Y(ori_ori_n433_));
  OR2        o0405(.A(n), .B(m), .Y(ori_ori_n434_));
  NO2        o0406(.A(ori_ori_n434_), .B(ori_ori_n155_), .Y(ori_ori_n435_));
  NO2        o0407(.A(ori_ori_n186_), .B(ori_ori_n150_), .Y(ori_ori_n436_));
  OAI210     o0408(.A0(ori_ori_n435_), .A1(ori_ori_n179_), .B0(ori_ori_n436_), .Y(ori_ori_n437_));
  INV        o0409(.A(ori_ori_n368_), .Y(ori_ori_n438_));
  NA3        o0410(.A(ori_ori_n438_), .B(ori_ori_n358_), .C(d), .Y(ori_ori_n439_));
  NO2        o0411(.A(ori_ori_n424_), .B(ori_ori_n49_), .Y(ori_ori_n440_));
  NO3        o0412(.A(ori_ori_n66_), .B(ori_ori_n113_), .C(e), .Y(ori_ori_n441_));
  NAi21      o0413(.An(k), .B(j), .Y(ori_ori_n442_));
  NA2        o0414(.A(ori_ori_n259_), .B(ori_ori_n442_), .Y(ori_ori_n443_));
  NA3        o0415(.A(ori_ori_n443_), .B(ori_ori_n441_), .C(ori_ori_n440_), .Y(ori_ori_n444_));
  NAi21      o0416(.An(e), .B(d), .Y(ori_ori_n445_));
  INV        o0417(.A(ori_ori_n445_), .Y(ori_ori_n446_));
  NO2        o0418(.A(ori_ori_n260_), .B(ori_ori_n218_), .Y(ori_ori_n447_));
  NA3        o0419(.A(ori_ori_n447_), .B(ori_ori_n446_), .C(ori_ori_n232_), .Y(ori_ori_n448_));
  NA4        o0420(.A(ori_ori_n448_), .B(ori_ori_n444_), .C(ori_ori_n439_), .D(ori_ori_n437_), .Y(ori_ori_n449_));
  NO2        o0421(.A(ori_ori_n334_), .B(ori_ori_n218_), .Y(ori_ori_n450_));
  NA2        o0422(.A(ori_ori_n450_), .B(ori_ori_n446_), .Y(ori_ori_n451_));
  NOi31      o0423(.An(n), .B(m), .C(k), .Y(ori_ori_n452_));
  AOI220     o0424(.A0(ori_ori_n452_), .A1(ori_ori_n383_), .B0(ori_ori_n226_), .B1(ori_ori_n50_), .Y(ori_ori_n453_));
  NAi31      o0425(.An(g), .B(f), .C(c), .Y(ori_ori_n454_));
  OR3        o0426(.A(ori_ori_n454_), .B(ori_ori_n453_), .C(e), .Y(ori_ori_n455_));
  NA3        o0427(.A(ori_ori_n455_), .B(ori_ori_n451_), .C(ori_ori_n312_), .Y(ori_ori_n456_));
  NO3        o0428(.A(ori_ori_n456_), .B(ori_ori_n449_), .C(ori_ori_n273_), .Y(ori_ori_n457_));
  NOi32      o0429(.An(c), .Bn(a), .C(b), .Y(ori_ori_n458_));
  NA2        o0430(.A(ori_ori_n458_), .B(ori_ori_n114_), .Y(ori_ori_n459_));
  INV        o0431(.A(ori_ori_n281_), .Y(ori_ori_n460_));
  AN2        o0432(.A(e), .B(d), .Y(ori_ori_n461_));
  NA2        o0433(.A(ori_ori_n461_), .B(ori_ori_n460_), .Y(ori_ori_n462_));
  INV        o0434(.A(ori_ori_n150_), .Y(ori_ori_n463_));
  NO2        o0435(.A(ori_ori_n132_), .B(ori_ori_n41_), .Y(ori_ori_n464_));
  NO2        o0436(.A(ori_ori_n66_), .B(e), .Y(ori_ori_n465_));
  NOi31      o0437(.An(j), .B(k), .C(i), .Y(ori_ori_n466_));
  NOi21      o0438(.An(ori_ori_n168_), .B(ori_ori_n466_), .Y(ori_ori_n467_));
  NA3        o0439(.A(ori_ori_n467_), .B(ori_ori_n268_), .C(ori_ori_n120_), .Y(ori_ori_n468_));
  NA2        o0440(.A(ori_ori_n468_), .B(ori_ori_n465_), .Y(ori_ori_n469_));
  AOI210     o0441(.A0(ori_ori_n469_), .A1(ori_ori_n462_), .B0(ori_ori_n459_), .Y(ori_ori_n470_));
  NO2        o0442(.A(ori_ori_n214_), .B(ori_ori_n209_), .Y(ori_ori_n471_));
  NOi21      o0443(.An(a), .B(b), .Y(ori_ori_n472_));
  NA3        o0444(.A(e), .B(d), .C(c), .Y(ori_ori_n473_));
  NAi21      o0445(.An(ori_ori_n473_), .B(ori_ori_n472_), .Y(ori_ori_n474_));
  NO2        o0446(.A(ori_ori_n423_), .B(ori_ori_n208_), .Y(ori_ori_n475_));
  NOi21      o0447(.An(ori_ori_n474_), .B(ori_ori_n475_), .Y(ori_ori_n476_));
  AOI210     o0448(.A0(ori_ori_n276_), .A1(ori_ori_n471_), .B0(ori_ori_n476_), .Y(ori_ori_n477_));
  NO4        o0449(.A(ori_ori_n191_), .B(ori_ori_n103_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n478_));
  NA2        o0450(.A(ori_ori_n378_), .B(ori_ori_n156_), .Y(ori_ori_n479_));
  OR2        o0451(.A(k), .B(j), .Y(ori_ori_n480_));
  NA2        o0452(.A(l), .B(k), .Y(ori_ori_n481_));
  NA3        o0453(.A(ori_ori_n481_), .B(ori_ori_n480_), .C(ori_ori_n226_), .Y(ori_ori_n482_));
  AOI210     o0454(.A0(ori_ori_n239_), .A1(ori_ori_n337_), .B0(ori_ori_n83_), .Y(ori_ori_n483_));
  NOi21      o0455(.An(ori_ori_n482_), .B(ori_ori_n483_), .Y(ori_ori_n484_));
  OR3        o0456(.A(ori_ori_n484_), .B(ori_ori_n146_), .C(ori_ori_n136_), .Y(ori_ori_n485_));
  NA3        o0457(.A(ori_ori_n284_), .B(ori_ori_n129_), .C(ori_ori_n127_), .Y(ori_ori_n486_));
  NO3        o0458(.A(ori_ori_n423_), .B(ori_ori_n91_), .C(ori_ori_n132_), .Y(ori_ori_n487_));
  NO2        o0459(.A(ori_ori_n487_), .B(ori_ori_n486_), .Y(ori_ori_n488_));
  NA3        o0460(.A(ori_ori_n488_), .B(ori_ori_n485_), .C(ori_ori_n479_), .Y(ori_ori_n489_));
  NO4        o0461(.A(ori_ori_n489_), .B(ori_ori_n478_), .C(ori_ori_n477_), .D(ori_ori_n470_), .Y(ori_ori_n490_));
  INV        o0462(.A(e), .Y(ori_ori_n491_));
  NO2        o0463(.A(ori_ori_n191_), .B(ori_ori_n56_), .Y(ori_ori_n492_));
  NAi31      o0464(.An(j), .B(l), .C(i), .Y(ori_ori_n493_));
  OAI210     o0465(.A0(ori_ori_n493_), .A1(ori_ori_n133_), .B0(ori_ori_n103_), .Y(ori_ori_n494_));
  NA3        o0466(.A(ori_ori_n494_), .B(ori_ori_n492_), .C(ori_ori_n491_), .Y(ori_ori_n495_));
  NO3        o0467(.A(ori_ori_n392_), .B(ori_ori_n343_), .C(ori_ori_n205_), .Y(ori_ori_n496_));
  NO2        o0468(.A(ori_ori_n392_), .B(ori_ori_n368_), .Y(ori_ori_n497_));
  NO4        o0469(.A(ori_ori_n497_), .B(ori_ori_n496_), .C(ori_ori_n188_), .D(ori_ori_n309_), .Y(ori_ori_n498_));
  NA3        o0470(.A(ori_ori_n498_), .B(ori_ori_n495_), .C(ori_ori_n248_), .Y(ori_ori_n499_));
  OAI210     o0471(.A0(ori_ori_n128_), .A1(ori_ori_n126_), .B0(n), .Y(ori_ori_n500_));
  NO2        o0472(.A(ori_ori_n500_), .B(ori_ori_n132_), .Y(ori_ori_n501_));
  XO2        o0473(.A(i), .B(h), .Y(ori_ori_n502_));
  NA3        o0474(.A(ori_ori_n502_), .B(ori_ori_n163_), .C(n), .Y(ori_ori_n503_));
  NAi41      o0475(.An(ori_ori_n301_), .B(ori_ori_n503_), .C(ori_ori_n453_), .D(ori_ori_n380_), .Y(ori_ori_n504_));
  NAi31      o0476(.An(c), .B(f), .C(d), .Y(ori_ori_n505_));
  AOI210     o0477(.A0(ori_ori_n285_), .A1(ori_ori_n199_), .B0(ori_ori_n505_), .Y(ori_ori_n506_));
  NOi21      o0478(.An(ori_ori_n81_), .B(ori_ori_n506_), .Y(ori_ori_n507_));
  NA3        o0479(.A(ori_ori_n376_), .B(ori_ori_n97_), .C(ori_ori_n96_), .Y(ori_ori_n508_));
  NA2        o0480(.A(ori_ori_n233_), .B(ori_ori_n109_), .Y(ori_ori_n509_));
  AOI210     o0481(.A0(ori_ori_n509_), .A1(ori_ori_n184_), .B0(ori_ori_n505_), .Y(ori_ori_n510_));
  NOi21      o0482(.An(ori_ori_n508_), .B(ori_ori_n510_), .Y(ori_ori_n511_));
  AO220      o0483(.A0(ori_ori_n293_), .A1(ori_ori_n271_), .B0(ori_ori_n169_), .B1(ori_ori_n67_), .Y(ori_ori_n512_));
  NA3        o0484(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n513_));
  NAi31      o0485(.An(ori_ori_n512_), .B(ori_ori_n511_), .C(ori_ori_n507_), .Y(ori_ori_n514_));
  NO2        o0486(.A(ori_ori_n514_), .B(ori_ori_n499_), .Y(ori_ori_n515_));
  NA4        o0487(.A(ori_ori_n515_), .B(ori_ori_n490_), .C(ori_ori_n457_), .D(ori_ori_n430_), .Y(ori11));
  NO2        o0488(.A(ori_ori_n71_), .B(f), .Y(ori_ori_n517_));
  NA2        o0489(.A(j), .B(g), .Y(ori_ori_n518_));
  NAi31      o0490(.An(i), .B(m), .C(l), .Y(ori_ori_n519_));
  NA3        o0491(.A(m), .B(k), .C(j), .Y(ori_ori_n520_));
  OAI220     o0492(.A0(ori_ori_n520_), .A1(ori_ori_n132_), .B0(ori_ori_n519_), .B1(ori_ori_n518_), .Y(ori_ori_n521_));
  NA2        o0493(.A(ori_ori_n521_), .B(ori_ori_n517_), .Y(ori_ori_n522_));
  NOi32      o0494(.An(e), .Bn(b), .C(f), .Y(ori_ori_n523_));
  NA2        o0495(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n524_));
  NO2        o0496(.A(ori_ori_n524_), .B(ori_ori_n303_), .Y(ori_ori_n525_));
  NAi31      o0497(.An(d), .B(e), .C(a), .Y(ori_ori_n526_));
  NO2        o0498(.A(ori_ori_n526_), .B(n), .Y(ori_ori_n527_));
  AOI220     o0499(.A0(ori_ori_n527_), .A1(ori_ori_n101_), .B0(ori_ori_n525_), .B1(ori_ori_n523_), .Y(ori_ori_n528_));
  NAi41      o0500(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n529_));
  AN2        o0501(.A(ori_ori_n529_), .B(ori_ori_n367_), .Y(ori_ori_n530_));
  NA2        o0502(.A(j), .B(i), .Y(ori_ori_n531_));
  NAi31      o0503(.An(n), .B(m), .C(k), .Y(ori_ori_n532_));
  NO3        o0504(.A(ori_ori_n532_), .B(ori_ori_n531_), .C(ori_ori_n113_), .Y(ori_ori_n533_));
  NO4        o0505(.A(n), .B(d), .C(ori_ori_n117_), .D(a), .Y(ori_ori_n534_));
  OR2        o0506(.A(n), .B(c), .Y(ori_ori_n535_));
  NO2        o0507(.A(ori_ori_n535_), .B(ori_ori_n152_), .Y(ori_ori_n536_));
  NO2        o0508(.A(ori_ori_n536_), .B(ori_ori_n534_), .Y(ori_ori_n537_));
  NOi32      o0509(.An(g), .Bn(f), .C(i), .Y(ori_ori_n538_));
  AOI220     o0510(.A0(ori_ori_n538_), .A1(ori_ori_n99_), .B0(ori_ori_n521_), .B1(f), .Y(ori_ori_n539_));
  NO2        o0511(.A(ori_ori_n281_), .B(ori_ori_n49_), .Y(ori_ori_n540_));
  NO2        o0512(.A(ori_ori_n539_), .B(ori_ori_n537_), .Y(ori_ori_n541_));
  INV        o0513(.A(ori_ori_n541_), .Y(ori_ori_n542_));
  NA2        o0514(.A(ori_ori_n142_), .B(ori_ori_n34_), .Y(ori_ori_n543_));
  OAI220     o0515(.A0(ori_ori_n543_), .A1(m), .B0(ori_ori_n524_), .B1(ori_ori_n239_), .Y(ori_ori_n544_));
  NOi41      o0516(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n545_));
  NAi32      o0517(.An(e), .Bn(b), .C(c), .Y(ori_ori_n546_));
  OR2        o0518(.A(ori_ori_n546_), .B(ori_ori_n83_), .Y(ori_ori_n547_));
  AN2        o0519(.A(ori_ori_n338_), .B(ori_ori_n323_), .Y(ori_ori_n548_));
  NA2        o0520(.A(ori_ori_n548_), .B(ori_ori_n547_), .Y(ori_ori_n549_));
  OA210      o0521(.A0(ori_ori_n549_), .A1(ori_ori_n545_), .B0(ori_ori_n544_), .Y(ori_ori_n550_));
  OAI220     o0522(.A0(ori_ori_n394_), .A1(ori_ori_n393_), .B0(ori_ori_n519_), .B1(ori_ori_n518_), .Y(ori_ori_n551_));
  NAi31      o0523(.An(d), .B(c), .C(a), .Y(ori_ori_n552_));
  NO2        o0524(.A(ori_ori_n552_), .B(n), .Y(ori_ori_n553_));
  NA3        o0525(.A(ori_ori_n553_), .B(ori_ori_n551_), .C(e), .Y(ori_ori_n554_));
  NO3        o0526(.A(ori_ori_n62_), .B(ori_ori_n49_), .C(ori_ori_n219_), .Y(ori_ori_n555_));
  NO2        o0527(.A(ori_ori_n236_), .B(ori_ori_n111_), .Y(ori_ori_n556_));
  OAI210     o0528(.A0(ori_ori_n555_), .A1(ori_ori_n395_), .B0(ori_ori_n556_), .Y(ori_ori_n557_));
  NA2        o0529(.A(ori_ori_n557_), .B(ori_ori_n554_), .Y(ori_ori_n558_));
  NO2        o0530(.A(ori_ori_n282_), .B(n), .Y(ori_ori_n559_));
  NO2        o0531(.A(ori_ori_n425_), .B(ori_ori_n559_), .Y(ori_ori_n560_));
  NA2        o0532(.A(ori_ori_n551_), .B(f), .Y(ori_ori_n561_));
  NAi21      o0533(.An(d), .B(b), .Y(ori_ori_n562_));
  NO2        o0534(.A(ori_ori_n562_), .B(ori_ori_n49_), .Y(ori_ori_n563_));
  NA2        o0535(.A(h), .B(f), .Y(ori_ori_n564_));
  NO2        o0536(.A(ori_ori_n564_), .B(ori_ori_n94_), .Y(ori_ori_n565_));
  NA2        o0537(.A(ori_ori_n565_), .B(ori_ori_n563_), .Y(ori_ori_n566_));
  OAI210     o0538(.A0(ori_ori_n561_), .A1(ori_ori_n560_), .B0(ori_ori_n566_), .Y(ori_ori_n567_));
  NO2        o0539(.A(ori_ori_n149_), .B(c), .Y(ori_ori_n568_));
  NA3        o0540(.A(f), .B(d), .C(b), .Y(ori_ori_n569_));
  NO4        o0541(.A(ori_ori_n569_), .B(ori_ori_n180_), .C(ori_ori_n177_), .D(g), .Y(ori_ori_n570_));
  NO4        o0542(.A(ori_ori_n570_), .B(ori_ori_n567_), .C(ori_ori_n558_), .D(ori_ori_n550_), .Y(ori_ori_n571_));
  AN4        o0543(.A(ori_ori_n571_), .B(ori_ori_n542_), .C(ori_ori_n528_), .D(ori_ori_n522_), .Y(ori_ori_n572_));
  INV        o0544(.A(k), .Y(ori_ori_n573_));
  NA3        o0545(.A(l), .B(ori_ori_n573_), .C(i), .Y(ori_ori_n574_));
  INV        o0546(.A(ori_ori_n574_), .Y(ori_ori_n575_));
  NAi32      o0547(.An(h), .Bn(f), .C(g), .Y(ori_ori_n576_));
  NAi41      o0548(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n577_));
  OAI210     o0549(.A0(ori_ori_n526_), .A1(n), .B0(ori_ori_n577_), .Y(ori_ori_n578_));
  NA2        o0550(.A(ori_ori_n578_), .B(m), .Y(ori_ori_n579_));
  NAi31      o0551(.An(h), .B(g), .C(f), .Y(ori_ori_n580_));
  OR3        o0552(.A(ori_ori_n580_), .B(ori_ori_n282_), .C(ori_ori_n49_), .Y(ori_ori_n581_));
  NA4        o0553(.A(ori_ori_n414_), .B(ori_ori_n122_), .C(ori_ori_n114_), .D(e), .Y(ori_ori_n582_));
  AN2        o0554(.A(ori_ori_n582_), .B(ori_ori_n581_), .Y(ori_ori_n583_));
  OA210      o0555(.A0(ori_ori_n579_), .A1(ori_ori_n576_), .B0(ori_ori_n583_), .Y(ori_ori_n584_));
  NO3        o0556(.A(ori_ori_n576_), .B(ori_ori_n71_), .C(ori_ori_n72_), .Y(ori_ori_n585_));
  NO4        o0557(.A(ori_ori_n580_), .B(ori_ori_n535_), .C(ori_ori_n152_), .D(ori_ori_n72_), .Y(ori_ori_n586_));
  OR2        o0558(.A(ori_ori_n586_), .B(ori_ori_n585_), .Y(ori_ori_n587_));
  NAi21      o0559(.An(ori_ori_n587_), .B(ori_ori_n584_), .Y(ori_ori_n588_));
  NAi31      o0560(.An(f), .B(h), .C(g), .Y(ori_ori_n589_));
  NOi32      o0561(.An(b), .Bn(a), .C(c), .Y(ori_ori_n590_));
  NOi32      o0562(.An(d), .Bn(a), .C(e), .Y(ori_ori_n591_));
  NA2        o0563(.A(ori_ori_n591_), .B(ori_ori_n114_), .Y(ori_ori_n592_));
  NO2        o0564(.A(n), .B(c), .Y(ori_ori_n593_));
  NA3        o0565(.A(ori_ori_n593_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n594_));
  NAi32      o0566(.An(n), .Bn(f), .C(m), .Y(ori_ori_n595_));
  NA3        o0567(.A(ori_ori_n595_), .B(ori_ori_n594_), .C(ori_ori_n592_), .Y(ori_ori_n596_));
  NOi32      o0568(.An(e), .Bn(a), .C(d), .Y(ori_ori_n597_));
  AOI210     o0569(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n597_), .Y(ori_ori_n598_));
  AOI210     o0570(.A0(ori_ori_n598_), .A1(ori_ori_n218_), .B0(ori_ori_n543_), .Y(ori_ori_n599_));
  NA2        o0571(.A(ori_ori_n599_), .B(ori_ori_n596_), .Y(ori_ori_n600_));
  OAI210     o0572(.A0(ori_ori_n255_), .A1(ori_ori_n86_), .B0(ori_ori_n600_), .Y(ori_ori_n601_));
  AOI210     o0573(.A0(ori_ori_n588_), .A1(ori_ori_n575_), .B0(ori_ori_n601_), .Y(ori_ori_n602_));
  NO3        o0574(.A(ori_ori_n321_), .B(ori_ori_n61_), .C(n), .Y(ori_ori_n603_));
  NA3        o0575(.A(ori_ori_n505_), .B(ori_ori_n175_), .C(ori_ori_n174_), .Y(ori_ori_n604_));
  NA2        o0576(.A(ori_ori_n454_), .B(ori_ori_n236_), .Y(ori_ori_n605_));
  OR2        o0577(.A(ori_ori_n605_), .B(ori_ori_n604_), .Y(ori_ori_n606_));
  NA2        o0578(.A(ori_ori_n606_), .B(ori_ori_n603_), .Y(ori_ori_n607_));
  NO2        o0579(.A(ori_ori_n607_), .B(ori_ori_n86_), .Y(ori_ori_n608_));
  NA3        o0580(.A(ori_ori_n545_), .B(ori_ori_n339_), .C(ori_ori_n46_), .Y(ori_ori_n609_));
  NOi32      o0581(.An(e), .Bn(c), .C(f), .Y(ori_ori_n610_));
  NOi21      o0582(.An(f), .B(g), .Y(ori_ori_n611_));
  NO2        o0583(.A(ori_ori_n611_), .B(ori_ori_n216_), .Y(ori_ori_n612_));
  AOI220     o0584(.A0(ori_ori_n612_), .A1(ori_ori_n388_), .B0(ori_ori_n610_), .B1(ori_ori_n179_), .Y(ori_ori_n613_));
  NA3        o0585(.A(ori_ori_n613_), .B(ori_ori_n609_), .C(ori_ori_n182_), .Y(ori_ori_n614_));
  AOI210     o0586(.A0(ori_ori_n530_), .A1(ori_ori_n392_), .B0(ori_ori_n302_), .Y(ori_ori_n615_));
  NOi21      o0587(.An(j), .B(l), .Y(ori_ori_n616_));
  NAi21      o0588(.An(k), .B(h), .Y(ori_ori_n617_));
  NO2        o0589(.A(ori_ori_n617_), .B(ori_ori_n270_), .Y(ori_ori_n618_));
  NOi31      o0590(.An(m), .B(n), .C(k), .Y(ori_ori_n619_));
  NA2        o0591(.A(ori_ori_n616_), .B(ori_ori_n619_), .Y(ori_ori_n620_));
  AOI210     o0592(.A0(ori_ori_n392_), .A1(ori_ori_n367_), .B0(ori_ori_n302_), .Y(ori_ori_n621_));
  NAi21      o0593(.An(ori_ori_n620_), .B(ori_ori_n621_), .Y(ori_ori_n622_));
  NO2        o0594(.A(ori_ori_n282_), .B(ori_ori_n49_), .Y(ori_ori_n623_));
  NO2        o0595(.A(ori_ori_n526_), .B(ori_ori_n49_), .Y(ori_ori_n624_));
  NA2        o0596(.A(ori_ori_n623_), .B(ori_ori_n565_), .Y(ori_ori_n625_));
  NA2        o0597(.A(ori_ori_n625_), .B(ori_ori_n622_), .Y(ori_ori_n626_));
  NA2        o0598(.A(ori_ori_n109_), .B(ori_ori_n36_), .Y(ori_ori_n627_));
  NO2        o0599(.A(k), .B(ori_ori_n219_), .Y(ori_ori_n628_));
  INV        o0600(.A(ori_ori_n358_), .Y(ori_ori_n629_));
  NO2        o0601(.A(ori_ori_n629_), .B(n), .Y(ori_ori_n630_));
  NAi31      o0602(.An(ori_ori_n627_), .B(ori_ori_n630_), .C(ori_ori_n628_), .Y(ori_ori_n631_));
  NO2        o0603(.A(ori_ori_n524_), .B(ori_ori_n180_), .Y(ori_ori_n632_));
  NA3        o0604(.A(ori_ori_n546_), .B(ori_ori_n278_), .C(ori_ori_n147_), .Y(ori_ori_n633_));
  NA2        o0605(.A(ori_ori_n502_), .B(ori_ori_n163_), .Y(ori_ori_n634_));
  NO3        o0606(.A(ori_ori_n389_), .B(ori_ori_n634_), .C(ori_ori_n86_), .Y(ori_ori_n635_));
  AOI210     o0607(.A0(ori_ori_n633_), .A1(ori_ori_n632_), .B0(ori_ori_n635_), .Y(ori_ori_n636_));
  AN3        o0608(.A(f), .B(d), .C(b), .Y(ori_ori_n637_));
  OAI210     o0609(.A0(ori_ori_n637_), .A1(ori_ori_n131_), .B0(n), .Y(ori_ori_n638_));
  NA3        o0610(.A(ori_ori_n502_), .B(ori_ori_n163_), .C(ori_ori_n219_), .Y(ori_ori_n639_));
  AOI210     o0611(.A0(ori_ori_n638_), .A1(ori_ori_n238_), .B0(ori_ori_n639_), .Y(ori_ori_n640_));
  NAi31      o0612(.An(m), .B(n), .C(k), .Y(ori_ori_n641_));
  INV        o0613(.A(ori_ori_n257_), .Y(ori_ori_n642_));
  OAI210     o0614(.A0(ori_ori_n642_), .A1(ori_ori_n640_), .B0(j), .Y(ori_ori_n643_));
  NA3        o0615(.A(ori_ori_n643_), .B(ori_ori_n636_), .C(ori_ori_n631_), .Y(ori_ori_n644_));
  NO4        o0616(.A(ori_ori_n644_), .B(ori_ori_n626_), .C(ori_ori_n614_), .D(ori_ori_n608_), .Y(ori_ori_n645_));
  NA2        o0617(.A(ori_ori_n376_), .B(ori_ori_n166_), .Y(ori_ori_n646_));
  NAi31      o0618(.An(g), .B(h), .C(f), .Y(ori_ori_n647_));
  OR3        o0619(.A(ori_ori_n647_), .B(ori_ori_n282_), .C(n), .Y(ori_ori_n648_));
  OA210      o0620(.A0(ori_ori_n526_), .A1(n), .B0(ori_ori_n577_), .Y(ori_ori_n649_));
  NA3        o0621(.A(ori_ori_n412_), .B(ori_ori_n122_), .C(ori_ori_n83_), .Y(ori_ori_n650_));
  OAI210     o0622(.A0(ori_ori_n649_), .A1(ori_ori_n90_), .B0(ori_ori_n650_), .Y(ori_ori_n651_));
  NOi21      o0623(.An(ori_ori_n648_), .B(ori_ori_n651_), .Y(ori_ori_n652_));
  AOI210     o0624(.A0(ori_ori_n652_), .A1(ori_ori_n646_), .B0(ori_ori_n520_), .Y(ori_ori_n653_));
  NO3        o0625(.A(g), .B(ori_ori_n218_), .C(ori_ori_n56_), .Y(ori_ori_n654_));
  NAi21      o0626(.An(h), .B(j), .Y(ori_ori_n655_));
  NO2        o0627(.A(ori_ori_n509_), .B(ori_ori_n86_), .Y(ori_ori_n656_));
  OAI210     o0628(.A0(ori_ori_n656_), .A1(ori_ori_n388_), .B0(ori_ori_n654_), .Y(ori_ori_n657_));
  OR2        o0629(.A(ori_ori_n71_), .B(ori_ori_n72_), .Y(ori_ori_n658_));
  NA3        o0630(.A(ori_ori_n517_), .B(ori_ori_n99_), .C(ori_ori_n98_), .Y(ori_ori_n659_));
  AN2        o0631(.A(h), .B(f), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n660_), .B(ori_ori_n37_), .Y(ori_ori_n661_));
  NA2        o0633(.A(ori_ori_n99_), .B(ori_ori_n46_), .Y(ori_ori_n662_));
  OAI220     o0634(.A0(ori_ori_n662_), .A1(ori_ori_n331_), .B0(ori_ori_n661_), .B1(ori_ori_n459_), .Y(ori_ori_n663_));
  AOI210     o0635(.A0(ori_ori_n562_), .A1(ori_ori_n424_), .B0(ori_ori_n49_), .Y(ori_ori_n664_));
  INV        o0636(.A(ori_ori_n663_), .Y(ori_ori_n665_));
  NA3        o0637(.A(ori_ori_n665_), .B(ori_ori_n659_), .C(ori_ori_n657_), .Y(ori_ori_n666_));
  NA2        o0638(.A(ori_ori_n133_), .B(ori_ori_n49_), .Y(ori_ori_n667_));
  AOI220     o0639(.A0(ori_ori_n667_), .A1(ori_ori_n523_), .B0(ori_ori_n358_), .B1(ori_ori_n114_), .Y(ori_ori_n668_));
  OA220      o0640(.A0(ori_ori_n668_), .A1(ori_ori_n543_), .B0(ori_ori_n356_), .B1(ori_ori_n112_), .Y(ori_ori_n669_));
  INV        o0641(.A(ori_ori_n669_), .Y(ori_ori_n670_));
  NO3        o0642(.A(ori_ori_n399_), .B(ori_ori_n196_), .C(ori_ori_n195_), .Y(ori_ori_n671_));
  NA2        o0643(.A(ori_ori_n671_), .B(ori_ori_n236_), .Y(ori_ori_n672_));
  NA3        o0644(.A(ori_ori_n672_), .B(ori_ori_n261_), .C(j), .Y(ori_ori_n673_));
  NO3        o0645(.A(ori_ori_n454_), .B(ori_ori_n177_), .C(i), .Y(ori_ori_n674_));
  NA2        o0646(.A(ori_ori_n458_), .B(ori_ori_n83_), .Y(ori_ori_n675_));
  NA3        o0647(.A(ori_ori_n673_), .B(ori_ori_n508_), .C(ori_ori_n397_), .Y(ori_ori_n676_));
  NO4        o0648(.A(ori_ori_n676_), .B(ori_ori_n670_), .C(ori_ori_n666_), .D(ori_ori_n653_), .Y(ori_ori_n677_));
  NA4        o0649(.A(ori_ori_n677_), .B(ori_ori_n645_), .C(ori_ori_n602_), .D(ori_ori_n572_), .Y(ori08));
  NO2        o0650(.A(k), .B(h), .Y(ori_ori_n679_));
  AO210      o0651(.A0(ori_ori_n259_), .A1(ori_ori_n442_), .B0(ori_ori_n679_), .Y(ori_ori_n680_));
  NO2        o0652(.A(ori_ori_n680_), .B(ori_ori_n300_), .Y(ori_ori_n681_));
  NA2        o0653(.A(ori_ori_n610_), .B(ori_ori_n83_), .Y(ori_ori_n682_));
  NA2        o0654(.A(ori_ori_n682_), .B(ori_ori_n454_), .Y(ori_ori_n683_));
  AOI210     o0655(.A0(ori_ori_n683_), .A1(ori_ori_n681_), .B0(ori_ori_n487_), .Y(ori_ori_n684_));
  NA2        o0656(.A(ori_ori_n83_), .B(ori_ori_n111_), .Y(ori_ori_n685_));
  NO2        o0657(.A(ori_ori_n685_), .B(ori_ori_n57_), .Y(ori_ori_n686_));
  NO4        o0658(.A(ori_ori_n374_), .B(ori_ori_n113_), .C(j), .D(ori_ori_n219_), .Y(ori_ori_n687_));
  NA2        o0659(.A(ori_ori_n687_), .B(ori_ori_n686_), .Y(ori_ori_n688_));
  AOI210     o0660(.A0(ori_ori_n569_), .A1(ori_ori_n159_), .B0(ori_ori_n83_), .Y(ori_ori_n689_));
  NA4        o0661(.A(ori_ori_n221_), .B(ori_ori_n142_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n690_));
  AN2        o0662(.A(l), .B(k), .Y(ori_ori_n691_));
  NA4        o0663(.A(ori_ori_n691_), .B(ori_ori_n109_), .C(ori_ori_n72_), .D(ori_ori_n219_), .Y(ori_ori_n692_));
  OAI210     o0664(.A0(ori_ori_n690_), .A1(g), .B0(ori_ori_n692_), .Y(ori_ori_n693_));
  NA2        o0665(.A(ori_ori_n693_), .B(ori_ori_n689_), .Y(ori_ori_n694_));
  NA4        o0666(.A(ori_ori_n694_), .B(ori_ori_n688_), .C(ori_ori_n684_), .D(ori_ori_n345_), .Y(ori_ori_n695_));
  NO2        o0667(.A(ori_ori_n38_), .B(ori_ori_n218_), .Y(ori_ori_n696_));
  AOI220     o0668(.A0(ori_ori_n612_), .A1(ori_ori_n344_), .B0(ori_ori_n696_), .B1(ori_ori_n559_), .Y(ori_ori_n697_));
  INV        o0669(.A(ori_ori_n697_), .Y(ori_ori_n698_));
  NO2        o0670(.A(ori_ori_n530_), .B(ori_ori_n35_), .Y(ori_ori_n699_));
  INV        o0671(.A(ori_ori_n699_), .Y(ori_ori_n700_));
  NO3        o0672(.A(ori_ori_n321_), .B(ori_ori_n132_), .C(ori_ori_n41_), .Y(ori_ori_n701_));
  NAi21      o0673(.An(ori_ori_n701_), .B(ori_ori_n692_), .Y(ori_ori_n702_));
  NA2        o0674(.A(ori_ori_n680_), .B(ori_ori_n137_), .Y(ori_ori_n703_));
  AOI220     o0675(.A0(ori_ori_n703_), .A1(ori_ori_n398_), .B0(ori_ori_n702_), .B1(ori_ori_n75_), .Y(ori_ori_n704_));
  OAI210     o0676(.A0(ori_ori_n700_), .A1(ori_ori_n86_), .B0(ori_ori_n704_), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n358_), .B(ori_ori_n43_), .Y(ori_ori_n706_));
  NA3        o0678(.A(ori_ori_n672_), .B(ori_ori_n333_), .C(ori_ori_n379_), .Y(ori_ori_n707_));
  NA3        o0679(.A(m), .B(l), .C(k), .Y(ori_ori_n708_));
  AOI210     o0680(.A0(ori_ori_n650_), .A1(ori_ori_n648_), .B0(ori_ori_n708_), .Y(ori_ori_n709_));
  NA3        o0681(.A(ori_ori_n114_), .B(k), .C(ori_ori_n86_), .Y(ori_ori_n710_));
  INV        o0682(.A(ori_ori_n709_), .Y(ori_ori_n711_));
  NA3        o0683(.A(ori_ori_n711_), .B(ori_ori_n707_), .C(ori_ori_n706_), .Y(ori_ori_n712_));
  NO4        o0684(.A(ori_ori_n712_), .B(ori_ori_n705_), .C(ori_ori_n698_), .D(ori_ori_n695_), .Y(ori_ori_n713_));
  NA2        o0685(.A(ori_ori_n612_), .B(ori_ori_n388_), .Y(ori_ori_n714_));
  NOi31      o0686(.An(g), .B(h), .C(f), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n624_), .B(ori_ori_n715_), .Y(ori_ori_n716_));
  AO210      o0688(.A0(ori_ori_n716_), .A1(ori_ori_n581_), .B0(ori_ori_n531_), .Y(ori_ori_n717_));
  NO3        o0689(.A(ori_ori_n392_), .B(ori_ori_n518_), .C(h), .Y(ori_ori_n718_));
  AOI210     o0690(.A0(ori_ori_n718_), .A1(ori_ori_n114_), .B0(ori_ori_n497_), .Y(ori_ori_n719_));
  NA4        o0691(.A(ori_ori_n719_), .B(ori_ori_n717_), .C(ori_ori_n714_), .D(ori_ori_n258_), .Y(ori_ori_n720_));
  NA2        o0692(.A(ori_ori_n691_), .B(ori_ori_n72_), .Y(ori_ori_n721_));
  NO4        o0693(.A(ori_ori_n671_), .B(ori_ori_n177_), .C(n), .D(i), .Y(ori_ori_n722_));
  NOi21      o0694(.An(h), .B(j), .Y(ori_ori_n723_));
  NA2        o0695(.A(ori_ori_n723_), .B(f), .Y(ori_ori_n724_));
  NO2        o0696(.A(ori_ori_n724_), .B(ori_ori_n252_), .Y(ori_ori_n725_));
  NO3        o0697(.A(ori_ori_n725_), .B(ori_ori_n722_), .C(ori_ori_n674_), .Y(ori_ori_n726_));
  OAI220     o0698(.A0(ori_ori_n726_), .A1(ori_ori_n721_), .B0(ori_ori_n583_), .B1(ori_ori_n62_), .Y(ori_ori_n727_));
  AOI210     o0699(.A0(ori_ori_n720_), .A1(l), .B0(ori_ori_n727_), .Y(ori_ori_n728_));
  NO2        o0700(.A(j), .B(i), .Y(ori_ori_n729_));
  NA3        o0701(.A(ori_ori_n729_), .B(ori_ori_n79_), .C(l), .Y(ori_ori_n730_));
  NA2        o0702(.A(ori_ori_n729_), .B(ori_ori_n33_), .Y(ori_ori_n731_));
  NA2        o0703(.A(ori_ori_n417_), .B(ori_ori_n122_), .Y(ori_ori_n732_));
  OA220      o0704(.A0(ori_ori_n732_), .A1(ori_ori_n731_), .B0(ori_ori_n730_), .B1(ori_ori_n579_), .Y(ori_ori_n733_));
  NO3        o0705(.A(ori_ori_n154_), .B(ori_ori_n49_), .C(ori_ori_n111_), .Y(ori_ori_n734_));
  NO2        o0706(.A(ori_ori_n716_), .B(ori_ori_n62_), .Y(ori_ori_n735_));
  INV        o0707(.A(j), .Y(ori_ori_n736_));
  NO3        o0708(.A(ori_ori_n300_), .B(ori_ori_n736_), .C(ori_ori_n40_), .Y(ori_ori_n737_));
  AOI210     o0709(.A0(ori_ori_n523_), .A1(n), .B0(ori_ori_n545_), .Y(ori_ori_n738_));
  NA2        o0710(.A(ori_ori_n738_), .B(ori_ori_n548_), .Y(ori_ori_n739_));
  AN3        o0711(.A(ori_ori_n739_), .B(ori_ori_n737_), .C(ori_ori_n98_), .Y(ori_ori_n740_));
  NO3        o0712(.A(ori_ori_n177_), .B(ori_ori_n387_), .C(ori_ori_n113_), .Y(ori_ori_n741_));
  AOI220     o0713(.A0(ori_ori_n741_), .A1(ori_ori_n253_), .B0(ori_ori_n605_), .B1(ori_ori_n311_), .Y(ori_ori_n742_));
  NAi31      o0714(.An(ori_ori_n598_), .B(ori_ori_n92_), .C(ori_ori_n83_), .Y(ori_ori_n743_));
  NA2        o0715(.A(ori_ori_n743_), .B(ori_ori_n742_), .Y(ori_ori_n744_));
  NO2        o0716(.A(ori_ori_n300_), .B(ori_ori_n137_), .Y(ori_ori_n745_));
  AOI220     o0717(.A0(ori_ori_n745_), .A1(ori_ori_n612_), .B0(ori_ori_n701_), .B1(ori_ori_n689_), .Y(ori_ori_n746_));
  NO2        o0718(.A(ori_ori_n708_), .B(ori_ori_n90_), .Y(ori_ori_n747_));
  NA2        o0719(.A(ori_ori_n747_), .B(ori_ori_n578_), .Y(ori_ori_n748_));
  NA2        o0720(.A(ori_ori_n748_), .B(ori_ori_n746_), .Y(ori_ori_n749_));
  OR4        o0721(.A(ori_ori_n749_), .B(ori_ori_n744_), .C(ori_ori_n740_), .D(ori_ori_n735_), .Y(ori_ori_n750_));
  NA3        o0722(.A(ori_ori_n738_), .B(ori_ori_n548_), .C(ori_ori_n547_), .Y(ori_ori_n751_));
  NA4        o0723(.A(ori_ori_n751_), .B(ori_ori_n221_), .C(ori_ori_n442_), .D(ori_ori_n34_), .Y(ori_ori_n752_));
  NO3        o0724(.A(ori_ori_n481_), .B(ori_ori_n431_), .C(j), .Y(ori_ori_n753_));
  OAI220     o0725(.A0(ori_ori_n690_), .A1(ori_ori_n682_), .B0(ori_ori_n331_), .B1(ori_ori_n38_), .Y(ori_ori_n754_));
  AOI210     o0726(.A0(ori_ori_n753_), .A1(ori_ori_n265_), .B0(ori_ori_n754_), .Y(ori_ori_n755_));
  NA3        o0727(.A(ori_ori_n538_), .B(ori_ori_n297_), .C(h), .Y(ori_ori_n756_));
  NO2        o0728(.A(ori_ori_n91_), .B(ori_ori_n47_), .Y(ori_ori_n757_));
  OAI220     o0729(.A0(ori_ori_n756_), .A1(ori_ori_n594_), .B0(ori_ori_n730_), .B1(ori_ori_n658_), .Y(ori_ori_n758_));
  AOI210     o0730(.A0(ori_ori_n757_), .A1(ori_ori_n630_), .B0(ori_ori_n758_), .Y(ori_ori_n759_));
  NA3        o0731(.A(ori_ori_n759_), .B(ori_ori_n755_), .C(ori_ori_n752_), .Y(ori_ori_n760_));
  NA2        o0732(.A(ori_ori_n747_), .B(ori_ori_n244_), .Y(ori_ori_n761_));
  NO2        o0733(.A(ori_ori_n649_), .B(ori_ori_n72_), .Y(ori_ori_n762_));
  AOI210     o0734(.A0(ori_ori_n753_), .A1(ori_ori_n762_), .B0(ori_ori_n335_), .Y(ori_ori_n763_));
  OAI210     o0735(.A0(ori_ori_n708_), .A1(ori_ori_n647_), .B0(ori_ori_n513_), .Y(ori_ori_n764_));
  NA3        o0736(.A(ori_ori_n256_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n765_));
  AOI220     o0737(.A0(ori_ori_n593_), .A1(ori_ori_n29_), .B0(ori_ori_n458_), .B1(ori_ori_n83_), .Y(ori_ori_n766_));
  NA2        o0738(.A(ori_ori_n766_), .B(ori_ori_n765_), .Y(ori_ori_n767_));
  NA2        o0739(.A(ori_ori_n767_), .B(ori_ori_n764_), .Y(ori_ori_n768_));
  NA3        o0740(.A(ori_ori_n768_), .B(ori_ori_n763_), .C(ori_ori_n761_), .Y(ori_ori_n769_));
  NOi41      o0741(.An(ori_ori_n733_), .B(ori_ori_n769_), .C(ori_ori_n760_), .D(ori_ori_n750_), .Y(ori_ori_n770_));
  OR3        o0742(.A(ori_ori_n690_), .B(ori_ori_n238_), .C(g), .Y(ori_ori_n771_));
  NO3        o0743(.A(ori_ori_n340_), .B(ori_ori_n302_), .C(ori_ori_n113_), .Y(ori_ori_n772_));
  NA2        o0744(.A(ori_ori_n772_), .B(ori_ori_n739_), .Y(ori_ori_n773_));
  NO3        o0745(.A(ori_ori_n518_), .B(ori_ori_n93_), .C(h), .Y(ori_ori_n774_));
  NA2        o0746(.A(ori_ori_n774_), .B(ori_ori_n686_), .Y(ori_ori_n775_));
  NA4        o0747(.A(ori_ori_n775_), .B(ori_ori_n773_), .C(ori_ori_n771_), .D(ori_ori_n400_), .Y(ori_ori_n776_));
  OR2        o0748(.A(ori_ori_n647_), .B(ori_ori_n91_), .Y(ori_ori_n777_));
  NOi31      o0749(.An(b), .B(d), .C(a), .Y(ori_ori_n778_));
  NO2        o0750(.A(ori_ori_n778_), .B(ori_ori_n591_), .Y(ori_ori_n779_));
  NO2        o0751(.A(ori_ori_n779_), .B(n), .Y(ori_ori_n780_));
  NO2        o0752(.A(ori_ori_n756_), .B(ori_ori_n592_), .Y(ori_ori_n781_));
  NO2        o0753(.A(ori_ori_n546_), .B(ori_ori_n83_), .Y(ori_ori_n782_));
  NO3        o0754(.A(ori_ori_n611_), .B(ori_ori_n329_), .C(ori_ori_n118_), .Y(ori_ori_n783_));
  NOi21      o0755(.An(ori_ori_n783_), .B(ori_ori_n164_), .Y(ori_ori_n784_));
  AOI210     o0756(.A0(ori_ori_n772_), .A1(ori_ori_n782_), .B0(ori_ori_n784_), .Y(ori_ori_n785_));
  OAI210     o0757(.A0(ori_ori_n690_), .A1(ori_ori_n389_), .B0(ori_ori_n785_), .Y(ori_ori_n786_));
  NO2        o0758(.A(ori_ori_n671_), .B(n), .Y(ori_ori_n787_));
  AOI220     o0759(.A0(ori_ori_n745_), .A1(ori_ori_n654_), .B0(ori_ori_n787_), .B1(ori_ori_n681_), .Y(ori_ori_n788_));
  NO2        o0760(.A(ori_ori_n326_), .B(ori_ori_n243_), .Y(ori_ori_n789_));
  OAI210     o0761(.A0(ori_ori_n95_), .A1(ori_ori_n92_), .B0(ori_ori_n789_), .Y(ori_ori_n790_));
  NA2        o0762(.A(ori_ori_n122_), .B(ori_ori_n83_), .Y(ori_ori_n791_));
  AOI210     o0763(.A0(ori_ori_n421_), .A1(ori_ori_n413_), .B0(ori_ori_n791_), .Y(ori_ori_n792_));
  NAi21      o0764(.An(ori_ori_n792_), .B(ori_ori_n790_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n279_), .B(i), .Y(ori_ori_n794_));
  OAI210     o0766(.A0(ori_ori_n586_), .A1(ori_ori_n585_), .B0(ori_ori_n359_), .Y(ori_ori_n795_));
  NAi31      o0767(.An(ori_ori_n793_), .B(ori_ori_n795_), .C(ori_ori_n788_), .Y(ori_ori_n796_));
  NO4        o0768(.A(ori_ori_n796_), .B(ori_ori_n786_), .C(ori_ori_n781_), .D(ori_ori_n776_), .Y(ori_ori_n797_));
  NA4        o0769(.A(ori_ori_n797_), .B(ori_ori_n770_), .C(ori_ori_n728_), .D(ori_ori_n713_), .Y(ori09));
  INV        o0770(.A(ori_ori_n123_), .Y(ori_ori_n799_));
  NA2        o0771(.A(f), .B(e), .Y(ori_ori_n800_));
  NO2        o0772(.A(ori_ori_n231_), .B(ori_ori_n113_), .Y(ori_ori_n801_));
  NA2        o0773(.A(ori_ori_n801_), .B(g), .Y(ori_ori_n802_));
  NA4        o0774(.A(ori_ori_n314_), .B(ori_ori_n467_), .C(ori_ori_n268_), .D(ori_ori_n120_), .Y(ori_ori_n803_));
  AOI210     o0775(.A0(ori_ori_n803_), .A1(g), .B0(ori_ori_n464_), .Y(ori_ori_n804_));
  AOI210     o0776(.A0(ori_ori_n804_), .A1(ori_ori_n802_), .B0(ori_ori_n800_), .Y(ori_ori_n805_));
  NA2        o0777(.A(ori_ori_n435_), .B(e), .Y(ori_ori_n806_));
  NO2        o0778(.A(ori_ori_n806_), .B(ori_ori_n505_), .Y(ori_ori_n807_));
  AOI210     o0779(.A0(ori_ori_n805_), .A1(ori_ori_n799_), .B0(ori_ori_n807_), .Y(ori_ori_n808_));
  NO2        o0780(.A(ori_ori_n208_), .B(ori_ori_n218_), .Y(ori_ori_n809_));
  NA3        o0781(.A(m), .B(l), .C(i), .Y(ori_ori_n810_));
  OAI220     o0782(.A0(ori_ori_n580_), .A1(ori_ori_n810_), .B0(ori_ori_n349_), .B1(ori_ori_n519_), .Y(ori_ori_n811_));
  NA4        o0783(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(g), .D(f), .Y(ori_ori_n812_));
  BUFFER     o0784(.A(ori_ori_n811_), .Y(ori_ori_n813_));
  OR2        o0785(.A(ori_ori_n813_), .B(ori_ori_n809_), .Y(ori_ori_n814_));
  NA3        o0786(.A(ori_ori_n777_), .B(ori_ori_n561_), .C(ori_ori_n513_), .Y(ori_ori_n815_));
  OA210      o0787(.A0(ori_ori_n815_), .A1(ori_ori_n814_), .B0(ori_ori_n780_), .Y(ori_ori_n816_));
  INV        o0788(.A(ori_ori_n338_), .Y(ori_ori_n817_));
  NO2        o0789(.A(ori_ori_n128_), .B(ori_ori_n126_), .Y(ori_ori_n818_));
  NOi31      o0790(.An(k), .B(m), .C(l), .Y(ori_ori_n819_));
  NO2        o0791(.A(ori_ori_n339_), .B(ori_ori_n819_), .Y(ori_ori_n820_));
  AOI210     o0792(.A0(ori_ori_n820_), .A1(ori_ori_n818_), .B0(ori_ori_n589_), .Y(ori_ori_n821_));
  NA2        o0793(.A(ori_ori_n765_), .B(ori_ori_n331_), .Y(ori_ori_n822_));
  NA2        o0794(.A(ori_ori_n341_), .B(ori_ori_n342_), .Y(ori_ori_n823_));
  OAI210     o0795(.A0(ori_ori_n208_), .A1(ori_ori_n218_), .B0(ori_ori_n823_), .Y(ori_ori_n824_));
  AOI220     o0796(.A0(ori_ori_n824_), .A1(ori_ori_n822_), .B0(ori_ori_n821_), .B1(ori_ori_n817_), .Y(ori_ori_n825_));
  NA2        o0797(.A(ori_ori_n680_), .B(ori_ori_n137_), .Y(ori_ori_n826_));
  NA3        o0798(.A(ori_ori_n826_), .B(ori_ori_n193_), .C(ori_ori_n31_), .Y(ori_ori_n827_));
  NA4        o0799(.A(ori_ori_n827_), .B(ori_ori_n825_), .C(ori_ori_n613_), .D(ori_ori_n81_), .Y(ori_ori_n828_));
  NO2        o0800(.A(ori_ori_n576_), .B(ori_ori_n493_), .Y(ori_ori_n829_));
  NA2        o0801(.A(ori_ori_n829_), .B(ori_ori_n193_), .Y(ori_ori_n830_));
  NOi21      o0802(.An(f), .B(d), .Y(ori_ori_n831_));
  NA2        o0803(.A(ori_ori_n831_), .B(m), .Y(ori_ori_n832_));
  NO2        o0804(.A(ori_ori_n832_), .B(ori_ori_n52_), .Y(ori_ori_n833_));
  NOi32      o0805(.An(g), .Bn(f), .C(d), .Y(ori_ori_n834_));
  NA4        o0806(.A(ori_ori_n834_), .B(ori_ori_n593_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n835_));
  NOi21      o0807(.An(ori_ori_n315_), .B(ori_ori_n835_), .Y(ori_ori_n836_));
  AOI210     o0808(.A0(ori_ori_n833_), .A1(ori_ori_n536_), .B0(ori_ori_n836_), .Y(ori_ori_n837_));
  NA2        o0809(.A(ori_ori_n268_), .B(ori_ori_n120_), .Y(ori_ori_n838_));
  AN2        o0810(.A(f), .B(d), .Y(ori_ori_n839_));
  NA3        o0811(.A(ori_ori_n472_), .B(ori_ori_n839_), .C(ori_ori_n83_), .Y(ori_ori_n840_));
  NO3        o0812(.A(ori_ori_n840_), .B(ori_ori_n72_), .C(ori_ori_n219_), .Y(ori_ori_n841_));
  NA2        o0813(.A(ori_ori_n838_), .B(ori_ori_n841_), .Y(ori_ori_n842_));
  NAi41      o0814(.An(ori_ori_n486_), .B(ori_ori_n842_), .C(ori_ori_n837_), .D(ori_ori_n830_), .Y(ori_ori_n843_));
  NO4        o0815(.A(ori_ori_n611_), .B(ori_ori_n133_), .C(ori_ori_n329_), .D(ori_ori_n155_), .Y(ori_ori_n844_));
  NO2        o0816(.A(ori_ori_n641_), .B(ori_ori_n329_), .Y(ori_ori_n845_));
  NO2        o0817(.A(ori_ori_n844_), .B(ori_ori_n240_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n591_), .B(ori_ori_n83_), .Y(ori_ori_n847_));
  NO2        o0819(.A(ori_ori_n823_), .B(ori_ori_n847_), .Y(ori_ori_n848_));
  NA3        o0820(.A(ori_ori_n163_), .B(ori_ori_n109_), .C(ori_ori_n108_), .Y(ori_ori_n849_));
  OAI220     o0821(.A0(ori_ori_n840_), .A1(ori_ori_n426_), .B0(ori_ori_n338_), .B1(ori_ori_n849_), .Y(ori_ori_n850_));
  NO3        o0822(.A(ori_ori_n850_), .B(ori_ori_n848_), .C(ori_ori_n309_), .Y(ori_ori_n851_));
  NA2        o0823(.A(c), .B(ori_ori_n117_), .Y(ori_ori_n852_));
  NO2        o0824(.A(ori_ori_n852_), .B(ori_ori_n404_), .Y(ori_ori_n853_));
  NA3        o0825(.A(ori_ori_n853_), .B(ori_ori_n504_), .C(f), .Y(ori_ori_n854_));
  OR2        o0826(.A(ori_ori_n647_), .B(ori_ori_n532_), .Y(ori_ori_n855_));
  INV        o0827(.A(ori_ori_n855_), .Y(ori_ori_n856_));
  NA2        o0828(.A(ori_ori_n779_), .B(ori_ori_n112_), .Y(ori_ori_n857_));
  NA2        o0829(.A(ori_ori_n857_), .B(ori_ori_n856_), .Y(ori_ori_n858_));
  NA4        o0830(.A(ori_ori_n858_), .B(ori_ori_n854_), .C(ori_ori_n851_), .D(ori_ori_n846_), .Y(ori_ori_n859_));
  NO4        o0831(.A(ori_ori_n859_), .B(ori_ori_n843_), .C(ori_ori_n828_), .D(ori_ori_n816_), .Y(ori_ori_n860_));
  NA2        o0832(.A(ori_ori_n113_), .B(j), .Y(ori_ori_n861_));
  NO2        o0833(.A(ori_ori_n331_), .B(ori_ori_n812_), .Y(ori_ori_n862_));
  NO2        o0834(.A(ori_ori_n137_), .B(ori_ori_n133_), .Y(ori_ori_n863_));
  NO2        o0835(.A(ori_ori_n236_), .B(ori_ori_n230_), .Y(ori_ori_n864_));
  AOI220     o0836(.A0(ori_ori_n864_), .A1(ori_ori_n233_), .B0(ori_ori_n307_), .B1(ori_ori_n863_), .Y(ori_ori_n865_));
  NO2        o0837(.A(ori_ori_n426_), .B(ori_ori_n800_), .Y(ori_ori_n866_));
  NA2        o0838(.A(ori_ori_n866_), .B(ori_ori_n553_), .Y(ori_ori_n867_));
  NA2        o0839(.A(ori_ori_n867_), .B(ori_ori_n865_), .Y(ori_ori_n868_));
  NA2        o0840(.A(e), .B(d), .Y(ori_ori_n869_));
  OAI220     o0841(.A0(ori_ori_n869_), .A1(c), .B0(ori_ori_n326_), .B1(d), .Y(ori_ori_n870_));
  NA3        o0842(.A(ori_ori_n870_), .B(ori_ori_n447_), .C(ori_ori_n502_), .Y(ori_ori_n871_));
  AOI210     o0843(.A0(ori_ori_n509_), .A1(ori_ori_n184_), .B0(ori_ori_n236_), .Y(ori_ori_n872_));
  AOI210     o0844(.A0(ori_ori_n612_), .A1(ori_ori_n344_), .B0(ori_ori_n872_), .Y(ori_ori_n873_));
  NA2        o0845(.A(ori_ori_n290_), .B(ori_ori_n168_), .Y(ori_ori_n874_));
  NA2        o0846(.A(ori_ori_n841_), .B(ori_ori_n874_), .Y(ori_ori_n875_));
  NA3        o0847(.A(ori_ori_n171_), .B(ori_ori_n84_), .C(ori_ori_n34_), .Y(ori_ori_n876_));
  NA4        o0848(.A(ori_ori_n876_), .B(ori_ori_n875_), .C(ori_ori_n873_), .D(ori_ori_n871_), .Y(ori_ori_n877_));
  NO3        o0849(.A(ori_ori_n877_), .B(ori_ori_n868_), .C(ori_ori_n862_), .Y(ori_ori_n878_));
  OR2        o0850(.A(ori_ori_n682_), .B(ori_ori_n222_), .Y(ori_ori_n879_));
  NO2        o0851(.A(ori_ori_n611_), .B(ori_ori_n61_), .Y(ori_ori_n880_));
  AOI220     o0852(.A0(ori_ori_n880_), .A1(ori_ori_n845_), .B0(ori_ori_n603_), .B1(ori_ori_n610_), .Y(ori_ori_n881_));
  OAI210     o0853(.A0(ori_ori_n806_), .A1(ori_ori_n174_), .B0(ori_ori_n881_), .Y(ori_ori_n882_));
  OAI210     o0854(.A0(ori_ori_n801_), .A1(ori_ori_n874_), .B0(ori_ori_n834_), .Y(ori_ori_n883_));
  NO2        o0855(.A(ori_ori_n883_), .B(ori_ori_n594_), .Y(ori_ori_n884_));
  AN2        o0856(.A(ori_ori_n822_), .B(ori_ori_n811_), .Y(ori_ori_n885_));
  NO3        o0857(.A(ori_ori_n885_), .B(ori_ori_n884_), .C(ori_ori_n882_), .Y(ori_ori_n886_));
  AO220      o0858(.A0(ori_ori_n447_), .A1(ori_ori_n723_), .B0(ori_ori_n179_), .B1(f), .Y(ori_ori_n887_));
  OAI210     o0859(.A0(ori_ori_n887_), .A1(ori_ori_n450_), .B0(ori_ori_n870_), .Y(ori_ori_n888_));
  NO2        o0860(.A(ori_ori_n433_), .B(ori_ori_n70_), .Y(ori_ori_n889_));
  OAI210     o0861(.A0(ori_ori_n815_), .A1(ori_ori_n889_), .B0(ori_ori_n686_), .Y(ori_ori_n890_));
  AN4        o0862(.A(ori_ori_n890_), .B(ori_ori_n888_), .C(ori_ori_n886_), .D(ori_ori_n879_), .Y(ori_ori_n891_));
  NA4        o0863(.A(ori_ori_n891_), .B(ori_ori_n878_), .C(ori_ori_n860_), .D(ori_ori_n808_), .Y(ori12));
  NO2        o0864(.A(ori_ori_n445_), .B(c), .Y(ori_ori_n893_));
  NO4        o0865(.A(ori_ori_n434_), .B(ori_ori_n259_), .C(ori_ori_n573_), .D(ori_ori_n219_), .Y(ori_ori_n894_));
  NA2        o0866(.A(ori_ori_n894_), .B(ori_ori_n893_), .Y(ori_ori_n895_));
  NA2        o0867(.A(ori_ori_n536_), .B(ori_ori_n889_), .Y(ori_ori_n896_));
  NO2        o0868(.A(ori_ori_n445_), .B(ori_ori_n117_), .Y(ori_ori_n897_));
  NO2        o0869(.A(ori_ori_n818_), .B(ori_ori_n349_), .Y(ori_ori_n898_));
  NO2        o0870(.A(ori_ori_n647_), .B(ori_ori_n374_), .Y(ori_ori_n899_));
  AOI220     o0871(.A0(ori_ori_n899_), .A1(ori_ori_n534_), .B0(ori_ori_n898_), .B1(ori_ori_n897_), .Y(ori_ori_n900_));
  NA3        o0872(.A(ori_ori_n900_), .B(ori_ori_n896_), .C(ori_ori_n895_), .Y(ori_ori_n901_));
  AOI210     o0873(.A0(ori_ori_n239_), .A1(ori_ori_n337_), .B0(ori_ori_n205_), .Y(ori_ori_n902_));
  OR2        o0874(.A(ori_ori_n902_), .B(ori_ori_n894_), .Y(ori_ori_n903_));
  AOI210     o0875(.A0(ori_ori_n334_), .A1(ori_ori_n385_), .B0(ori_ori_n219_), .Y(ori_ori_n904_));
  OAI210     o0876(.A0(ori_ori_n904_), .A1(ori_ori_n903_), .B0(ori_ori_n399_), .Y(ori_ori_n905_));
  NO2        o0877(.A(ori_ori_n627_), .B(ori_ori_n270_), .Y(ori_ori_n906_));
  NO2        o0878(.A(ori_ori_n580_), .B(ori_ori_n810_), .Y(ori_ori_n907_));
  AOI220     o0879(.A0(ori_ori_n907_), .A1(ori_ori_n559_), .B0(ori_ori_n789_), .B1(ori_ori_n906_), .Y(ori_ori_n908_));
  NO2        o0880(.A(ori_ori_n154_), .B(ori_ori_n243_), .Y(ori_ori_n909_));
  NA3        o0881(.A(ori_ori_n909_), .B(ori_ori_n246_), .C(i), .Y(ori_ori_n910_));
  NA3        o0882(.A(ori_ori_n910_), .B(ori_ori_n908_), .C(ori_ori_n905_), .Y(ori_ori_n911_));
  OR2        o0883(.A(ori_ori_n327_), .B(ori_ori_n897_), .Y(ori_ori_n912_));
  NA2        o0884(.A(ori_ori_n912_), .B(ori_ori_n350_), .Y(ori_ori_n913_));
  NO3        o0885(.A(ori_ori_n133_), .B(ori_ori_n155_), .C(ori_ori_n219_), .Y(ori_ori_n914_));
  NA2        o0886(.A(ori_ori_n914_), .B(ori_ori_n523_), .Y(ori_ori_n915_));
  NA4        o0887(.A(ori_ori_n435_), .B(ori_ori_n432_), .C(ori_ori_n185_), .D(g), .Y(ori_ori_n916_));
  NA3        o0888(.A(ori_ori_n916_), .B(ori_ori_n915_), .C(ori_ori_n913_), .Y(ori_ori_n917_));
  NO3        o0889(.A(ori_ori_n652_), .B(ori_ori_n91_), .C(ori_ori_n45_), .Y(ori_ori_n918_));
  NO4        o0890(.A(ori_ori_n918_), .B(ori_ori_n917_), .C(ori_ori_n911_), .D(ori_ori_n901_), .Y(ori_ori_n919_));
  NO2        o0891(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n920_));
  INV        o0892(.A(ori_ori_n71_), .Y(ori_ori_n921_));
  NA2        o0893(.A(ori_ori_n546_), .B(ori_ori_n147_), .Y(ori_ori_n922_));
  NOi21      o0894(.An(ori_ori_n34_), .B(ori_ori_n641_), .Y(ori_ori_n923_));
  AOI220     o0895(.A0(ori_ori_n923_), .A1(ori_ori_n922_), .B0(ori_ori_n921_), .B1(ori_ori_n920_), .Y(ori_ori_n924_));
  OAI210     o0896(.A0(ori_ori_n257_), .A1(ori_ori_n45_), .B0(ori_ori_n924_), .Y(ori_ori_n925_));
  INV        o0897(.A(ori_ori_n325_), .Y(ori_ori_n926_));
  NO2        o0898(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n927_));
  NO2        o0899(.A(ori_ori_n500_), .B(ori_ori_n302_), .Y(ori_ori_n928_));
  INV        o0900(.A(ori_ori_n928_), .Y(ori_ori_n929_));
  NO2        o0901(.A(ori_ori_n929_), .B(ori_ori_n147_), .Y(ori_ori_n930_));
  INV        o0902(.A(ori_ori_n361_), .Y(ori_ori_n931_));
  NO4        o0903(.A(ori_ori_n931_), .B(ori_ori_n930_), .C(ori_ori_n926_), .D(ori_ori_n925_), .Y(ori_ori_n932_));
  NA2        o0904(.A(ori_ori_n344_), .B(g), .Y(ori_ori_n933_));
  NA2        o0905(.A(ori_ori_n166_), .B(i), .Y(ori_ori_n934_));
  NO2        o0906(.A(ori_ori_n934_), .B(ori_ori_n91_), .Y(ori_ori_n935_));
  AOI210     o0907(.A0(ori_ori_n415_), .A1(ori_ori_n37_), .B0(ori_ori_n935_), .Y(ori_ori_n936_));
  NO2        o0908(.A(ori_ori_n147_), .B(ori_ori_n83_), .Y(ori_ori_n937_));
  OR2        o0909(.A(ori_ori_n937_), .B(ori_ori_n545_), .Y(ori_ori_n938_));
  NA2        o0910(.A(ori_ori_n546_), .B(ori_ori_n377_), .Y(ori_ori_n939_));
  AOI210     o0911(.A0(ori_ori_n939_), .A1(n), .B0(ori_ori_n938_), .Y(ori_ori_n940_));
  OAI220     o0912(.A0(ori_ori_n940_), .A1(ori_ori_n933_), .B0(ori_ori_n936_), .B1(ori_ori_n331_), .Y(ori_ori_n941_));
  NA3        o0913(.A(ori_ori_n341_), .B(ori_ori_n616_), .C(i), .Y(ori_ori_n942_));
  OAI210     o0914(.A0(ori_ori_n433_), .A1(ori_ori_n314_), .B0(ori_ori_n942_), .Y(ori_ori_n943_));
  NA2        o0915(.A(ori_ori_n943_), .B(ori_ori_n664_), .Y(ori_ori_n944_));
  NA3        o0916(.A(ori_ori_n328_), .B(ori_ori_n119_), .C(g), .Y(ori_ori_n945_));
  AOI210     o0917(.A0(ori_ori_n661_), .A1(ori_ori_n945_), .B0(m), .Y(ori_ori_n946_));
  OAI210     o0918(.A0(ori_ori_n946_), .A1(ori_ori_n898_), .B0(ori_ori_n327_), .Y(ori_ori_n947_));
  NA2        o0919(.A(ori_ori_n675_), .B(ori_ori_n847_), .Y(ori_ori_n948_));
  INV        o0920(.A(ori_ori_n812_), .Y(ori_ori_n949_));
  NA2        o0921(.A(ori_ori_n949_), .B(ori_ori_n948_), .Y(ori_ori_n950_));
  NA3        o0922(.A(ori_ori_n950_), .B(ori_ori_n947_), .C(ori_ori_n944_), .Y(ori_ori_n951_));
  NO2        o0923(.A(ori_ori_n374_), .B(ori_ori_n90_), .Y(ori_ori_n952_));
  OAI210     o0924(.A0(ori_ori_n952_), .A1(ori_ori_n906_), .B0(ori_ori_n244_), .Y(ori_ori_n953_));
  NA2        o0925(.A(ori_ori_n651_), .B(ori_ori_n87_), .Y(ori_ori_n954_));
  NO2        o0926(.A(ori_ori_n453_), .B(ori_ori_n219_), .Y(ori_ori_n955_));
  AOI220     o0927(.A0(ori_ori_n955_), .A1(ori_ori_n378_), .B0(ori_ori_n912_), .B1(ori_ori_n223_), .Y(ori_ori_n956_));
  NA2        o0928(.A(ori_ori_n578_), .B(ori_ori_n89_), .Y(ori_ori_n957_));
  NA4        o0929(.A(ori_ori_n957_), .B(ori_ori_n956_), .C(ori_ori_n954_), .D(ori_ori_n953_), .Y(ori_ori_n958_));
  AOI210     o0930(.A0(ori_ori_n416_), .A1(ori_ori_n408_), .B0(ori_ori_n791_), .Y(ori_ori_n959_));
  OAI210     o0931(.A0(ori_ori_n364_), .A1(ori_ori_n363_), .B0(ori_ori_n110_), .Y(ori_ori_n960_));
  AOI210     o0932(.A0(ori_ori_n960_), .A1(ori_ori_n527_), .B0(ori_ori_n959_), .Y(ori_ori_n961_));
  NA2        o0933(.A(ori_ori_n946_), .B(ori_ori_n897_), .Y(ori_ori_n962_));
  NO3        o0934(.A(ori_ori_n861_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n963_));
  AOI220     o0935(.A0(ori_ori_n963_), .A1(ori_ori_n615_), .B0(ori_ori_n632_), .B1(ori_ori_n523_), .Y(ori_ori_n964_));
  NA3        o0936(.A(ori_ori_n964_), .B(ori_ori_n962_), .C(ori_ori_n961_), .Y(ori_ori_n965_));
  NO4        o0937(.A(ori_ori_n965_), .B(ori_ori_n958_), .C(ori_ori_n951_), .D(ori_ori_n941_), .Y(ori_ori_n966_));
  NAi31      o0938(.An(ori_ori_n143_), .B(ori_ori_n417_), .C(n), .Y(ori_ori_n967_));
  NO3        o0939(.A(ori_ori_n126_), .B(ori_ori_n339_), .C(ori_ori_n819_), .Y(ori_ori_n968_));
  NO2        o0940(.A(ori_ori_n968_), .B(ori_ori_n967_), .Y(ori_ori_n969_));
  NO3        o0941(.A(ori_ori_n279_), .B(ori_ori_n143_), .C(ori_ori_n404_), .Y(ori_ori_n970_));
  AOI210     o0942(.A0(ori_ori_n970_), .A1(ori_ori_n494_), .B0(ori_ori_n969_), .Y(ori_ori_n971_));
  NA2        o0943(.A(ori_ori_n487_), .B(i), .Y(ori_ori_n972_));
  NA2        o0944(.A(ori_ori_n972_), .B(ori_ori_n971_), .Y(ori_ori_n973_));
  NA2        o0945(.A(ori_ori_n236_), .B(ori_ori_n175_), .Y(ori_ori_n974_));
  NO3        o0946(.A(ori_ori_n311_), .B(ori_ori_n435_), .C(ori_ori_n179_), .Y(ori_ori_n975_));
  NOi31      o0947(.An(ori_ori_n974_), .B(ori_ori_n975_), .C(ori_ori_n219_), .Y(ori_ori_n976_));
  NAi21      o0948(.An(ori_ori_n546_), .B(ori_ori_n955_), .Y(ori_ori_n977_));
  NA2        o0949(.A(ori_ori_n478_), .B(g), .Y(ori_ori_n978_));
  NA2        o0950(.A(ori_ori_n978_), .B(ori_ori_n977_), .Y(ori_ori_n979_));
  OAI220     o0951(.A0(ori_ori_n967_), .A1(ori_ori_n239_), .B0(ori_ori_n942_), .B1(ori_ori_n592_), .Y(ori_ori_n980_));
  NO2        o0952(.A(ori_ori_n648_), .B(ori_ori_n374_), .Y(ori_ori_n981_));
  NA2        o0953(.A(ori_ori_n902_), .B(ori_ori_n893_), .Y(ori_ori_n982_));
  OAI220     o0954(.A0(ori_ori_n899_), .A1(ori_ori_n907_), .B0(ori_ori_n536_), .B1(ori_ori_n425_), .Y(ori_ori_n983_));
  NA3        o0955(.A(ori_ori_n983_), .B(ori_ori_n982_), .C(ori_ori_n609_), .Y(ori_ori_n984_));
  OAI210     o0956(.A0(ori_ori_n902_), .A1(ori_ori_n894_), .B0(ori_ori_n974_), .Y(ori_ori_n985_));
  NA3        o0957(.A(ori_ori_n939_), .B(ori_ori_n483_), .C(ori_ori_n46_), .Y(ori_ori_n986_));
  NA3        o0958(.A(ori_ori_n986_), .B(ori_ori_n985_), .C(ori_ori_n280_), .Y(ori_ori_n987_));
  OR4        o0959(.A(ori_ori_n987_), .B(ori_ori_n984_), .C(ori_ori_n981_), .D(ori_ori_n980_), .Y(ori_ori_n988_));
  NO4        o0960(.A(ori_ori_n988_), .B(ori_ori_n979_), .C(ori_ori_n976_), .D(ori_ori_n973_), .Y(ori_ori_n989_));
  NA4        o0961(.A(ori_ori_n989_), .B(ori_ori_n966_), .C(ori_ori_n932_), .D(ori_ori_n919_), .Y(ori13));
  NAi32      o0962(.An(d), .Bn(c), .C(e), .Y(ori_ori_n991_));
  NA2        o0963(.A(ori_ori_n142_), .B(ori_ori_n45_), .Y(ori_ori_n992_));
  NA2        o0964(.A(ori_ori_n407_), .B(ori_ori_n218_), .Y(ori_ori_n993_));
  AN2        o0965(.A(d), .B(c), .Y(ori_ori_n994_));
  NA2        o0966(.A(ori_ori_n994_), .B(ori_ori_n117_), .Y(ori_ori_n995_));
  NO2        o0967(.A(j), .B(ori_ori_n45_), .Y(ori_ori_n996_));
  NA2        o0968(.A(ori_ori_n618_), .B(ori_ori_n996_), .Y(ori_ori_n997_));
  NOi41      o0969(.An(n), .B(m), .C(i), .D(h), .Y(ori_ori_n998_));
  OR3        o0970(.A(e), .B(d), .C(c), .Y(ori_ori_n999_));
  NA3        o0971(.A(k), .B(j), .C(i), .Y(ori_ori_n1000_));
  NO3        o0972(.A(ori_ori_n1000_), .B(ori_ori_n310_), .C(ori_ori_n90_), .Y(ori_ori_n1001_));
  NOi21      o0973(.An(ori_ori_n1001_), .B(ori_ori_n999_), .Y(ori_ori_n1002_));
  NA3        o0974(.A(ori_ori_n461_), .B(ori_ori_n333_), .C(ori_ori_n56_), .Y(ori_ori_n1003_));
  NO2        o0975(.A(ori_ori_n1003_), .B(ori_ori_n997_), .Y(ori_ori_n1004_));
  NO3        o0976(.A(ori_ori_n1003_), .B(ori_ori_n576_), .C(ori_ori_n442_), .Y(ori_ori_n1005_));
  NO2        o0977(.A(f), .B(c), .Y(ori_ori_n1006_));
  NOi21      o0978(.An(ori_ori_n1006_), .B(ori_ori_n434_), .Y(ori_ori_n1007_));
  NA2        o0979(.A(ori_ori_n1007_), .B(ori_ori_n59_), .Y(ori_ori_n1008_));
  OR2        o0980(.A(k), .B(i), .Y(ori_ori_n1009_));
  NO3        o0981(.A(ori_ori_n1009_), .B(ori_ori_n249_), .C(l), .Y(ori_ori_n1010_));
  NOi31      o0982(.An(ori_ori_n1010_), .B(ori_ori_n1008_), .C(j), .Y(ori_ori_n1011_));
  OR3        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1005_), .C(ori_ori_n1004_), .Y(ori_ori_n1012_));
  OR2        o0984(.A(ori_ori_n1012_), .B(ori_ori_n1002_), .Y(ori02));
  OR2        o0985(.A(l), .B(k), .Y(ori_ori_n1014_));
  OR3        o0986(.A(h), .B(g), .C(f), .Y(ori_ori_n1015_));
  OR3        o0987(.A(n), .B(m), .C(i), .Y(ori_ori_n1016_));
  NO4        o0988(.A(ori_ori_n1016_), .B(ori_ori_n1015_), .C(ori_ori_n1014_), .D(ori_ori_n999_), .Y(ori_ori_n1017_));
  AN3        o0989(.A(g), .B(f), .C(c), .Y(ori_ori_n1018_));
  NO3        o0990(.A(ori_ori_n1003_), .B(ori_ori_n992_), .C(ori_ori_n576_), .Y(ori_ori_n1019_));
  INV        o0991(.A(ori_ori_n1019_), .Y(ori_ori_n1020_));
  NA3        o0992(.A(l), .B(k), .C(j), .Y(ori_ori_n1021_));
  NA2        o0993(.A(i), .B(h), .Y(ori_ori_n1022_));
  NO3        o0994(.A(ori_ori_n1022_), .B(ori_ori_n1021_), .C(ori_ori_n133_), .Y(ori_ori_n1023_));
  NO3        o0995(.A(ori_ori_n144_), .B(ori_ori_n288_), .C(ori_ori_n219_), .Y(ori_ori_n1024_));
  NA3        o0996(.A(c), .B(b), .C(a), .Y(ori_ori_n1025_));
  INV        o0997(.A(ori_ori_n1004_), .Y(ori_ori_n1026_));
  AN2        o0998(.A(ori_ori_n1026_), .B(ori_ori_n1020_), .Y(ori_ori_n1027_));
  NAi21      o0999(.An(ori_ori_n1017_), .B(ori_ori_n1027_), .Y(ori03));
  NO2        o1000(.A(ori_ori_n519_), .B(ori_ori_n589_), .Y(ori_ori_n1029_));
  NA4        o1001(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(g), .D(ori_ori_n218_), .Y(ori_ori_n1030_));
  NA2        o1002(.A(ori_ori_n365_), .B(ori_ori_n1030_), .Y(ori_ori_n1031_));
  NO3        o1003(.A(ori_ori_n1031_), .B(ori_ori_n1029_), .C(ori_ori_n960_), .Y(ori_ori_n1032_));
  NO3        o1004(.A(ori_ori_n824_), .B(ori_ori_n813_), .C(ori_ori_n696_), .Y(ori_ori_n1033_));
  OAI220     o1005(.A0(ori_ori_n1033_), .A1(ori_ori_n675_), .B0(ori_ori_n1032_), .B1(ori_ori_n577_), .Y(ori_ori_n1034_));
  NO2        o1006(.A(ori_ori_n791_), .B(ori_ori_n418_), .Y(ori_ori_n1035_));
  NOi31      o1007(.An(m), .B(n), .C(f), .Y(ori_ori_n1036_));
  NA2        o1008(.A(ori_ori_n1036_), .B(ori_ori_n51_), .Y(ori_ori_n1037_));
  AN2        o1009(.A(e), .B(c), .Y(ori_ori_n1038_));
  NA2        o1010(.A(ori_ori_n1038_), .B(a), .Y(ori_ori_n1039_));
  OAI220     o1011(.A0(ori_ori_n1039_), .A1(ori_ori_n1037_), .B0(ori_ori_n855_), .B1(ori_ori_n424_), .Y(ori_ori_n1040_));
  NA2        o1012(.A(ori_ori_n502_), .B(l), .Y(ori_ori_n1041_));
  NO3        o1013(.A(ori_ori_n1040_), .B(ori_ori_n1035_), .C(ori_ori_n959_), .Y(ori_ori_n1042_));
  NO2        o1014(.A(ori_ori_n288_), .B(a), .Y(ori_ori_n1043_));
  NO2        o1015(.A(ori_ori_n1022_), .B(ori_ori_n481_), .Y(ori_ori_n1044_));
  NO2        o1016(.A(ori_ori_n86_), .B(g), .Y(ori_ori_n1045_));
  AOI210     o1017(.A0(ori_ori_n1045_), .A1(ori_ori_n1044_), .B0(ori_ori_n1010_), .Y(ori_ori_n1046_));
  OR2        o1018(.A(ori_ori_n1046_), .B(ori_ori_n1008_), .Y(ori_ori_n1047_));
  NA2        o1019(.A(ori_ori_n1047_), .B(ori_ori_n1042_), .Y(ori_ori_n1048_));
  NO4        o1020(.A(ori_ori_n1048_), .B(ori_ori_n1034_), .C(ori_ori_n793_), .D(ori_ori_n558_), .Y(ori_ori_n1049_));
  NA2        o1021(.A(c), .B(b), .Y(ori_ori_n1050_));
  NO2        o1022(.A(ori_ori_n685_), .B(ori_ori_n1050_), .Y(ori_ori_n1051_));
  OAI210     o1023(.A0(ori_ori_n832_), .A1(ori_ori_n804_), .B0(ori_ori_n411_), .Y(ori_ori_n1052_));
  OAI210     o1024(.A0(ori_ori_n1052_), .A1(ori_ori_n833_), .B0(ori_ori_n1051_), .Y(ori_ori_n1053_));
  NAi21      o1025(.An(ori_ori_n419_), .B(ori_ori_n1051_), .Y(ori_ori_n1054_));
  OAI210     o1026(.A0(ori_ori_n540_), .A1(ori_ori_n39_), .B0(ori_ori_n1043_), .Y(ori_ori_n1055_));
  NA2        o1027(.A(ori_ori_n1055_), .B(ori_ori_n1054_), .Y(ori_ori_n1056_));
  NA2        o1028(.A(ori_ori_n268_), .B(ori_ori_n120_), .Y(ori_ori_n1057_));
  OAI210     o1029(.A0(ori_ori_n1057_), .A1(ori_ori_n292_), .B0(g), .Y(ori_ori_n1058_));
  NAi21      o1030(.An(f), .B(d), .Y(ori_ori_n1059_));
  NO2        o1031(.A(ori_ori_n1059_), .B(ori_ori_n1025_), .Y(ori_ori_n1060_));
  INV        o1032(.A(ori_ori_n1060_), .Y(ori_ori_n1061_));
  AOI210     o1033(.A0(ori_ori_n1058_), .A1(ori_ori_n298_), .B0(ori_ori_n1061_), .Y(ori_ori_n1062_));
  AOI210     o1034(.A0(ori_ori_n1062_), .A1(ori_ori_n114_), .B0(ori_ori_n1056_), .Y(ori_ori_n1063_));
  NA2        o1035(.A(ori_ori_n464_), .B(ori_ori_n463_), .Y(ori_ori_n1064_));
  NO2        o1036(.A(ori_ori_n186_), .B(ori_ori_n243_), .Y(ori_ori_n1065_));
  NA2        o1037(.A(ori_ori_n1065_), .B(m), .Y(ori_ori_n1066_));
  NA2        o1038(.A(ori_ori_n1041_), .B(ori_ori_n467_), .Y(ori_ori_n1067_));
  OAI210     o1039(.A0(ori_ori_n1067_), .A1(ori_ori_n315_), .B0(ori_ori_n465_), .Y(ori_ori_n1068_));
  AOI210     o1040(.A0(ori_ori_n1068_), .A1(ori_ori_n1064_), .B0(ori_ori_n1066_), .Y(ori_ori_n1069_));
  NA2        o1041(.A(ori_ori_n553_), .B(ori_ori_n406_), .Y(ori_ori_n1070_));
  NA2        o1042(.A(ori_ori_n438_), .B(ori_ori_n1060_), .Y(ori_ori_n1071_));
  NO2        o1043(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n1072_));
  NA2        o1044(.A(ori_ori_n1065_), .B(ori_ori_n427_), .Y(ori_ori_n1073_));
  NAi41      o1045(.An(ori_ori_n1072_), .B(ori_ori_n1073_), .C(ori_ori_n1071_), .D(ori_ori_n1070_), .Y(ori_ori_n1074_));
  NO2        o1046(.A(ori_ori_n1074_), .B(ori_ori_n1069_), .Y(ori_ori_n1075_));
  NA4        o1047(.A(ori_ori_n1075_), .B(ori_ori_n1063_), .C(ori_ori_n1053_), .D(ori_ori_n1049_), .Y(ori00));
  AOI210     o1048(.A0(ori_ori_n866_), .A1(ori_ori_n909_), .B0(ori_ori_n1035_), .Y(ori_ori_n1077_));
  INV        o1049(.A(ori_ori_n1019_), .Y(ori_ori_n1078_));
  NA3        o1050(.A(ori_ori_n1078_), .B(ori_ori_n1077_), .C(ori_ori_n961_), .Y(ori_ori_n1079_));
  NA2        o1051(.A(ori_ori_n504_), .B(f), .Y(ori_ori_n1080_));
  OAI210     o1052(.A0(ori_ori_n968_), .A1(ori_ori_n40_), .B0(ori_ori_n634_), .Y(ori_ori_n1081_));
  NA3        o1053(.A(ori_ori_n1081_), .B(ori_ori_n264_), .C(n), .Y(ori_ori_n1082_));
  AOI210     o1054(.A0(ori_ori_n1082_), .A1(ori_ori_n1080_), .B0(ori_ori_n995_), .Y(ori_ori_n1083_));
  NO3        o1055(.A(ori_ori_n1083_), .B(ori_ori_n1079_), .C(ori_ori_n1002_), .Y(ori_ori_n1084_));
  INV        o1056(.A(ori_ori_n1072_), .Y(ori_ori_n1085_));
  NO4        o1057(.A(ori_ori_n484_), .B(ori_ori_n352_), .C(ori_ori_n1050_), .D(ori_ori_n59_), .Y(ori_ori_n1086_));
  NA3        o1058(.A(ori_ori_n379_), .B(ori_ori_n226_), .C(g), .Y(ori_ori_n1087_));
  OR2        o1059(.A(ori_ori_n380_), .B(ori_ori_n136_), .Y(ori_ori_n1088_));
  NO2        o1060(.A(h), .B(g), .Y(ori_ori_n1089_));
  OAI220     o1061(.A0(ori_ori_n519_), .A1(ori_ori_n589_), .B0(ori_ori_n91_), .B1(ori_ori_n90_), .Y(ori_ori_n1090_));
  AOI220     o1062(.A0(ori_ori_n1090_), .A1(ori_ori_n527_), .B0(ori_ori_n914_), .B1(ori_ori_n568_), .Y(ori_ori_n1091_));
  AOI220     o1063(.A0(ori_ori_n322_), .A1(ori_ori_n253_), .B0(ori_ori_n181_), .B1(ori_ori_n151_), .Y(ori_ori_n1092_));
  NA3        o1064(.A(ori_ori_n1092_), .B(ori_ori_n1091_), .C(ori_ori_n1088_), .Y(ori_ori_n1093_));
  NO3        o1065(.A(ori_ori_n1093_), .B(ori_ori_n1086_), .C(ori_ori_n273_), .Y(ori_ori_n1094_));
  AOI210     o1066(.A0(ori_ori_n253_), .A1(ori_ori_n344_), .B0(ori_ori_n570_), .Y(ori_ori_n1095_));
  NA2        o1067(.A(ori_ori_n1095_), .B(ori_ori_n157_), .Y(ori_ori_n1096_));
  NO2        o1068(.A(ori_ori_n245_), .B(ori_ori_n185_), .Y(ori_ori_n1097_));
  NA2        o1069(.A(ori_ori_n1097_), .B(ori_ori_n425_), .Y(ori_ori_n1098_));
  NAi31      o1070(.An(ori_ori_n189_), .B(ori_ori_n829_), .C(ori_ori_n461_), .Y(ori_ori_n1099_));
  NA2        o1071(.A(ori_ori_n1099_), .B(ori_ori_n1098_), .Y(ori_ori_n1100_));
  NO4        o1072(.A(ori_ori_n1017_), .B(ori_ori_n1100_), .C(ori_ori_n1096_), .D(ori_ori_n512_), .Y(ori_ori_n1101_));
  AN3        o1073(.A(ori_ori_n1101_), .B(ori_ori_n1094_), .C(ori_ori_n1085_), .Y(ori_ori_n1102_));
  NA2        o1074(.A(ori_ori_n527_), .B(ori_ori_n101_), .Y(ori_ori_n1103_));
  NA3        o1075(.A(ori_ori_n1036_), .B(ori_ori_n597_), .C(ori_ori_n460_), .Y(ori_ori_n1104_));
  NA4        o1076(.A(ori_ori_n1104_), .B(ori_ori_n554_), .C(ori_ori_n1103_), .D(ori_ori_n247_), .Y(ori_ori_n1105_));
  NA2        o1077(.A(ori_ori_n1031_), .B(ori_ori_n527_), .Y(ori_ori_n1106_));
  NA4        o1078(.A(ori_ori_n637_), .B(ori_ori_n210_), .C(ori_ori_n226_), .D(ori_ori_n166_), .Y(ori_ori_n1107_));
  NA2        o1079(.A(ori_ori_n1107_), .B(ori_ori_n1106_), .Y(ori_ori_n1108_));
  OAI210     o1080(.A0(ori_ori_n459_), .A1(ori_ori_n121_), .B0(ori_ori_n835_), .Y(ori_ori_n1109_));
  AOI220     o1081(.A0(ori_ori_n1109_), .A1(ori_ori_n1067_), .B0(ori_ori_n553_), .B1(ori_ori_n406_), .Y(ori_ori_n1110_));
  NA2        o1082(.A(n), .B(e), .Y(ori_ori_n1111_));
  NO2        o1083(.A(ori_ori_n1111_), .B(ori_ori_n149_), .Y(ori_ori_n1112_));
  OAI210     o1084(.A0(ori_ori_n353_), .A1(ori_ori_n316_), .B0(ori_ori_n440_), .Y(ori_ori_n1113_));
  NA2        o1085(.A(ori_ori_n1113_), .B(ori_ori_n1110_), .Y(ori_ori_n1114_));
  AOI210     o1086(.A0(ori_ori_n1112_), .A1(ori_ori_n821_), .B0(ori_ori_n792_), .Y(ori_ori_n1115_));
  AOI220     o1087(.A0(ori_ori_n923_), .A1(ori_ori_n568_), .B0(ori_ori_n637_), .B1(ori_ori_n250_), .Y(ori_ori_n1116_));
  NO2        o1088(.A(ori_ori_n68_), .B(h), .Y(ori_ori_n1117_));
  NA3        o1089(.A(ori_ori_n1116_), .B(ori_ori_n1115_), .C(ori_ori_n837_), .Y(ori_ori_n1118_));
  NO4        o1090(.A(ori_ori_n1118_), .B(ori_ori_n1114_), .C(ori_ori_n1108_), .D(ori_ori_n1105_), .Y(ori_ori_n1119_));
  NA2        o1091(.A(ori_ori_n805_), .B(ori_ori_n734_), .Y(ori_ori_n1120_));
  NA4        o1092(.A(ori_ori_n1120_), .B(ori_ori_n1119_), .C(ori_ori_n1102_), .D(ori_ori_n1084_), .Y(ori01));
  NO2        o1093(.A(ori_ori_n475_), .B(ori_ori_n286_), .Y(ori_ori_n1122_));
  NA2        o1094(.A(ori_ori_n390_), .B(i), .Y(ori_ori_n1123_));
  NA3        o1095(.A(ori_ori_n1123_), .B(ori_ori_n1122_), .C(ori_ori_n982_), .Y(ori_ori_n1124_));
  NA2        o1096(.A(ori_ori_n578_), .B(ori_ori_n89_), .Y(ori_ori_n1125_));
  NA2        o1097(.A(ori_ori_n546_), .B(ori_ori_n278_), .Y(ori_ori_n1126_));
  NA2        o1098(.A(ori_ori_n928_), .B(ori_ori_n1126_), .Y(ori_ori_n1127_));
  NA4        o1099(.A(ori_ori_n1127_), .B(ori_ori_n1125_), .C(ori_ori_n881_), .D(ori_ori_n332_), .Y(ori_ori_n1128_));
  NA2        o1100(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1129_));
  NA2        o1101(.A(ori_ori_n691_), .B(ori_ori_n96_), .Y(ori_ori_n1130_));
  NO2        o1102(.A(ori_ori_n1130_), .B(ori_ori_n1129_), .Y(ori_ori_n1131_));
  OAI210     o1103(.A0(ori_ori_n756_), .A1(ori_ori_n592_), .B0(ori_ori_n1107_), .Y(ori_ori_n1132_));
  AOI210     o1104(.A0(ori_ori_n1131_), .A1(ori_ori_n623_), .B0(ori_ori_n1132_), .Y(ori_ori_n1133_));
  INV        o1105(.A(ori_ori_n119_), .Y(ori_ori_n1134_));
  OR2        o1106(.A(ori_ori_n649_), .B(ori_ori_n365_), .Y(ori_ori_n1135_));
  NAi41      o1107(.An(ori_ori_n165_), .B(ori_ori_n1135_), .C(ori_ori_n1133_), .D(ori_ori_n865_), .Y(ori_ori_n1136_));
  NO2        o1108(.A(ori_ori_n663_), .B(ori_ori_n506_), .Y(ori_ori_n1137_));
  OR2        o1109(.A(ori_ori_n199_), .B(ori_ori_n197_), .Y(ori_ori_n1138_));
  NA3        o1110(.A(ori_ori_n1138_), .B(ori_ori_n1137_), .C(ori_ori_n139_), .Y(ori_ori_n1139_));
  NO4        o1111(.A(ori_ori_n1139_), .B(ori_ori_n1136_), .C(ori_ori_n1128_), .D(ori_ori_n1124_), .Y(ori_ori_n1140_));
  INV        o1112(.A(ori_ori_n1087_), .Y(ori_ori_n1141_));
  OAI210     o1113(.A0(ori_ori_n1141_), .A1(ori_ori_n304_), .B0(ori_ori_n523_), .Y(ori_ori_n1142_));
  NA2        o1114(.A(ori_ori_n530_), .B(ori_ori_n392_), .Y(ori_ori_n1143_));
  NOi21      o1115(.An(ori_ori_n555_), .B(ori_ori_n573_), .Y(ori_ori_n1144_));
  NA2        o1116(.A(ori_ori_n1144_), .B(ori_ori_n1143_), .Y(ori_ori_n1145_));
  AOI210     o1117(.A0(ori_ori_n208_), .A1(ori_ori_n88_), .B0(ori_ori_n218_), .Y(ori_ori_n1146_));
  OAI210     o1118(.A0(ori_ori_n780_), .A1(ori_ori_n425_), .B0(ori_ori_n1146_), .Y(ori_ori_n1147_));
  AN3        o1119(.A(m), .B(l), .C(k), .Y(ori_ori_n1148_));
  OAI210     o1120(.A0(ori_ori_n355_), .A1(ori_ori_n34_), .B0(ori_ori_n1148_), .Y(ori_ori_n1149_));
  NA2        o1121(.A(ori_ori_n207_), .B(ori_ori_n34_), .Y(ori_ori_n1150_));
  AO210      o1122(.A0(ori_ori_n1150_), .A1(ori_ori_n1149_), .B0(ori_ori_n331_), .Y(ori_ori_n1151_));
  NA4        o1123(.A(ori_ori_n1151_), .B(ori_ori_n1147_), .C(ori_ori_n1145_), .D(ori_ori_n1142_), .Y(ori_ori_n1152_));
  NA2        o1124(.A(ori_ori_n587_), .B(ori_ori_n119_), .Y(ori_ori_n1153_));
  OAI210     o1125(.A0(ori_ori_n1134_), .A1(ori_ori_n584_), .B0(ori_ori_n1153_), .Y(ori_ori_n1154_));
  NA2        o1126(.A(ori_ori_n285_), .B(ori_ori_n199_), .Y(ori_ori_n1155_));
  NA2        o1127(.A(ori_ori_n1155_), .B(ori_ori_n654_), .Y(ori_ori_n1156_));
  NO3        o1128(.A(ori_ori_n791_), .B(ori_ori_n208_), .C(ori_ori_n404_), .Y(ori_ori_n1157_));
  INV        o1129(.A(ori_ori_n1157_), .Y(ori_ori_n1158_));
  NA2        o1130(.A(ori_ori_n1131_), .B(ori_ori_n664_), .Y(ori_ori_n1159_));
  NA4        o1131(.A(ori_ori_n1159_), .B(ori_ori_n1158_), .C(ori_ori_n1156_), .D(ori_ori_n759_), .Y(ori_ori_n1160_));
  NO3        o1132(.A(ori_ori_n1160_), .B(ori_ori_n1154_), .C(ori_ori_n1152_), .Y(ori_ori_n1161_));
  NA3        o1133(.A(ori_ori_n593_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1162_));
  NO2        o1134(.A(ori_ori_n1162_), .B(ori_ori_n208_), .Y(ori_ori_n1163_));
  AOI210     o1135(.A0(ori_ori_n501_), .A1(ori_ori_n58_), .B0(ori_ori_n1163_), .Y(ori_ori_n1164_));
  NO2        o1136(.A(ori_ori_n211_), .B(ori_ori_n112_), .Y(ori_ori_n1165_));
  INV        o1137(.A(ori_ori_n1165_), .Y(ori_ori_n1166_));
  NA3        o1138(.A(ori_ori_n1166_), .B(ori_ori_n1164_), .C(ori_ori_n733_), .Y(ori_ori_n1167_));
  NO2        o1139(.A(ori_ori_n934_), .B(ori_ori_n238_), .Y(ori_ori_n1168_));
  NA2        o1140(.A(ori_ori_n565_), .B(ori_ori_n563_), .Y(ori_ori_n1169_));
  NO3        o1141(.A(ori_ori_n78_), .B(ori_ori_n302_), .C(ori_ori_n45_), .Y(ori_ori_n1170_));
  NA2        o1142(.A(ori_ori_n1170_), .B(ori_ori_n545_), .Y(ori_ori_n1171_));
  NA2        o1143(.A(ori_ori_n1171_), .B(ori_ori_n1169_), .Y(ori_ori_n1172_));
  NO2        o1144(.A(ori_ori_n365_), .B(ori_ori_n71_), .Y(ori_ori_n1173_));
  INV        o1145(.A(ori_ori_n1173_), .Y(ori_ori_n1174_));
  NA2        o1146(.A(ori_ori_n1170_), .B(ori_ori_n782_), .Y(ori_ori_n1175_));
  NA3        o1147(.A(ori_ori_n1175_), .B(ori_ori_n1174_), .C(ori_ori_n382_), .Y(ori_ori_n1176_));
  NO3        o1148(.A(ori_ori_n1176_), .B(ori_ori_n1172_), .C(ori_ori_n1167_), .Y(ori_ori_n1177_));
  NO2        o1149(.A(ori_ori_n132_), .B(ori_ori_n45_), .Y(ori_ori_n1178_));
  NO2        o1150(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1179_));
  AO220      o1151(.A0(ori_ori_n1179_), .A1(ori_ori_n612_), .B0(ori_ori_n1178_), .B1(ori_ori_n689_), .Y(ori_ori_n1180_));
  NA2        o1152(.A(ori_ori_n1180_), .B(ori_ori_n339_), .Y(ori_ori_n1181_));
  INV        o1153(.A(ori_ori_n136_), .Y(ori_ori_n1182_));
  NO3        o1154(.A(ori_ori_n1022_), .B(ori_ori_n180_), .C(ori_ori_n86_), .Y(ori_ori_n1183_));
  AOI220     o1155(.A0(ori_ori_n1183_), .A1(ori_ori_n1182_), .B0(ori_ori_n1170_), .B1(ori_ori_n937_), .Y(ori_ori_n1184_));
  NA2        o1156(.A(ori_ori_n1184_), .B(ori_ori_n1181_), .Y(ori_ori_n1185_));
  NO2        o1157(.A(ori_ori_n605_), .B(ori_ori_n604_), .Y(ori_ori_n1186_));
  NO4        o1158(.A(ori_ori_n1022_), .B(ori_ori_n1186_), .C(ori_ori_n178_), .D(ori_ori_n86_), .Y(ori_ori_n1187_));
  NO3        o1159(.A(ori_ori_n1187_), .B(ori_ori_n1185_), .C(ori_ori_n626_), .Y(ori_ori_n1188_));
  NA4        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1177_), .C(ori_ori_n1161_), .D(ori_ori_n1140_), .Y(ori06));
  NO2        o1161(.A(ori_ori_n405_), .B(ori_ori_n552_), .Y(ori_ori_n1190_));
  NA2        o1162(.A(ori_ori_n274_), .B(ori_ori_n1190_), .Y(ori_ori_n1191_));
  NO2        o1163(.A(ori_ori_n230_), .B(ori_ori_n103_), .Y(ori_ori_n1192_));
  OAI210     o1164(.A0(ori_ori_n1192_), .A1(ori_ori_n1183_), .B0(ori_ori_n378_), .Y(ori_ori_n1193_));
  NO3        o1165(.A(ori_ori_n590_), .B(ori_ori_n778_), .C(ori_ori_n591_), .Y(ori_ori_n1194_));
  OR2        o1166(.A(ori_ori_n1194_), .B(ori_ori_n855_), .Y(ori_ori_n1195_));
  NA3        o1167(.A(ori_ori_n1195_), .B(ori_ori_n1193_), .C(ori_ori_n1191_), .Y(ori_ori_n1196_));
  NO3        o1168(.A(ori_ori_n1196_), .B(ori_ori_n1172_), .C(ori_ori_n263_), .Y(ori_ori_n1197_));
  NO2        o1169(.A(ori_ori_n302_), .B(ori_ori_n45_), .Y(ori_ori_n1198_));
  AOI210     o1170(.A0(ori_ori_n1198_), .A1(ori_ori_n938_), .B0(ori_ori_n1168_), .Y(ori_ori_n1199_));
  AOI210     o1171(.A0(ori_ori_n1198_), .A1(ori_ori_n549_), .B0(ori_ori_n1180_), .Y(ori_ori_n1200_));
  AOI210     o1172(.A0(ori_ori_n1200_), .A1(ori_ori_n1199_), .B0(ori_ori_n337_), .Y(ori_ori_n1201_));
  OAI210     o1173(.A0(ori_ori_n88_), .A1(ori_ori_n40_), .B0(ori_ori_n662_), .Y(ori_ori_n1202_));
  NA2        o1174(.A(ori_ori_n1202_), .B(ori_ori_n630_), .Y(ori_ori_n1203_));
  NO2        o1175(.A(ori_ori_n509_), .B(ori_ori_n175_), .Y(ori_ori_n1204_));
  NOi21      o1176(.An(ori_ori_n138_), .B(ori_ori_n45_), .Y(ori_ori_n1205_));
  NO2        o1177(.A(ori_ori_n598_), .B(ori_ori_n1037_), .Y(ori_ori_n1206_));
  OAI210     o1178(.A0(ori_ori_n454_), .A1(ori_ori_n254_), .B0(ori_ori_n876_), .Y(ori_ori_n1207_));
  NO4        o1179(.A(ori_ori_n1207_), .B(ori_ori_n1206_), .C(ori_ori_n1205_), .D(ori_ori_n1204_), .Y(ori_ori_n1208_));
  NA2        o1180(.A(ori_ori_n1208_), .B(ori_ori_n1203_), .Y(ori_ori_n1209_));
  AN2        o1181(.A(ori_ori_n923_), .B(ori_ori_n633_), .Y(ori_ori_n1210_));
  NO3        o1182(.A(ori_ori_n1210_), .B(ori_ori_n1209_), .C(ori_ori_n1201_), .Y(ori_ori_n1211_));
  NO2        o1183(.A(ori_ori_n710_), .B(ori_ori_n47_), .Y(ori_ori_n1212_));
  NA2        o1184(.A(ori_ori_n358_), .B(ori_ori_n1212_), .Y(ori_ori_n1213_));
  NO3        o1185(.A(ori_ori_n249_), .B(ori_ori_n103_), .C(ori_ori_n288_), .Y(ori_ori_n1214_));
  OAI220     o1186(.A0(ori_ori_n682_), .A1(ori_ori_n254_), .B0(ori_ori_n505_), .B1(ori_ori_n509_), .Y(ori_ori_n1215_));
  INV        o1187(.A(k), .Y(ori_ori_n1216_));
  NO3        o1188(.A(ori_ori_n1216_), .B(ori_ori_n589_), .C(j), .Y(ori_ori_n1217_));
  NOi21      o1189(.An(ori_ori_n1217_), .B(ori_ori_n658_), .Y(ori_ori_n1218_));
  NO4        o1190(.A(ori_ori_n1218_), .B(ori_ori_n1215_), .C(ori_ori_n1214_), .D(ori_ori_n1040_), .Y(ori_ori_n1219_));
  NA3        o1191(.A(ori_ori_n766_), .B(ori_ori_n765_), .C(ori_ori_n847_), .Y(ori_ori_n1220_));
  NAi31      o1192(.An(ori_ori_n724_), .B(ori_ori_n1220_), .C(ori_ori_n207_), .Y(ori_ori_n1221_));
  NA4        o1193(.A(ori_ori_n1221_), .B(ori_ori_n1219_), .C(ori_ori_n1213_), .D(ori_ori_n1116_), .Y(ori_ori_n1222_));
  AOI210     o1194(.A0(ori_ori_n565_), .A1(ori_ori_n440_), .B0(ori_ori_n369_), .Y(ori_ori_n1223_));
  NA2        o1195(.A(ori_ori_n1217_), .B(ori_ori_n762_), .Y(ori_ori_n1224_));
  NA2        o1196(.A(ori_ori_n1224_), .B(ori_ori_n1223_), .Y(ori_ori_n1225_));
  AN2        o1197(.A(ori_ori_n894_), .B(ori_ori_n893_), .Y(ori_ori_n1226_));
  NO3        o1198(.A(ori_ori_n1226_), .B(ori_ori_n497_), .C(ori_ori_n478_), .Y(ori_ori_n1227_));
  NA2        o1199(.A(ori_ori_n1227_), .B(ori_ori_n1175_), .Y(ori_ori_n1228_));
  NAi21      o1200(.An(j), .B(i), .Y(ori_ori_n1229_));
  NO4        o1201(.A(ori_ori_n1186_), .B(ori_ori_n1229_), .C(ori_ori_n434_), .D(ori_ori_n241_), .Y(ori_ori_n1230_));
  NO4        o1202(.A(ori_ori_n1230_), .B(ori_ori_n1228_), .C(ori_ori_n1225_), .D(ori_ori_n1222_), .Y(ori_ori_n1231_));
  NA4        o1203(.A(ori_ori_n1231_), .B(ori_ori_n1211_), .C(ori_ori_n1197_), .D(ori_ori_n1188_), .Y(ori07));
  NOi21      o1204(.An(j), .B(k), .Y(ori_ori_n1233_));
  NA4        o1205(.A(ori_ori_n183_), .B(ori_ori_n109_), .C(ori_ori_n1233_), .D(f), .Y(ori_ori_n1234_));
  NAi32      o1206(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1235_));
  NO3        o1207(.A(ori_ori_n1235_), .B(g), .C(f), .Y(ori_ori_n1236_));
  INV        o1208(.A(ori_ori_n1236_), .Y(ori_ori_n1237_));
  NAi21      o1209(.An(f), .B(c), .Y(ori_ori_n1238_));
  OR2        o1210(.A(e), .B(d), .Y(ori_ori_n1239_));
  NO2        o1211(.A(ori_ori_n617_), .B(ori_ori_n326_), .Y(ori_ori_n1240_));
  NA3        o1212(.A(ori_ori_n1240_), .B(ori_ori_n996_), .C(ori_ori_n183_), .Y(ori_ori_n1241_));
  NOi31      o1213(.An(n), .B(m), .C(b), .Y(ori_ori_n1242_));
  NA3        o1214(.A(ori_ori_n1241_), .B(ori_ori_n1237_), .C(ori_ori_n1234_), .Y(ori_ori_n1243_));
  NOi41      o1215(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1244_));
  NO2        o1216(.A(ori_ori_n1000_), .B(ori_ori_n310_), .Y(ori_ori_n1245_));
  NA2        o1217(.A(ori_ori_n533_), .B(ori_ori_n79_), .Y(ori_ori_n1246_));
  NA2        o1218(.A(ori_ori_n1117_), .B(ori_ori_n296_), .Y(ori_ori_n1247_));
  NA2        o1219(.A(ori_ori_n1247_), .B(ori_ori_n1246_), .Y(ori_ori_n1248_));
  NO2        o1220(.A(ori_ori_n1248_), .B(ori_ori_n1243_), .Y(ori_ori_n1249_));
  NO3        o1221(.A(e), .B(d), .C(c), .Y(ori_ori_n1250_));
  NO2        o1222(.A(ori_ori_n133_), .B(ori_ori_n219_), .Y(ori_ori_n1251_));
  NA2        o1223(.A(ori_ori_n1251_), .B(ori_ori_n1250_), .Y(ori_ori_n1252_));
  INV        o1224(.A(ori_ori_n1252_), .Y(ori_ori_n1253_));
  BUFFER     o1225(.A(h), .Y(ori_ori_n1254_));
  NO3        o1226(.A(n), .B(m), .C(i), .Y(ori_ori_n1255_));
  OAI210     o1227(.A0(ori_ori_n1038_), .A1(ori_ori_n160_), .B0(ori_ori_n1255_), .Y(ori_ori_n1256_));
  NO2        o1228(.A(ori_ori_n1256_), .B(ori_ori_n1254_), .Y(ori_ori_n1257_));
  NA3        o1229(.A(ori_ori_n679_), .B(ori_ori_n667_), .C(ori_ori_n113_), .Y(ori_ori_n1258_));
  NO2        o1230(.A(ori_ori_n1258_), .B(ori_ori_n45_), .Y(ori_ori_n1259_));
  NO2        o1231(.A(l), .B(k), .Y(ori_ori_n1260_));
  NO3        o1232(.A(ori_ori_n434_), .B(d), .C(c), .Y(ori_ori_n1261_));
  NO3        o1233(.A(ori_ori_n1259_), .B(ori_ori_n1257_), .C(ori_ori_n1253_), .Y(ori_ori_n1262_));
  NO2        o1234(.A(ori_ori_n150_), .B(h), .Y(ori_ori_n1263_));
  NO2        o1235(.A(ori_ori_n1009_), .B(l), .Y(ori_ori_n1264_));
  NO2        o1236(.A(g), .B(c), .Y(ori_ori_n1265_));
  NA3        o1237(.A(ori_ori_n1265_), .B(ori_ori_n144_), .C(ori_ori_n190_), .Y(ori_ori_n1266_));
  NO2        o1238(.A(ori_ori_n1266_), .B(ori_ori_n1264_), .Y(ori_ori_n1267_));
  NA2        o1239(.A(ori_ori_n1267_), .B(ori_ori_n183_), .Y(ori_ori_n1268_));
  NO2        o1240(.A(ori_ori_n445_), .B(a), .Y(ori_ori_n1269_));
  NA2        o1241(.A(ori_ori_n1269_), .B(ori_ori_n114_), .Y(ori_ori_n1270_));
  INV        o1242(.A(h), .Y(ori_ori_n1271_));
  NA2        o1243(.A(ori_ori_n140_), .B(ori_ori_n226_), .Y(ori_ori_n1272_));
  NO2        o1244(.A(ori_ori_n1272_), .B(ori_ori_n1380_), .Y(ori_ori_n1273_));
  NO2        o1245(.A(ori_ori_n731_), .B(ori_ori_n191_), .Y(ori_ori_n1274_));
  NOi31      o1246(.An(m), .B(n), .C(b), .Y(ori_ori_n1275_));
  NOi31      o1247(.An(f), .B(d), .C(c), .Y(ori_ori_n1276_));
  NA2        o1248(.A(ori_ori_n1276_), .B(ori_ori_n1275_), .Y(ori_ori_n1277_));
  INV        o1249(.A(ori_ori_n1277_), .Y(ori_ori_n1278_));
  NO3        o1250(.A(ori_ori_n1278_), .B(ori_ori_n1274_), .C(ori_ori_n1273_), .Y(ori_ori_n1279_));
  NA2        o1251(.A(ori_ori_n1018_), .B(ori_ori_n461_), .Y(ori_ori_n1280_));
  NO2        o1252(.A(ori_ori_n1280_), .B(ori_ori_n434_), .Y(ori_ori_n1281_));
  NO3        o1253(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1282_));
  NO2        o1254(.A(ori_ori_n998_), .B(ori_ori_n1281_), .Y(ori_ori_n1283_));
  AN4        o1255(.A(ori_ori_n1283_), .B(ori_ori_n1279_), .C(ori_ori_n1270_), .D(ori_ori_n1268_), .Y(ori_ori_n1284_));
  NA2        o1256(.A(ori_ori_n1242_), .B(ori_ori_n375_), .Y(ori_ori_n1285_));
  INV        o1257(.A(ori_ori_n1285_), .Y(ori_ori_n1286_));
  NA2        o1258(.A(ori_ori_n1261_), .B(ori_ori_n220_), .Y(ori_ori_n1287_));
  INV        o1259(.A(ori_ori_n1023_), .Y(ori_ori_n1288_));
  NAi31      o1260(.An(ori_ori_n1286_), .B(ori_ori_n1288_), .C(ori_ori_n1287_), .Y(ori_ori_n1289_));
  NO4        o1261(.A(ori_ori_n133_), .B(g), .C(f), .D(e), .Y(ori_ori_n1290_));
  NA2        o1262(.A(ori_ori_n30_), .B(h), .Y(ori_ori_n1291_));
  NO2        o1263(.A(ori_ori_n1291_), .B(ori_ori_n1016_), .Y(ori_ori_n1292_));
  NA2        o1264(.A(ori_ori_n1244_), .B(ori_ori_n1260_), .Y(ori_ori_n1293_));
  INV        o1265(.A(ori_ori_n1293_), .Y(ori_ori_n1294_));
  OR3        o1266(.A(ori_ori_n532_), .B(ori_ori_n531_), .C(ori_ori_n113_), .Y(ori_ori_n1295_));
  NA2        o1267(.A(ori_ori_n1036_), .B(ori_ori_n404_), .Y(ori_ori_n1296_));
  NO2        o1268(.A(ori_ori_n1296_), .B(ori_ori_n432_), .Y(ori_ori_n1297_));
  AO210      o1269(.A0(ori_ori_n1297_), .A1(ori_ori_n117_), .B0(ori_ori_n1294_), .Y(ori_ori_n1298_));
  NO3        o1270(.A(ori_ori_n1298_), .B(ori_ori_n1292_), .C(ori_ori_n1289_), .Y(ori_ori_n1299_));
  NA4        o1271(.A(ori_ori_n1299_), .B(ori_ori_n1284_), .C(ori_ori_n1262_), .D(ori_ori_n1249_), .Y(ori_ori_n1300_));
  NO2        o1272(.A(ori_ori_n1050_), .B(ori_ori_n111_), .Y(ori_ori_n1301_));
  NO2        o1273(.A(ori_ori_n387_), .B(j), .Y(ori_ori_n1302_));
  NA2        o1274(.A(ori_ori_n1282_), .B(ori_ori_n1036_), .Y(ori_ori_n1303_));
  NAi41      o1275(.An(ori_ori_n1271_), .B(ori_ori_n1007_), .C(ori_ori_n172_), .D(ori_ori_n153_), .Y(ori_ori_n1304_));
  NA2        o1276(.A(ori_ori_n1304_), .B(ori_ori_n1303_), .Y(ori_ori_n1305_));
  NA2        o1277(.A(ori_ori_n1302_), .B(ori_ori_n162_), .Y(ori_ori_n1306_));
  INV        o1278(.A(ori_ori_n1306_), .Y(ori_ori_n1307_));
  NO2        o1279(.A(ori_ori_n1307_), .B(ori_ori_n1305_), .Y(ori_ori_n1308_));
  INV        o1280(.A(ori_ori_n49_), .Y(ori_ori_n1309_));
  AOI220     o1281(.A0(ori_ori_n1309_), .A1(ori_ori_n1089_), .B0(ori_ori_n794_), .B1(ori_ori_n198_), .Y(ori_ori_n1310_));
  INV        o1282(.A(ori_ori_n1310_), .Y(ori_ori_n1311_));
  NO2        o1283(.A(ori_ori_n655_), .B(ori_ori_n180_), .Y(ori_ori_n1312_));
  NO2        o1284(.A(ori_ori_n1312_), .B(ori_ori_n1311_), .Y(ori_ori_n1313_));
  NO3        o1285(.A(ori_ori_n1025_), .B(ori_ori_n1239_), .C(ori_ori_n49_), .Y(ori_ori_n1314_));
  NO2        o1286(.A(ori_ori_n1016_), .B(h), .Y(ori_ori_n1315_));
  NA3        o1287(.A(ori_ori_n1315_), .B(d), .C(ori_ori_n993_), .Y(ori_ori_n1316_));
  INV        o1288(.A(ori_ori_n1316_), .Y(ori_ori_n1317_));
  NA3        o1289(.A(ori_ori_n1301_), .B(ori_ori_n461_), .C(f), .Y(ori_ori_n1318_));
  INV        o1290(.A(ori_ori_n183_), .Y(ori_ori_n1319_));
  NO2        o1291(.A(ori_ori_n1379_), .B(ori_ori_n1318_), .Y(ori_ori_n1320_));
  NO2        o1292(.A(ori_ori_n1229_), .B(ori_ori_n178_), .Y(ori_ori_n1321_));
  NOi21      o1293(.An(d), .B(f), .Y(ori_ori_n1322_));
  NO2        o1294(.A(ori_ori_n1322_), .B(ori_ori_n40_), .Y(ori_ori_n1323_));
  NA2        o1295(.A(ori_ori_n1323_), .B(ori_ori_n1321_), .Y(ori_ori_n1324_));
  INV        o1296(.A(ori_ori_n1324_), .Y(ori_ori_n1325_));
  NO3        o1297(.A(ori_ori_n1325_), .B(ori_ori_n1320_), .C(ori_ori_n1317_), .Y(ori_ori_n1326_));
  NA3        o1298(.A(ori_ori_n1326_), .B(ori_ori_n1313_), .C(ori_ori_n1308_), .Y(ori_ori_n1327_));
  NO2        o1299(.A(ori_ori_n1006_), .B(ori_ori_n40_), .Y(ori_ori_n1328_));
  INV        o1300(.A(ori_ori_n302_), .Y(ori_ori_n1329_));
  OAI210     o1301(.A0(ori_ori_n1329_), .A1(ori_ori_n1328_), .B0(ori_ori_n1245_), .Y(ori_ori_n1330_));
  OAI210     o1302(.A0(ori_ori_n1290_), .A1(ori_ori_n1242_), .B0(ori_ori_n852_), .Y(ori_ori_n1331_));
  NO2        o1303(.A(ori_ori_n991_), .B(ori_ori_n133_), .Y(ori_ori_n1332_));
  NA2        o1304(.A(ori_ori_n1332_), .B(ori_ori_n611_), .Y(ori_ori_n1333_));
  NA3        o1305(.A(ori_ori_n1333_), .B(ori_ori_n1331_), .C(ori_ori_n1330_), .Y(ori_ori_n1334_));
  NA2        o1306(.A(ori_ori_n1265_), .B(ori_ori_n1322_), .Y(ori_ori_n1335_));
  NO2        o1307(.A(ori_ori_n1335_), .B(m), .Y(ori_ori_n1336_));
  NO2        o1308(.A(ori_ori_n154_), .B(ori_ori_n185_), .Y(ori_ori_n1337_));
  OAI210     o1309(.A0(ori_ori_n1337_), .A1(ori_ori_n111_), .B0(ori_ori_n1275_), .Y(ori_ori_n1338_));
  INV        o1310(.A(ori_ori_n1338_), .Y(ori_ori_n1339_));
  NO3        o1311(.A(ori_ori_n1339_), .B(ori_ori_n1336_), .C(ori_ori_n1334_), .Y(ori_ori_n1340_));
  NO2        o1312(.A(ori_ori_n1238_), .B(e), .Y(ori_ori_n1341_));
  NA2        o1313(.A(ori_ori_n1341_), .B(ori_ori_n402_), .Y(ori_ori_n1342_));
  BUFFER     o1314(.A(ori_ori_n133_), .Y(ori_ori_n1343_));
  NO2        o1315(.A(ori_ori_n1343_), .B(ori_ori_n1342_), .Y(ori_ori_n1344_));
  NO2        o1316(.A(ori_ori_n1295_), .B(ori_ori_n349_), .Y(ori_ori_n1345_));
  NO2        o1317(.A(ori_ori_n1345_), .B(ori_ori_n1344_), .Y(ori_ori_n1346_));
  NO2        o1318(.A(ori_ori_n185_), .B(c), .Y(ori_ori_n1347_));
  NA2        o1319(.A(ori_ori_n1347_), .B(ori_ori_n183_), .Y(ori_ori_n1348_));
  AOI220     o1320(.A0(ori_ori_n1348_), .A1(ori_ori_n1008_), .B0(ori_ori_n524_), .B1(ori_ori_n363_), .Y(ori_ori_n1349_));
  NO2        o1321(.A(ori_ori_n1261_), .B(ori_ori_n1314_), .Y(ori_ori_n1350_));
  INV        o1322(.A(ori_ori_n1045_), .Y(ori_ori_n1351_));
  OAI220     o1323(.A0(ori_ori_n1351_), .A1(ori_ori_n69_), .B0(ori_ori_n1350_), .B1(ori_ori_n218_), .Y(ori_ori_n1352_));
  AOI210     o1324(.A0(ori_ori_n869_), .A1(ori_ori_n414_), .B0(ori_ori_n105_), .Y(ori_ori_n1353_));
  OR2        o1325(.A(ori_ori_n1353_), .B(ori_ori_n531_), .Y(ori_ori_n1354_));
  NO2        o1326(.A(ori_ori_n1354_), .B(ori_ori_n178_), .Y(ori_ori_n1355_));
  NA2        o1327(.A(ori_ori_n1024_), .B(ori_ori_n226_), .Y(ori_ori_n1356_));
  NO2        o1328(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1357_));
  INV        o1329(.A(ori_ori_n480_), .Y(ori_ori_n1358_));
  NA2        o1330(.A(ori_ori_n1358_), .B(ori_ori_n1357_), .Y(ori_ori_n1359_));
  NO2        o1331(.A(ori_ori_n259_), .B(g), .Y(ori_ori_n1360_));
  NO2        o1332(.A(m), .B(i), .Y(ori_ori_n1361_));
  BUFFER     o1333(.A(ori_ori_n1361_), .Y(ori_ori_n1362_));
  AOI220     o1334(.A0(ori_ori_n1362_), .A1(ori_ori_n1263_), .B0(ori_ori_n1007_), .B1(ori_ori_n1360_), .Y(ori_ori_n1363_));
  NA3        o1335(.A(ori_ori_n1363_), .B(ori_ori_n1359_), .C(ori_ori_n1356_), .Y(ori_ori_n1364_));
  NO4        o1336(.A(ori_ori_n1364_), .B(ori_ori_n1355_), .C(ori_ori_n1352_), .D(ori_ori_n1349_), .Y(ori_ori_n1365_));
  NA3        o1337(.A(ori_ori_n1365_), .B(ori_ori_n1346_), .C(ori_ori_n1340_), .Y(ori_ori_n1366_));
  NA3        o1338(.A(ori_ori_n927_), .B(ori_ori_n140_), .C(ori_ori_n46_), .Y(ori_ori_n1367_));
  INV        o1339(.A(ori_ori_n1341_), .Y(ori_ori_n1368_));
  NO2        o1340(.A(ori_ori_n1368_), .B(ori_ori_n1319_), .Y(ori_ori_n1369_));
  INV        o1341(.A(ori_ori_n1369_), .Y(ori_ori_n1370_));
  NO2        o1342(.A(ori_ori_n1296_), .B(d), .Y(ori_ori_n1371_));
  INV        o1343(.A(ori_ori_n1371_), .Y(ori_ori_n1372_));
  NA3        o1344(.A(ori_ori_n1372_), .B(ori_ori_n1370_), .C(ori_ori_n1367_), .Y(ori_ori_n1373_));
  OR4        o1345(.A(ori_ori_n1373_), .B(ori_ori_n1366_), .C(ori_ori_n1327_), .D(ori_ori_n1300_), .Y(ori04));
  INV        o1346(.A(ori_ori_n1005_), .Y(ori_ori_n1375_));
  NA3        o1347(.A(ori_ori_n1375_), .B(ori_ori_n1047_), .C(ori_ori_n1027_), .Y(ori05));
  INV        o1348(.A(ori_ori_n114_), .Y(ori_ori_n1379_));
  INV        o1349(.A(h), .Y(ori_ori_n1380_));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  INV        m0010(.A(h), .Y(mai_mai_n39_));
  NAi21      m0011(.An(j), .B(l), .Y(mai_mai_n40_));
  NAi32      m0012(.An(n), .Bn(g), .C(m), .Y(mai_mai_n41_));
  NO3        m0013(.A(mai_mai_n41_), .B(mai_mai_n40_), .C(mai_mai_n39_), .Y(mai_mai_n42_));
  NAi31      m0014(.An(n), .B(m), .C(l), .Y(mai_mai_n43_));
  INV        m0015(.A(i), .Y(mai_mai_n44_));
  AN2        m0016(.A(h), .B(g), .Y(mai_mai_n45_));
  NA2        m0017(.A(mai_mai_n45_), .B(mai_mai_n44_), .Y(mai_mai_n46_));
  NO2        m0018(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n47_));
  NAi21      m0019(.An(n), .B(m), .Y(mai_mai_n48_));
  NOi32      m0020(.An(k), .Bn(h), .C(l), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(g), .Y(mai_mai_n50_));
  INV        m0022(.A(mai_mai_n50_), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n48_), .Y(mai_mai_n52_));
  NO3        m0024(.A(mai_mai_n52_), .B(mai_mai_n47_), .C(mai_mai_n42_), .Y(mai_mai_n53_));
  NO2        m0025(.A(mai_mai_n53_), .B(mai_mai_n32_), .Y(mai_mai_n54_));
  INV        m0026(.A(c), .Y(mai_mai_n55_));
  NA2        m0027(.A(e), .B(b), .Y(mai_mai_n56_));
  NO2        m0028(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  INV        m0029(.A(d), .Y(mai_mai_n58_));
  NAi21      m0030(.An(i), .B(h), .Y(mai_mai_n59_));
  NAi31      m0031(.An(i), .B(l), .C(j), .Y(mai_mai_n60_));
  NAi41      m0032(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n61_));
  NA2        m0033(.A(g), .B(f), .Y(mai_mai_n62_));
  NO2        m0034(.A(mai_mai_n62_), .B(mai_mai_n61_), .Y(mai_mai_n63_));
  NAi21      m0035(.An(i), .B(j), .Y(mai_mai_n64_));
  NAi32      m0036(.An(n), .Bn(k), .C(m), .Y(mai_mai_n65_));
  NO2        m0037(.A(mai_mai_n65_), .B(mai_mai_n64_), .Y(mai_mai_n66_));
  NAi31      m0038(.An(l), .B(m), .C(k), .Y(mai_mai_n67_));
  NAi21      m0039(.An(e), .B(h), .Y(mai_mai_n68_));
  NAi41      m0040(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n69_));
  NA2        m0041(.A(mai_mai_n66_), .B(mai_mai_n63_), .Y(mai_mai_n70_));
  INV        m0042(.A(m), .Y(mai_mai_n71_));
  NOi21      m0043(.An(k), .B(l), .Y(mai_mai_n72_));
  NA2        m0044(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n73_));
  AN4        m0045(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n74_));
  NOi31      m0046(.An(h), .B(g), .C(f), .Y(mai_mai_n75_));
  NA2        m0047(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  NAi32      m0048(.An(m), .Bn(k), .C(j), .Y(mai_mai_n77_));
  NOi32      m0049(.An(h), .Bn(g), .C(f), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n74_), .Y(mai_mai_n79_));
  OA220      m0051(.A0(mai_mai_n79_), .A1(mai_mai_n77_), .B0(mai_mai_n76_), .B1(mai_mai_n73_), .Y(mai_mai_n80_));
  NA2        m0052(.A(mai_mai_n80_), .B(mai_mai_n70_), .Y(mai_mai_n81_));
  INV        m0053(.A(n), .Y(mai_mai_n82_));
  NOi32      m0054(.An(e), .Bn(b), .C(d), .Y(mai_mai_n83_));
  NA2        m0055(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  INV        m0056(.A(j), .Y(mai_mai_n85_));
  AN3        m0057(.A(m), .B(k), .C(i), .Y(mai_mai_n86_));
  NA3        m0058(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(g), .Y(mai_mai_n87_));
  NAi32      m0059(.An(g), .Bn(f), .C(h), .Y(mai_mai_n88_));
  NAi31      m0060(.An(j), .B(m), .C(l), .Y(mai_mai_n89_));
  NO2        m0061(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n90_));
  NA2        m0062(.A(m), .B(l), .Y(mai_mai_n91_));
  NAi31      m0063(.An(k), .B(j), .C(g), .Y(mai_mai_n92_));
  NO3        m0064(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(f), .Y(mai_mai_n93_));
  AN2        m0065(.A(j), .B(g), .Y(mai_mai_n94_));
  NOi32      m0066(.An(m), .Bn(l), .C(i), .Y(mai_mai_n95_));
  NOi21      m0067(.An(g), .B(i), .Y(mai_mai_n96_));
  NOi32      m0068(.An(m), .Bn(j), .C(k), .Y(mai_mai_n97_));
  AOI220     m0069(.A0(mai_mai_n97_), .A1(mai_mai_n96_), .B0(mai_mai_n95_), .B1(mai_mai_n94_), .Y(mai_mai_n98_));
  NO2        m0070(.A(mai_mai_n98_), .B(f), .Y(mai_mai_n99_));
  NO3        m0071(.A(mai_mai_n99_), .B(mai_mai_n93_), .C(mai_mai_n90_), .Y(mai_mai_n100_));
  NAi41      m0072(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n101_));
  AN2        m0073(.A(e), .B(b), .Y(mai_mai_n102_));
  NOi31      m0074(.An(c), .B(h), .C(f), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NO2        m0076(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n105_));
  NOi21      m0077(.An(g), .B(f), .Y(mai_mai_n106_));
  NOi21      m0078(.An(i), .B(h), .Y(mai_mai_n107_));
  NA3        m0079(.A(mai_mai_n107_), .B(mai_mai_n106_), .C(mai_mai_n36_), .Y(mai_mai_n108_));
  INV        m0080(.A(a), .Y(mai_mai_n109_));
  NA2        m0081(.A(mai_mai_n102_), .B(mai_mai_n109_), .Y(mai_mai_n110_));
  INV        m0082(.A(l), .Y(mai_mai_n111_));
  NOi21      m0083(.An(m), .B(n), .Y(mai_mai_n112_));
  AN2        m0084(.A(k), .B(h), .Y(mai_mai_n113_));
  NO2        m0085(.A(mai_mai_n108_), .B(mai_mai_n84_), .Y(mai_mai_n114_));
  INV        m0086(.A(b), .Y(mai_mai_n115_));
  NA2        m0087(.A(l), .B(j), .Y(mai_mai_n116_));
  AN2        m0088(.A(k), .B(i), .Y(mai_mai_n117_));
  NA2        m0089(.A(mai_mai_n117_), .B(mai_mai_n116_), .Y(mai_mai_n118_));
  NA2        m0090(.A(g), .B(e), .Y(mai_mai_n119_));
  NOi32      m0091(.An(c), .Bn(a), .C(d), .Y(mai_mai_n120_));
  NA2        m0092(.A(mai_mai_n120_), .B(mai_mai_n112_), .Y(mai_mai_n121_));
  NO4        m0093(.A(mai_mai_n121_), .B(mai_mai_n119_), .C(mai_mai_n118_), .D(mai_mai_n115_), .Y(mai_mai_n122_));
  NO3        m0094(.A(mai_mai_n122_), .B(mai_mai_n114_), .C(mai_mai_n105_), .Y(mai_mai_n123_));
  OAI210     m0095(.A0(mai_mai_n100_), .A1(mai_mai_n84_), .B0(mai_mai_n123_), .Y(mai_mai_n124_));
  NOi31      m0096(.An(k), .B(m), .C(j), .Y(mai_mai_n125_));
  NA3        m0097(.A(mai_mai_n125_), .B(mai_mai_n75_), .C(mai_mai_n74_), .Y(mai_mai_n126_));
  NOi31      m0098(.An(k), .B(m), .C(i), .Y(mai_mai_n127_));
  NA3        m0099(.A(mai_mai_n127_), .B(mai_mai_n78_), .C(mai_mai_n74_), .Y(mai_mai_n128_));
  NA2        m0100(.A(mai_mai_n128_), .B(mai_mai_n126_), .Y(mai_mai_n129_));
  NOi32      m0101(.An(f), .Bn(b), .C(e), .Y(mai_mai_n130_));
  NAi21      m0102(.An(g), .B(h), .Y(mai_mai_n131_));
  NAi21      m0103(.An(m), .B(n), .Y(mai_mai_n132_));
  NAi21      m0104(.An(j), .B(k), .Y(mai_mai_n133_));
  NO3        m0105(.A(mai_mai_n133_), .B(mai_mai_n132_), .C(mai_mai_n131_), .Y(mai_mai_n134_));
  NAi41      m0106(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n135_));
  NAi31      m0107(.An(j), .B(k), .C(h), .Y(mai_mai_n136_));
  NA2        m0108(.A(mai_mai_n134_), .B(mai_mai_n130_), .Y(mai_mai_n137_));
  NO2        m0109(.A(k), .B(j), .Y(mai_mai_n138_));
  NO2        m0110(.A(mai_mai_n138_), .B(mai_mai_n132_), .Y(mai_mai_n139_));
  AN2        m0111(.A(k), .B(j), .Y(mai_mai_n140_));
  NAi21      m0112(.An(c), .B(b), .Y(mai_mai_n141_));
  NA2        m0113(.A(f), .B(d), .Y(mai_mai_n142_));
  NO4        m0114(.A(mai_mai_n142_), .B(mai_mai_n141_), .C(mai_mai_n140_), .D(mai_mai_n131_), .Y(mai_mai_n143_));
  NAi31      m0115(.An(f), .B(e), .C(b), .Y(mai_mai_n144_));
  NA2        m0116(.A(mai_mai_n143_), .B(mai_mai_n139_), .Y(mai_mai_n145_));
  NA2        m0117(.A(d), .B(b), .Y(mai_mai_n146_));
  NAi21      m0118(.An(e), .B(f), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NA2        m0120(.A(b), .B(a), .Y(mai_mai_n149_));
  NAi21      m0121(.An(e), .B(g), .Y(mai_mai_n150_));
  NAi21      m0122(.An(c), .B(d), .Y(mai_mai_n151_));
  NAi31      m0123(.An(l), .B(k), .C(h), .Y(mai_mai_n152_));
  NO2        m0124(.A(mai_mai_n132_), .B(mai_mai_n152_), .Y(mai_mai_n153_));
  NAi31      m0125(.An(mai_mai_n129_), .B(mai_mai_n145_), .C(mai_mai_n137_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(b), .Y(mai_mai_n155_));
  NOi21      m0127(.An(g), .B(d), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  NOi21      m0129(.An(h), .B(i), .Y(mai_mai_n158_));
  NOi21      m0130(.An(k), .B(m), .Y(mai_mai_n159_));
  NA3        m0131(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n160_));
  NOi21      m0132(.An(h), .B(g), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n162_));
  NA2        m0134(.A(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  NAi31      m0135(.An(l), .B(j), .C(h), .Y(mai_mai_n164_));
  NO2        m0136(.A(mai_mai_n164_), .B(mai_mai_n48_), .Y(mai_mai_n165_));
  NA2        m0137(.A(mai_mai_n165_), .B(mai_mai_n63_), .Y(mai_mai_n166_));
  NOi32      m0138(.An(n), .Bn(k), .C(m), .Y(mai_mai_n167_));
  NA2        m0139(.A(l), .B(i), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  OAI210     m0141(.A0(mai_mai_n169_), .A1(mai_mai_n163_), .B0(mai_mai_n166_), .Y(mai_mai_n170_));
  NAi31      m0142(.An(d), .B(f), .C(c), .Y(mai_mai_n171_));
  NAi31      m0143(.An(e), .B(f), .C(c), .Y(mai_mai_n172_));
  NA2        m0144(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  NA2        m0145(.A(j), .B(h), .Y(mai_mai_n174_));
  OR3        m0146(.A(n), .B(m), .C(k), .Y(mai_mai_n175_));
  NO2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NAi32      m0148(.An(m), .Bn(k), .C(n), .Y(mai_mai_n177_));
  NO2        m0149(.A(mai_mai_n177_), .B(mai_mai_n174_), .Y(mai_mai_n178_));
  AOI220     m0150(.A0(mai_mai_n178_), .A1(mai_mai_n157_), .B0(mai_mai_n176_), .B1(mai_mai_n173_), .Y(mai_mai_n179_));
  NO2        m0151(.A(n), .B(m), .Y(mai_mai_n180_));
  NA2        m0152(.A(mai_mai_n180_), .B(mai_mai_n49_), .Y(mai_mai_n181_));
  NAi21      m0153(.An(f), .B(e), .Y(mai_mai_n182_));
  NA2        m0154(.A(d), .B(c), .Y(mai_mai_n183_));
  NO2        m0155(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  NOi21      m0156(.An(mai_mai_n184_), .B(mai_mai_n181_), .Y(mai_mai_n185_));
  NAi21      m0157(.An(d), .B(c), .Y(mai_mai_n186_));
  NAi31      m0158(.An(m), .B(n), .C(b), .Y(mai_mai_n187_));
  NA2        m0159(.A(k), .B(i), .Y(mai_mai_n188_));
  NAi21      m0160(.An(h), .B(f), .Y(mai_mai_n189_));
  NO2        m0161(.A(mai_mai_n189_), .B(mai_mai_n188_), .Y(mai_mai_n190_));
  NO2        m0162(.A(mai_mai_n187_), .B(mai_mai_n151_), .Y(mai_mai_n191_));
  NA2        m0163(.A(mai_mai_n191_), .B(mai_mai_n190_), .Y(mai_mai_n192_));
  NOi32      m0164(.An(f), .Bn(c), .C(d), .Y(mai_mai_n193_));
  NOi32      m0165(.An(f), .Bn(c), .C(e), .Y(mai_mai_n194_));
  NO2        m0166(.A(mai_mai_n194_), .B(mai_mai_n193_), .Y(mai_mai_n195_));
  NO3        m0167(.A(n), .B(m), .C(j), .Y(mai_mai_n196_));
  NA2        m0168(.A(mai_mai_n196_), .B(mai_mai_n113_), .Y(mai_mai_n197_));
  AO210      m0169(.A0(mai_mai_n197_), .A1(mai_mai_n181_), .B0(mai_mai_n195_), .Y(mai_mai_n198_));
  NAi41      m0170(.An(mai_mai_n185_), .B(mai_mai_n198_), .C(mai_mai_n192_), .D(mai_mai_n179_), .Y(mai_mai_n199_));
  OR3        m0171(.A(mai_mai_n199_), .B(mai_mai_n170_), .C(mai_mai_n154_), .Y(mai_mai_n200_));
  NO4        m0172(.A(mai_mai_n200_), .B(mai_mai_n124_), .C(mai_mai_n81_), .D(mai_mai_n54_), .Y(mai_mai_n201_));
  NA3        m0173(.A(m), .B(mai_mai_n111_), .C(j), .Y(mai_mai_n202_));
  NAi31      m0174(.An(n), .B(h), .C(g), .Y(mai_mai_n203_));
  NO2        m0175(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  NOi32      m0176(.An(m), .Bn(k), .C(l), .Y(mai_mai_n205_));
  NA3        m0177(.A(mai_mai_n205_), .B(mai_mai_n85_), .C(g), .Y(mai_mai_n206_));
  NO2        m0178(.A(mai_mai_n206_), .B(n), .Y(mai_mai_n207_));
  NOi21      m0179(.An(k), .B(j), .Y(mai_mai_n208_));
  NA4        m0180(.A(mai_mai_n208_), .B(mai_mai_n112_), .C(i), .D(g), .Y(mai_mai_n209_));
  AN2        m0181(.A(i), .B(g), .Y(mai_mai_n210_));
  INV        m0182(.A(mai_mai_n209_), .Y(mai_mai_n211_));
  NAi41      m0183(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n212_));
  INV        m0184(.A(mai_mai_n212_), .Y(mai_mai_n213_));
  INV        m0185(.A(f), .Y(mai_mai_n214_));
  INV        m0186(.A(g), .Y(mai_mai_n215_));
  NOi31      m0187(.An(i), .B(j), .C(h), .Y(mai_mai_n216_));
  NOi21      m0188(.An(l), .B(m), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  NO3        m0190(.A(mai_mai_n218_), .B(mai_mai_n215_), .C(mai_mai_n214_), .Y(mai_mai_n219_));
  NA2        m0191(.A(mai_mai_n219_), .B(mai_mai_n213_), .Y(mai_mai_n220_));
  OAI210     m0192(.A0(mai_mai_n209_), .A1(mai_mai_n32_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  NOi21      m0193(.An(n), .B(m), .Y(mai_mai_n222_));
  NOi32      m0194(.An(l), .Bn(i), .C(j), .Y(mai_mai_n223_));
  NA2        m0195(.A(mai_mai_n223_), .B(mai_mai_n222_), .Y(mai_mai_n224_));
  OA220      m0196(.A0(mai_mai_n224_), .A1(mai_mai_n104_), .B0(mai_mai_n77_), .B1(mai_mai_n76_), .Y(mai_mai_n225_));
  NAi21      m0197(.An(j), .B(h), .Y(mai_mai_n226_));
  XN2        m0198(.A(i), .B(h), .Y(mai_mai_n227_));
  NA2        m0199(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  NOi31      m0200(.An(k), .B(n), .C(m), .Y(mai_mai_n229_));
  NOi31      m0201(.An(mai_mai_n229_), .B(mai_mai_n183_), .C(mai_mai_n182_), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n230_), .B(mai_mai_n228_), .Y(mai_mai_n231_));
  NAi31      m0203(.An(f), .B(e), .C(c), .Y(mai_mai_n232_));
  NO4        m0204(.A(mai_mai_n232_), .B(mai_mai_n175_), .C(mai_mai_n174_), .D(mai_mai_n58_), .Y(mai_mai_n233_));
  NA3        m0205(.A(e), .B(c), .C(b), .Y(mai_mai_n234_));
  NAi32      m0206(.An(m), .Bn(i), .C(k), .Y(mai_mai_n235_));
  INV        m0207(.A(k), .Y(mai_mai_n236_));
  INV        m0208(.A(mai_mai_n233_), .Y(mai_mai_n237_));
  NAi21      m0209(.An(n), .B(a), .Y(mai_mai_n238_));
  NO2        m0210(.A(mai_mai_n238_), .B(mai_mai_n146_), .Y(mai_mai_n239_));
  NAi41      m0211(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n240_), .B(e), .Y(mai_mai_n241_));
  NO3        m0213(.A(mai_mai_n147_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n242_));
  OAI210     m0214(.A0(mai_mai_n242_), .A1(mai_mai_n241_), .B0(mai_mai_n239_), .Y(mai_mai_n243_));
  AN4        m0215(.A(mai_mai_n243_), .B(mai_mai_n237_), .C(mai_mai_n231_), .D(mai_mai_n225_), .Y(mai_mai_n244_));
  OR2        m0216(.A(h), .B(g), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n245_), .B(mai_mai_n101_), .Y(mai_mai_n246_));
  NA2        m0218(.A(mai_mai_n246_), .B(mai_mai_n130_), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n159_), .B(mai_mai_n107_), .Y(mai_mai_n248_));
  NO2        m0220(.A(n), .B(a), .Y(mai_mai_n249_));
  NAi31      m0221(.An(mai_mai_n240_), .B(mai_mai_n249_), .C(mai_mai_n102_), .Y(mai_mai_n250_));
  NAi21      m0222(.An(h), .B(i), .Y(mai_mai_n251_));
  NA2        m0223(.A(mai_mai_n180_), .B(k), .Y(mai_mai_n252_));
  NO2        m0224(.A(mai_mai_n252_), .B(mai_mai_n251_), .Y(mai_mai_n253_));
  NA2        m0225(.A(mai_mai_n253_), .B(mai_mai_n193_), .Y(mai_mai_n254_));
  NA3        m0226(.A(mai_mai_n254_), .B(mai_mai_n250_), .C(mai_mai_n247_), .Y(mai_mai_n255_));
  NOi21      m0227(.An(g), .B(e), .Y(mai_mai_n256_));
  NO2        m0228(.A(mai_mai_n69_), .B(mai_mai_n71_), .Y(mai_mai_n257_));
  NOi32      m0229(.An(l), .Bn(j), .C(i), .Y(mai_mai_n258_));
  AOI210     m0230(.A0(mai_mai_n72_), .A1(mai_mai_n85_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n251_), .B(mai_mai_n43_), .Y(mai_mai_n260_));
  NAi21      m0232(.An(f), .B(g), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n261_), .B(mai_mai_n61_), .Y(mai_mai_n262_));
  NO2        m0234(.A(mai_mai_n65_), .B(mai_mai_n116_), .Y(mai_mai_n263_));
  AOI220     m0235(.A0(mai_mai_n263_), .A1(mai_mai_n262_), .B0(mai_mai_n260_), .B1(mai_mai_n63_), .Y(mai_mai_n264_));
  INV        m0236(.A(mai_mai_n264_), .Y(mai_mai_n265_));
  NO3        m0237(.A(mai_mai_n133_), .B(mai_mai_n48_), .C(mai_mai_n44_), .Y(mai_mai_n266_));
  NOi41      m0238(.An(mai_mai_n244_), .B(mai_mai_n265_), .C(mai_mai_n255_), .D(mai_mai_n221_), .Y(mai_mai_n267_));
  NO3        m0239(.A(mai_mai_n204_), .B(mai_mai_n47_), .C(mai_mai_n42_), .Y(mai_mai_n268_));
  NO2        m0240(.A(mai_mai_n268_), .B(mai_mai_n110_), .Y(mai_mai_n269_));
  NA3        m0241(.A(mai_mai_n58_), .B(c), .C(b), .Y(mai_mai_n270_));
  NAi21      m0242(.An(h), .B(g), .Y(mai_mai_n271_));
  NO2        m0243(.A(mai_mai_n248_), .B(mai_mai_n261_), .Y(mai_mai_n272_));
  NAi31      m0244(.An(g), .B(k), .C(h), .Y(mai_mai_n273_));
  NO3        m0245(.A(mai_mai_n132_), .B(mai_mai_n273_), .C(l), .Y(mai_mai_n274_));
  NAi31      m0246(.An(e), .B(d), .C(a), .Y(mai_mai_n275_));
  NA2        m0247(.A(mai_mai_n274_), .B(mai_mai_n130_), .Y(mai_mai_n276_));
  INV        m0248(.A(mai_mai_n276_), .Y(mai_mai_n277_));
  NA3        m0249(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(mai_mai_n82_), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n278_), .B(mai_mai_n195_), .Y(mai_mai_n279_));
  INV        m0251(.A(mai_mai_n279_), .Y(mai_mai_n280_));
  NA3        m0252(.A(e), .B(c), .C(b), .Y(mai_mai_n281_));
  NAi32      m0253(.An(k), .Bn(i), .C(j), .Y(mai_mai_n282_));
  NAi21      m0254(.An(l), .B(k), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n283_), .B(mai_mai_n48_), .Y(mai_mai_n284_));
  NOi21      m0256(.An(l), .B(j), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n161_), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  NA3        m0258(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(g), .Y(mai_mai_n287_));
  OR3        m0259(.A(mai_mai_n69_), .B(mai_mai_n71_), .C(e), .Y(mai_mai_n288_));
  AOI210     m0260(.A0(mai_mai_n287_), .A1(mai_mai_n286_), .B0(mai_mai_n288_), .Y(mai_mai_n289_));
  INV        m0261(.A(mai_mai_n289_), .Y(mai_mai_n290_));
  NAi32      m0262(.An(j), .Bn(h), .C(i), .Y(mai_mai_n291_));
  NAi21      m0263(.An(m), .B(l), .Y(mai_mai_n292_));
  NO3        m0264(.A(mai_mai_n292_), .B(mai_mai_n291_), .C(mai_mai_n82_), .Y(mai_mai_n293_));
  NA2        m0265(.A(h), .B(g), .Y(mai_mai_n294_));
  NA2        m0266(.A(mai_mai_n167_), .B(mai_mai_n44_), .Y(mai_mai_n295_));
  NO2        m0267(.A(mai_mai_n295_), .B(mai_mai_n294_), .Y(mai_mai_n296_));
  OAI210     m0268(.A0(mai_mai_n296_), .A1(mai_mai_n293_), .B0(mai_mai_n162_), .Y(mai_mai_n297_));
  NA3        m0269(.A(mai_mai_n297_), .B(mai_mai_n290_), .C(mai_mai_n280_), .Y(mai_mai_n298_));
  NO2        m0270(.A(mai_mai_n144_), .B(d), .Y(mai_mai_n299_));
  NA2        m0271(.A(mai_mai_n299_), .B(mai_mai_n52_), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n301_));
  NAi32      m0273(.An(n), .Bn(m), .C(l), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n302_), .B(mai_mai_n291_), .Y(mai_mai_n303_));
  NA2        m0275(.A(mai_mai_n303_), .B(mai_mai_n184_), .Y(mai_mai_n304_));
  NAi31      m0276(.An(k), .B(l), .C(j), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n304_), .B(mai_mai_n300_), .Y(mai_mai_n306_));
  NO4        m0278(.A(mai_mai_n306_), .B(mai_mai_n298_), .C(mai_mai_n277_), .D(mai_mai_n269_), .Y(mai_mai_n307_));
  NA2        m0279(.A(mai_mai_n253_), .B(mai_mai_n194_), .Y(mai_mai_n308_));
  NAi21      m0280(.An(m), .B(k), .Y(mai_mai_n309_));
  NO2        m0281(.A(mai_mai_n227_), .B(mai_mai_n309_), .Y(mai_mai_n310_));
  NAi41      m0282(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n311_));
  NO2        m0283(.A(mai_mai_n311_), .B(mai_mai_n150_), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n312_), .B(mai_mai_n310_), .Y(mai_mai_n313_));
  NAi31      m0285(.An(i), .B(l), .C(h), .Y(mai_mai_n314_));
  NO4        m0286(.A(mai_mai_n314_), .B(mai_mai_n150_), .C(mai_mai_n69_), .D(mai_mai_n71_), .Y(mai_mai_n315_));
  NA2        m0287(.A(e), .B(c), .Y(mai_mai_n316_));
  NO3        m0288(.A(mai_mai_n316_), .B(n), .C(d), .Y(mai_mai_n317_));
  NOi21      m0289(.An(f), .B(h), .Y(mai_mai_n318_));
  NA2        m0290(.A(mai_mai_n318_), .B(mai_mai_n117_), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n319_), .B(mai_mai_n215_), .Y(mai_mai_n320_));
  NAi31      m0292(.An(d), .B(e), .C(b), .Y(mai_mai_n321_));
  NO2        m0293(.A(mai_mai_n132_), .B(mai_mai_n321_), .Y(mai_mai_n322_));
  NA2        m0294(.A(mai_mai_n322_), .B(mai_mai_n320_), .Y(mai_mai_n323_));
  NAi41      m0295(.An(mai_mai_n315_), .B(mai_mai_n323_), .C(mai_mai_n313_), .D(mai_mai_n308_), .Y(mai_mai_n324_));
  NO4        m0296(.A(mai_mai_n311_), .B(mai_mai_n77_), .C(mai_mai_n68_), .D(mai_mai_n215_), .Y(mai_mai_n325_));
  NA2        m0297(.A(mai_mai_n249_), .B(mai_mai_n102_), .Y(mai_mai_n326_));
  OR2        m0298(.A(mai_mai_n326_), .B(mai_mai_n206_), .Y(mai_mai_n327_));
  NOi31      m0299(.An(l), .B(n), .C(m), .Y(mai_mai_n328_));
  NA2        m0300(.A(mai_mai_n328_), .B(mai_mai_n216_), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n329_), .B(mai_mai_n195_), .Y(mai_mai_n330_));
  NAi32      m0302(.An(mai_mai_n330_), .Bn(mai_mai_n325_), .C(mai_mai_n327_), .Y(mai_mai_n331_));
  NAi32      m0303(.An(m), .Bn(j), .C(k), .Y(mai_mai_n332_));
  NAi41      m0304(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n333_));
  OAI210     m0305(.A0(mai_mai_n212_), .A1(mai_mai_n332_), .B0(mai_mai_n333_), .Y(mai_mai_n334_));
  NOi31      m0306(.An(j), .B(m), .C(k), .Y(mai_mai_n335_));
  NO2        m0307(.A(mai_mai_n125_), .B(mai_mai_n335_), .Y(mai_mai_n336_));
  AN3        m0308(.A(h), .B(g), .C(f), .Y(mai_mai_n337_));
  NAi31      m0309(.An(mai_mai_n336_), .B(mai_mai_n337_), .C(mai_mai_n334_), .Y(mai_mai_n338_));
  NOi32      m0310(.An(m), .Bn(j), .C(l), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n339_), .B(mai_mai_n95_), .Y(mai_mai_n340_));
  NAi32      m0312(.An(mai_mai_n340_), .Bn(mai_mai_n203_), .C(mai_mai_n299_), .Y(mai_mai_n341_));
  NO2        m0313(.A(mai_mai_n292_), .B(mai_mai_n291_), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n218_), .B(g), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n155_), .B(mai_mai_n82_), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n344_), .B(mai_mai_n343_), .Y(mai_mai_n345_));
  NA2        m0317(.A(mai_mai_n235_), .B(mai_mai_n77_), .Y(mai_mai_n346_));
  NA3        m0318(.A(mai_mai_n346_), .B(mai_mai_n337_), .C(mai_mai_n213_), .Y(mai_mai_n347_));
  NA4        m0319(.A(mai_mai_n347_), .B(mai_mai_n345_), .C(mai_mai_n341_), .D(mai_mai_n338_), .Y(mai_mai_n348_));
  NA3        m0320(.A(h), .B(g), .C(f), .Y(mai_mai_n349_));
  NOi32      m0321(.An(j), .Bn(g), .C(i), .Y(mai_mai_n350_));
  NA3        m0322(.A(mai_mai_n350_), .B(mai_mai_n283_), .C(mai_mai_n112_), .Y(mai_mai_n351_));
  AO210      m0323(.A0(mai_mai_n110_), .A1(mai_mai_n32_), .B0(mai_mai_n351_), .Y(mai_mai_n352_));
  NOi32      m0324(.An(e), .Bn(b), .C(a), .Y(mai_mai_n353_));
  AN2        m0325(.A(l), .B(j), .Y(mai_mai_n354_));
  NO2        m0326(.A(mai_mai_n309_), .B(mai_mai_n354_), .Y(mai_mai_n355_));
  NO3        m0327(.A(mai_mai_n311_), .B(mai_mai_n68_), .C(mai_mai_n215_), .Y(mai_mai_n356_));
  NA2        m0328(.A(mai_mai_n209_), .B(mai_mai_n35_), .Y(mai_mai_n357_));
  AOI220     m0329(.A0(mai_mai_n357_), .A1(mai_mai_n353_), .B0(mai_mai_n356_), .B1(mai_mai_n355_), .Y(mai_mai_n358_));
  NA2        m0330(.A(mai_mai_n210_), .B(k), .Y(mai_mai_n359_));
  NA3        m0331(.A(m), .B(mai_mai_n111_), .C(mai_mai_n214_), .Y(mai_mai_n360_));
  NAi41      m0332(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n361_));
  NA2        m0333(.A(mai_mai_n50_), .B(mai_mai_n112_), .Y(mai_mai_n362_));
  NA2        m0334(.A(mai_mai_n358_), .B(mai_mai_n352_), .Y(mai_mai_n363_));
  NO4        m0335(.A(mai_mai_n363_), .B(mai_mai_n348_), .C(mai_mai_n331_), .D(mai_mai_n324_), .Y(mai_mai_n364_));
  NA4        m0336(.A(mai_mai_n364_), .B(mai_mai_n307_), .C(mai_mai_n267_), .D(mai_mai_n201_), .Y(mai10));
  NA3        m0337(.A(m), .B(k), .C(i), .Y(mai_mai_n366_));
  NO3        m0338(.A(mai_mai_n366_), .B(j), .C(mai_mai_n215_), .Y(mai_mai_n367_));
  NOi21      m0339(.An(e), .B(f), .Y(mai_mai_n368_));
  NO4        m0340(.A(mai_mai_n151_), .B(mai_mai_n368_), .C(n), .D(mai_mai_n109_), .Y(mai_mai_n369_));
  NAi31      m0341(.An(b), .B(f), .C(c), .Y(mai_mai_n370_));
  INV        m0342(.A(mai_mai_n370_), .Y(mai_mai_n371_));
  NOi32      m0343(.An(k), .Bn(h), .C(j), .Y(mai_mai_n372_));
  NA2        m0344(.A(mai_mai_n372_), .B(mai_mai_n222_), .Y(mai_mai_n373_));
  NA2        m0345(.A(mai_mai_n160_), .B(mai_mai_n373_), .Y(mai_mai_n374_));
  AOI220     m0346(.A0(mai_mai_n374_), .A1(mai_mai_n371_), .B0(mai_mai_n369_), .B1(mai_mai_n367_), .Y(mai_mai_n375_));
  AN2        m0347(.A(j), .B(h), .Y(mai_mai_n376_));
  NO3        m0348(.A(n), .B(m), .C(k), .Y(mai_mai_n377_));
  NA2        m0349(.A(mai_mai_n377_), .B(mai_mai_n376_), .Y(mai_mai_n378_));
  NO3        m0350(.A(mai_mai_n378_), .B(mai_mai_n151_), .C(mai_mai_n214_), .Y(mai_mai_n379_));
  OR2        m0351(.A(m), .B(k), .Y(mai_mai_n380_));
  NO2        m0352(.A(mai_mai_n174_), .B(mai_mai_n380_), .Y(mai_mai_n381_));
  NA4        m0353(.A(n), .B(f), .C(c), .D(mai_mai_n115_), .Y(mai_mai_n382_));
  NOi21      m0354(.An(mai_mai_n381_), .B(mai_mai_n382_), .Y(mai_mai_n383_));
  NOi32      m0355(.An(d), .Bn(a), .C(c), .Y(mai_mai_n384_));
  NA2        m0356(.A(mai_mai_n384_), .B(mai_mai_n182_), .Y(mai_mai_n385_));
  NAi21      m0357(.An(i), .B(g), .Y(mai_mai_n386_));
  NAi31      m0358(.An(k), .B(m), .C(j), .Y(mai_mai_n387_));
  NO3        m0359(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(n), .Y(mai_mai_n388_));
  NOi21      m0360(.An(mai_mai_n388_), .B(mai_mai_n385_), .Y(mai_mai_n389_));
  NO3        m0361(.A(mai_mai_n389_), .B(mai_mai_n383_), .C(mai_mai_n379_), .Y(mai_mai_n390_));
  NO2        m0362(.A(mai_mai_n382_), .B(mai_mai_n292_), .Y(mai_mai_n391_));
  NOi32      m0363(.An(f), .Bn(d), .C(c), .Y(mai_mai_n392_));
  AOI220     m0364(.A0(mai_mai_n392_), .A1(mai_mai_n303_), .B0(mai_mai_n391_), .B1(mai_mai_n216_), .Y(mai_mai_n393_));
  NA3        m0365(.A(mai_mai_n393_), .B(mai_mai_n390_), .C(mai_mai_n375_), .Y(mai_mai_n394_));
  NO2        m0366(.A(mai_mai_n58_), .B(mai_mai_n115_), .Y(mai_mai_n395_));
  NA2        m0367(.A(mai_mai_n249_), .B(mai_mai_n395_), .Y(mai_mai_n396_));
  INV        m0368(.A(e), .Y(mai_mai_n397_));
  NA2        m0369(.A(mai_mai_n45_), .B(e), .Y(mai_mai_n398_));
  OAI220     m0370(.A0(mai_mai_n398_), .A1(mai_mai_n202_), .B0(mai_mai_n206_), .B1(mai_mai_n397_), .Y(mai_mai_n399_));
  AN2        m0371(.A(g), .B(e), .Y(mai_mai_n400_));
  NO2        m0372(.A(mai_mai_n87_), .B(mai_mai_n397_), .Y(mai_mai_n401_));
  NO2        m0373(.A(mai_mai_n98_), .B(mai_mai_n397_), .Y(mai_mai_n402_));
  NO3        m0374(.A(mai_mai_n402_), .B(mai_mai_n401_), .C(mai_mai_n399_), .Y(mai_mai_n403_));
  NOi21      m0375(.An(g), .B(h), .Y(mai_mai_n404_));
  AN3        m0376(.A(m), .B(l), .C(i), .Y(mai_mai_n405_));
  NA3        m0377(.A(mai_mai_n405_), .B(mai_mai_n404_), .C(e), .Y(mai_mai_n406_));
  AN3        m0378(.A(h), .B(g), .C(e), .Y(mai_mai_n407_));
  NA2        m0379(.A(mai_mai_n407_), .B(mai_mai_n95_), .Y(mai_mai_n408_));
  AN2        m0380(.A(mai_mai_n408_), .B(mai_mai_n406_), .Y(mai_mai_n409_));
  AOI210     m0381(.A0(mai_mai_n409_), .A1(mai_mai_n403_), .B0(mai_mai_n396_), .Y(mai_mai_n410_));
  NA3        m0382(.A(mai_mai_n384_), .B(mai_mai_n182_), .C(mai_mai_n82_), .Y(mai_mai_n411_));
  NAi31      m0383(.An(b), .B(c), .C(a), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n412_), .B(n), .Y(mai_mai_n413_));
  NA2        m0385(.A(mai_mai_n50_), .B(m), .Y(mai_mai_n414_));
  NO2        m0386(.A(mai_mai_n414_), .B(mai_mai_n147_), .Y(mai_mai_n415_));
  NA2        m0387(.A(mai_mai_n415_), .B(mai_mai_n413_), .Y(mai_mai_n416_));
  INV        m0388(.A(mai_mai_n416_), .Y(mai_mai_n417_));
  NO3        m0389(.A(mai_mai_n417_), .B(mai_mai_n410_), .C(mai_mai_n394_), .Y(mai_mai_n418_));
  NA2        m0390(.A(i), .B(g), .Y(mai_mai_n419_));
  NO3        m0391(.A(mai_mai_n275_), .B(mai_mai_n419_), .C(c), .Y(mai_mai_n420_));
  NOi21      m0392(.An(a), .B(n), .Y(mai_mai_n421_));
  NOi21      m0393(.An(d), .B(c), .Y(mai_mai_n422_));
  NA2        m0394(.A(mai_mai_n422_), .B(mai_mai_n421_), .Y(mai_mai_n423_));
  NA3        m0395(.A(i), .B(g), .C(f), .Y(mai_mai_n424_));
  OR2        m0396(.A(mai_mai_n424_), .B(mai_mai_n67_), .Y(mai_mai_n425_));
  NA3        m0397(.A(mai_mai_n405_), .B(mai_mai_n404_), .C(mai_mai_n182_), .Y(mai_mai_n426_));
  AOI210     m0398(.A0(mai_mai_n426_), .A1(mai_mai_n425_), .B0(mai_mai_n423_), .Y(mai_mai_n427_));
  AOI210     m0399(.A0(mai_mai_n420_), .A1(mai_mai_n284_), .B0(mai_mai_n427_), .Y(mai_mai_n428_));
  OR2        m0400(.A(n), .B(m), .Y(mai_mai_n429_));
  NO2        m0401(.A(mai_mai_n429_), .B(mai_mai_n152_), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n183_), .B(mai_mai_n147_), .Y(mai_mai_n431_));
  OAI210     m0403(.A0(mai_mai_n430_), .A1(mai_mai_n176_), .B0(mai_mai_n431_), .Y(mai_mai_n432_));
  INV        m0404(.A(mai_mai_n362_), .Y(mai_mai_n433_));
  NA3        m0405(.A(mai_mai_n433_), .B(mai_mai_n353_), .C(d), .Y(mai_mai_n434_));
  NO2        m0406(.A(mai_mai_n412_), .B(mai_mai_n48_), .Y(mai_mai_n435_));
  NO3        m0407(.A(mai_mai_n62_), .B(mai_mai_n111_), .C(e), .Y(mai_mai_n436_));
  NAi21      m0408(.An(k), .B(j), .Y(mai_mai_n437_));
  NA2        m0409(.A(mai_mai_n251_), .B(mai_mai_n437_), .Y(mai_mai_n438_));
  NA3        m0410(.A(mai_mai_n438_), .B(mai_mai_n436_), .C(mai_mai_n435_), .Y(mai_mai_n439_));
  NAi21      m0411(.An(e), .B(d), .Y(mai_mai_n440_));
  INV        m0412(.A(mai_mai_n440_), .Y(mai_mai_n441_));
  NO2        m0413(.A(mai_mai_n252_), .B(mai_mai_n214_), .Y(mai_mai_n442_));
  NA3        m0414(.A(mai_mai_n442_), .B(mai_mai_n441_), .C(mai_mai_n228_), .Y(mai_mai_n443_));
  NA4        m0415(.A(mai_mai_n443_), .B(mai_mai_n439_), .C(mai_mai_n434_), .D(mai_mai_n432_), .Y(mai_mai_n444_));
  NO2        m0416(.A(mai_mai_n329_), .B(mai_mai_n214_), .Y(mai_mai_n445_));
  NA2        m0417(.A(mai_mai_n445_), .B(mai_mai_n441_), .Y(mai_mai_n446_));
  NOi31      m0418(.An(n), .B(m), .C(k), .Y(mai_mai_n447_));
  AOI220     m0419(.A0(mai_mai_n447_), .A1(mai_mai_n376_), .B0(mai_mai_n222_), .B1(mai_mai_n49_), .Y(mai_mai_n448_));
  NAi31      m0420(.An(g), .B(f), .C(c), .Y(mai_mai_n449_));
  OR3        m0421(.A(mai_mai_n449_), .B(mai_mai_n448_), .C(e), .Y(mai_mai_n450_));
  NA3        m0422(.A(mai_mai_n450_), .B(mai_mai_n446_), .C(mai_mai_n304_), .Y(mai_mai_n451_));
  NOi41      m0423(.An(mai_mai_n428_), .B(mai_mai_n451_), .C(mai_mai_n444_), .D(mai_mai_n265_), .Y(mai_mai_n452_));
  NOi32      m0424(.An(c), .Bn(a), .C(b), .Y(mai_mai_n453_));
  NA2        m0425(.A(mai_mai_n453_), .B(mai_mai_n112_), .Y(mai_mai_n454_));
  INV        m0426(.A(mai_mai_n273_), .Y(mai_mai_n455_));
  AN2        m0427(.A(e), .B(d), .Y(mai_mai_n456_));
  NA2        m0428(.A(mai_mai_n456_), .B(mai_mai_n455_), .Y(mai_mai_n457_));
  INV        m0429(.A(mai_mai_n147_), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n131_), .B(mai_mai_n40_), .Y(mai_mai_n459_));
  NO2        m0431(.A(mai_mai_n62_), .B(e), .Y(mai_mai_n460_));
  NA4        m0432(.A(mai_mai_n314_), .B(mai_mai_n164_), .C(mai_mai_n259_), .D(mai_mai_n118_), .Y(mai_mai_n461_));
  AOI220     m0433(.A0(mai_mai_n461_), .A1(mai_mai_n460_), .B0(mai_mai_n459_), .B1(mai_mai_n458_), .Y(mai_mai_n462_));
  AOI210     m0434(.A0(mai_mai_n462_), .A1(mai_mai_n457_), .B0(mai_mai_n454_), .Y(mai_mai_n463_));
  NO2        m0435(.A(mai_mai_n211_), .B(mai_mai_n207_), .Y(mai_mai_n464_));
  NOi21      m0436(.An(a), .B(b), .Y(mai_mai_n465_));
  NA3        m0437(.A(e), .B(d), .C(c), .Y(mai_mai_n466_));
  NAi21      m0438(.An(mai_mai_n466_), .B(mai_mai_n465_), .Y(mai_mai_n467_));
  NO2        m0439(.A(mai_mai_n411_), .B(mai_mai_n206_), .Y(mai_mai_n468_));
  NOi21      m0440(.An(mai_mai_n467_), .B(mai_mai_n468_), .Y(mai_mai_n469_));
  AOI210     m0441(.A0(mai_mai_n268_), .A1(mai_mai_n464_), .B0(mai_mai_n469_), .Y(mai_mai_n470_));
  NO4        m0442(.A(mai_mai_n189_), .B(mai_mai_n101_), .C(mai_mai_n55_), .D(b), .Y(mai_mai_n471_));
  NA2        m0443(.A(mai_mai_n371_), .B(mai_mai_n153_), .Y(mai_mai_n472_));
  OR2        m0444(.A(k), .B(j), .Y(mai_mai_n473_));
  NA2        m0445(.A(l), .B(k), .Y(mai_mai_n474_));
  AOI210     m0446(.A0(mai_mai_n235_), .A1(mai_mai_n332_), .B0(mai_mai_n82_), .Y(mai_mai_n475_));
  NA2        m0447(.A(mai_mai_n128_), .B(mai_mai_n126_), .Y(mai_mai_n476_));
  NA2        m0448(.A(mai_mai_n384_), .B(mai_mai_n112_), .Y(mai_mai_n477_));
  NO4        m0449(.A(mai_mai_n477_), .B(mai_mai_n92_), .C(mai_mai_n111_), .D(e), .Y(mai_mai_n478_));
  NO3        m0450(.A(mai_mai_n411_), .B(mai_mai_n89_), .C(mai_mai_n131_), .Y(mai_mai_n479_));
  NO4        m0451(.A(mai_mai_n479_), .B(mai_mai_n478_), .C(mai_mai_n476_), .D(mai_mai_n315_), .Y(mai_mai_n480_));
  NA2        m0452(.A(mai_mai_n480_), .B(mai_mai_n472_), .Y(mai_mai_n481_));
  NO4        m0453(.A(mai_mai_n481_), .B(mai_mai_n471_), .C(mai_mai_n470_), .D(mai_mai_n463_), .Y(mai_mai_n482_));
  NA2        m0454(.A(mai_mai_n66_), .B(mai_mai_n63_), .Y(mai_mai_n483_));
  NOi21      m0455(.An(d), .B(e), .Y(mai_mai_n484_));
  NAi31      m0456(.An(j), .B(l), .C(i), .Y(mai_mai_n485_));
  OAI210     m0457(.A0(mai_mai_n485_), .A1(mai_mai_n132_), .B0(mai_mai_n101_), .Y(mai_mai_n486_));
  NO3        m0458(.A(mai_mai_n385_), .B(mai_mai_n340_), .C(mai_mai_n203_), .Y(mai_mai_n487_));
  NO2        m0459(.A(mai_mai_n385_), .B(mai_mai_n362_), .Y(mai_mai_n488_));
  NO4        m0460(.A(mai_mai_n488_), .B(mai_mai_n487_), .C(mai_mai_n185_), .D(mai_mai_n301_), .Y(mai_mai_n489_));
  NA3        m0461(.A(mai_mai_n489_), .B(mai_mai_n483_), .C(mai_mai_n244_), .Y(mai_mai_n490_));
  OAI210     m0462(.A0(mai_mai_n127_), .A1(mai_mai_n125_), .B0(n), .Y(mai_mai_n491_));
  NO2        m0463(.A(mai_mai_n491_), .B(mai_mai_n131_), .Y(mai_mai_n492_));
  OA210      m0464(.A0(mai_mai_n246_), .A1(mai_mai_n492_), .B0(mai_mai_n194_), .Y(mai_mai_n493_));
  XO2        m0465(.A(i), .B(h), .Y(mai_mai_n494_));
  NA3        m0466(.A(mai_mai_n494_), .B(mai_mai_n159_), .C(n), .Y(mai_mai_n495_));
  NAi41      m0467(.An(mai_mai_n293_), .B(mai_mai_n495_), .C(mai_mai_n448_), .D(mai_mai_n373_), .Y(mai_mai_n496_));
  NOi32      m0468(.An(mai_mai_n496_), .Bn(mai_mai_n460_), .C(mai_mai_n270_), .Y(mai_mai_n497_));
  NAi31      m0469(.An(c), .B(f), .C(d), .Y(mai_mai_n498_));
  AOI210     m0470(.A0(mai_mai_n278_), .A1(mai_mai_n197_), .B0(mai_mai_n498_), .Y(mai_mai_n499_));
  NOi21      m0471(.An(mai_mai_n80_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NA3        m0472(.A(mai_mai_n369_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n501_));
  NA2        m0473(.A(mai_mai_n229_), .B(mai_mai_n107_), .Y(mai_mai_n502_));
  AOI210     m0474(.A0(mai_mai_n502_), .A1(mai_mai_n181_), .B0(mai_mai_n498_), .Y(mai_mai_n503_));
  AOI210     m0475(.A0(mai_mai_n351_), .A1(mai_mai_n35_), .B0(mai_mai_n467_), .Y(mai_mai_n504_));
  NOi31      m0476(.An(mai_mai_n501_), .B(mai_mai_n504_), .C(mai_mai_n503_), .Y(mai_mai_n505_));
  AN2        m0477(.A(mai_mai_n165_), .B(mai_mai_n63_), .Y(mai_mai_n506_));
  NA3        m0478(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n507_));
  NO2        m0479(.A(mai_mai_n507_), .B(mai_mai_n423_), .Y(mai_mai_n508_));
  NO2        m0480(.A(mai_mai_n508_), .B(mai_mai_n289_), .Y(mai_mai_n509_));
  NAi41      m0481(.An(mai_mai_n506_), .B(mai_mai_n509_), .C(mai_mai_n505_), .D(mai_mai_n500_), .Y(mai_mai_n510_));
  NO4        m0482(.A(mai_mai_n510_), .B(mai_mai_n497_), .C(mai_mai_n493_), .D(mai_mai_n490_), .Y(mai_mai_n511_));
  NA4        m0483(.A(mai_mai_n511_), .B(mai_mai_n482_), .C(mai_mai_n452_), .D(mai_mai_n418_), .Y(mai11));
  NO2        m0484(.A(mai_mai_n69_), .B(f), .Y(mai_mai_n513_));
  NA2        m0485(.A(j), .B(g), .Y(mai_mai_n514_));
  NAi31      m0486(.An(i), .B(m), .C(l), .Y(mai_mai_n515_));
  NA3        m0487(.A(m), .B(k), .C(j), .Y(mai_mai_n516_));
  OAI220     m0488(.A0(mai_mai_n516_), .A1(mai_mai_n131_), .B0(mai_mai_n515_), .B1(mai_mai_n514_), .Y(mai_mai_n517_));
  NA2        m0489(.A(mai_mai_n517_), .B(mai_mai_n513_), .Y(mai_mai_n518_));
  NOi32      m0490(.An(e), .Bn(b), .C(f), .Y(mai_mai_n519_));
  NA2        m0491(.A(mai_mai_n258_), .B(mai_mai_n112_), .Y(mai_mai_n520_));
  NA2        m0492(.A(mai_mai_n45_), .B(j), .Y(mai_mai_n521_));
  NO2        m0493(.A(mai_mai_n521_), .B(mai_mai_n295_), .Y(mai_mai_n522_));
  NAi31      m0494(.An(d), .B(e), .C(a), .Y(mai_mai_n523_));
  NO2        m0495(.A(mai_mai_n523_), .B(n), .Y(mai_mai_n524_));
  AOI220     m0496(.A0(mai_mai_n524_), .A1(mai_mai_n99_), .B0(mai_mai_n522_), .B1(mai_mai_n519_), .Y(mai_mai_n525_));
  NAi41      m0497(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n526_));
  AN2        m0498(.A(mai_mai_n526_), .B(mai_mai_n361_), .Y(mai_mai_n527_));
  AOI210     m0499(.A0(mai_mai_n527_), .A1(mai_mai_n385_), .B0(mai_mai_n271_), .Y(mai_mai_n528_));
  NA2        m0500(.A(j), .B(i), .Y(mai_mai_n529_));
  NAi31      m0501(.An(n), .B(m), .C(k), .Y(mai_mai_n530_));
  NO3        m0502(.A(mai_mai_n530_), .B(mai_mai_n529_), .C(mai_mai_n111_), .Y(mai_mai_n531_));
  NO4        m0503(.A(n), .B(d), .C(mai_mai_n115_), .D(a), .Y(mai_mai_n532_));
  OR2        m0504(.A(n), .B(c), .Y(mai_mai_n533_));
  NO2        m0505(.A(mai_mai_n533_), .B(mai_mai_n149_), .Y(mai_mai_n534_));
  NO2        m0506(.A(mai_mai_n534_), .B(mai_mai_n532_), .Y(mai_mai_n535_));
  NOi32      m0507(.An(g), .Bn(f), .C(i), .Y(mai_mai_n536_));
  NA2        m0508(.A(mai_mai_n517_), .B(f), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n273_), .B(mai_mai_n48_), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n537_), .B(mai_mai_n535_), .Y(mai_mai_n539_));
  AOI210     m0511(.A0(mai_mai_n531_), .A1(mai_mai_n528_), .B0(mai_mai_n539_), .Y(mai_mai_n540_));
  NA2        m0512(.A(mai_mai_n140_), .B(mai_mai_n34_), .Y(mai_mai_n541_));
  OAI220     m0513(.A0(mai_mai_n541_), .A1(m), .B0(mai_mai_n521_), .B1(mai_mai_n235_), .Y(mai_mai_n542_));
  NOi41      m0514(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n543_));
  NAi32      m0515(.An(e), .Bn(b), .C(c), .Y(mai_mai_n544_));
  OR2        m0516(.A(mai_mai_n544_), .B(mai_mai_n82_), .Y(mai_mai_n545_));
  AN2        m0517(.A(mai_mai_n333_), .B(mai_mai_n311_), .Y(mai_mai_n546_));
  NA2        m0518(.A(mai_mai_n546_), .B(mai_mai_n545_), .Y(mai_mai_n547_));
  OA210      m0519(.A0(mai_mai_n547_), .A1(mai_mai_n543_), .B0(mai_mai_n542_), .Y(mai_mai_n548_));
  OAI220     m0520(.A0(mai_mai_n387_), .A1(mai_mai_n386_), .B0(mai_mai_n515_), .B1(mai_mai_n514_), .Y(mai_mai_n549_));
  NO3        m0521(.A(mai_mai_n60_), .B(mai_mai_n48_), .C(mai_mai_n215_), .Y(mai_mai_n550_));
  NO2        m0522(.A(mai_mai_n232_), .B(mai_mai_n109_), .Y(mai_mai_n551_));
  OAI210     m0523(.A0(mai_mai_n550_), .A1(mai_mai_n388_), .B0(mai_mai_n551_), .Y(mai_mai_n552_));
  INV        m0524(.A(mai_mai_n552_), .Y(mai_mai_n553_));
  NO2        m0525(.A(mai_mai_n275_), .B(n), .Y(mai_mai_n554_));
  NO2        m0526(.A(mai_mai_n413_), .B(mai_mai_n554_), .Y(mai_mai_n555_));
  NA2        m0527(.A(mai_mai_n549_), .B(f), .Y(mai_mai_n556_));
  NAi32      m0528(.An(d), .Bn(a), .C(b), .Y(mai_mai_n557_));
  NA2        m0529(.A(h), .B(f), .Y(mai_mai_n558_));
  NO2        m0530(.A(mai_mai_n558_), .B(mai_mai_n92_), .Y(mai_mai_n559_));
  NO3        m0531(.A(mai_mai_n177_), .B(mai_mai_n174_), .C(g), .Y(mai_mai_n560_));
  NA2        m0532(.A(mai_mai_n560_), .B(mai_mai_n57_), .Y(mai_mai_n561_));
  OAI210     m0533(.A0(mai_mai_n556_), .A1(mai_mai_n555_), .B0(mai_mai_n561_), .Y(mai_mai_n562_));
  AN3        m0534(.A(j), .B(h), .C(g), .Y(mai_mai_n563_));
  NO2        m0535(.A(mai_mai_n146_), .B(c), .Y(mai_mai_n564_));
  NA3        m0536(.A(mai_mai_n564_), .B(mai_mai_n563_), .C(mai_mai_n447_), .Y(mai_mai_n565_));
  NA3        m0537(.A(f), .B(d), .C(b), .Y(mai_mai_n566_));
  NO4        m0538(.A(mai_mai_n566_), .B(mai_mai_n177_), .C(mai_mai_n174_), .D(g), .Y(mai_mai_n567_));
  NAi21      m0539(.An(mai_mai_n567_), .B(mai_mai_n565_), .Y(mai_mai_n568_));
  NO4        m0540(.A(mai_mai_n568_), .B(mai_mai_n562_), .C(mai_mai_n553_), .D(mai_mai_n548_), .Y(mai_mai_n569_));
  AN4        m0541(.A(mai_mai_n569_), .B(mai_mai_n540_), .C(mai_mai_n525_), .D(mai_mai_n518_), .Y(mai_mai_n570_));
  INV        m0542(.A(k), .Y(mai_mai_n571_));
  NA3        m0543(.A(l), .B(mai_mai_n571_), .C(i), .Y(mai_mai_n572_));
  INV        m0544(.A(mai_mai_n572_), .Y(mai_mai_n573_));
  NA4        m0545(.A(mai_mai_n384_), .B(mai_mai_n404_), .C(mai_mai_n182_), .D(mai_mai_n112_), .Y(mai_mai_n574_));
  NAi32      m0546(.An(h), .Bn(f), .C(g), .Y(mai_mai_n575_));
  NAi41      m0547(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n576_));
  OAI210     m0548(.A0(mai_mai_n523_), .A1(n), .B0(mai_mai_n576_), .Y(mai_mai_n577_));
  NA2        m0549(.A(mai_mai_n577_), .B(m), .Y(mai_mai_n578_));
  NAi31      m0550(.An(h), .B(g), .C(f), .Y(mai_mai_n579_));
  OR2        m0551(.A(mai_mai_n578_), .B(mai_mai_n575_), .Y(mai_mai_n580_));
  NA2        m0552(.A(mai_mai_n580_), .B(mai_mai_n574_), .Y(mai_mai_n581_));
  NAi31      m0553(.An(f), .B(h), .C(g), .Y(mai_mai_n582_));
  NO4        m0554(.A(mai_mai_n305_), .B(mai_mai_n582_), .C(mai_mai_n69_), .D(mai_mai_n71_), .Y(mai_mai_n583_));
  NOi32      m0555(.An(b), .Bn(a), .C(c), .Y(mai_mai_n584_));
  NOi32      m0556(.An(d), .Bn(a), .C(e), .Y(mai_mai_n585_));
  NA2        m0557(.A(mai_mai_n585_), .B(mai_mai_n112_), .Y(mai_mai_n586_));
  NO2        m0558(.A(n), .B(c), .Y(mai_mai_n587_));
  NAi32      m0559(.An(n), .Bn(f), .C(m), .Y(mai_mai_n588_));
  NOi32      m0560(.An(e), .Bn(a), .C(d), .Y(mai_mai_n589_));
  AOI210     m0561(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n589_), .Y(mai_mai_n590_));
  NO2        m0562(.A(mai_mai_n590_), .B(mai_mai_n541_), .Y(mai_mai_n591_));
  AOI210     m0563(.A0(mai_mai_n591_), .A1(mai_mai_n1499_), .B0(mai_mai_n583_), .Y(mai_mai_n592_));
  INV        m0564(.A(mai_mai_n592_), .Y(mai_mai_n593_));
  AOI210     m0565(.A0(mai_mai_n581_), .A1(mai_mai_n573_), .B0(mai_mai_n593_), .Y(mai_mai_n594_));
  NO3        m0566(.A(mai_mai_n309_), .B(mai_mai_n59_), .C(n), .Y(mai_mai_n595_));
  NA3        m0567(.A(mai_mai_n498_), .B(mai_mai_n172_), .C(mai_mai_n171_), .Y(mai_mai_n596_));
  NA2        m0568(.A(mai_mai_n449_), .B(mai_mai_n232_), .Y(mai_mai_n597_));
  OR2        m0569(.A(mai_mai_n597_), .B(mai_mai_n596_), .Y(mai_mai_n598_));
  NA2        m0570(.A(mai_mai_n72_), .B(mai_mai_n112_), .Y(mai_mai_n599_));
  NO2        m0571(.A(mai_mai_n599_), .B(mai_mai_n44_), .Y(mai_mai_n600_));
  AOI220     m0572(.A0(mai_mai_n600_), .A1(mai_mai_n528_), .B0(mai_mai_n598_), .B1(mai_mai_n595_), .Y(mai_mai_n601_));
  NO2        m0573(.A(mai_mai_n601_), .B(mai_mai_n85_), .Y(mai_mai_n602_));
  NOi32      m0574(.An(e), .Bn(c), .C(f), .Y(mai_mai_n603_));
  NOi21      m0575(.An(f), .B(g), .Y(mai_mai_n604_));
  NO2        m0576(.A(mai_mai_n604_), .B(mai_mai_n212_), .Y(mai_mai_n605_));
  AOI220     m0577(.A0(mai_mai_n605_), .A1(mai_mai_n381_), .B0(mai_mai_n603_), .B1(mai_mai_n176_), .Y(mai_mai_n606_));
  NA2        m0578(.A(mai_mai_n606_), .B(mai_mai_n179_), .Y(mai_mai_n607_));
  AOI210     m0579(.A0(mai_mai_n527_), .A1(mai_mai_n385_), .B0(mai_mai_n294_), .Y(mai_mai_n608_));
  NA2        m0580(.A(mai_mai_n608_), .B(mai_mai_n263_), .Y(mai_mai_n609_));
  NOi21      m0581(.An(j), .B(l), .Y(mai_mai_n610_));
  NAi21      m0582(.An(k), .B(h), .Y(mai_mai_n611_));
  NO2        m0583(.A(mai_mai_n611_), .B(mai_mai_n261_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n610_), .Y(mai_mai_n613_));
  OR2        m0585(.A(mai_mai_n613_), .B(mai_mai_n578_), .Y(mai_mai_n614_));
  NOi31      m0586(.An(m), .B(n), .C(k), .Y(mai_mai_n615_));
  NA2        m0587(.A(mai_mai_n610_), .B(mai_mai_n615_), .Y(mai_mai_n616_));
  NO2        m0588(.A(mai_mai_n275_), .B(mai_mai_n48_), .Y(mai_mai_n617_));
  NO2        m0589(.A(mai_mai_n305_), .B(mai_mai_n582_), .Y(mai_mai_n618_));
  NO2        m0590(.A(mai_mai_n523_), .B(mai_mai_n48_), .Y(mai_mai_n619_));
  AOI220     m0591(.A0(mai_mai_n619_), .A1(mai_mai_n618_), .B0(mai_mai_n617_), .B1(mai_mai_n559_), .Y(mai_mai_n620_));
  NA3        m0592(.A(mai_mai_n620_), .B(mai_mai_n614_), .C(mai_mai_n609_), .Y(mai_mai_n621_));
  NA2        m0593(.A(mai_mai_n107_), .B(mai_mai_n36_), .Y(mai_mai_n622_));
  NO2        m0594(.A(k), .B(mai_mai_n215_), .Y(mai_mai_n623_));
  INV        m0595(.A(mai_mai_n353_), .Y(mai_mai_n624_));
  NO2        m0596(.A(mai_mai_n624_), .B(n), .Y(mai_mai_n625_));
  NAi31      m0597(.An(mai_mai_n622_), .B(mai_mai_n625_), .C(mai_mai_n623_), .Y(mai_mai_n626_));
  NO2        m0598(.A(mai_mai_n521_), .B(mai_mai_n177_), .Y(mai_mai_n627_));
  NA3        m0599(.A(mai_mai_n544_), .B(mai_mai_n270_), .C(mai_mai_n144_), .Y(mai_mai_n628_));
  NA2        m0600(.A(mai_mai_n494_), .B(mai_mai_n159_), .Y(mai_mai_n629_));
  NO3        m0601(.A(mai_mai_n382_), .B(mai_mai_n629_), .C(mai_mai_n85_), .Y(mai_mai_n630_));
  AOI210     m0602(.A0(mai_mai_n628_), .A1(mai_mai_n627_), .B0(mai_mai_n630_), .Y(mai_mai_n631_));
  AN3        m0603(.A(f), .B(d), .C(b), .Y(mai_mai_n632_));
  OAI210     m0604(.A0(mai_mai_n632_), .A1(mai_mai_n130_), .B0(n), .Y(mai_mai_n633_));
  NA3        m0605(.A(mai_mai_n494_), .B(mai_mai_n159_), .C(mai_mai_n215_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(mai_mai_n633_), .A1(mai_mai_n234_), .B0(mai_mai_n634_), .Y(mai_mai_n635_));
  NAi31      m0607(.An(m), .B(n), .C(k), .Y(mai_mai_n636_));
  OR2        m0608(.A(mai_mai_n135_), .B(mai_mai_n59_), .Y(mai_mai_n637_));
  OAI210     m0609(.A0(mai_mai_n637_), .A1(mai_mai_n636_), .B0(mai_mai_n250_), .Y(mai_mai_n638_));
  OAI210     m0610(.A0(mai_mai_n638_), .A1(mai_mai_n635_), .B0(j), .Y(mai_mai_n639_));
  NA3        m0611(.A(mai_mai_n639_), .B(mai_mai_n631_), .C(mai_mai_n626_), .Y(mai_mai_n640_));
  NO4        m0612(.A(mai_mai_n640_), .B(mai_mai_n621_), .C(mai_mai_n607_), .D(mai_mai_n602_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n369_), .B(mai_mai_n161_), .Y(mai_mai_n642_));
  NAi31      m0614(.An(g), .B(h), .C(f), .Y(mai_mai_n643_));
  OA210      m0615(.A0(mai_mai_n523_), .A1(n), .B0(mai_mai_n576_), .Y(mai_mai_n644_));
  NO2        m0616(.A(mai_mai_n644_), .B(mai_mai_n88_), .Y(mai_mai_n645_));
  INV        m0617(.A(mai_mai_n645_), .Y(mai_mai_n646_));
  AOI210     m0618(.A0(mai_mai_n646_), .A1(mai_mai_n642_), .B0(mai_mai_n516_), .Y(mai_mai_n647_));
  NO3        m0619(.A(g), .B(mai_mai_n214_), .C(mai_mai_n55_), .Y(mai_mai_n648_));
  NAi21      m0620(.An(h), .B(j), .Y(mai_mai_n649_));
  NA2        m0621(.A(mai_mai_n381_), .B(mai_mai_n648_), .Y(mai_mai_n650_));
  OR2        m0622(.A(mai_mai_n69_), .B(mai_mai_n71_), .Y(mai_mai_n651_));
  NA2        m0623(.A(mai_mai_n584_), .B(mai_mai_n337_), .Y(mai_mai_n652_));
  OA220      m0624(.A0(mai_mai_n616_), .A1(mai_mai_n652_), .B0(mai_mai_n613_), .B1(mai_mai_n651_), .Y(mai_mai_n653_));
  AN2        m0625(.A(h), .B(f), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n654_), .B(mai_mai_n37_), .Y(mai_mai_n655_));
  NA2        m0627(.A(mai_mai_n97_), .B(mai_mai_n45_), .Y(mai_mai_n656_));
  OAI220     m0628(.A0(mai_mai_n656_), .A1(mai_mai_n326_), .B0(mai_mai_n655_), .B1(mai_mai_n454_), .Y(mai_mai_n657_));
  AOI210     m0629(.A0(mai_mai_n557_), .A1(mai_mai_n412_), .B0(mai_mai_n48_), .Y(mai_mai_n658_));
  OAI220     m0630(.A0(mai_mai_n579_), .A1(mai_mai_n572_), .B0(mai_mai_n319_), .B1(mai_mai_n514_), .Y(mai_mai_n659_));
  AOI210     m0631(.A0(mai_mai_n659_), .A1(mai_mai_n658_), .B0(mai_mai_n657_), .Y(mai_mai_n660_));
  NA3        m0632(.A(mai_mai_n660_), .B(mai_mai_n653_), .C(mai_mai_n650_), .Y(mai_mai_n661_));
  NO2        m0633(.A(mai_mai_n251_), .B(f), .Y(mai_mai_n662_));
  NO2        m0634(.A(mai_mai_n604_), .B(mai_mai_n59_), .Y(mai_mai_n663_));
  NO3        m0635(.A(mai_mai_n663_), .B(mai_mai_n662_), .C(mai_mai_n34_), .Y(mai_mai_n664_));
  NA2        m0636(.A(mai_mai_n322_), .B(mai_mai_n140_), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n132_), .B(mai_mai_n48_), .Y(mai_mai_n666_));
  OR2        m0638(.A(mai_mai_n351_), .B(mai_mai_n110_), .Y(mai_mai_n667_));
  OAI210     m0639(.A0(mai_mai_n665_), .A1(mai_mai_n664_), .B0(mai_mai_n667_), .Y(mai_mai_n668_));
  NO3        m0640(.A(mai_mai_n392_), .B(mai_mai_n194_), .C(mai_mai_n193_), .Y(mai_mai_n669_));
  NA2        m0641(.A(mai_mai_n669_), .B(mai_mai_n232_), .Y(mai_mai_n670_));
  NA3        m0642(.A(mai_mai_n670_), .B(mai_mai_n253_), .C(j), .Y(mai_mai_n671_));
  NO3        m0643(.A(mai_mai_n449_), .B(mai_mai_n174_), .C(i), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n453_), .B(mai_mai_n82_), .Y(mai_mai_n673_));
  NO4        m0645(.A(mai_mai_n516_), .B(mai_mai_n673_), .C(mai_mai_n131_), .D(mai_mai_n214_), .Y(mai_mai_n674_));
  INV        m0646(.A(mai_mai_n674_), .Y(mai_mai_n675_));
  NA4        m0647(.A(mai_mai_n675_), .B(mai_mai_n671_), .C(mai_mai_n501_), .D(mai_mai_n390_), .Y(mai_mai_n676_));
  NO4        m0648(.A(mai_mai_n676_), .B(mai_mai_n668_), .C(mai_mai_n661_), .D(mai_mai_n647_), .Y(mai_mai_n677_));
  NA4        m0649(.A(mai_mai_n677_), .B(mai_mai_n641_), .C(mai_mai_n594_), .D(mai_mai_n570_), .Y(mai08));
  NO2        m0650(.A(k), .B(h), .Y(mai_mai_n679_));
  AO210      m0651(.A0(mai_mai_n251_), .A1(mai_mai_n437_), .B0(mai_mai_n679_), .Y(mai_mai_n680_));
  NO2        m0652(.A(mai_mai_n680_), .B(mai_mai_n292_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n603_), .B(mai_mai_n82_), .Y(mai_mai_n682_));
  NA2        m0654(.A(mai_mai_n682_), .B(mai_mai_n449_), .Y(mai_mai_n683_));
  AOI210     m0655(.A0(mai_mai_n683_), .A1(mai_mai_n681_), .B0(mai_mai_n479_), .Y(mai_mai_n684_));
  NA2        m0656(.A(mai_mai_n82_), .B(mai_mai_n109_), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n685_), .B(mai_mai_n56_), .Y(mai_mai_n686_));
  NO4        m0658(.A(mai_mai_n366_), .B(mai_mai_n111_), .C(j), .D(mai_mai_n215_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n566_), .B(mai_mai_n234_), .Y(mai_mai_n688_));
  AOI220     m0660(.A0(mai_mai_n688_), .A1(mai_mai_n343_), .B0(mai_mai_n687_), .B1(mai_mai_n686_), .Y(mai_mai_n689_));
  AOI210     m0661(.A0(mai_mai_n566_), .A1(mai_mai_n155_), .B0(mai_mai_n82_), .Y(mai_mai_n690_));
  NA4        m0662(.A(mai_mai_n217_), .B(mai_mai_n140_), .C(mai_mai_n44_), .D(h), .Y(mai_mai_n691_));
  AN2        m0663(.A(l), .B(k), .Y(mai_mai_n692_));
  NA3        m0664(.A(mai_mai_n689_), .B(mai_mai_n684_), .C(mai_mai_n345_), .Y(mai_mai_n693_));
  AN2        m0665(.A(mai_mai_n524_), .B(mai_mai_n93_), .Y(mai_mai_n694_));
  NO4        m0666(.A(mai_mai_n174_), .B(mai_mai_n380_), .C(mai_mai_n111_), .D(g), .Y(mai_mai_n695_));
  AOI210     m0667(.A0(mai_mai_n695_), .A1(mai_mai_n688_), .B0(mai_mai_n508_), .Y(mai_mai_n696_));
  NO2        m0668(.A(mai_mai_n38_), .B(mai_mai_n214_), .Y(mai_mai_n697_));
  AOI220     m0669(.A0(mai_mai_n605_), .A1(mai_mai_n342_), .B0(mai_mai_n697_), .B1(mai_mai_n554_), .Y(mai_mai_n698_));
  NAi31      m0670(.An(mai_mai_n694_), .B(mai_mai_n698_), .C(mai_mai_n696_), .Y(mai_mai_n699_));
  OAI210     m0671(.A0(mai_mai_n544_), .A1(mai_mai_n46_), .B0(mai_mai_n637_), .Y(mai_mai_n700_));
  NO2        m0672(.A(mai_mai_n474_), .B(mai_mai_n132_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n701_), .B(mai_mai_n700_), .Y(mai_mai_n702_));
  NO3        m0674(.A(mai_mai_n309_), .B(mai_mai_n131_), .C(mai_mai_n40_), .Y(mai_mai_n703_));
  BUFFER     m0675(.A(mai_mai_n703_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n680_), .B(mai_mai_n136_), .Y(mai_mai_n705_));
  AOI220     m0677(.A0(mai_mai_n705_), .A1(mai_mai_n391_), .B0(mai_mai_n704_), .B1(mai_mai_n74_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n702_), .B(mai_mai_n706_), .Y(mai_mai_n707_));
  NA3        m0679(.A(mai_mai_n670_), .B(mai_mai_n328_), .C(mai_mai_n372_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n692_), .B(mai_mai_n222_), .Y(mai_mai_n709_));
  NO2        m0681(.A(mai_mai_n709_), .B(mai_mai_n321_), .Y(mai_mai_n710_));
  AOI210     m0682(.A0(mai_mai_n710_), .A1(mai_mai_n662_), .B0(mai_mai_n478_), .Y(mai_mai_n711_));
  NA3        m0683(.A(m), .B(l), .C(k), .Y(mai_mai_n712_));
  NO2        m0684(.A(mai_mai_n526_), .B(mai_mai_n271_), .Y(mai_mai_n713_));
  NOi21      m0685(.An(mai_mai_n713_), .B(mai_mai_n520_), .Y(mai_mai_n714_));
  NA4        m0686(.A(mai_mai_n112_), .B(l), .C(k), .D(mai_mai_n85_), .Y(mai_mai_n715_));
  NA3        m0687(.A(mai_mai_n120_), .B(mai_mai_n400_), .C(i), .Y(mai_mai_n716_));
  NO2        m0688(.A(mai_mai_n716_), .B(mai_mai_n715_), .Y(mai_mai_n717_));
  NO2        m0689(.A(mai_mai_n717_), .B(mai_mai_n714_), .Y(mai_mai_n718_));
  NA3        m0690(.A(mai_mai_n718_), .B(mai_mai_n711_), .C(mai_mai_n708_), .Y(mai_mai_n719_));
  NO4        m0691(.A(mai_mai_n719_), .B(mai_mai_n707_), .C(mai_mai_n699_), .D(mai_mai_n693_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n605_), .B(mai_mai_n381_), .Y(mai_mai_n721_));
  NOi31      m0693(.An(g), .B(h), .C(f), .Y(mai_mai_n722_));
  NA2        m0694(.A(mai_mai_n619_), .B(mai_mai_n722_), .Y(mai_mai_n723_));
  OR2        m0695(.A(mai_mai_n723_), .B(mai_mai_n529_), .Y(mai_mai_n724_));
  NO3        m0696(.A(mai_mai_n385_), .B(mai_mai_n514_), .C(h), .Y(mai_mai_n725_));
  AOI210     m0697(.A0(mai_mai_n725_), .A1(mai_mai_n112_), .B0(mai_mai_n488_), .Y(mai_mai_n726_));
  NA4        m0698(.A(mai_mai_n726_), .B(mai_mai_n724_), .C(mai_mai_n721_), .D(mai_mai_n250_), .Y(mai_mai_n727_));
  NA2        m0699(.A(mai_mai_n692_), .B(mai_mai_n71_), .Y(mai_mai_n728_));
  NO4        m0700(.A(mai_mai_n669_), .B(mai_mai_n174_), .C(n), .D(i), .Y(mai_mai_n729_));
  NOi21      m0701(.An(h), .B(j), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n730_), .B(f), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n729_), .B(mai_mai_n672_), .Y(mai_mai_n732_));
  NO2        m0704(.A(mai_mai_n732_), .B(mai_mai_n728_), .Y(mai_mai_n733_));
  AOI210     m0705(.A0(mai_mai_n727_), .A1(l), .B0(mai_mai_n733_), .Y(mai_mai_n734_));
  NO2        m0706(.A(j), .B(i), .Y(mai_mai_n735_));
  NA3        m0707(.A(mai_mai_n735_), .B(mai_mai_n78_), .C(l), .Y(mai_mai_n736_));
  NA2        m0708(.A(mai_mai_n735_), .B(mai_mai_n33_), .Y(mai_mai_n737_));
  OR2        m0709(.A(mai_mai_n736_), .B(mai_mai_n578_), .Y(mai_mai_n738_));
  NO3        m0710(.A(mai_mai_n151_), .B(mai_mai_n48_), .C(mai_mai_n109_), .Y(mai_mai_n739_));
  NO3        m0711(.A(mai_mai_n533_), .B(mai_mai_n149_), .C(mai_mai_n71_), .Y(mai_mai_n740_));
  NO3        m0712(.A(mai_mai_n474_), .B(mai_mai_n424_), .C(j), .Y(mai_mai_n741_));
  OAI210     m0713(.A0(mai_mai_n740_), .A1(mai_mai_n739_), .B0(mai_mai_n741_), .Y(mai_mai_n742_));
  OAI210     m0714(.A0(mai_mai_n723_), .A1(mai_mai_n60_), .B0(mai_mai_n742_), .Y(mai_mai_n743_));
  NA2        m0715(.A(k), .B(j), .Y(mai_mai_n744_));
  NO3        m0716(.A(mai_mai_n292_), .B(mai_mai_n744_), .C(mai_mai_n39_), .Y(mai_mai_n745_));
  AOI210     m0717(.A0(mai_mai_n519_), .A1(n), .B0(mai_mai_n543_), .Y(mai_mai_n746_));
  NA2        m0718(.A(mai_mai_n746_), .B(mai_mai_n546_), .Y(mai_mai_n747_));
  AN3        m0719(.A(mai_mai_n747_), .B(mai_mai_n745_), .C(mai_mai_n96_), .Y(mai_mai_n748_));
  NA2        m0720(.A(mai_mai_n597_), .B(mai_mai_n303_), .Y(mai_mai_n749_));
  NAi31      m0721(.An(mai_mai_n590_), .B(mai_mai_n90_), .C(mai_mai_n82_), .Y(mai_mai_n750_));
  NA2        m0722(.A(mai_mai_n750_), .B(mai_mai_n749_), .Y(mai_mai_n751_));
  NO2        m0723(.A(mai_mai_n292_), .B(mai_mai_n136_), .Y(mai_mai_n752_));
  AOI220     m0724(.A0(mai_mai_n752_), .A1(mai_mai_n605_), .B0(mai_mai_n703_), .B1(mai_mai_n690_), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n712_), .B(mai_mai_n88_), .Y(mai_mai_n754_));
  NA2        m0726(.A(mai_mai_n754_), .B(mai_mai_n577_), .Y(mai_mai_n755_));
  NO2        m0727(.A(mai_mai_n579_), .B(mai_mai_n116_), .Y(mai_mai_n756_));
  OAI210     m0728(.A0(mai_mai_n756_), .A1(mai_mai_n741_), .B0(mai_mai_n658_), .Y(mai_mai_n757_));
  NA3        m0729(.A(mai_mai_n757_), .B(mai_mai_n755_), .C(mai_mai_n753_), .Y(mai_mai_n758_));
  OR4        m0730(.A(mai_mai_n758_), .B(mai_mai_n751_), .C(mai_mai_n748_), .D(mai_mai_n743_), .Y(mai_mai_n759_));
  NA3        m0731(.A(mai_mai_n746_), .B(mai_mai_n546_), .C(mai_mai_n545_), .Y(mai_mai_n760_));
  NA4        m0732(.A(mai_mai_n760_), .B(mai_mai_n217_), .C(mai_mai_n437_), .D(mai_mai_n34_), .Y(mai_mai_n761_));
  NO4        m0733(.A(mai_mai_n474_), .B(mai_mai_n419_), .C(j), .D(f), .Y(mai_mai_n762_));
  OAI220     m0734(.A0(mai_mai_n691_), .A1(mai_mai_n682_), .B0(mai_mai_n326_), .B1(mai_mai_n38_), .Y(mai_mai_n763_));
  AOI210     m0735(.A0(mai_mai_n762_), .A1(mai_mai_n257_), .B0(mai_mai_n763_), .Y(mai_mai_n764_));
  NA3        m0736(.A(mai_mai_n536_), .B(mai_mai_n285_), .C(h), .Y(mai_mai_n765_));
  NOi21      m0737(.An(mai_mai_n658_), .B(mai_mai_n765_), .Y(mai_mai_n766_));
  NO2        m0738(.A(mai_mai_n89_), .B(mai_mai_n46_), .Y(mai_mai_n767_));
  NO2        m0739(.A(mai_mai_n736_), .B(mai_mai_n651_), .Y(mai_mai_n768_));
  AOI210     m0740(.A0(mai_mai_n767_), .A1(mai_mai_n625_), .B0(mai_mai_n768_), .Y(mai_mai_n769_));
  NAi41      m0741(.An(mai_mai_n766_), .B(mai_mai_n769_), .C(mai_mai_n764_), .D(mai_mai_n761_), .Y(mai_mai_n770_));
  BUFFER     m0742(.A(mai_mai_n93_), .Y(mai_mai_n771_));
  NA2        m0743(.A(mai_mai_n771_), .B(mai_mai_n239_), .Y(mai_mai_n772_));
  NO2        m0744(.A(mai_mai_n644_), .B(mai_mai_n71_), .Y(mai_mai_n773_));
  AOI210     m0745(.A0(mai_mai_n762_), .A1(mai_mai_n773_), .B0(mai_mai_n330_), .Y(mai_mai_n774_));
  OAI210     m0746(.A0(mai_mai_n712_), .A1(mai_mai_n643_), .B0(mai_mai_n507_), .Y(mai_mai_n775_));
  NA3        m0747(.A(mai_mai_n249_), .B(mai_mai_n58_), .C(b), .Y(mai_mai_n776_));
  AOI220     m0748(.A0(mai_mai_n587_), .A1(mai_mai_n29_), .B0(mai_mai_n453_), .B1(mai_mai_n82_), .Y(mai_mai_n777_));
  NA2        m0749(.A(mai_mai_n777_), .B(mai_mai_n776_), .Y(mai_mai_n778_));
  NO2        m0750(.A(mai_mai_n765_), .B(mai_mai_n477_), .Y(mai_mai_n779_));
  AOI210     m0751(.A0(mai_mai_n778_), .A1(mai_mai_n775_), .B0(mai_mai_n779_), .Y(mai_mai_n780_));
  NA3        m0752(.A(mai_mai_n780_), .B(mai_mai_n774_), .C(mai_mai_n772_), .Y(mai_mai_n781_));
  NOi41      m0753(.An(mai_mai_n738_), .B(mai_mai_n781_), .C(mai_mai_n770_), .D(mai_mai_n759_), .Y(mai_mai_n782_));
  NO3        m0754(.A(mai_mai_n336_), .B(mai_mai_n294_), .C(mai_mai_n111_), .Y(mai_mai_n783_));
  NA2        m0755(.A(mai_mai_n783_), .B(mai_mai_n747_), .Y(mai_mai_n784_));
  NA2        m0756(.A(mai_mai_n45_), .B(mai_mai_n55_), .Y(mai_mai_n785_));
  NO3        m0757(.A(mai_mai_n785_), .B(mai_mai_n737_), .C(mai_mai_n275_), .Y(mai_mai_n786_));
  NO3        m0758(.A(mai_mai_n514_), .B(mai_mai_n91_), .C(h), .Y(mai_mai_n787_));
  AOI210     m0759(.A0(mai_mai_n787_), .A1(mai_mai_n686_), .B0(mai_mai_n786_), .Y(mai_mai_n788_));
  NA3        m0760(.A(mai_mai_n788_), .B(mai_mai_n784_), .C(mai_mai_n393_), .Y(mai_mai_n789_));
  OR2        m0761(.A(mai_mai_n643_), .B(mai_mai_n89_), .Y(mai_mai_n790_));
  NOi31      m0762(.An(b), .B(d), .C(a), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n791_), .B(mai_mai_n585_), .Y(mai_mai_n792_));
  NO2        m0764(.A(mai_mai_n792_), .B(n), .Y(mai_mai_n793_));
  NOi21      m0765(.An(mai_mai_n777_), .B(mai_mai_n793_), .Y(mai_mai_n794_));
  NO2        m0766(.A(mai_mai_n794_), .B(mai_mai_n790_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n669_), .B(n), .Y(mai_mai_n796_));
  AOI220     m0768(.A0(mai_mai_n752_), .A1(mai_mai_n648_), .B0(mai_mai_n796_), .B1(mai_mai_n681_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n316_), .B(mai_mai_n238_), .Y(mai_mai_n798_));
  OAI210     m0770(.A0(mai_mai_n93_), .A1(mai_mai_n90_), .B0(mai_mai_n798_), .Y(mai_mai_n799_));
  NA2        m0771(.A(mai_mai_n120_), .B(mai_mai_n82_), .Y(mai_mai_n800_));
  INV        m0772(.A(mai_mai_n799_), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n710_), .B(mai_mai_n34_), .Y(mai_mai_n802_));
  NAi21      m0774(.An(mai_mai_n715_), .B(mai_mai_n420_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n271_), .B(i), .Y(mai_mai_n804_));
  NA2        m0776(.A(mai_mai_n695_), .B(mai_mai_n344_), .Y(mai_mai_n805_));
  AN2        m0777(.A(mai_mai_n805_), .B(mai_mai_n803_), .Y(mai_mai_n806_));
  NAi41      m0778(.An(mai_mai_n801_), .B(mai_mai_n806_), .C(mai_mai_n802_), .D(mai_mai_n797_), .Y(mai_mai_n807_));
  NO3        m0779(.A(mai_mai_n807_), .B(mai_mai_n795_), .C(mai_mai_n789_), .Y(mai_mai_n808_));
  NA4        m0780(.A(mai_mai_n808_), .B(mai_mai_n782_), .C(mai_mai_n734_), .D(mai_mai_n720_), .Y(mai09));
  INV        m0781(.A(mai_mai_n121_), .Y(mai_mai_n810_));
  NA2        m0782(.A(f), .B(e), .Y(mai_mai_n811_));
  NO2        m0783(.A(mai_mai_n227_), .B(mai_mai_n111_), .Y(mai_mai_n812_));
  NA2        m0784(.A(mai_mai_n812_), .B(g), .Y(mai_mai_n813_));
  NA4        m0785(.A(mai_mai_n305_), .B(mai_mai_n164_), .C(mai_mai_n259_), .D(mai_mai_n118_), .Y(mai_mai_n814_));
  AOI210     m0786(.A0(mai_mai_n814_), .A1(g), .B0(mai_mai_n459_), .Y(mai_mai_n815_));
  AOI210     m0787(.A0(mai_mai_n815_), .A1(mai_mai_n813_), .B0(mai_mai_n811_), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n430_), .B(e), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n817_), .B(mai_mai_n498_), .Y(mai_mai_n818_));
  AOI210     m0790(.A0(mai_mai_n816_), .A1(mai_mai_n810_), .B0(mai_mai_n818_), .Y(mai_mai_n819_));
  NA3        m0791(.A(m), .B(l), .C(i), .Y(mai_mai_n820_));
  OAI220     m0792(.A0(mai_mai_n579_), .A1(mai_mai_n820_), .B0(mai_mai_n349_), .B1(mai_mai_n515_), .Y(mai_mai_n821_));
  NA4        m0793(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(g), .D(f), .Y(mai_mai_n822_));
  NAi31      m0794(.An(mai_mai_n821_), .B(mai_mai_n822_), .C(mai_mai_n425_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n790_), .B(mai_mai_n556_), .Y(mai_mai_n824_));
  OA210      m0796(.A0(mai_mai_n824_), .A1(mai_mai_n823_), .B0(mai_mai_n793_), .Y(mai_mai_n825_));
  INV        m0797(.A(mai_mai_n333_), .Y(mai_mai_n826_));
  NO2        m0798(.A(mai_mai_n127_), .B(mai_mai_n125_), .Y(mai_mai_n827_));
  INV        m0799(.A(mai_mai_n335_), .Y(mai_mai_n828_));
  AOI210     m0800(.A0(mai_mai_n828_), .A1(mai_mai_n827_), .B0(mai_mai_n582_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n776_), .B(mai_mai_n326_), .Y(mai_mai_n830_));
  NA2        m0802(.A(mai_mai_n337_), .B(mai_mai_n339_), .Y(mai_mai_n831_));
  OAI210     m0803(.A0(mai_mai_n206_), .A1(mai_mai_n214_), .B0(mai_mai_n831_), .Y(mai_mai_n832_));
  AOI220     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n830_), .B0(mai_mai_n829_), .B1(mai_mai_n826_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n168_), .B(mai_mai_n113_), .Y(mai_mai_n834_));
  NA3        m0806(.A(mai_mai_n834_), .B(mai_mai_n680_), .C(mai_mai_n136_), .Y(mai_mai_n835_));
  NA3        m0807(.A(mai_mai_n835_), .B(mai_mai_n191_), .C(mai_mai_n31_), .Y(mai_mai_n836_));
  NA4        m0808(.A(mai_mai_n836_), .B(mai_mai_n833_), .C(mai_mai_n606_), .D(mai_mai_n80_), .Y(mai_mai_n837_));
  NOi21      m0809(.An(f), .B(d), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n838_), .B(m), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n839_), .B(mai_mai_n51_), .Y(mai_mai_n840_));
  NOi32      m0812(.An(g), .Bn(f), .C(d), .Y(mai_mai_n841_));
  NA4        m0813(.A(mai_mai_n841_), .B(mai_mai_n587_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n840_), .B(mai_mai_n534_), .Y(mai_mai_n843_));
  NA3        m0815(.A(mai_mai_n305_), .B(mai_mai_n259_), .C(mai_mai_n118_), .Y(mai_mai_n844_));
  AN2        m0816(.A(f), .B(d), .Y(mai_mai_n845_));
  NA3        m0817(.A(mai_mai_n465_), .B(mai_mai_n845_), .C(mai_mai_n82_), .Y(mai_mai_n846_));
  NO3        m0818(.A(mai_mai_n846_), .B(mai_mai_n71_), .C(mai_mai_n215_), .Y(mai_mai_n847_));
  NO2        m0819(.A(mai_mai_n282_), .B(mai_mai_n55_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n844_), .B(mai_mai_n847_), .Y(mai_mai_n849_));
  NAi31      m0821(.An(mai_mai_n476_), .B(mai_mai_n849_), .C(mai_mai_n843_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n636_), .B(mai_mai_n321_), .Y(mai_mai_n851_));
  AN2        m0823(.A(mai_mai_n851_), .B(mai_mai_n662_), .Y(mai_mai_n852_));
  INV        m0824(.A(mai_mai_n852_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n585_), .B(mai_mai_n82_), .Y(mai_mai_n854_));
  NO2        m0826(.A(mai_mai_n831_), .B(mai_mai_n854_), .Y(mai_mai_n855_));
  NA3        m0827(.A(mai_mai_n159_), .B(mai_mai_n107_), .C(mai_mai_n106_), .Y(mai_mai_n856_));
  OAI220     m0828(.A0(mai_mai_n846_), .A1(mai_mai_n414_), .B0(mai_mai_n333_), .B1(mai_mai_n856_), .Y(mai_mai_n857_));
  NOi41      m0829(.An(mai_mai_n225_), .B(mai_mai_n857_), .C(mai_mai_n855_), .D(mai_mai_n301_), .Y(mai_mai_n858_));
  NA2        m0830(.A(c), .B(mai_mai_n115_), .Y(mai_mai_n859_));
  NO2        m0831(.A(mai_mai_n859_), .B(mai_mai_n397_), .Y(mai_mai_n860_));
  NA3        m0832(.A(mai_mai_n860_), .B(mai_mai_n496_), .C(f), .Y(mai_mai_n861_));
  OR2        m0833(.A(mai_mai_n643_), .B(mai_mai_n530_), .Y(mai_mai_n862_));
  INV        m0834(.A(mai_mai_n862_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n792_), .B(mai_mai_n110_), .Y(mai_mai_n864_));
  NA2        m0836(.A(mai_mai_n864_), .B(mai_mai_n863_), .Y(mai_mai_n865_));
  NA4        m0837(.A(mai_mai_n865_), .B(mai_mai_n861_), .C(mai_mai_n858_), .D(mai_mai_n853_), .Y(mai_mai_n866_));
  NO4        m0838(.A(mai_mai_n866_), .B(mai_mai_n850_), .C(mai_mai_n837_), .D(mai_mai_n825_), .Y(mai_mai_n867_));
  OR2        m0839(.A(mai_mai_n846_), .B(mai_mai_n71_), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n812_), .B(g), .Y(mai_mai_n869_));
  AOI210     m0841(.A0(mai_mai_n869_), .A1(mai_mai_n286_), .B0(mai_mai_n868_), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n136_), .B(mai_mai_n132_), .Y(mai_mai_n871_));
  NO2        m0843(.A(mai_mai_n232_), .B(mai_mai_n226_), .Y(mai_mai_n872_));
  AOI220     m0844(.A0(mai_mai_n872_), .A1(mai_mai_n229_), .B0(mai_mai_n299_), .B1(mai_mai_n871_), .Y(mai_mai_n873_));
  NO2        m0845(.A(mai_mai_n414_), .B(mai_mai_n811_), .Y(mai_mai_n874_));
  INV        m0846(.A(mai_mai_n873_), .Y(mai_mai_n875_));
  NA2        m0847(.A(e), .B(d), .Y(mai_mai_n876_));
  OAI220     m0848(.A0(mai_mai_n876_), .A1(c), .B0(mai_mai_n316_), .B1(d), .Y(mai_mai_n877_));
  NA3        m0849(.A(mai_mai_n877_), .B(mai_mai_n442_), .C(mai_mai_n494_), .Y(mai_mai_n878_));
  AOI210     m0850(.A0(mai_mai_n502_), .A1(mai_mai_n181_), .B0(mai_mai_n232_), .Y(mai_mai_n879_));
  AOI210     m0851(.A0(mai_mai_n605_), .A1(mai_mai_n342_), .B0(mai_mai_n879_), .Y(mai_mai_n880_));
  NA3        m0852(.A(mai_mai_n167_), .B(mai_mai_n83_), .C(mai_mai_n34_), .Y(mai_mai_n881_));
  NA3        m0853(.A(mai_mai_n881_), .B(mai_mai_n880_), .C(mai_mai_n878_), .Y(mai_mai_n882_));
  NO3        m0854(.A(mai_mai_n882_), .B(mai_mai_n875_), .C(mai_mai_n870_), .Y(mai_mai_n883_));
  NA2        m0855(.A(mai_mai_n826_), .B(mai_mai_n31_), .Y(mai_mai_n884_));
  AO210      m0856(.A0(mai_mai_n884_), .A1(mai_mai_n682_), .B0(mai_mai_n218_), .Y(mai_mai_n885_));
  OAI220     m0857(.A0(mai_mai_n604_), .A1(mai_mai_n59_), .B0(mai_mai_n294_), .B1(j), .Y(mai_mai_n886_));
  AOI220     m0858(.A0(mai_mai_n886_), .A1(mai_mai_n851_), .B0(mai_mai_n595_), .B1(mai_mai_n603_), .Y(mai_mai_n887_));
  OAI210     m0859(.A0(mai_mai_n817_), .A1(mai_mai_n171_), .B0(mai_mai_n887_), .Y(mai_mai_n888_));
  AOI210     m0860(.A0(mai_mai_n117_), .A1(mai_mai_n116_), .B0(mai_mai_n258_), .Y(mai_mai_n889_));
  NO2        m0861(.A(mai_mai_n889_), .B(mai_mai_n842_), .Y(mai_mai_n890_));
  AO210      m0862(.A0(mai_mai_n830_), .A1(mai_mai_n821_), .B0(mai_mai_n890_), .Y(mai_mai_n891_));
  NOi31      m0863(.An(mai_mai_n534_), .B(mai_mai_n839_), .C(mai_mai_n286_), .Y(mai_mai_n892_));
  NO3        m0864(.A(mai_mai_n892_), .B(mai_mai_n891_), .C(mai_mai_n888_), .Y(mai_mai_n893_));
  AO220      m0865(.A0(mai_mai_n442_), .A1(mai_mai_n730_), .B0(mai_mai_n176_), .B1(f), .Y(mai_mai_n894_));
  OAI210     m0866(.A0(mai_mai_n894_), .A1(mai_mai_n445_), .B0(mai_mai_n877_), .Y(mai_mai_n895_));
  NA2        m0867(.A(mai_mai_n824_), .B(mai_mai_n686_), .Y(mai_mai_n896_));
  AN4        m0868(.A(mai_mai_n896_), .B(mai_mai_n895_), .C(mai_mai_n893_), .D(mai_mai_n885_), .Y(mai_mai_n897_));
  NA4        m0869(.A(mai_mai_n897_), .B(mai_mai_n883_), .C(mai_mai_n867_), .D(mai_mai_n819_), .Y(mai12));
  NO2        m0870(.A(mai_mai_n440_), .B(c), .Y(mai_mai_n899_));
  NO4        m0871(.A(mai_mai_n429_), .B(mai_mai_n251_), .C(mai_mai_n571_), .D(mai_mai_n215_), .Y(mai_mai_n900_));
  NA2        m0872(.A(mai_mai_n900_), .B(mai_mai_n899_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n440_), .B(mai_mai_n115_), .Y(mai_mai_n902_));
  NO2        m0874(.A(mai_mai_n827_), .B(mai_mai_n349_), .Y(mai_mai_n903_));
  NO2        m0875(.A(mai_mai_n643_), .B(mai_mai_n366_), .Y(mai_mai_n904_));
  AOI220     m0876(.A0(mai_mai_n904_), .A1(mai_mai_n532_), .B0(mai_mai_n903_), .B1(mai_mai_n902_), .Y(mai_mai_n905_));
  NA3        m0877(.A(mai_mai_n905_), .B(mai_mai_n901_), .C(mai_mai_n428_), .Y(mai_mai_n906_));
  AOI210     m0878(.A0(mai_mai_n235_), .A1(mai_mai_n332_), .B0(mai_mai_n203_), .Y(mai_mai_n907_));
  OR2        m0879(.A(mai_mai_n907_), .B(mai_mai_n900_), .Y(mai_mai_n908_));
  AOI210     m0880(.A0(mai_mai_n329_), .A1(mai_mai_n378_), .B0(mai_mai_n215_), .Y(mai_mai_n909_));
  OAI210     m0881(.A0(mai_mai_n909_), .A1(mai_mai_n908_), .B0(mai_mai_n392_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n622_), .B(mai_mai_n261_), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n579_), .B(mai_mai_n820_), .Y(mai_mai_n912_));
  AOI220     m0884(.A0(mai_mai_n912_), .A1(mai_mai_n554_), .B0(mai_mai_n798_), .B1(mai_mai_n911_), .Y(mai_mai_n913_));
  NO2        m0885(.A(mai_mai_n151_), .B(mai_mai_n238_), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n913_), .B(mai_mai_n910_), .Y(mai_mai_n915_));
  BUFFER     m0887(.A(mai_mai_n317_), .Y(mai_mai_n916_));
  NO3        m0888(.A(mai_mai_n132_), .B(mai_mai_n152_), .C(mai_mai_n215_), .Y(mai_mai_n917_));
  NA2        m0889(.A(mai_mai_n917_), .B(mai_mai_n519_), .Y(mai_mai_n918_));
  NA4        m0890(.A(mai_mai_n430_), .B(mai_mai_n422_), .C(mai_mai_n182_), .D(g), .Y(mai_mai_n919_));
  NA2        m0891(.A(mai_mai_n919_), .B(mai_mai_n918_), .Y(mai_mai_n920_));
  NO3        m0892(.A(mai_mai_n920_), .B(mai_mai_n915_), .C(mai_mai_n906_), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n360_), .B(mai_mai_n359_), .Y(mai_mai_n922_));
  INV        m0894(.A(mai_mai_n576_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n544_), .B(mai_mai_n144_), .Y(mai_mai_n924_));
  NOi21      m0896(.An(mai_mai_n34_), .B(mai_mai_n636_), .Y(mai_mai_n925_));
  AOI220     m0897(.A0(mai_mai_n925_), .A1(mai_mai_n924_), .B0(mai_mai_n923_), .B1(mai_mai_n922_), .Y(mai_mai_n926_));
  OAI210     m0898(.A0(mai_mai_n250_), .A1(mai_mai_n44_), .B0(mai_mai_n926_), .Y(mai_mai_n927_));
  NA2        m0899(.A(mai_mai_n420_), .B(mai_mai_n263_), .Y(mai_mai_n928_));
  NO3        m0900(.A(mai_mai_n800_), .B(mai_mai_n87_), .C(mai_mai_n397_), .Y(mai_mai_n929_));
  NAi31      m0901(.An(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n313_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n48_), .B(mai_mai_n44_), .Y(mai_mai_n931_));
  NO2        m0903(.A(mai_mai_n491_), .B(mai_mai_n294_), .Y(mai_mai_n932_));
  INV        m0904(.A(mai_mai_n932_), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n933_), .B(mai_mai_n144_), .Y(mai_mai_n934_));
  NA2        m0906(.A(mai_mai_n615_), .B(mai_mai_n354_), .Y(mai_mai_n935_));
  OAI210     m0907(.A0(mai_mai_n716_), .A1(mai_mai_n935_), .B0(mai_mai_n358_), .Y(mai_mai_n936_));
  NO4        m0908(.A(mai_mai_n936_), .B(mai_mai_n934_), .C(mai_mai_n930_), .D(mai_mai_n927_), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n342_), .B(g), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n161_), .B(i), .Y(mai_mai_n939_));
  NA2        m0911(.A(mai_mai_n45_), .B(i), .Y(mai_mai_n940_));
  NO2        m0912(.A(mai_mai_n940_), .B(mai_mai_n202_), .Y(mai_mai_n941_));
  INV        m0913(.A(mai_mai_n941_), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n544_), .B(mai_mai_n370_), .Y(mai_mai_n943_));
  AOI210     m0915(.A0(mai_mai_n943_), .A1(n), .B0(mai_mai_n543_), .Y(mai_mai_n944_));
  OAI220     m0916(.A0(mai_mai_n944_), .A1(mai_mai_n938_), .B0(mai_mai_n942_), .B1(mai_mai_n326_), .Y(mai_mai_n945_));
  NO2        m0917(.A(mai_mai_n643_), .B(mai_mai_n485_), .Y(mai_mai_n946_));
  NA3        m0918(.A(mai_mai_n337_), .B(mai_mai_n610_), .C(i), .Y(mai_mai_n947_));
  OAI210     m0919(.A0(mai_mai_n424_), .A1(mai_mai_n305_), .B0(mai_mai_n947_), .Y(mai_mai_n948_));
  OAI220     m0920(.A0(mai_mai_n948_), .A1(mai_mai_n946_), .B0(mai_mai_n658_), .B1(mai_mai_n740_), .Y(mai_mai_n949_));
  NA2        m0921(.A(mai_mai_n589_), .B(mai_mai_n112_), .Y(mai_mai_n950_));
  OR3        m0922(.A(mai_mai_n305_), .B(mai_mai_n419_), .C(f), .Y(mai_mai_n951_));
  NA3        m0923(.A(mai_mai_n610_), .B(mai_mai_n78_), .C(i), .Y(mai_mai_n952_));
  OA220      m0924(.A0(mai_mai_n952_), .A1(mai_mai_n950_), .B0(mai_mai_n951_), .B1(mai_mai_n578_), .Y(mai_mai_n953_));
  NA3        m0925(.A(mai_mai_n318_), .B(mai_mai_n117_), .C(g), .Y(mai_mai_n954_));
  AOI210     m0926(.A0(mai_mai_n655_), .A1(mai_mai_n954_), .B0(m), .Y(mai_mai_n955_));
  OAI210     m0927(.A0(mai_mai_n955_), .A1(mai_mai_n903_), .B0(mai_mai_n317_), .Y(mai_mai_n956_));
  NA2        m0928(.A(mai_mai_n673_), .B(mai_mai_n854_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n822_), .B(mai_mai_n425_), .Y(mai_mai_n958_));
  NA2        m0930(.A(mai_mai_n223_), .B(mai_mai_n75_), .Y(mai_mai_n959_));
  NA3        m0931(.A(mai_mai_n959_), .B(mai_mai_n952_), .C(mai_mai_n951_), .Y(mai_mai_n960_));
  AOI220     m0932(.A0(mai_mai_n960_), .A1(mai_mai_n257_), .B0(mai_mai_n958_), .B1(mai_mai_n957_), .Y(mai_mai_n961_));
  NA4        m0933(.A(mai_mai_n961_), .B(mai_mai_n956_), .C(mai_mai_n953_), .D(mai_mai_n949_), .Y(mai_mai_n962_));
  NA2        m0934(.A(mai_mai_n645_), .B(mai_mai_n86_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n448_), .B(mai_mai_n215_), .Y(mai_mai_n964_));
  AOI220     m0936(.A0(mai_mai_n964_), .A1(mai_mai_n371_), .B0(mai_mai_n916_), .B1(mai_mai_n219_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n904_), .B(mai_mai_n914_), .Y(mai_mai_n966_));
  NA3        m0938(.A(mai_mai_n966_), .B(mai_mai_n965_), .C(mai_mai_n963_), .Y(mai_mai_n967_));
  OAI210     m0939(.A0(mai_mai_n958_), .A1(mai_mai_n912_), .B0(mai_mai_n532_), .Y(mai_mai_n968_));
  OAI210     m0940(.A0(mai_mai_n360_), .A1(mai_mai_n359_), .B0(mai_mai_n108_), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n969_), .B(mai_mai_n524_), .Y(mai_mai_n970_));
  NA2        m0942(.A(mai_mai_n955_), .B(mai_mai_n902_), .Y(mai_mai_n971_));
  NA2        m0943(.A(mai_mai_n627_), .B(mai_mai_n519_), .Y(mai_mai_n972_));
  NA4        m0944(.A(mai_mai_n972_), .B(mai_mai_n971_), .C(mai_mai_n970_), .D(mai_mai_n968_), .Y(mai_mai_n973_));
  NO4        m0945(.A(mai_mai_n973_), .B(mai_mai_n967_), .C(mai_mai_n962_), .D(mai_mai_n945_), .Y(mai_mai_n974_));
  NAi31      m0946(.An(mai_mai_n141_), .B(mai_mai_n407_), .C(n), .Y(mai_mai_n975_));
  NO2        m0947(.A(mai_mai_n125_), .B(mai_mai_n335_), .Y(mai_mai_n976_));
  NO2        m0948(.A(mai_mai_n976_), .B(mai_mai_n975_), .Y(mai_mai_n977_));
  NO3        m0949(.A(mai_mai_n271_), .B(mai_mai_n141_), .C(mai_mai_n397_), .Y(mai_mai_n978_));
  AOI210     m0950(.A0(mai_mai_n978_), .A1(mai_mai_n486_), .B0(mai_mai_n977_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n479_), .B(i), .Y(mai_mai_n980_));
  NA2        m0952(.A(mai_mai_n980_), .B(mai_mai_n979_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n232_), .B(mai_mai_n172_), .Y(mai_mai_n982_));
  NO3        m0954(.A(mai_mai_n303_), .B(mai_mai_n430_), .C(mai_mai_n176_), .Y(mai_mai_n983_));
  NOi31      m0955(.An(mai_mai_n982_), .B(mai_mai_n983_), .C(mai_mai_n215_), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n423_), .B(mai_mai_n854_), .Y(mai_mai_n985_));
  NO3        m0957(.A(mai_mai_n424_), .B(mai_mai_n305_), .C(mai_mai_n71_), .Y(mai_mai_n986_));
  AOI220     m0958(.A0(mai_mai_n986_), .A1(mai_mai_n985_), .B0(mai_mai_n471_), .B1(g), .Y(mai_mai_n987_));
  INV        m0959(.A(mai_mai_n987_), .Y(mai_mai_n988_));
  OAI220     m0960(.A0(mai_mai_n975_), .A1(mai_mai_n235_), .B0(mai_mai_n947_), .B1(mai_mai_n586_), .Y(mai_mai_n989_));
  NA2        m0961(.A(mai_mai_n907_), .B(mai_mai_n899_), .Y(mai_mai_n990_));
  NO3        m0962(.A(mai_mai_n533_), .B(mai_mai_n149_), .C(mai_mai_n214_), .Y(mai_mai_n991_));
  OAI210     m0963(.A0(mai_mai_n991_), .A1(mai_mai_n513_), .B0(mai_mai_n367_), .Y(mai_mai_n992_));
  OAI220     m0964(.A0(mai_mai_n904_), .A1(mai_mai_n912_), .B0(mai_mai_n534_), .B1(mai_mai_n413_), .Y(mai_mai_n993_));
  NA3        m0965(.A(mai_mai_n993_), .B(mai_mai_n992_), .C(mai_mai_n990_), .Y(mai_mai_n994_));
  OAI210     m0966(.A0(mai_mai_n907_), .A1(mai_mai_n900_), .B0(mai_mai_n982_), .Y(mai_mai_n995_));
  NA3        m0967(.A(mai_mai_n943_), .B(mai_mai_n475_), .C(mai_mai_n45_), .Y(mai_mai_n996_));
  AOI210     m0968(.A0(mai_mai_n369_), .A1(mai_mai_n367_), .B0(mai_mai_n325_), .Y(mai_mai_n997_));
  NA3        m0969(.A(mai_mai_n997_), .B(mai_mai_n996_), .C(mai_mai_n995_), .Y(mai_mai_n998_));
  OR3        m0970(.A(mai_mai_n998_), .B(mai_mai_n994_), .C(mai_mai_n989_), .Y(mai_mai_n999_));
  NO4        m0971(.A(mai_mai_n999_), .B(mai_mai_n988_), .C(mai_mai_n984_), .D(mai_mai_n981_), .Y(mai_mai_n1000_));
  NA4        m0972(.A(mai_mai_n1000_), .B(mai_mai_n974_), .C(mai_mai_n937_), .D(mai_mai_n921_), .Y(mai13));
  INV        m0973(.A(mai_mai_n45_), .Y(mai_mai_n1002_));
  AN2        m0974(.A(c), .B(b), .Y(mai_mai_n1003_));
  NA3        m0975(.A(mai_mai_n249_), .B(mai_mai_n1003_), .C(m), .Y(mai_mai_n1004_));
  NA2        m0976(.A(mai_mai_n484_), .B(f), .Y(mai_mai_n1005_));
  NO4        m0977(.A(mai_mai_n1005_), .B(mai_mai_n1004_), .C(mai_mai_n1002_), .D(mai_mai_n572_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n263_), .B(mai_mai_n1003_), .Y(mai_mai_n1007_));
  NO3        m0979(.A(mai_mai_n1007_), .B(mai_mai_n1005_), .C(mai_mai_n939_), .Y(mai_mai_n1008_));
  NAi32      m0980(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1009_));
  NA2        m0981(.A(mai_mai_n140_), .B(mai_mai_n44_), .Y(mai_mai_n1010_));
  NO4        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1009_), .C(mai_mai_n579_), .D(mai_mai_n302_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n649_), .B(mai_mai_n226_), .Y(mai_mai_n1012_));
  NA2        m0984(.A(mai_mai_n400_), .B(mai_mai_n214_), .Y(mai_mai_n1013_));
  AN2        m0985(.A(d), .B(c), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n1014_), .B(mai_mai_n115_), .Y(mai_mai_n1015_));
  NO4        m0987(.A(mai_mai_n1015_), .B(mai_mai_n1013_), .C(mai_mai_n177_), .D(mai_mai_n168_), .Y(mai_mai_n1016_));
  NA2        m0988(.A(mai_mai_n484_), .B(c), .Y(mai_mai_n1017_));
  NO4        m0989(.A(mai_mai_n1010_), .B(mai_mai_n575_), .C(mai_mai_n1017_), .D(mai_mai_n302_), .Y(mai_mai_n1018_));
  AO210      m0990(.A0(mai_mai_n1016_), .A1(mai_mai_n1012_), .B0(mai_mai_n1018_), .Y(mai_mai_n1019_));
  OR4        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1011_), .C(mai_mai_n1008_), .D(mai_mai_n1006_), .Y(mai_mai_n1020_));
  NAi32      m0992(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1021_));
  NO2        m0993(.A(mai_mai_n1021_), .B(mai_mai_n146_), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n1022_), .B(g), .Y(mai_mai_n1023_));
  OR3        m0995(.A(mai_mai_n226_), .B(mai_mai_n177_), .C(mai_mai_n168_), .Y(mai_mai_n1024_));
  NO2        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1023_), .Y(mai_mai_n1025_));
  NO2        m0997(.A(mai_mai_n1017_), .B(mai_mai_n302_), .Y(mai_mai_n1026_));
  NO2        m0998(.A(j), .B(mai_mai_n44_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n612_), .B(mai_mai_n1027_), .Y(mai_mai_n1028_));
  NOi21      m1000(.An(mai_mai_n1026_), .B(mai_mai_n1028_), .Y(mai_mai_n1029_));
  NO2        m1001(.A(mai_mai_n744_), .B(mai_mai_n111_), .Y(mai_mai_n1030_));
  NOi41      m1002(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1030_), .Y(mai_mai_n1032_));
  NO2        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1023_), .Y(mai_mai_n1033_));
  OR3        m1005(.A(e), .B(d), .C(c), .Y(mai_mai_n1034_));
  NA3        m1006(.A(k), .B(j), .C(i), .Y(mai_mai_n1035_));
  NO3        m1007(.A(mai_mai_n1035_), .B(mai_mai_n302_), .C(mai_mai_n88_), .Y(mai_mai_n1036_));
  NOi21      m1008(.An(mai_mai_n1036_), .B(mai_mai_n1034_), .Y(mai_mai_n1037_));
  OR4        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1033_), .C(mai_mai_n1029_), .D(mai_mai_n1025_), .Y(mai_mai_n1038_));
  NA3        m1010(.A(mai_mai_n456_), .B(mai_mai_n328_), .C(mai_mai_n55_), .Y(mai_mai_n1039_));
  NO2        m1011(.A(mai_mai_n1039_), .B(mai_mai_n1028_), .Y(mai_mai_n1040_));
  NO4        m1012(.A(mai_mai_n1039_), .B(mai_mai_n575_), .C(mai_mai_n437_), .D(mai_mai_n44_), .Y(mai_mai_n1041_));
  NO2        m1013(.A(f), .B(c), .Y(mai_mai_n1042_));
  NOi21      m1014(.An(mai_mai_n1042_), .B(mai_mai_n429_), .Y(mai_mai_n1043_));
  NA2        m1015(.A(mai_mai_n1043_), .B(mai_mai_n58_), .Y(mai_mai_n1044_));
  OR2        m1016(.A(k), .B(i), .Y(mai_mai_n1045_));
  NO3        m1017(.A(mai_mai_n1045_), .B(mai_mai_n245_), .C(l), .Y(mai_mai_n1046_));
  NOi31      m1018(.An(mai_mai_n1046_), .B(mai_mai_n1044_), .C(j), .Y(mai_mai_n1047_));
  OR3        m1019(.A(mai_mai_n1047_), .B(mai_mai_n1041_), .C(mai_mai_n1040_), .Y(mai_mai_n1048_));
  OR3        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1038_), .C(mai_mai_n1020_), .Y(mai02));
  OR2        m1021(.A(l), .B(k), .Y(mai_mai_n1050_));
  OR3        m1022(.A(h), .B(g), .C(f), .Y(mai_mai_n1051_));
  OR3        m1023(.A(n), .B(m), .C(i), .Y(mai_mai_n1052_));
  NO4        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1051_), .C(mai_mai_n1050_), .D(mai_mai_n1034_), .Y(mai_mai_n1053_));
  NOi31      m1025(.An(e), .B(d), .C(c), .Y(mai_mai_n1054_));
  AOI210     m1026(.A0(mai_mai_n1036_), .A1(mai_mai_n1054_), .B0(mai_mai_n1011_), .Y(mai_mai_n1055_));
  AN3        m1027(.A(g), .B(f), .C(c), .Y(mai_mai_n1056_));
  NA3        m1028(.A(mai_mai_n1056_), .B(mai_mai_n456_), .C(h), .Y(mai_mai_n1057_));
  OR2        m1029(.A(mai_mai_n1035_), .B(mai_mai_n302_), .Y(mai_mai_n1058_));
  OR2        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1057_), .Y(mai_mai_n1059_));
  NO3        m1031(.A(mai_mai_n1039_), .B(mai_mai_n1010_), .C(mai_mai_n575_), .Y(mai_mai_n1060_));
  NO2        m1032(.A(mai_mai_n1060_), .B(mai_mai_n1025_), .Y(mai_mai_n1061_));
  NA3        m1033(.A(l), .B(k), .C(j), .Y(mai_mai_n1062_));
  NA2        m1034(.A(i), .B(h), .Y(mai_mai_n1063_));
  NO3        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1062_), .C(mai_mai_n132_), .Y(mai_mai_n1064_));
  NO3        m1036(.A(mai_mai_n142_), .B(mai_mai_n281_), .C(mai_mai_n215_), .Y(mai_mai_n1065_));
  AOI210     m1037(.A0(mai_mai_n1065_), .A1(mai_mai_n1064_), .B0(mai_mai_n1029_), .Y(mai_mai_n1066_));
  NA3        m1038(.A(c), .B(b), .C(a), .Y(mai_mai_n1067_));
  NO3        m1039(.A(mai_mai_n1067_), .B(mai_mai_n876_), .C(mai_mai_n214_), .Y(mai_mai_n1068_));
  NO4        m1040(.A(mai_mai_n1035_), .B(mai_mai_n294_), .C(mai_mai_n48_), .D(mai_mai_n111_), .Y(mai_mai_n1069_));
  AOI210     m1041(.A0(mai_mai_n1069_), .A1(mai_mai_n1068_), .B0(mai_mai_n1040_), .Y(mai_mai_n1070_));
  AN4        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1066_), .C(mai_mai_n1061_), .D(mai_mai_n1059_), .Y(mai_mai_n1071_));
  NO2        m1043(.A(mai_mai_n1015_), .B(mai_mai_n1013_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n1032_), .B(mai_mai_n1024_), .Y(mai_mai_n1073_));
  AOI210     m1045(.A0(mai_mai_n1073_), .A1(mai_mai_n1072_), .B0(mai_mai_n1006_), .Y(mai_mai_n1074_));
  NAi41      m1046(.An(mai_mai_n1053_), .B(mai_mai_n1074_), .C(mai_mai_n1071_), .D(mai_mai_n1055_), .Y(mai03));
  NO2        m1047(.A(mai_mai_n515_), .B(mai_mai_n582_), .Y(mai_mai_n1076_));
  NA4        m1048(.A(mai_mai_n563_), .B(m), .C(mai_mai_n111_), .D(mai_mai_n214_), .Y(mai_mai_n1077_));
  INV        m1049(.A(mai_mai_n1077_), .Y(mai_mai_n1078_));
  NO3        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1076_), .C(mai_mai_n969_), .Y(mai_mai_n1079_));
  NOi41      m1051(.An(mai_mai_n790_), .B(mai_mai_n832_), .C(mai_mai_n823_), .D(mai_mai_n697_), .Y(mai_mai_n1080_));
  OAI220     m1052(.A0(mai_mai_n1080_), .A1(mai_mai_n673_), .B0(mai_mai_n1079_), .B1(mai_mai_n576_), .Y(mai_mai_n1081_));
  NOi31      m1053(.An(i), .B(k), .C(j), .Y(mai_mai_n1082_));
  NA4        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1054_), .C(mai_mai_n337_), .D(mai_mai_n328_), .Y(mai_mai_n1083_));
  INV        m1055(.A(mai_mai_n1083_), .Y(mai_mai_n1084_));
  NOi31      m1056(.An(m), .B(n), .C(f), .Y(mai_mai_n1085_));
  NA2        m1057(.A(mai_mai_n1085_), .B(mai_mai_n50_), .Y(mai_mai_n1086_));
  AN2        m1058(.A(e), .B(c), .Y(mai_mai_n1087_));
  NO2        m1059(.A(mai_mai_n862_), .B(mai_mai_n412_), .Y(mai_mai_n1088_));
  NA2        m1060(.A(mai_mai_n494_), .B(l), .Y(mai_mai_n1089_));
  NOi31      m1061(.An(mai_mai_n841_), .B(mai_mai_n1004_), .C(mai_mai_n1089_), .Y(mai_mai_n1090_));
  NO3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1088_), .C(mai_mai_n1084_), .Y(mai_mai_n1091_));
  NO2        m1063(.A(mai_mai_n281_), .B(a), .Y(mai_mai_n1092_));
  INV        m1064(.A(mai_mai_n1011_), .Y(mai_mai_n1093_));
  NO2        m1065(.A(mai_mai_n1063_), .B(mai_mai_n474_), .Y(mai_mai_n1094_));
  NO2        m1066(.A(mai_mai_n85_), .B(g), .Y(mai_mai_n1095_));
  AOI210     m1067(.A0(mai_mai_n1095_), .A1(mai_mai_n1094_), .B0(mai_mai_n1046_), .Y(mai_mai_n1096_));
  OR2        m1068(.A(mai_mai_n1096_), .B(mai_mai_n1044_), .Y(mai_mai_n1097_));
  NA3        m1069(.A(mai_mai_n1097_), .B(mai_mai_n1093_), .C(mai_mai_n1091_), .Y(mai_mai_n1098_));
  NO4        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1081_), .C(mai_mai_n801_), .D(mai_mai_n553_), .Y(mai_mai_n1099_));
  NA2        m1071(.A(c), .B(b), .Y(mai_mai_n1100_));
  NO2        m1072(.A(mai_mai_n685_), .B(mai_mai_n1100_), .Y(mai_mai_n1101_));
  OAI210     m1073(.A0(mai_mai_n839_), .A1(mai_mai_n815_), .B0(mai_mai_n403_), .Y(mai_mai_n1102_));
  OAI210     m1074(.A0(mai_mai_n1102_), .A1(mai_mai_n840_), .B0(mai_mai_n1101_), .Y(mai_mai_n1103_));
  NAi21      m1075(.An(mai_mai_n409_), .B(mai_mai_n1101_), .Y(mai_mai_n1104_));
  NA3        m1076(.A(mai_mai_n413_), .B(mai_mai_n549_), .C(f), .Y(mai_mai_n1105_));
  NA2        m1077(.A(mai_mai_n538_), .B(mai_mai_n1092_), .Y(mai_mai_n1106_));
  NA3        m1078(.A(mai_mai_n1106_), .B(mai_mai_n1105_), .C(mai_mai_n1104_), .Y(mai_mai_n1107_));
  NAi21      m1079(.An(f), .B(d), .Y(mai_mai_n1108_));
  NO2        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1067_), .Y(mai_mai_n1109_));
  INV        m1081(.A(mai_mai_n1107_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n183_), .B(mai_mai_n238_), .Y(mai_mai_n1111_));
  NA2        m1083(.A(mai_mai_n1111_), .B(m), .Y(mai_mai_n1112_));
  NA3        m1084(.A(mai_mai_n889_), .B(mai_mai_n1089_), .C(mai_mai_n164_), .Y(mai_mai_n1113_));
  NA2        m1085(.A(mai_mai_n1113_), .B(mai_mai_n460_), .Y(mai_mai_n1114_));
  NO2        m1086(.A(mai_mai_n1114_), .B(mai_mai_n1112_), .Y(mai_mai_n1115_));
  NA2        m1087(.A(mai_mai_n158_), .B(mai_mai_n33_), .Y(mai_mai_n1116_));
  AOI210     m1088(.A0(mai_mai_n935_), .A1(mai_mai_n1116_), .B0(mai_mai_n215_), .Y(mai_mai_n1117_));
  OAI210     m1089(.A0(mai_mai_n1117_), .A1(mai_mai_n433_), .B0(mai_mai_n1109_), .Y(mai_mai_n1118_));
  NO2        m1090(.A(mai_mai_n362_), .B(mai_mai_n361_), .Y(mai_mai_n1119_));
  INV        m1091(.A(mai_mai_n929_), .Y(mai_mai_n1120_));
  NAi31      m1092(.An(mai_mai_n1119_), .B(mai_mai_n1120_), .C(mai_mai_n1118_), .Y(mai_mai_n1121_));
  NO2        m1093(.A(mai_mai_n1121_), .B(mai_mai_n1115_), .Y(mai_mai_n1122_));
  NA4        m1094(.A(mai_mai_n1122_), .B(mai_mai_n1110_), .C(mai_mai_n1103_), .D(mai_mai_n1099_), .Y(mai00));
  AOI210     m1095(.A0(mai_mai_n293_), .A1(mai_mai_n215_), .B0(mai_mai_n274_), .Y(mai_mai_n1124_));
  NO2        m1096(.A(mai_mai_n1124_), .B(mai_mai_n566_), .Y(mai_mai_n1125_));
  AOI210     m1097(.A0(mai_mai_n874_), .A1(mai_mai_n914_), .B0(mai_mai_n1084_), .Y(mai_mai_n1126_));
  NO3        m1098(.A(mai_mai_n1060_), .B(mai_mai_n929_), .C(mai_mai_n694_), .Y(mai_mai_n1127_));
  NA3        m1099(.A(mai_mai_n1127_), .B(mai_mai_n1126_), .C(mai_mai_n970_), .Y(mai_mai_n1128_));
  NA2        m1100(.A(mai_mai_n496_), .B(f), .Y(mai_mai_n1129_));
  INV        m1101(.A(mai_mai_n629_), .Y(mai_mai_n1130_));
  NA3        m1102(.A(mai_mai_n1130_), .B(mai_mai_n256_), .C(n), .Y(mai_mai_n1131_));
  AOI210     m1103(.A0(mai_mai_n1131_), .A1(mai_mai_n1129_), .B0(mai_mai_n1015_), .Y(mai_mai_n1132_));
  NO4        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1128_), .C(mai_mai_n1125_), .D(mai_mai_n1038_), .Y(mai_mai_n1133_));
  NA3        m1105(.A(mai_mai_n167_), .B(mai_mai_n45_), .C(mai_mai_n44_), .Y(mai_mai_n1134_));
  NA3        m1106(.A(d), .B(mai_mai_n55_), .C(b), .Y(mai_mai_n1135_));
  NOi31      m1107(.An(n), .B(m), .C(i), .Y(mai_mai_n1136_));
  NA3        m1108(.A(mai_mai_n1136_), .B(mai_mai_n632_), .C(mai_mai_n50_), .Y(mai_mai_n1137_));
  OAI210     m1109(.A0(mai_mai_n1135_), .A1(mai_mai_n1134_), .B0(mai_mai_n1137_), .Y(mai_mai_n1138_));
  INV        m1110(.A(mai_mai_n565_), .Y(mai_mai_n1139_));
  NO3        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1138_), .C(mai_mai_n892_), .Y(mai_mai_n1140_));
  NA3        m1112(.A(mai_mai_n372_), .B(mai_mai_n222_), .C(g), .Y(mai_mai_n1141_));
  OR2        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1135_), .Y(mai_mai_n1142_));
  NO2        m1114(.A(h), .B(g), .Y(mai_mai_n1143_));
  NA4        m1115(.A(mai_mai_n486_), .B(mai_mai_n456_), .C(mai_mai_n1143_), .D(mai_mai_n1003_), .Y(mai_mai_n1144_));
  OAI220     m1116(.A0(mai_mai_n515_), .A1(mai_mai_n582_), .B0(mai_mai_n89_), .B1(mai_mai_n88_), .Y(mai_mai_n1145_));
  AOI220     m1117(.A0(mai_mai_n1145_), .A1(mai_mai_n524_), .B0(mai_mai_n917_), .B1(mai_mai_n564_), .Y(mai_mai_n1146_));
  NA3        m1118(.A(mai_mai_n1146_), .B(mai_mai_n1144_), .C(mai_mai_n1142_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n1147_), .B(mai_mai_n265_), .Y(mai_mai_n1148_));
  INV        m1120(.A(mai_mai_n315_), .Y(mai_mai_n1149_));
  INV        m1121(.A(mai_mai_n567_), .Y(mai_mai_n1150_));
  NA2        m1122(.A(mai_mai_n1150_), .B(mai_mai_n1149_), .Y(mai_mai_n1151_));
  NA3        m1123(.A(mai_mai_n180_), .B(mai_mai_n111_), .C(g), .Y(mai_mai_n1152_));
  NA3        m1124(.A(mai_mai_n456_), .B(mai_mai_n39_), .C(f), .Y(mai_mai_n1153_));
  NOi31      m1125(.An(mai_mai_n848_), .B(mai_mai_n1153_), .C(mai_mai_n1152_), .Y(mai_mai_n1154_));
  NO2        m1126(.A(mai_mai_n273_), .B(mai_mai_n71_), .Y(mai_mai_n1155_));
  NO3        m1127(.A(mai_mai_n412_), .B(mai_mai_n811_), .C(n), .Y(mai_mai_n1156_));
  AOI210     m1128(.A0(mai_mai_n1156_), .A1(mai_mai_n1155_), .B0(mai_mai_n1053_), .Y(mai_mai_n1157_));
  NAi31      m1129(.An(mai_mai_n1018_), .B(mai_mai_n1157_), .C(mai_mai_n70_), .Y(mai_mai_n1158_));
  NO4        m1130(.A(mai_mai_n1158_), .B(mai_mai_n1154_), .C(mai_mai_n1151_), .D(mai_mai_n506_), .Y(mai_mai_n1159_));
  AN3        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1148_), .C(mai_mai_n1140_), .Y(mai_mai_n1160_));
  NA2        m1132(.A(mai_mai_n524_), .B(mai_mai_n99_), .Y(mai_mai_n1161_));
  NA3        m1133(.A(mai_mai_n1085_), .B(mai_mai_n589_), .C(mai_mai_n455_), .Y(mai_mai_n1162_));
  NA3        m1134(.A(mai_mai_n1162_), .B(mai_mai_n1161_), .C(mai_mai_n243_), .Y(mai_mai_n1163_));
  NA2        m1135(.A(mai_mai_n1078_), .B(mai_mai_n524_), .Y(mai_mai_n1164_));
  NA4        m1136(.A(mai_mai_n632_), .B(mai_mai_n208_), .C(mai_mai_n222_), .D(mai_mai_n161_), .Y(mai_mai_n1165_));
  NA3        m1137(.A(mai_mai_n1165_), .B(mai_mai_n1164_), .C(mai_mai_n290_), .Y(mai_mai_n1166_));
  OAI210     m1138(.A0(mai_mai_n454_), .A1(mai_mai_n119_), .B0(mai_mai_n842_), .Y(mai_mai_n1167_));
  NA2        m1139(.A(mai_mai_n1167_), .B(mai_mai_n1113_), .Y(mai_mai_n1168_));
  OR4        m1140(.A(mai_mai_n1015_), .B(mai_mai_n271_), .C(mai_mai_n224_), .D(e), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n218_), .B(mai_mai_n215_), .Y(mai_mai_n1170_));
  NA2        m1142(.A(n), .B(e), .Y(mai_mai_n1171_));
  NO2        m1143(.A(mai_mai_n1171_), .B(mai_mai_n146_), .Y(mai_mai_n1172_));
  AOI220     m1144(.A0(mai_mai_n1172_), .A1(mai_mai_n272_), .B0(mai_mai_n826_), .B1(mai_mai_n1170_), .Y(mai_mai_n1173_));
  NA3        m1145(.A(mai_mai_n1173_), .B(mai_mai_n1169_), .C(mai_mai_n1168_), .Y(mai_mai_n1174_));
  NA2        m1146(.A(mai_mai_n1172_), .B(mai_mai_n829_), .Y(mai_mai_n1175_));
  AOI220     m1147(.A0(mai_mai_n925_), .A1(mai_mai_n564_), .B0(mai_mai_n632_), .B1(mai_mai_n246_), .Y(mai_mai_n1176_));
  NO2        m1148(.A(mai_mai_n64_), .B(h), .Y(mai_mai_n1177_));
  NO3        m1149(.A(mai_mai_n1015_), .B(mai_mai_n1013_), .C(mai_mai_n709_), .Y(mai_mai_n1178_));
  NO2        m1150(.A(mai_mai_n1050_), .B(mai_mai_n132_), .Y(mai_mai_n1179_));
  AN2        m1151(.A(mai_mai_n1179_), .B(mai_mai_n1065_), .Y(mai_mai_n1180_));
  OAI210     m1152(.A0(mai_mai_n1180_), .A1(mai_mai_n1178_), .B0(mai_mai_n1177_), .Y(mai_mai_n1181_));
  NA4        m1153(.A(mai_mai_n1181_), .B(mai_mai_n1176_), .C(mai_mai_n1175_), .D(mai_mai_n843_), .Y(mai_mai_n1182_));
  NO4        m1154(.A(mai_mai_n1182_), .B(mai_mai_n1174_), .C(mai_mai_n1166_), .D(mai_mai_n1163_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n816_), .B(mai_mai_n739_), .Y(mai_mai_n1184_));
  NA4        m1156(.A(mai_mai_n1184_), .B(mai_mai_n1183_), .C(mai_mai_n1160_), .D(mai_mai_n1133_), .Y(mai01));
  AN2        m1157(.A(mai_mai_n992_), .B(mai_mai_n990_), .Y(mai_mai_n1186_));
  NO4        m1158(.A(mai_mai_n786_), .B(mai_mai_n779_), .C(mai_mai_n468_), .D(mai_mai_n279_), .Y(mai_mai_n1187_));
  NA2        m1159(.A(mai_mai_n383_), .B(i), .Y(mai_mai_n1188_));
  NA3        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1187_), .C(mai_mai_n1186_), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n544_), .B(mai_mai_n270_), .Y(mai_mai_n1190_));
  NA2        m1162(.A(mai_mai_n932_), .B(mai_mai_n1190_), .Y(mai_mai_n1191_));
  NA3        m1163(.A(mai_mai_n1191_), .B(mai_mai_n887_), .C(mai_mai_n327_), .Y(mai_mai_n1192_));
  INV        m1164(.A(mai_mai_n117_), .Y(mai_mai_n1193_));
  OR2        m1165(.A(mai_mai_n1193_), .B(mai_mai_n574_), .Y(mai_mai_n1194_));
  NA3        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1165_), .C(mai_mai_n873_), .Y(mai_mai_n1195_));
  NO3        m1167(.A(mai_mai_n766_), .B(mai_mai_n657_), .C(mai_mai_n499_), .Y(mai_mai_n1196_));
  NA3        m1168(.A(mai_mai_n692_), .B(mai_mai_n94_), .C(mai_mai_n44_), .Y(mai_mai_n1197_));
  OA220      m1169(.A0(mai_mai_n1197_), .A1(mai_mai_n651_), .B0(mai_mai_n197_), .B1(mai_mai_n195_), .Y(mai_mai_n1198_));
  NA3        m1170(.A(mai_mai_n1198_), .B(mai_mai_n1196_), .C(mai_mai_n137_), .Y(mai_mai_n1199_));
  NO4        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1195_), .C(mai_mai_n1192_), .D(mai_mai_n1189_), .Y(mai_mai_n1200_));
  NA2        m1172(.A(mai_mai_n296_), .B(mai_mai_n519_), .Y(mai_mai_n1201_));
  NA2        m1173(.A(mai_mai_n527_), .B(mai_mai_n385_), .Y(mai_mai_n1202_));
  NOi21      m1174(.An(mai_mai_n550_), .B(mai_mai_n571_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n1203_), .B(mai_mai_n1202_), .Y(mai_mai_n1204_));
  AOI210     m1176(.A0(mai_mai_n206_), .A1(mai_mai_n87_), .B0(mai_mai_n214_), .Y(mai_mai_n1205_));
  OAI210     m1177(.A0(mai_mai_n793_), .A1(mai_mai_n413_), .B0(mai_mai_n1205_), .Y(mai_mai_n1206_));
  AN3        m1178(.A(m), .B(l), .C(k), .Y(mai_mai_n1207_));
  OAI210     m1179(.A0(mai_mai_n350_), .A1(mai_mai_n34_), .B0(mai_mai_n1207_), .Y(mai_mai_n1208_));
  OR2        m1180(.A(mai_mai_n1208_), .B(mai_mai_n326_), .Y(mai_mai_n1209_));
  NA4        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1206_), .C(mai_mai_n1204_), .D(mai_mai_n1201_), .Y(mai_mai_n1210_));
  INV        m1182(.A(mai_mai_n583_), .Y(mai_mai_n1211_));
  OAI210     m1183(.A0(mai_mai_n1193_), .A1(mai_mai_n580_), .B0(mai_mai_n1211_), .Y(mai_mai_n1212_));
  NA2        m1184(.A(mai_mai_n278_), .B(mai_mai_n197_), .Y(mai_mai_n1213_));
  NA2        m1185(.A(mai_mai_n1213_), .B(mai_mai_n648_), .Y(mai_mai_n1214_));
  INV        m1186(.A(mai_mai_n929_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n320_), .B(mai_mai_n658_), .Y(mai_mai_n1216_));
  NA4        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1215_), .C(mai_mai_n1214_), .D(mai_mai_n769_), .Y(mai_mai_n1217_));
  NO3        m1189(.A(mai_mai_n1217_), .B(mai_mai_n1212_), .C(mai_mai_n1210_), .Y(mai_mai_n1218_));
  NA2        m1190(.A(mai_mai_n492_), .B(mai_mai_n57_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n1197_), .B(mai_mai_n950_), .Y(mai_mai_n1220_));
  NO2        m1192(.A(mai_mai_n209_), .B(mai_mai_n110_), .Y(mai_mai_n1221_));
  NO3        m1193(.A(mai_mai_n1221_), .B(mai_mai_n1220_), .C(mai_mai_n1138_), .Y(mai_mai_n1222_));
  NA3        m1194(.A(mai_mai_n1222_), .B(mai_mai_n1219_), .C(mai_mai_n738_), .Y(mai_mai_n1223_));
  NO2        m1195(.A(mai_mai_n939_), .B(mai_mai_n234_), .Y(mai_mai_n1224_));
  NO2        m1196(.A(mai_mai_n940_), .B(mai_mai_n546_), .Y(mai_mai_n1225_));
  OAI210     m1197(.A0(mai_mai_n1225_), .A1(mai_mai_n1224_), .B0(mai_mai_n335_), .Y(mai_mai_n1226_));
  INV        m1198(.A(mai_mai_n653_), .Y(mai_mai_n1227_));
  OR2        m1199(.A(mai_mai_n1141_), .B(mai_mai_n1135_), .Y(mai_mai_n1228_));
  NA2        m1200(.A(mai_mai_n1228_), .B(mai_mai_n375_), .Y(mai_mai_n1229_));
  NOi41      m1201(.An(mai_mai_n1226_), .B(mai_mai_n1229_), .C(mai_mai_n1227_), .D(mai_mai_n1223_), .Y(mai_mai_n1230_));
  NO2        m1202(.A(mai_mai_n131_), .B(mai_mai_n44_), .Y(mai_mai_n1231_));
  NO2        m1203(.A(mai_mai_n44_), .B(mai_mai_n39_), .Y(mai_mai_n1232_));
  AO220      m1204(.A0(mai_mai_n1232_), .A1(mai_mai_n605_), .B0(mai_mai_n1231_), .B1(mai_mai_n690_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n1233_), .B(mai_mai_n335_), .Y(mai_mai_n1234_));
  NO3        m1206(.A(mai_mai_n1063_), .B(mai_mai_n177_), .C(mai_mai_n85_), .Y(mai_mai_n1235_));
  INV        m1207(.A(mai_mai_n1234_), .Y(mai_mai_n1236_));
  NO2        m1208(.A(mai_mai_n597_), .B(mai_mai_n596_), .Y(mai_mai_n1237_));
  NO4        m1209(.A(mai_mai_n1063_), .B(mai_mai_n1237_), .C(mai_mai_n175_), .D(mai_mai_n85_), .Y(mai_mai_n1238_));
  NO3        m1210(.A(mai_mai_n1238_), .B(mai_mai_n1236_), .C(mai_mai_n621_), .Y(mai_mai_n1239_));
  NA4        m1211(.A(mai_mai_n1239_), .B(mai_mai_n1230_), .C(mai_mai_n1218_), .D(mai_mai_n1200_), .Y(mai06));
  NO2        m1212(.A(mai_mai_n226_), .B(mai_mai_n101_), .Y(mai_mai_n1241_));
  OAI210     m1213(.A0(mai_mai_n1241_), .A1(mai_mai_n1235_), .B0(mai_mai_n371_), .Y(mai_mai_n1242_));
  NO3        m1214(.A(mai_mai_n584_), .B(mai_mai_n791_), .C(mai_mai_n585_), .Y(mai_mai_n1243_));
  OR2        m1215(.A(mai_mai_n1243_), .B(mai_mai_n862_), .Y(mai_mai_n1244_));
  NA3        m1216(.A(mai_mai_n1244_), .B(mai_mai_n1242_), .C(mai_mai_n1226_), .Y(mai_mai_n1245_));
  NO3        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1227_), .C(mai_mai_n255_), .Y(mai_mai_n1246_));
  NO2        m1218(.A(mai_mai_n294_), .B(mai_mai_n44_), .Y(mai_mai_n1247_));
  AOI210     m1219(.A0(mai_mai_n1247_), .A1(mai_mai_n543_), .B0(mai_mai_n1224_), .Y(mai_mai_n1248_));
  AOI210     m1220(.A0(mai_mai_n1247_), .A1(mai_mai_n547_), .B0(mai_mai_n1233_), .Y(mai_mai_n1249_));
  AOI210     m1221(.A0(mai_mai_n1249_), .A1(mai_mai_n1248_), .B0(mai_mai_n332_), .Y(mai_mai_n1250_));
  OAI210     m1222(.A0(mai_mai_n87_), .A1(mai_mai_n39_), .B0(mai_mai_n656_), .Y(mai_mai_n1251_));
  NA2        m1223(.A(mai_mai_n1251_), .B(mai_mai_n625_), .Y(mai_mai_n1252_));
  NO2        m1224(.A(mai_mai_n502_), .B(mai_mai_n172_), .Y(mai_mai_n1253_));
  NO2        m1225(.A(mai_mai_n590_), .B(mai_mai_n1086_), .Y(mai_mai_n1254_));
  OAI210     m1226(.A0(mai_mai_n449_), .A1(mai_mai_n248_), .B0(mai_mai_n881_), .Y(mai_mai_n1255_));
  NO3        m1227(.A(mai_mai_n1255_), .B(mai_mai_n1254_), .C(mai_mai_n1253_), .Y(mai_mai_n1256_));
  INV        m1228(.A(mai_mai_n583_), .Y(mai_mai_n1257_));
  NA3        m1229(.A(mai_mai_n1257_), .B(mai_mai_n1256_), .C(mai_mai_n1252_), .Y(mai_mai_n1258_));
  NO2        m1230(.A(mai_mai_n731_), .B(mai_mai_n359_), .Y(mai_mai_n1259_));
  NO3        m1231(.A(mai_mai_n658_), .B(mai_mai_n740_), .C(mai_mai_n617_), .Y(mai_mai_n1260_));
  NOi21      m1232(.An(mai_mai_n1259_), .B(mai_mai_n1260_), .Y(mai_mai_n1261_));
  AN2        m1233(.A(mai_mai_n925_), .B(mai_mai_n628_), .Y(mai_mai_n1262_));
  NO4        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1261_), .C(mai_mai_n1258_), .D(mai_mai_n1250_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n785_), .B(mai_mai_n275_), .Y(mai_mai_n1264_));
  OAI220     m1236(.A0(mai_mai_n715_), .A1(mai_mai_n46_), .B0(mai_mai_n226_), .B1(mai_mai_n599_), .Y(mai_mai_n1265_));
  OAI210     m1237(.A0(mai_mai_n275_), .A1(c), .B0(mai_mai_n624_), .Y(mai_mai_n1266_));
  AOI220     m1238(.A0(mai_mai_n1266_), .A1(mai_mai_n1265_), .B0(mai_mai_n1264_), .B1(mai_mai_n266_), .Y(mai_mai_n1267_));
  OAI220     m1239(.A0(mai_mai_n682_), .A1(mai_mai_n248_), .B0(mai_mai_n498_), .B1(mai_mai_n502_), .Y(mai_mai_n1268_));
  OAI210     m1240(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1269_));
  NO3        m1241(.A(mai_mai_n1269_), .B(mai_mai_n582_), .C(j), .Y(mai_mai_n1270_));
  NOi21      m1242(.An(mai_mai_n1270_), .B(mai_mai_n651_), .Y(mai_mai_n1271_));
  NO3        m1243(.A(mai_mai_n1271_), .B(mai_mai_n1268_), .C(mai_mai_n1088_), .Y(mai_mai_n1272_));
  NA3        m1244(.A(mai_mai_n777_), .B(mai_mai_n776_), .C(mai_mai_n423_), .Y(mai_mai_n1273_));
  NAi31      m1245(.An(mai_mai_n731_), .B(mai_mai_n1273_), .C(mai_mai_n205_), .Y(mai_mai_n1274_));
  NA4        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1272_), .C(mai_mai_n1267_), .D(mai_mai_n1176_), .Y(mai_mai_n1275_));
  NOi31      m1247(.An(mai_mai_n1243_), .B(mai_mai_n453_), .C(mai_mai_n384_), .Y(mai_mai_n1276_));
  OR3        m1248(.A(mai_mai_n1276_), .B(mai_mai_n765_), .C(mai_mai_n530_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n559_), .B(mai_mai_n435_), .Y(mai_mai_n1278_));
  NA2        m1250(.A(mai_mai_n1270_), .B(mai_mai_n773_), .Y(mai_mai_n1279_));
  NA3        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1278_), .C(mai_mai_n1277_), .Y(mai_mai_n1280_));
  NA2        m1252(.A(mai_mai_n1259_), .B(mai_mai_n739_), .Y(mai_mai_n1281_));
  AN2        m1253(.A(mai_mai_n900_), .B(mai_mai_n899_), .Y(mai_mai_n1282_));
  NO4        m1254(.A(mai_mai_n1282_), .B(mai_mai_n852_), .C(mai_mai_n488_), .D(mai_mai_n471_), .Y(mai_mai_n1283_));
  NA2        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1281_), .Y(mai_mai_n1284_));
  NAi21      m1256(.An(j), .B(i), .Y(mai_mai_n1285_));
  NO4        m1257(.A(mai_mai_n1237_), .B(mai_mai_n1285_), .C(mai_mai_n429_), .D(mai_mai_n236_), .Y(mai_mai_n1286_));
  NO4        m1258(.A(mai_mai_n1286_), .B(mai_mai_n1284_), .C(mai_mai_n1280_), .D(mai_mai_n1275_), .Y(mai_mai_n1287_));
  NA4        m1259(.A(mai_mai_n1287_), .B(mai_mai_n1263_), .C(mai_mai_n1246_), .D(mai_mai_n1239_), .Y(mai07));
  NOi21      m1260(.An(j), .B(k), .Y(mai_mai_n1289_));
  NA4        m1261(.A(mai_mai_n180_), .B(mai_mai_n107_), .C(mai_mai_n1289_), .D(f), .Y(mai_mai_n1290_));
  NAi32      m1262(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1291_));
  NO3        m1263(.A(mai_mai_n1291_), .B(g), .C(f), .Y(mai_mai_n1292_));
  OAI210     m1264(.A0(mai_mai_n314_), .A1(mai_mai_n473_), .B0(mai_mai_n1292_), .Y(mai_mai_n1293_));
  NAi21      m1265(.An(f), .B(c), .Y(mai_mai_n1294_));
  OR2        m1266(.A(e), .B(d), .Y(mai_mai_n1295_));
  OAI220     m1267(.A0(mai_mai_n1295_), .A1(mai_mai_n1294_), .B0(mai_mai_n611_), .B1(mai_mai_n316_), .Y(mai_mai_n1296_));
  NA3        m1268(.A(mai_mai_n1296_), .B(mai_mai_n1027_), .C(mai_mai_n180_), .Y(mai_mai_n1297_));
  NOi31      m1269(.An(n), .B(m), .C(b), .Y(mai_mai_n1298_));
  NO3        m1270(.A(mai_mai_n132_), .B(mai_mai_n437_), .C(h), .Y(mai_mai_n1299_));
  NA3        m1271(.A(mai_mai_n1297_), .B(mai_mai_n1293_), .C(mai_mai_n1290_), .Y(mai_mai_n1300_));
  NOi41      m1272(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1301_));
  NOi21      m1273(.An(h), .B(k), .Y(mai_mai_n1302_));
  NO2        m1274(.A(k), .B(i), .Y(mai_mai_n1303_));
  NA3        m1275(.A(mai_mai_n1303_), .B(mai_mai_n872_), .C(mai_mai_n180_), .Y(mai_mai_n1304_));
  NA2        m1276(.A(mai_mai_n85_), .B(mai_mai_n44_), .Y(mai_mai_n1305_));
  NO2        m1277(.A(mai_mai_n1021_), .B(mai_mai_n429_), .Y(mai_mai_n1306_));
  NA3        m1278(.A(mai_mai_n1306_), .B(mai_mai_n1305_), .C(mai_mai_n215_), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n1035_), .B(mai_mai_n302_), .Y(mai_mai_n1308_));
  NA2        m1280(.A(mai_mai_n531_), .B(mai_mai_n78_), .Y(mai_mai_n1309_));
  NA2        m1281(.A(mai_mai_n1177_), .B(mai_mai_n284_), .Y(mai_mai_n1310_));
  NA4        m1282(.A(mai_mai_n1310_), .B(mai_mai_n1309_), .C(mai_mai_n1307_), .D(mai_mai_n1304_), .Y(mai_mai_n1311_));
  NO2        m1283(.A(mai_mai_n1311_), .B(mai_mai_n1300_), .Y(mai_mai_n1312_));
  NO3        m1284(.A(e), .B(d), .C(c), .Y(mai_mai_n1313_));
  OAI210     m1285(.A0(mai_mai_n132_), .A1(mai_mai_n215_), .B0(mai_mai_n588_), .Y(mai_mai_n1314_));
  NA2        m1286(.A(mai_mai_n1314_), .B(mai_mai_n1313_), .Y(mai_mai_n1315_));
  NO2        m1287(.A(mai_mai_n1315_), .B(c), .Y(mai_mai_n1316_));
  OR2        m1288(.A(h), .B(f), .Y(mai_mai_n1317_));
  NO3        m1289(.A(n), .B(m), .C(i), .Y(mai_mai_n1318_));
  OAI210     m1290(.A0(mai_mai_n1087_), .A1(mai_mai_n156_), .B0(mai_mai_n1318_), .Y(mai_mai_n1319_));
  NO2        m1291(.A(mai_mai_n1319_), .B(mai_mai_n1317_), .Y(mai_mai_n1320_));
  NA3        m1292(.A(mai_mai_n679_), .B(mai_mai_n666_), .C(mai_mai_n111_), .Y(mai_mai_n1321_));
  NO2        m1293(.A(mai_mai_n1321_), .B(mai_mai_n44_), .Y(mai_mai_n1322_));
  NA2        m1294(.A(mai_mai_n1318_), .B(mai_mai_n623_), .Y(mai_mai_n1323_));
  NO2        m1295(.A(l), .B(k), .Y(mai_mai_n1324_));
  NOi41      m1296(.An(mai_mai_n536_), .B(mai_mai_n1324_), .C(mai_mai_n466_), .D(mai_mai_n429_), .Y(mai_mai_n1325_));
  NO3        m1297(.A(mai_mai_n429_), .B(d), .C(c), .Y(mai_mai_n1326_));
  NO4        m1298(.A(mai_mai_n1325_), .B(mai_mai_n1322_), .C(mai_mai_n1320_), .D(mai_mai_n1316_), .Y(mai_mai_n1327_));
  NO2        m1299(.A(mai_mai_n147_), .B(h), .Y(mai_mai_n1328_));
  NO2        m1300(.A(mai_mai_n1045_), .B(l), .Y(mai_mai_n1329_));
  NO2        m1301(.A(g), .B(c), .Y(mai_mai_n1330_));
  NA3        m1302(.A(mai_mai_n1330_), .B(mai_mai_n142_), .C(mai_mai_n188_), .Y(mai_mai_n1331_));
  NO2        m1303(.A(mai_mai_n1331_), .B(mai_mai_n1329_), .Y(mai_mai_n1332_));
  NA2        m1304(.A(mai_mai_n1332_), .B(mai_mai_n180_), .Y(mai_mai_n1333_));
  NA2        m1305(.A(mai_mai_n1302_), .B(mai_mai_n1045_), .Y(mai_mai_n1334_));
  NO2        m1306(.A(mai_mai_n440_), .B(a), .Y(mai_mai_n1335_));
  NA3        m1307(.A(mai_mai_n1335_), .B(mai_mai_n1334_), .C(mai_mai_n112_), .Y(mai_mai_n1336_));
  NO2        m1308(.A(i), .B(h), .Y(mai_mai_n1337_));
  NA2        m1309(.A(mai_mai_n1108_), .B(h), .Y(mai_mai_n1338_));
  NA2        m1310(.A(mai_mai_n138_), .B(mai_mai_n222_), .Y(mai_mai_n1339_));
  NO2        m1311(.A(mai_mai_n1339_), .B(mai_mai_n1338_), .Y(mai_mai_n1340_));
  NO2        m1312(.A(mai_mai_n737_), .B(mai_mai_n189_), .Y(mai_mai_n1341_));
  NOi31      m1313(.An(m), .B(n), .C(b), .Y(mai_mai_n1342_));
  NOi31      m1314(.An(f), .B(d), .C(c), .Y(mai_mai_n1343_));
  NA2        m1315(.A(mai_mai_n1343_), .B(mai_mai_n1342_), .Y(mai_mai_n1344_));
  INV        m1316(.A(mai_mai_n1344_), .Y(mai_mai_n1345_));
  NO3        m1317(.A(mai_mai_n1345_), .B(mai_mai_n1341_), .C(mai_mai_n1340_), .Y(mai_mai_n1346_));
  NA2        m1318(.A(mai_mai_n1056_), .B(mai_mai_n456_), .Y(mai_mai_n1347_));
  NO4        m1319(.A(mai_mai_n1347_), .B(mai_mai_n1030_), .C(mai_mai_n429_), .D(mai_mai_n44_), .Y(mai_mai_n1348_));
  OAI210     m1320(.A0(mai_mai_n183_), .A1(mai_mai_n514_), .B0(mai_mai_n1031_), .Y(mai_mai_n1349_));
  NO3        m1321(.A(mai_mai_n40_), .B(i), .C(h), .Y(mai_mai_n1350_));
  INV        m1322(.A(mai_mai_n1349_), .Y(mai_mai_n1351_));
  NO2        m1323(.A(mai_mai_n1351_), .B(mai_mai_n1348_), .Y(mai_mai_n1352_));
  AN4        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1346_), .C(mai_mai_n1336_), .D(mai_mai_n1333_), .Y(mai_mai_n1353_));
  NA2        m1325(.A(mai_mai_n1298_), .B(mai_mai_n368_), .Y(mai_mai_n1354_));
  NO2        m1326(.A(mai_mai_n1354_), .B(mai_mai_n1012_), .Y(mai_mai_n1355_));
  NA2        m1327(.A(mai_mai_n1326_), .B(mai_mai_n216_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n189_), .B(b), .Y(mai_mai_n1357_));
  AOI220     m1329(.A0(mai_mai_n1136_), .A1(mai_mai_n1357_), .B0(mai_mai_n1064_), .B1(mai_mai_n1347_), .Y(mai_mai_n1358_));
  NAi31      m1330(.An(mai_mai_n1355_), .B(mai_mai_n1358_), .C(mai_mai_n1356_), .Y(mai_mai_n1359_));
  NO4        m1331(.A(mai_mai_n132_), .B(g), .C(f), .D(e), .Y(mai_mai_n1360_));
  NA3        m1332(.A(mai_mai_n1303_), .B(mai_mai_n285_), .C(h), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n196_), .B(mai_mai_n96_), .Y(mai_mai_n1362_));
  OR2        m1334(.A(e), .B(a), .Y(mai_mai_n1363_));
  NO2        m1335(.A(mai_mai_n1295_), .B(mai_mai_n1294_), .Y(mai_mai_n1364_));
  AOI210     m1336(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1364_), .Y(mai_mai_n1365_));
  NO2        m1337(.A(mai_mai_n1365_), .B(mai_mai_n1052_), .Y(mai_mai_n1366_));
  NA2        m1338(.A(mai_mai_n1301_), .B(mai_mai_n1324_), .Y(mai_mai_n1367_));
  INV        m1339(.A(mai_mai_n1367_), .Y(mai_mai_n1368_));
  OR3        m1340(.A(mai_mai_n530_), .B(mai_mai_n529_), .C(mai_mai_n111_), .Y(mai_mai_n1369_));
  NA2        m1341(.A(mai_mai_n1085_), .B(mai_mai_n397_), .Y(mai_mai_n1370_));
  NO2        m1342(.A(mai_mai_n1370_), .B(mai_mai_n422_), .Y(mai_mai_n1371_));
  AO210      m1343(.A0(mai_mai_n1371_), .A1(mai_mai_n115_), .B0(mai_mai_n1368_), .Y(mai_mai_n1372_));
  NO3        m1344(.A(mai_mai_n1372_), .B(mai_mai_n1366_), .C(mai_mai_n1359_), .Y(mai_mai_n1373_));
  NA4        m1345(.A(mai_mai_n1373_), .B(mai_mai_n1353_), .C(mai_mai_n1327_), .D(mai_mai_n1312_), .Y(mai_mai_n1374_));
  NO2        m1346(.A(mai_mai_n1100_), .B(mai_mai_n109_), .Y(mai_mai_n1375_));
  NA2        m1347(.A(mai_mai_n368_), .B(mai_mai_n55_), .Y(mai_mai_n1376_));
  AOI210     m1348(.A0(mai_mai_n1376_), .A1(mai_mai_n1021_), .B0(mai_mai_n1323_), .Y(mai_mai_n1377_));
  NA2        m1349(.A(mai_mai_n216_), .B(mai_mai_n180_), .Y(mai_mai_n1378_));
  AOI210     m1350(.A0(mai_mai_n1378_), .A1(mai_mai_n1152_), .B0(mai_mai_n1376_), .Y(mai_mai_n1379_));
  NO2        m1351(.A(mai_mai_n1057_), .B(mai_mai_n1052_), .Y(mai_mai_n1380_));
  NO3        m1352(.A(mai_mai_n1380_), .B(mai_mai_n1379_), .C(mai_mai_n1377_), .Y(mai_mai_n1381_));
  NO2        m1353(.A(mai_mai_n380_), .B(j), .Y(mai_mai_n1382_));
  NA3        m1354(.A(mai_mai_n1350_), .B(mai_mai_n1295_), .C(mai_mai_n1085_), .Y(mai_mai_n1383_));
  NAi41      m1355(.An(mai_mai_n1337_), .B(mai_mai_n1043_), .C(mai_mai_n168_), .D(mai_mai_n150_), .Y(mai_mai_n1384_));
  NA2        m1356(.A(mai_mai_n1384_), .B(mai_mai_n1383_), .Y(mai_mai_n1385_));
  NA3        m1357(.A(g), .B(mai_mai_n1382_), .C(mai_mai_n158_), .Y(mai_mai_n1386_));
  INV        m1358(.A(mai_mai_n1386_), .Y(mai_mai_n1387_));
  NO3        m1359(.A(mai_mai_n731_), .B(mai_mai_n175_), .C(mai_mai_n400_), .Y(mai_mai_n1388_));
  NO3        m1360(.A(mai_mai_n1388_), .B(mai_mai_n1387_), .C(mai_mai_n1385_), .Y(mai_mai_n1389_));
  AOI210     m1361(.A0(mai_mai_n1378_), .A1(mai_mai_n1362_), .B0(mai_mai_n1021_), .Y(mai_mai_n1390_));
  OR2        m1362(.A(n), .B(i), .Y(mai_mai_n1391_));
  OAI210     m1363(.A0(mai_mai_n1391_), .A1(mai_mai_n1042_), .B0(mai_mai_n48_), .Y(mai_mai_n1392_));
  AOI220     m1364(.A0(mai_mai_n1392_), .A1(mai_mai_n1143_), .B0(mai_mai_n804_), .B1(mai_mai_n196_), .Y(mai_mai_n1393_));
  INV        m1365(.A(mai_mai_n1393_), .Y(mai_mai_n1394_));
  OAI220     m1366(.A0(mai_mai_n649_), .A1(g), .B0(mai_mai_n226_), .B1(c), .Y(mai_mai_n1395_));
  AOI210     m1367(.A0(mai_mai_n1357_), .A1(mai_mai_n40_), .B0(mai_mai_n1395_), .Y(mai_mai_n1396_));
  NO2        m1368(.A(mai_mai_n132_), .B(l), .Y(mai_mai_n1397_));
  NO2        m1369(.A(mai_mai_n226_), .B(k), .Y(mai_mai_n1398_));
  OAI210     m1370(.A0(mai_mai_n1398_), .A1(mai_mai_n1337_), .B0(mai_mai_n1397_), .Y(mai_mai_n1399_));
  OAI220     m1371(.A0(mai_mai_n1399_), .A1(mai_mai_n31_), .B0(mai_mai_n1396_), .B1(mai_mai_n177_), .Y(mai_mai_n1400_));
  NO3        m1372(.A(mai_mai_n1369_), .B(mai_mai_n456_), .C(mai_mai_n349_), .Y(mai_mai_n1401_));
  NO4        m1373(.A(mai_mai_n1401_), .B(mai_mai_n1400_), .C(mai_mai_n1394_), .D(mai_mai_n1390_), .Y(mai_mai_n1402_));
  NO3        m1374(.A(mai_mai_n1067_), .B(mai_mai_n1295_), .C(mai_mai_n48_), .Y(mai_mai_n1403_));
  NO2        m1375(.A(mai_mai_n1052_), .B(h), .Y(mai_mai_n1404_));
  NA3        m1376(.A(mai_mai_n1404_), .B(d), .C(mai_mai_n1013_), .Y(mai_mai_n1405_));
  NO2        m1377(.A(mai_mai_n1405_), .B(c), .Y(mai_mai_n1406_));
  NA3        m1378(.A(mai_mai_n1375_), .B(mai_mai_n456_), .C(f), .Y(mai_mai_n1407_));
  NA2        m1379(.A(mai_mai_n180_), .B(mai_mai_n111_), .Y(mai_mai_n1408_));
  NO2        m1380(.A(mai_mai_n1289_), .B(mai_mai_n41_), .Y(mai_mai_n1409_));
  AOI210     m1381(.A0(mai_mai_n112_), .A1(mai_mai_n39_), .B0(mai_mai_n1409_), .Y(mai_mai_n1410_));
  NO2        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1407_), .Y(mai_mai_n1411_));
  NO2        m1383(.A(mai_mai_n1285_), .B(mai_mai_n175_), .Y(mai_mai_n1412_));
  NOi21      m1384(.An(d), .B(f), .Y(mai_mai_n1413_));
  NO3        m1385(.A(mai_mai_n1343_), .B(mai_mai_n1413_), .C(mai_mai_n39_), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1414_), .B(mai_mai_n1412_), .Y(mai_mai_n1415_));
  NO2        m1387(.A(mai_mai_n1295_), .B(f), .Y(mai_mai_n1416_));
  NA2        m1388(.A(mai_mai_n1335_), .B(mai_mai_n1409_), .Y(mai_mai_n1417_));
  NA2        m1389(.A(mai_mai_n1417_), .B(mai_mai_n1415_), .Y(mai_mai_n1418_));
  NO3        m1390(.A(mai_mai_n1418_), .B(mai_mai_n1411_), .C(mai_mai_n1406_), .Y(mai_mai_n1419_));
  NA4        m1391(.A(mai_mai_n1419_), .B(mai_mai_n1402_), .C(mai_mai_n1389_), .D(mai_mai_n1381_), .Y(mai_mai_n1420_));
  NO3        m1392(.A(mai_mai_n1056_), .B(mai_mai_n1042_), .C(mai_mai_n39_), .Y(mai_mai_n1421_));
  NO2        m1393(.A(mai_mai_n456_), .B(mai_mai_n294_), .Y(mai_mai_n1422_));
  OAI210     m1394(.A0(mai_mai_n1422_), .A1(mai_mai_n1421_), .B0(mai_mai_n1308_), .Y(mai_mai_n1423_));
  OAI210     m1395(.A0(mai_mai_n1360_), .A1(mai_mai_n1298_), .B0(mai_mai_n859_), .Y(mai_mai_n1424_));
  NO2        m1396(.A(mai_mai_n1009_), .B(mai_mai_n132_), .Y(mai_mai_n1425_));
  NA2        m1397(.A(mai_mai_n1425_), .B(mai_mai_n604_), .Y(mai_mai_n1426_));
  NA3        m1398(.A(mai_mai_n1426_), .B(mai_mai_n1424_), .C(mai_mai_n1423_), .Y(mai_mai_n1427_));
  NA2        m1399(.A(mai_mai_n1330_), .B(mai_mai_n1413_), .Y(mai_mai_n1428_));
  NO2        m1400(.A(mai_mai_n1428_), .B(m), .Y(mai_mai_n1429_));
  NO2        m1401(.A(mai_mai_n151_), .B(mai_mai_n182_), .Y(mai_mai_n1430_));
  OAI210     m1402(.A0(mai_mai_n1430_), .A1(mai_mai_n109_), .B0(mai_mai_n1342_), .Y(mai_mai_n1431_));
  INV        m1403(.A(mai_mai_n1431_), .Y(mai_mai_n1432_));
  NO3        m1404(.A(mai_mai_n1432_), .B(mai_mai_n1429_), .C(mai_mai_n1427_), .Y(mai_mai_n1433_));
  NO2        m1405(.A(mai_mai_n1294_), .B(e), .Y(mai_mai_n1434_));
  NA2        m1406(.A(mai_mai_n1434_), .B(mai_mai_n395_), .Y(mai_mai_n1435_));
  OAI210     m1407(.A0(mai_mai_n1416_), .A1(mai_mai_n1095_), .B0(mai_mai_n615_), .Y(mai_mai_n1436_));
  OR3        m1408(.A(mai_mai_n1398_), .B(mai_mai_n1177_), .C(mai_mai_n132_), .Y(mai_mai_n1437_));
  OAI220     m1409(.A0(mai_mai_n1437_), .A1(mai_mai_n1435_), .B0(mai_mai_n1436_), .B1(mai_mai_n431_), .Y(mai_mai_n1438_));
  INV        m1410(.A(mai_mai_n1438_), .Y(mai_mai_n1439_));
  NO2        m1411(.A(mai_mai_n182_), .B(c), .Y(mai_mai_n1440_));
  OAI210     m1412(.A0(mai_mai_n1440_), .A1(mai_mai_n1434_), .B0(mai_mai_n180_), .Y(mai_mai_n1441_));
  AOI220     m1413(.A0(mai_mai_n1441_), .A1(mai_mai_n1044_), .B0(mai_mai_n521_), .B1(mai_mai_n359_), .Y(mai_mai_n1442_));
  NA2        m1414(.A(mai_mai_n529_), .B(g), .Y(mai_mai_n1443_));
  AOI210     m1415(.A0(mai_mai_n1443_), .A1(mai_mai_n1326_), .B0(mai_mai_n1403_), .Y(mai_mai_n1444_));
  NO2        m1416(.A(mai_mai_n1363_), .B(f), .Y(mai_mai_n1445_));
  NA2        m1417(.A(mai_mai_n1095_), .B(a), .Y(mai_mai_n1446_));
  OAI220     m1418(.A0(mai_mai_n1446_), .A1(mai_mai_n65_), .B0(mai_mai_n1444_), .B1(mai_mai_n214_), .Y(mai_mai_n1447_));
  AOI210     m1419(.A0(mai_mai_n876_), .A1(mai_mai_n404_), .B0(mai_mai_n103_), .Y(mai_mai_n1448_));
  OR2        m1420(.A(mai_mai_n1448_), .B(mai_mai_n529_), .Y(mai_mai_n1449_));
  NA2        m1421(.A(mai_mai_n1445_), .B(mai_mai_n1305_), .Y(mai_mai_n1450_));
  OAI220     m1422(.A0(mai_mai_n1450_), .A1(mai_mai_n48_), .B0(mai_mai_n1449_), .B1(mai_mai_n175_), .Y(mai_mai_n1451_));
  NA4        m1423(.A(mai_mai_n1065_), .B(mai_mai_n1062_), .C(mai_mai_n222_), .D(mai_mai_n64_), .Y(mai_mai_n1452_));
  NA2        m1424(.A(mai_mai_n1299_), .B(mai_mai_n183_), .Y(mai_mai_n1453_));
  NO2        m1425(.A(mai_mai_n48_), .B(l), .Y(mai_mai_n1454_));
  OAI210     m1426(.A0(mai_mai_n1363_), .A1(mai_mai_n838_), .B0(mai_mai_n473_), .Y(mai_mai_n1455_));
  OAI210     m1427(.A0(mai_mai_n1455_), .A1(mai_mai_n1068_), .B0(mai_mai_n1454_), .Y(mai_mai_n1456_));
  NO2        m1428(.A(mai_mai_n251_), .B(g), .Y(mai_mai_n1457_));
  NO2        m1429(.A(m), .B(i), .Y(mai_mai_n1458_));
  BUFFER     m1430(.A(mai_mai_n1458_), .Y(mai_mai_n1459_));
  AOI220     m1431(.A0(mai_mai_n1459_), .A1(mai_mai_n1328_), .B0(mai_mai_n1043_), .B1(mai_mai_n1457_), .Y(mai_mai_n1460_));
  NA4        m1432(.A(mai_mai_n1460_), .B(mai_mai_n1456_), .C(mai_mai_n1453_), .D(mai_mai_n1452_), .Y(mai_mai_n1461_));
  NO4        m1433(.A(mai_mai_n1461_), .B(mai_mai_n1451_), .C(mai_mai_n1447_), .D(mai_mai_n1442_), .Y(mai_mai_n1462_));
  NA3        m1434(.A(mai_mai_n1462_), .B(mai_mai_n1439_), .C(mai_mai_n1433_), .Y(mai_mai_n1463_));
  NA3        m1435(.A(mai_mai_n931_), .B(mai_mai_n138_), .C(mai_mai_n45_), .Y(mai_mai_n1464_));
  AOI210     m1436(.A0(mai_mai_n148_), .A1(c), .B0(mai_mai_n1464_), .Y(mai_mai_n1465_));
  INV        m1437(.A(mai_mai_n186_), .Y(mai_mai_n1466_));
  NA2        m1438(.A(mai_mai_n1466_), .B(mai_mai_n1404_), .Y(mai_mai_n1467_));
  OR2        m1439(.A(mai_mai_n133_), .B(mai_mai_n1354_), .Y(mai_mai_n1468_));
  NO2        m1440(.A(mai_mai_n68_), .B(c), .Y(mai_mai_n1469_));
  NA2        m1441(.A(mai_mai_n1412_), .B(mai_mai_n1469_), .Y(mai_mai_n1470_));
  NA3        m1442(.A(mai_mai_n1470_), .B(mai_mai_n1468_), .C(mai_mai_n1467_), .Y(mai_mai_n1471_));
  NO2        m1443(.A(mai_mai_n1471_), .B(mai_mai_n1465_), .Y(mai_mai_n1472_));
  AOI210     m1444(.A0(mai_mai_n156_), .A1(mai_mai_n55_), .B0(mai_mai_n1434_), .Y(mai_mai_n1473_));
  NO2        m1445(.A(mai_mai_n1473_), .B(mai_mai_n1408_), .Y(mai_mai_n1474_));
  NOi21      m1446(.An(mai_mai_n1299_), .B(e), .Y(mai_mai_n1475_));
  NO2        m1447(.A(mai_mai_n1475_), .B(mai_mai_n1474_), .Y(mai_mai_n1476_));
  AN2        m1448(.A(mai_mai_n1065_), .B(mai_mai_n1050_), .Y(mai_mai_n1477_));
  NA2        m1449(.A(mai_mai_n1027_), .B(mai_mai_n159_), .Y(mai_mai_n1478_));
  NOi31      m1450(.An(mai_mai_n30_), .B(mai_mai_n1478_), .C(n), .Y(mai_mai_n1479_));
  AOI210     m1451(.A0(mai_mai_n1477_), .A1(mai_mai_n1136_), .B0(mai_mai_n1479_), .Y(mai_mai_n1480_));
  NO2        m1452(.A(mai_mai_n1407_), .B(mai_mai_n65_), .Y(mai_mai_n1481_));
  NA2        m1453(.A(mai_mai_n58_), .B(a), .Y(mai_mai_n1482_));
  NO2        m1454(.A(mai_mai_n1303_), .B(mai_mai_n117_), .Y(mai_mai_n1483_));
  OAI220     m1455(.A0(mai_mai_n1483_), .A1(mai_mai_n1354_), .B0(mai_mai_n1370_), .B1(mai_mai_n1482_), .Y(mai_mai_n1484_));
  NO2        m1456(.A(mai_mai_n1484_), .B(mai_mai_n1481_), .Y(mai_mai_n1485_));
  NA4        m1457(.A(mai_mai_n1485_), .B(mai_mai_n1480_), .C(mai_mai_n1476_), .D(mai_mai_n1472_), .Y(mai_mai_n1486_));
  OR4        m1458(.A(mai_mai_n1486_), .B(mai_mai_n1463_), .C(mai_mai_n1420_), .D(mai_mai_n1374_), .Y(mai04));
  NOi31      m1459(.An(mai_mai_n1360_), .B(mai_mai_n1361_), .C(mai_mai_n1015_), .Y(mai_mai_n1488_));
  NA2        m1460(.A(mai_mai_n1416_), .B(mai_mai_n804_), .Y(mai_mai_n1489_));
  NO3        m1461(.A(mai_mai_n1489_), .B(mai_mai_n1004_), .C(mai_mai_n474_), .Y(mai_mai_n1490_));
  OR3        m1462(.A(mai_mai_n1490_), .B(mai_mai_n1488_), .C(mai_mai_n1033_), .Y(mai_mai_n1491_));
  NO2        m1463(.A(mai_mai_n1305_), .B(mai_mai_n88_), .Y(mai_mai_n1492_));
  AOI210     m1464(.A0(mai_mai_n1492_), .A1(mai_mai_n1026_), .B0(mai_mai_n1154_), .Y(mai_mai_n1493_));
  NA2        m1465(.A(mai_mai_n1493_), .B(mai_mai_n1181_), .Y(mai_mai_n1494_));
  NO4        m1466(.A(mai_mai_n1494_), .B(mai_mai_n1491_), .C(mai_mai_n1041_), .D(mai_mai_n1020_), .Y(mai_mai_n1495_));
  NA4        m1467(.A(mai_mai_n1495_), .B(mai_mai_n1097_), .C(mai_mai_n1083_), .D(mai_mai_n1071_), .Y(mai05));
  INV        m1468(.A(mai_mai_n588_), .Y(mai_mai_n1499_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NA2        u0033(.A(l), .B(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NA2        u0066(.A(m), .B(l), .Y(men_men_n95_));
  NAi31      u0067(.An(k), .B(j), .C(g), .Y(men_men_n96_));
  NO3        u0068(.A(men_men_n96_), .B(men_men_n95_), .C(f), .Y(men_men_n97_));
  AN2        u0069(.A(j), .B(g), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(l), .C(i), .Y(men_men_n99_));
  BUFFER     u0071(.A(g), .Y(men_men_n100_));
  NOi32      u0072(.An(m), .Bn(j), .C(k), .Y(men_men_n101_));
  NO2        u0073(.A(men_men_n97_), .B(men_men_n92_), .Y(men_men_n102_));
  NAi41      u0074(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n103_));
  AN2        u0075(.A(e), .B(b), .Y(men_men_n104_));
  NOi31      u0076(.An(c), .B(h), .C(f), .Y(men_men_n105_));
  NA2        u0077(.A(men_men_n105_), .B(men_men_n104_), .Y(men_men_n106_));
  NO2        u0078(.A(men_men_n106_), .B(men_men_n103_), .Y(men_men_n107_));
  NOi21      u0079(.An(i), .B(h), .Y(men_men_n108_));
  INV        u0080(.A(a), .Y(men_men_n109_));
  NA2        u0081(.A(men_men_n104_), .B(men_men_n109_), .Y(men_men_n110_));
  INV        u0082(.A(l), .Y(men_men_n111_));
  NOi21      u0083(.An(m), .B(n), .Y(men_men_n112_));
  AN2        u0084(.A(k), .B(h), .Y(men_men_n113_));
  INV        u0085(.A(b), .Y(men_men_n114_));
  NA2        u0086(.A(l), .B(j), .Y(men_men_n115_));
  AN2        u0087(.A(k), .B(i), .Y(men_men_n116_));
  NA2        u0088(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NA2        u0089(.A(g), .B(e), .Y(men_men_n118_));
  NOi32      u0090(.An(c), .Bn(a), .C(d), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n112_), .Y(men_men_n120_));
  NO4        u0092(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n117_), .D(men_men_n114_), .Y(men_men_n121_));
  NO2        u0093(.A(men_men_n121_), .B(men_men_n107_), .Y(men_men_n122_));
  OAI210     u0094(.A0(men_men_n102_), .A1(men_men_n88_), .B0(men_men_n122_), .Y(men_men_n123_));
  NOi31      u0095(.An(k), .B(m), .C(j), .Y(men_men_n124_));
  NOi31      u0096(.An(k), .B(m), .C(i), .Y(men_men_n125_));
  NOi32      u0097(.An(f), .Bn(b), .C(e), .Y(men_men_n126_));
  NAi21      u0098(.An(g), .B(h), .Y(men_men_n127_));
  NAi21      u0099(.An(m), .B(n), .Y(men_men_n128_));
  NAi21      u0100(.An(j), .B(k), .Y(men_men_n129_));
  NAi41      u0101(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n130_));
  NAi31      u0102(.An(j), .B(k), .C(h), .Y(men_men_n131_));
  NO3        u0103(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n132_));
  INV        u0104(.A(men_men_n132_), .Y(men_men_n133_));
  NO2        u0105(.A(k), .B(j), .Y(men_men_n134_));
  AN2        u0106(.A(k), .B(j), .Y(men_men_n135_));
  NAi21      u0107(.An(c), .B(b), .Y(men_men_n136_));
  NA2        u0108(.A(f), .B(d), .Y(men_men_n137_));
  NA2        u0109(.A(h), .B(c), .Y(men_men_n138_));
  NAi31      u0110(.An(f), .B(e), .C(b), .Y(men_men_n139_));
  NA2        u0111(.A(d), .B(b), .Y(men_men_n140_));
  NAi21      u0112(.An(e), .B(f), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n142_));
  NA2        u0114(.A(b), .B(a), .Y(men_men_n143_));
  NAi21      u0115(.An(c), .B(d), .Y(men_men_n144_));
  NAi31      u0116(.An(l), .B(k), .C(h), .Y(men_men_n145_));
  NO2        u0117(.A(men_men_n128_), .B(men_men_n145_), .Y(men_men_n146_));
  NA2        u0118(.A(men_men_n146_), .B(men_men_n142_), .Y(men_men_n147_));
  NA2        u0119(.A(men_men_n147_), .B(men_men_n133_), .Y(men_men_n148_));
  NAi31      u0120(.An(e), .B(f), .C(b), .Y(men_men_n149_));
  NOi21      u0121(.An(g), .B(d), .Y(men_men_n150_));
  NO2        u0122(.A(men_men_n150_), .B(men_men_n149_), .Y(men_men_n151_));
  NOi21      u0123(.An(h), .B(i), .Y(men_men_n152_));
  NOi21      u0124(.An(k), .B(m), .Y(men_men_n153_));
  NA3        u0125(.A(men_men_n153_), .B(men_men_n152_), .C(n), .Y(men_men_n154_));
  NOi21      u0126(.An(men_men_n151_), .B(men_men_n154_), .Y(men_men_n155_));
  NOi21      u0127(.An(h), .B(g), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n137_), .B(men_men_n136_), .Y(men_men_n157_));
  NA2        u0129(.A(men_men_n157_), .B(men_men_n156_), .Y(men_men_n158_));
  NAi31      u0130(.An(l), .B(j), .C(h), .Y(men_men_n159_));
  NOi32      u0131(.An(n), .Bn(k), .C(m), .Y(men_men_n160_));
  NA2        u0132(.A(l), .B(i), .Y(men_men_n161_));
  NA2        u0133(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NO2        u0134(.A(men_men_n162_), .B(men_men_n158_), .Y(men_men_n163_));
  NAi31      u0135(.An(d), .B(f), .C(c), .Y(men_men_n164_));
  NAi31      u0136(.An(e), .B(f), .C(c), .Y(men_men_n165_));
  NA2        u0137(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  NA2        u0138(.A(j), .B(h), .Y(men_men_n167_));
  OR3        u0139(.A(n), .B(m), .C(k), .Y(men_men_n168_));
  NO2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NAi32      u0141(.An(m), .Bn(k), .C(n), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n170_), .B(men_men_n167_), .Y(men_men_n171_));
  AOI220     u0143(.A0(men_men_n171_), .A1(men_men_n151_), .B0(men_men_n169_), .B1(men_men_n166_), .Y(men_men_n172_));
  NO2        u0144(.A(n), .B(m), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n50_), .Y(men_men_n174_));
  NAi21      u0146(.An(f), .B(e), .Y(men_men_n175_));
  NA2        u0147(.A(d), .B(c), .Y(men_men_n176_));
  NAi21      u0148(.An(d), .B(c), .Y(men_men_n177_));
  NAi31      u0149(.An(m), .B(n), .C(b), .Y(men_men_n178_));
  NAi21      u0150(.An(h), .B(f), .Y(men_men_n179_));
  NO2        u0151(.A(men_men_n178_), .B(men_men_n144_), .Y(men_men_n180_));
  NOi32      u0152(.An(f), .Bn(c), .C(d), .Y(men_men_n181_));
  NOi32      u0153(.An(f), .Bn(c), .C(e), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  NO3        u0155(.A(n), .B(m), .C(j), .Y(men_men_n184_));
  NA2        u0156(.A(men_men_n184_), .B(men_men_n113_), .Y(men_men_n185_));
  AO210      u0157(.A0(men_men_n185_), .A1(men_men_n174_), .B0(men_men_n183_), .Y(men_men_n186_));
  NA2        u0158(.A(men_men_n186_), .B(men_men_n172_), .Y(men_men_n187_));
  OR4        u0159(.A(men_men_n187_), .B(men_men_n163_), .C(men_men_n155_), .D(men_men_n148_), .Y(men_men_n188_));
  NO4        u0160(.A(men_men_n188_), .B(men_men_n123_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n189_));
  NA3        u0161(.A(m), .B(men_men_n111_), .C(j), .Y(men_men_n190_));
  NAi31      u0162(.An(n), .B(h), .C(g), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi32      u0164(.An(m), .Bn(k), .C(l), .Y(men_men_n193_));
  NA3        u0165(.A(men_men_n193_), .B(men_men_n89_), .C(g), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(n), .Y(men_men_n195_));
  AN2        u0167(.A(i), .B(g), .Y(men_men_n196_));
  NA3        u0168(.A(men_men_n76_), .B(men_men_n196_), .C(men_men_n112_), .Y(men_men_n197_));
  INV        u0169(.A(men_men_n197_), .Y(men_men_n198_));
  NO3        u0170(.A(men_men_n198_), .B(men_men_n195_), .C(men_men_n192_), .Y(men_men_n199_));
  NAi41      u0171(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n200_));
  INV        u0172(.A(f), .Y(men_men_n201_));
  INV        u0173(.A(g), .Y(men_men_n202_));
  NOi31      u0174(.An(i), .B(j), .C(h), .Y(men_men_n203_));
  NOi21      u0175(.An(l), .B(m), .Y(men_men_n204_));
  NA2        u0176(.A(men_men_n204_), .B(men_men_n203_), .Y(men_men_n205_));
  NO3        u0177(.A(men_men_n205_), .B(men_men_n202_), .C(men_men_n201_), .Y(men_men_n206_));
  NO2        u0178(.A(men_men_n199_), .B(men_men_n32_), .Y(men_men_n207_));
  NOi21      u0179(.An(n), .B(m), .Y(men_men_n208_));
  NOi32      u0180(.An(l), .Bn(i), .C(j), .Y(men_men_n209_));
  NA2        u0181(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  OA220      u0182(.A0(men_men_n210_), .A1(men_men_n106_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n211_));
  NAi21      u0183(.An(j), .B(h), .Y(men_men_n212_));
  XN2        u0184(.A(i), .B(h), .Y(men_men_n213_));
  NA2        u0185(.A(men_men_n213_), .B(men_men_n212_), .Y(men_men_n214_));
  NOi31      u0186(.An(k), .B(n), .C(m), .Y(men_men_n215_));
  NOi31      u0187(.An(men_men_n215_), .B(men_men_n176_), .C(men_men_n175_), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n214_), .Y(men_men_n217_));
  NAi31      u0189(.An(f), .B(e), .C(c), .Y(men_men_n218_));
  NO4        u0190(.A(men_men_n218_), .B(men_men_n168_), .C(men_men_n167_), .D(men_men_n59_), .Y(men_men_n219_));
  NA4        u0191(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n220_));
  NAi32      u0192(.An(m), .Bn(i), .C(k), .Y(men_men_n221_));
  NO3        u0193(.A(men_men_n221_), .B(men_men_n93_), .C(men_men_n220_), .Y(men_men_n222_));
  INV        u0194(.A(k), .Y(men_men_n223_));
  NO2        u0195(.A(men_men_n222_), .B(men_men_n219_), .Y(men_men_n224_));
  NAi21      u0196(.An(n), .B(a), .Y(men_men_n225_));
  NO2        u0197(.A(men_men_n225_), .B(men_men_n140_), .Y(men_men_n226_));
  NAi41      u0198(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n227_));
  NO2        u0199(.A(men_men_n227_), .B(e), .Y(men_men_n228_));
  NO3        u0200(.A(men_men_n141_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n229_));
  OAI210     u0201(.A0(men_men_n229_), .A1(men_men_n228_), .B0(men_men_n226_), .Y(men_men_n230_));
  AN4        u0202(.A(men_men_n230_), .B(men_men_n224_), .C(men_men_n217_), .D(men_men_n211_), .Y(men_men_n231_));
  OR2        u0203(.A(h), .B(g), .Y(men_men_n232_));
  NAi41      u0204(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n233_));
  NO2        u0205(.A(men_men_n233_), .B(men_men_n201_), .Y(men_men_n234_));
  NA2        u0206(.A(men_men_n153_), .B(men_men_n108_), .Y(men_men_n235_));
  NAi21      u0207(.An(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  NO2        u0208(.A(n), .B(a), .Y(men_men_n237_));
  NAi31      u0209(.An(men_men_n227_), .B(men_men_n237_), .C(men_men_n104_), .Y(men_men_n238_));
  AN2        u0210(.A(men_men_n238_), .B(men_men_n236_), .Y(men_men_n239_));
  NAi21      u0211(.An(h), .B(i), .Y(men_men_n240_));
  NA2        u0212(.A(men_men_n173_), .B(k), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n240_), .Y(men_men_n242_));
  NA2        u0214(.A(men_men_n242_), .B(men_men_n181_), .Y(men_men_n243_));
  NA2        u0215(.A(men_men_n243_), .B(men_men_n239_), .Y(men_men_n244_));
  NOi21      u0216(.An(g), .B(e), .Y(men_men_n245_));
  NO2        u0217(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n246_));
  NA2        u0218(.A(men_men_n246_), .B(men_men_n245_), .Y(men_men_n247_));
  NOi32      u0219(.An(l), .Bn(j), .C(i), .Y(men_men_n248_));
  AOI210     u0220(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n248_), .Y(men_men_n249_));
  NAi21      u0221(.An(f), .B(g), .Y(men_men_n250_));
  NO2        u0222(.A(men_men_n250_), .B(men_men_n65_), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n69_), .B(men_men_n115_), .Y(men_men_n252_));
  NA2        u0224(.A(men_men_n252_), .B(men_men_n251_), .Y(men_men_n253_));
  OAI210     u0225(.A0(men_men_n249_), .A1(men_men_n247_), .B0(men_men_n253_), .Y(men_men_n254_));
  NO3        u0226(.A(men_men_n129_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n255_));
  NOi41      u0227(.An(men_men_n231_), .B(men_men_n254_), .C(men_men_n244_), .D(men_men_n207_), .Y(men_men_n256_));
  NO4        u0228(.A(men_men_n192_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n257_), .B(men_men_n110_), .Y(men_men_n258_));
  NA3        u0230(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n259_));
  NAi21      u0231(.An(h), .B(g), .Y(men_men_n260_));
  OR4        u0232(.A(men_men_n260_), .B(men_men_n259_), .C(men_men_n210_), .D(e), .Y(men_men_n261_));
  NO2        u0233(.A(men_men_n235_), .B(men_men_n250_), .Y(men_men_n262_));
  NAi31      u0234(.An(g), .B(k), .C(h), .Y(men_men_n263_));
  NO3        u0235(.A(men_men_n128_), .B(men_men_n263_), .C(l), .Y(men_men_n264_));
  NAi31      u0236(.An(e), .B(d), .C(a), .Y(men_men_n265_));
  NA2        u0237(.A(men_men_n264_), .B(men_men_n126_), .Y(men_men_n266_));
  NA2        u0238(.A(men_men_n266_), .B(men_men_n261_), .Y(men_men_n267_));
  NA4        u0239(.A(men_men_n153_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n115_), .Y(men_men_n268_));
  NA3        u0240(.A(men_men_n153_), .B(men_men_n152_), .C(men_men_n86_), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n269_), .B(men_men_n183_), .Y(men_men_n270_));
  NOi21      u0242(.An(men_men_n268_), .B(men_men_n270_), .Y(men_men_n271_));
  NA3        u0243(.A(e), .B(c), .C(b), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n60_), .B(men_men_n272_), .Y(men_men_n273_));
  NAi32      u0245(.An(k), .Bn(i), .C(j), .Y(men_men_n274_));
  NAi31      u0246(.An(h), .B(l), .C(i), .Y(men_men_n275_));
  NA3        u0247(.A(men_men_n275_), .B(men_men_n274_), .C(men_men_n159_), .Y(men_men_n276_));
  NOi21      u0248(.An(men_men_n276_), .B(men_men_n49_), .Y(men_men_n277_));
  OAI210     u0249(.A0(men_men_n251_), .A1(men_men_n273_), .B0(men_men_n277_), .Y(men_men_n278_));
  NAi21      u0250(.An(l), .B(k), .Y(men_men_n279_));
  NO2        u0251(.A(men_men_n279_), .B(men_men_n49_), .Y(men_men_n280_));
  NOi21      u0252(.An(l), .B(j), .Y(men_men_n281_));
  NA2        u0253(.A(men_men_n156_), .B(men_men_n281_), .Y(men_men_n282_));
  NA3        u0254(.A(men_men_n116_), .B(men_men_n115_), .C(g), .Y(men_men_n283_));
  OR3        u0255(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n284_));
  AOI210     u0256(.A0(men_men_n283_), .A1(men_men_n282_), .B0(men_men_n284_), .Y(men_men_n285_));
  INV        u0257(.A(men_men_n285_), .Y(men_men_n286_));
  NAi32      u0258(.An(j), .Bn(h), .C(i), .Y(men_men_n287_));
  NAi21      u0259(.An(m), .B(l), .Y(men_men_n288_));
  NO3        u0260(.A(men_men_n288_), .B(men_men_n287_), .C(men_men_n86_), .Y(men_men_n289_));
  NA2        u0261(.A(h), .B(g), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n289_), .B(men_men_n157_), .Y(men_men_n291_));
  NA4        u0263(.A(men_men_n291_), .B(men_men_n286_), .C(men_men_n278_), .D(men_men_n271_), .Y(men_men_n292_));
  NO2        u0264(.A(men_men_n139_), .B(d), .Y(men_men_n293_));
  NA2        u0265(.A(men_men_n293_), .B(men_men_n53_), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n106_), .B(men_men_n103_), .Y(men_men_n295_));
  NAi32      u0267(.An(n), .Bn(m), .C(l), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n296_), .B(men_men_n287_), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n120_), .B(men_men_n114_), .Y(men_men_n298_));
  NAi31      u0270(.An(k), .B(l), .C(j), .Y(men_men_n299_));
  OAI210     u0271(.A0(men_men_n279_), .A1(j), .B0(men_men_n299_), .Y(men_men_n300_));
  NOi21      u0272(.An(men_men_n300_), .B(men_men_n118_), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n301_), .B(men_men_n298_), .Y(men_men_n302_));
  NA2        u0274(.A(men_men_n302_), .B(men_men_n294_), .Y(men_men_n303_));
  NO4        u0275(.A(men_men_n303_), .B(men_men_n292_), .C(men_men_n267_), .D(men_men_n258_), .Y(men_men_n304_));
  NA2        u0276(.A(men_men_n242_), .B(men_men_n182_), .Y(men_men_n305_));
  NAi21      u0277(.An(m), .B(k), .Y(men_men_n306_));
  NO2        u0278(.A(men_men_n213_), .B(men_men_n306_), .Y(men_men_n307_));
  NAi41      u0279(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n308_));
  NAi31      u0280(.An(i), .B(l), .C(h), .Y(men_men_n309_));
  NO4        u0281(.A(men_men_n309_), .B(e), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n310_));
  NA2        u0282(.A(e), .B(c), .Y(men_men_n311_));
  NO3        u0283(.A(men_men_n311_), .B(n), .C(d), .Y(men_men_n312_));
  NOi21      u0284(.An(f), .B(h), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n116_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n314_), .B(men_men_n202_), .Y(men_men_n315_));
  NAi31      u0287(.An(d), .B(e), .C(b), .Y(men_men_n316_));
  NO2        u0288(.A(men_men_n128_), .B(men_men_n316_), .Y(men_men_n317_));
  NA2        u0289(.A(men_men_n317_), .B(men_men_n315_), .Y(men_men_n318_));
  NAi31      u0290(.An(men_men_n310_), .B(men_men_n318_), .C(men_men_n305_), .Y(men_men_n319_));
  NO4        u0291(.A(men_men_n308_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n202_), .Y(men_men_n320_));
  NA2        u0292(.A(men_men_n237_), .B(men_men_n104_), .Y(men_men_n321_));
  OR2        u0293(.A(men_men_n321_), .B(men_men_n194_), .Y(men_men_n322_));
  NOi31      u0294(.An(l), .B(n), .C(m), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n203_), .Y(men_men_n324_));
  NO2        u0296(.A(men_men_n324_), .B(men_men_n183_), .Y(men_men_n325_));
  NAi32      u0297(.An(men_men_n325_), .Bn(men_men_n320_), .C(men_men_n322_), .Y(men_men_n326_));
  NAi32      u0298(.An(m), .Bn(j), .C(k), .Y(men_men_n327_));
  NAi41      u0299(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n328_));
  OAI210     u0300(.A0(men_men_n200_), .A1(men_men_n327_), .B0(men_men_n328_), .Y(men_men_n329_));
  NOi31      u0301(.An(j), .B(m), .C(k), .Y(men_men_n330_));
  NO2        u0302(.A(men_men_n124_), .B(men_men_n330_), .Y(men_men_n331_));
  AN3        u0303(.A(h), .B(g), .C(f), .Y(men_men_n332_));
  NAi31      u0304(.An(men_men_n331_), .B(men_men_n332_), .C(men_men_n329_), .Y(men_men_n333_));
  NOi32      u0305(.An(m), .Bn(j), .C(l), .Y(men_men_n334_));
  NO2        u0306(.A(men_men_n334_), .B(men_men_n99_), .Y(men_men_n335_));
  NAi32      u0307(.An(men_men_n335_), .Bn(men_men_n191_), .C(men_men_n293_), .Y(men_men_n336_));
  NO2        u0308(.A(men_men_n288_), .B(men_men_n287_), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n205_), .B(g), .Y(men_men_n338_));
  NO2        u0310(.A(men_men_n149_), .B(men_men_n86_), .Y(men_men_n339_));
  AOI220     u0311(.A0(men_men_n339_), .A1(men_men_n338_), .B0(men_men_n234_), .B1(men_men_n337_), .Y(men_men_n340_));
  NA3        u0312(.A(men_men_n340_), .B(men_men_n336_), .C(men_men_n333_), .Y(men_men_n341_));
  NA3        u0313(.A(h), .B(g), .C(f), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n342_), .B(men_men_n77_), .Y(men_men_n343_));
  NA2        u0315(.A(men_men_n328_), .B(men_men_n200_), .Y(men_men_n344_));
  NA2        u0316(.A(men_men_n156_), .B(e), .Y(men_men_n345_));
  NO2        u0317(.A(men_men_n345_), .B(men_men_n41_), .Y(men_men_n346_));
  AOI220     u0318(.A0(men_men_n346_), .A1(men_men_n298_), .B0(men_men_n344_), .B1(men_men_n343_), .Y(men_men_n347_));
  NOi32      u0319(.An(j), .Bn(g), .C(i), .Y(men_men_n348_));
  NA3        u0320(.A(men_men_n348_), .B(men_men_n279_), .C(men_men_n112_), .Y(men_men_n349_));
  NOi32      u0321(.An(e), .Bn(b), .C(a), .Y(men_men_n350_));
  AN2        u0322(.A(l), .B(j), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n306_), .B(men_men_n351_), .Y(men_men_n352_));
  NO3        u0324(.A(men_men_n308_), .B(men_men_n72_), .C(men_men_n202_), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n197_), .B(men_men_n35_), .Y(men_men_n354_));
  AOI220     u0326(.A0(men_men_n354_), .A1(men_men_n350_), .B0(men_men_n353_), .B1(men_men_n352_), .Y(men_men_n355_));
  NO2        u0327(.A(men_men_n316_), .B(n), .Y(men_men_n356_));
  NA2        u0328(.A(men_men_n196_), .B(k), .Y(men_men_n357_));
  NA3        u0329(.A(m), .B(men_men_n111_), .C(men_men_n201_), .Y(men_men_n358_));
  NA4        u0330(.A(men_men_n193_), .B(men_men_n89_), .C(g), .D(men_men_n201_), .Y(men_men_n359_));
  OAI210     u0331(.A0(men_men_n358_), .A1(men_men_n357_), .B0(men_men_n359_), .Y(men_men_n360_));
  NAi41      u0332(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n361_));
  NA2        u0333(.A(men_men_n51_), .B(men_men_n112_), .Y(men_men_n362_));
  NO2        u0334(.A(men_men_n362_), .B(men_men_n361_), .Y(men_men_n363_));
  AOI220     u0335(.A0(men_men_n363_), .A1(b), .B0(men_men_n360_), .B1(men_men_n356_), .Y(men_men_n364_));
  NA3        u0336(.A(men_men_n364_), .B(men_men_n355_), .C(men_men_n347_), .Y(men_men_n365_));
  NO4        u0337(.A(men_men_n365_), .B(men_men_n341_), .C(men_men_n326_), .D(men_men_n319_), .Y(men_men_n366_));
  NA4        u0338(.A(men_men_n366_), .B(men_men_n304_), .C(men_men_n256_), .D(men_men_n189_), .Y(men10));
  NA3        u0339(.A(m), .B(k), .C(i), .Y(men_men_n368_));
  NO3        u0340(.A(men_men_n368_), .B(j), .C(men_men_n202_), .Y(men_men_n369_));
  NOi21      u0341(.An(e), .B(f), .Y(men_men_n370_));
  NO4        u0342(.A(men_men_n144_), .B(men_men_n370_), .C(n), .D(men_men_n109_), .Y(men_men_n371_));
  NAi31      u0343(.An(b), .B(f), .C(c), .Y(men_men_n372_));
  INV        u0344(.A(men_men_n372_), .Y(men_men_n373_));
  NOi32      u0345(.An(k), .Bn(h), .C(j), .Y(men_men_n374_));
  NA2        u0346(.A(men_men_n374_), .B(men_men_n208_), .Y(men_men_n375_));
  NA2        u0347(.A(men_men_n154_), .B(men_men_n375_), .Y(men_men_n376_));
  AOI220     u0348(.A0(men_men_n376_), .A1(men_men_n373_), .B0(men_men_n371_), .B1(men_men_n369_), .Y(men_men_n377_));
  AN2        u0349(.A(j), .B(h), .Y(men_men_n378_));
  NO3        u0350(.A(n), .B(m), .C(k), .Y(men_men_n379_));
  NA2        u0351(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n380_));
  NO3        u0352(.A(men_men_n380_), .B(men_men_n144_), .C(men_men_n201_), .Y(men_men_n381_));
  OR2        u0353(.A(m), .B(k), .Y(men_men_n382_));
  NO2        u0354(.A(men_men_n167_), .B(men_men_n382_), .Y(men_men_n383_));
  NA4        u0355(.A(n), .B(f), .C(c), .D(men_men_n114_), .Y(men_men_n384_));
  NOi21      u0356(.An(men_men_n383_), .B(men_men_n384_), .Y(men_men_n385_));
  NOi32      u0357(.An(d), .Bn(a), .C(c), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n386_), .B(men_men_n175_), .Y(men_men_n387_));
  NAi21      u0359(.An(i), .B(g), .Y(men_men_n388_));
  NAi31      u0360(.An(k), .B(m), .C(j), .Y(men_men_n389_));
  NO2        u0361(.A(men_men_n385_), .B(men_men_n381_), .Y(men_men_n390_));
  NO2        u0362(.A(men_men_n384_), .B(men_men_n288_), .Y(men_men_n391_));
  NOi32      u0363(.An(f), .Bn(d), .C(c), .Y(men_men_n392_));
  AOI220     u0364(.A0(men_men_n392_), .A1(men_men_n297_), .B0(men_men_n391_), .B1(men_men_n203_), .Y(men_men_n393_));
  NA3        u0365(.A(men_men_n393_), .B(men_men_n390_), .C(men_men_n377_), .Y(men_men_n394_));
  NO2        u0366(.A(men_men_n59_), .B(men_men_n114_), .Y(men_men_n395_));
  NA2        u0367(.A(men_men_n237_), .B(men_men_n395_), .Y(men_men_n396_));
  INV        u0368(.A(e), .Y(men_men_n397_));
  NA2        u0369(.A(men_men_n46_), .B(e), .Y(men_men_n398_));
  OAI220     u0370(.A0(men_men_n398_), .A1(men_men_n190_), .B0(men_men_n194_), .B1(men_men_n397_), .Y(men_men_n399_));
  AN2        u0371(.A(g), .B(e), .Y(men_men_n400_));
  NA3        u0372(.A(men_men_n400_), .B(men_men_n193_), .C(i), .Y(men_men_n401_));
  INV        u0373(.A(men_men_n401_), .Y(men_men_n402_));
  NO2        u0374(.A(men_men_n402_), .B(men_men_n399_), .Y(men_men_n403_));
  NOi32      u0375(.An(h), .Bn(e), .C(g), .Y(men_men_n404_));
  NA3        u0376(.A(men_men_n404_), .B(men_men_n281_), .C(m), .Y(men_men_n405_));
  NOi21      u0377(.An(g), .B(h), .Y(men_men_n406_));
  AN3        u0378(.A(m), .B(l), .C(i), .Y(men_men_n407_));
  NA3        u0379(.A(men_men_n407_), .B(men_men_n406_), .C(e), .Y(men_men_n408_));
  AN3        u0380(.A(h), .B(g), .C(e), .Y(men_men_n409_));
  NA2        u0381(.A(men_men_n409_), .B(men_men_n99_), .Y(men_men_n410_));
  AN3        u0382(.A(men_men_n410_), .B(men_men_n408_), .C(men_men_n405_), .Y(men_men_n411_));
  AOI210     u0383(.A0(men_men_n411_), .A1(men_men_n403_), .B0(men_men_n396_), .Y(men_men_n412_));
  NA3        u0384(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n413_), .B(men_men_n396_), .Y(men_men_n414_));
  NAi31      u0386(.An(b), .B(c), .C(a), .Y(men_men_n415_));
  NO2        u0387(.A(men_men_n415_), .B(n), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n51_), .B(m), .Y(men_men_n417_));
  NO2        u0389(.A(men_men_n417_), .B(men_men_n141_), .Y(men_men_n418_));
  NA2        u0390(.A(men_men_n418_), .B(men_men_n416_), .Y(men_men_n419_));
  INV        u0391(.A(men_men_n419_), .Y(men_men_n420_));
  NO4        u0392(.A(men_men_n420_), .B(men_men_n414_), .C(men_men_n412_), .D(men_men_n394_), .Y(men_men_n421_));
  NA2        u0393(.A(i), .B(g), .Y(men_men_n422_));
  NO3        u0394(.A(men_men_n265_), .B(men_men_n422_), .C(c), .Y(men_men_n423_));
  NOi21      u0395(.An(a), .B(n), .Y(men_men_n424_));
  NOi21      u0396(.An(d), .B(c), .Y(men_men_n425_));
  NA2        u0397(.A(men_men_n425_), .B(men_men_n424_), .Y(men_men_n426_));
  NA3        u0398(.A(i), .B(g), .C(f), .Y(men_men_n427_));
  OR2        u0399(.A(men_men_n427_), .B(men_men_n71_), .Y(men_men_n428_));
  NA3        u0400(.A(men_men_n407_), .B(men_men_n406_), .C(men_men_n175_), .Y(men_men_n429_));
  AOI210     u0401(.A0(men_men_n429_), .A1(men_men_n428_), .B0(men_men_n426_), .Y(men_men_n430_));
  AOI210     u0402(.A0(men_men_n423_), .A1(men_men_n280_), .B0(men_men_n430_), .Y(men_men_n431_));
  OR2        u0403(.A(n), .B(m), .Y(men_men_n432_));
  NO2        u0404(.A(men_men_n432_), .B(men_men_n145_), .Y(men_men_n433_));
  NO2        u0405(.A(men_men_n176_), .B(men_men_n141_), .Y(men_men_n434_));
  OAI210     u0406(.A0(men_men_n433_), .A1(men_men_n169_), .B0(men_men_n434_), .Y(men_men_n435_));
  INV        u0407(.A(men_men_n362_), .Y(men_men_n436_));
  NA3        u0408(.A(men_men_n436_), .B(men_men_n350_), .C(d), .Y(men_men_n437_));
  NO2        u0409(.A(men_men_n415_), .B(men_men_n49_), .Y(men_men_n438_));
  NAi21      u0410(.An(k), .B(j), .Y(men_men_n439_));
  NAi21      u0411(.An(e), .B(d), .Y(men_men_n440_));
  INV        u0412(.A(men_men_n440_), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n241_), .B(men_men_n201_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n442_), .B(men_men_n441_), .C(men_men_n214_), .Y(men_men_n443_));
  NA3        u0415(.A(men_men_n443_), .B(men_men_n437_), .C(men_men_n435_), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n324_), .B(men_men_n201_), .Y(men_men_n445_));
  NA2        u0417(.A(men_men_n445_), .B(men_men_n441_), .Y(men_men_n446_));
  NOi31      u0418(.An(n), .B(m), .C(k), .Y(men_men_n447_));
  AOI220     u0419(.A0(men_men_n447_), .A1(men_men_n378_), .B0(men_men_n208_), .B1(men_men_n50_), .Y(men_men_n448_));
  NAi31      u0420(.An(g), .B(f), .C(c), .Y(men_men_n449_));
  INV        u0421(.A(men_men_n446_), .Y(men_men_n450_));
  NOi41      u0422(.An(men_men_n431_), .B(men_men_n450_), .C(men_men_n444_), .D(men_men_n254_), .Y(men_men_n451_));
  NOi32      u0423(.An(c), .Bn(a), .C(b), .Y(men_men_n452_));
  NA2        u0424(.A(men_men_n452_), .B(men_men_n112_), .Y(men_men_n453_));
  INV        u0425(.A(men_men_n263_), .Y(men_men_n454_));
  AN2        u0426(.A(e), .B(d), .Y(men_men_n455_));
  NA2        u0427(.A(men_men_n455_), .B(men_men_n454_), .Y(men_men_n456_));
  INV        u0428(.A(men_men_n141_), .Y(men_men_n457_));
  NO2        u0429(.A(men_men_n127_), .B(men_men_n41_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n66_), .B(e), .Y(men_men_n459_));
  NOi31      u0431(.An(j), .B(k), .C(i), .Y(men_men_n460_));
  NOi21      u0432(.An(men_men_n159_), .B(men_men_n460_), .Y(men_men_n461_));
  NA4        u0433(.A(men_men_n309_), .B(men_men_n461_), .C(men_men_n249_), .D(men_men_n117_), .Y(men_men_n462_));
  AOI220     u0434(.A0(men_men_n462_), .A1(men_men_n459_), .B0(men_men_n458_), .B1(men_men_n457_), .Y(men_men_n463_));
  AOI210     u0435(.A0(men_men_n463_), .A1(men_men_n456_), .B0(men_men_n453_), .Y(men_men_n464_));
  NOi21      u0436(.An(a), .B(b), .Y(men_men_n465_));
  NA3        u0437(.A(e), .B(d), .C(c), .Y(men_men_n466_));
  NAi21      u0438(.An(men_men_n466_), .B(men_men_n465_), .Y(men_men_n467_));
  AOI210     u0439(.A0(men_men_n257_), .A1(men_men_n197_), .B0(men_men_n467_), .Y(men_men_n468_));
  NO4        u0440(.A(men_men_n179_), .B(men_men_n103_), .C(men_men_n56_), .D(b), .Y(men_men_n469_));
  NA2        u0441(.A(men_men_n373_), .B(men_men_n146_), .Y(men_men_n470_));
  OR2        u0442(.A(k), .B(j), .Y(men_men_n471_));
  NA2        u0443(.A(l), .B(k), .Y(men_men_n472_));
  NA3        u0444(.A(men_men_n472_), .B(men_men_n471_), .C(men_men_n208_), .Y(men_men_n473_));
  AOI210     u0445(.A0(men_men_n221_), .A1(men_men_n327_), .B0(men_men_n86_), .Y(men_men_n474_));
  NOi21      u0446(.An(men_men_n473_), .B(men_men_n474_), .Y(men_men_n475_));
  OR3        u0447(.A(men_men_n475_), .B(men_men_n138_), .C(men_men_n130_), .Y(men_men_n476_));
  INV        u0448(.A(men_men_n268_), .Y(men_men_n477_));
  NA2        u0449(.A(men_men_n386_), .B(men_men_n112_), .Y(men_men_n478_));
  NO4        u0450(.A(men_men_n478_), .B(men_men_n96_), .C(men_men_n111_), .D(e), .Y(men_men_n479_));
  NO3        u0451(.A(men_men_n479_), .B(men_men_n477_), .C(men_men_n310_), .Y(men_men_n480_));
  NA3        u0452(.A(men_men_n480_), .B(men_men_n476_), .C(men_men_n470_), .Y(men_men_n481_));
  NO4        u0453(.A(men_men_n481_), .B(men_men_n469_), .C(men_men_n468_), .D(men_men_n464_), .Y(men_men_n482_));
  NA2        u0454(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n483_));
  NOi21      u0455(.An(d), .B(e), .Y(men_men_n484_));
  NO2        u0456(.A(men_men_n179_), .B(men_men_n56_), .Y(men_men_n485_));
  NAi31      u0457(.An(j), .B(l), .C(i), .Y(men_men_n486_));
  OAI210     u0458(.A0(men_men_n486_), .A1(men_men_n128_), .B0(men_men_n103_), .Y(men_men_n487_));
  NA3        u0459(.A(men_men_n487_), .B(men_men_n485_), .C(men_men_n484_), .Y(men_men_n488_));
  NO3        u0460(.A(men_men_n387_), .B(men_men_n335_), .C(men_men_n191_), .Y(men_men_n489_));
  NO2        u0461(.A(men_men_n387_), .B(men_men_n362_), .Y(men_men_n490_));
  NO3        u0462(.A(men_men_n490_), .B(men_men_n489_), .C(men_men_n295_), .Y(men_men_n491_));
  NA4        u0463(.A(men_men_n491_), .B(men_men_n488_), .C(men_men_n483_), .D(men_men_n231_), .Y(men_men_n492_));
  OAI210     u0464(.A0(men_men_n125_), .A1(men_men_n124_), .B0(n), .Y(men_men_n493_));
  NO2        u0465(.A(men_men_n493_), .B(men_men_n127_), .Y(men_men_n494_));
  OA210      u0466(.A0(men_men_n289_), .A1(men_men_n494_), .B0(men_men_n182_), .Y(men_men_n495_));
  XO2        u0467(.A(i), .B(h), .Y(men_men_n496_));
  NA3        u0468(.A(men_men_n496_), .B(men_men_n153_), .C(n), .Y(men_men_n497_));
  NAi41      u0469(.An(men_men_n289_), .B(men_men_n497_), .C(men_men_n448_), .D(men_men_n375_), .Y(men_men_n498_));
  NOi32      u0470(.An(men_men_n498_), .Bn(men_men_n459_), .C(men_men_n259_), .Y(men_men_n499_));
  NAi31      u0471(.An(c), .B(f), .C(d), .Y(men_men_n500_));
  AOI210     u0472(.A0(men_men_n269_), .A1(men_men_n185_), .B0(men_men_n500_), .Y(men_men_n501_));
  NOi21      u0473(.An(men_men_n84_), .B(men_men_n501_), .Y(men_men_n502_));
  NA2        u0474(.A(men_men_n215_), .B(men_men_n108_), .Y(men_men_n503_));
  AOI210     u0475(.A0(men_men_n503_), .A1(men_men_n174_), .B0(men_men_n500_), .Y(men_men_n504_));
  AOI210     u0476(.A0(men_men_n349_), .A1(men_men_n35_), .B0(men_men_n467_), .Y(men_men_n505_));
  NO2        u0477(.A(men_men_n505_), .B(men_men_n504_), .Y(men_men_n506_));
  AN2        u0478(.A(men_men_n277_), .B(men_men_n251_), .Y(men_men_n507_));
  NA3        u0479(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n508_));
  NO2        u0480(.A(men_men_n508_), .B(men_men_n426_), .Y(men_men_n509_));
  NO2        u0481(.A(men_men_n509_), .B(men_men_n285_), .Y(men_men_n510_));
  NAi41      u0482(.An(men_men_n507_), .B(men_men_n510_), .C(men_men_n506_), .D(men_men_n502_), .Y(men_men_n511_));
  NO4        u0483(.A(men_men_n511_), .B(men_men_n499_), .C(men_men_n495_), .D(men_men_n492_), .Y(men_men_n512_));
  NA4        u0484(.A(men_men_n512_), .B(men_men_n482_), .C(men_men_n451_), .D(men_men_n421_), .Y(men11));
  NO2        u0485(.A(men_men_n73_), .B(f), .Y(men_men_n514_));
  NA2        u0486(.A(j), .B(g), .Y(men_men_n515_));
  NAi31      u0487(.An(i), .B(m), .C(l), .Y(men_men_n516_));
  NA3        u0488(.A(m), .B(k), .C(j), .Y(men_men_n517_));
  OAI220     u0489(.A0(men_men_n517_), .A1(men_men_n127_), .B0(men_men_n516_), .B1(men_men_n515_), .Y(men_men_n518_));
  NA2        u0490(.A(men_men_n518_), .B(men_men_n514_), .Y(men_men_n519_));
  NOi32      u0491(.An(e), .Bn(b), .C(f), .Y(men_men_n520_));
  NA2        u0492(.A(men_men_n248_), .B(men_men_n112_), .Y(men_men_n521_));
  NA2        u0493(.A(men_men_n46_), .B(j), .Y(men_men_n522_));
  NAi31      u0494(.An(d), .B(e), .C(a), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n523_), .B(n), .Y(men_men_n524_));
  NAi41      u0496(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n525_));
  AN2        u0497(.A(men_men_n525_), .B(men_men_n361_), .Y(men_men_n526_));
  AOI210     u0498(.A0(men_men_n526_), .A1(men_men_n387_), .B0(men_men_n260_), .Y(men_men_n527_));
  NA2        u0499(.A(j), .B(i), .Y(men_men_n528_));
  NAi31      u0500(.An(n), .B(m), .C(k), .Y(men_men_n529_));
  NO3        u0501(.A(men_men_n529_), .B(men_men_n528_), .C(men_men_n111_), .Y(men_men_n530_));
  NO4        u0502(.A(n), .B(d), .C(men_men_n114_), .D(a), .Y(men_men_n531_));
  OR2        u0503(.A(n), .B(c), .Y(men_men_n532_));
  NO2        u0504(.A(men_men_n532_), .B(men_men_n143_), .Y(men_men_n533_));
  NO2        u0505(.A(men_men_n533_), .B(men_men_n531_), .Y(men_men_n534_));
  NOi32      u0506(.An(g), .Bn(f), .C(i), .Y(men_men_n535_));
  AOI220     u0507(.A0(men_men_n535_), .A1(men_men_n101_), .B0(men_men_n518_), .B1(f), .Y(men_men_n536_));
  NO2        u0508(.A(men_men_n263_), .B(men_men_n49_), .Y(men_men_n537_));
  NO2        u0509(.A(men_men_n536_), .B(men_men_n534_), .Y(men_men_n538_));
  AOI210     u0510(.A0(men_men_n530_), .A1(men_men_n527_), .B0(men_men_n538_), .Y(men_men_n539_));
  NA2        u0511(.A(men_men_n135_), .B(men_men_n34_), .Y(men_men_n540_));
  OAI220     u0512(.A0(men_men_n540_), .A1(m), .B0(men_men_n522_), .B1(men_men_n221_), .Y(men_men_n541_));
  NOi41      u0513(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n542_));
  NAi32      u0514(.An(e), .Bn(b), .C(c), .Y(men_men_n543_));
  OR2        u0515(.A(men_men_n543_), .B(men_men_n86_), .Y(men_men_n544_));
  AN2        u0516(.A(men_men_n328_), .B(men_men_n308_), .Y(men_men_n545_));
  NA2        u0517(.A(men_men_n545_), .B(men_men_n544_), .Y(men_men_n546_));
  OA210      u0518(.A0(men_men_n546_), .A1(men_men_n542_), .B0(men_men_n541_), .Y(men_men_n547_));
  OAI220     u0519(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n516_), .B1(men_men_n515_), .Y(men_men_n548_));
  NAi31      u0520(.An(d), .B(c), .C(a), .Y(men_men_n549_));
  NO2        u0521(.A(men_men_n549_), .B(n), .Y(men_men_n550_));
  NA3        u0522(.A(men_men_n550_), .B(men_men_n548_), .C(e), .Y(men_men_n551_));
  INV        u0523(.A(men_men_n551_), .Y(men_men_n552_));
  NO2        u0524(.A(men_men_n265_), .B(n), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n416_), .B(men_men_n553_), .Y(men_men_n554_));
  NA2        u0526(.A(men_men_n548_), .B(f), .Y(men_men_n555_));
  NAi32      u0527(.An(d), .Bn(a), .C(b), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n556_), .B(men_men_n49_), .Y(men_men_n557_));
  NA2        u0529(.A(h), .B(f), .Y(men_men_n558_));
  NO2        u0530(.A(men_men_n558_), .B(men_men_n96_), .Y(men_men_n559_));
  NO3        u0531(.A(men_men_n170_), .B(men_men_n167_), .C(g), .Y(men_men_n560_));
  AOI220     u0532(.A0(men_men_n560_), .A1(men_men_n58_), .B0(men_men_n559_), .B1(men_men_n557_), .Y(men_men_n561_));
  OAI210     u0533(.A0(men_men_n555_), .A1(men_men_n554_), .B0(men_men_n561_), .Y(men_men_n562_));
  AN3        u0534(.A(j), .B(h), .C(g), .Y(men_men_n563_));
  NO2        u0535(.A(men_men_n140_), .B(c), .Y(men_men_n564_));
  NA3        u0536(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n447_), .Y(men_men_n565_));
  NA3        u0537(.A(f), .B(d), .C(b), .Y(men_men_n566_));
  INV        u0538(.A(men_men_n565_), .Y(men_men_n567_));
  NO4        u0539(.A(men_men_n567_), .B(men_men_n562_), .C(men_men_n552_), .D(men_men_n547_), .Y(men_men_n568_));
  AN3        u0540(.A(men_men_n568_), .B(men_men_n539_), .C(men_men_n519_), .Y(men_men_n569_));
  INV        u0541(.A(k), .Y(men_men_n570_));
  NA3        u0542(.A(l), .B(men_men_n570_), .C(i), .Y(men_men_n571_));
  INV        u0543(.A(men_men_n571_), .Y(men_men_n572_));
  NA4        u0544(.A(men_men_n386_), .B(men_men_n406_), .C(men_men_n175_), .D(men_men_n112_), .Y(men_men_n573_));
  NAi32      u0545(.An(h), .Bn(f), .C(g), .Y(men_men_n574_));
  NAi41      u0546(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n575_));
  OAI210     u0547(.A0(men_men_n523_), .A1(n), .B0(men_men_n575_), .Y(men_men_n576_));
  NA2        u0548(.A(men_men_n576_), .B(m), .Y(men_men_n577_));
  NAi31      u0549(.An(h), .B(g), .C(f), .Y(men_men_n578_));
  OR3        u0550(.A(men_men_n578_), .B(men_men_n265_), .C(men_men_n49_), .Y(men_men_n579_));
  NA4        u0551(.A(men_men_n406_), .B(men_men_n119_), .C(men_men_n112_), .D(e), .Y(men_men_n580_));
  AN2        u0552(.A(men_men_n580_), .B(men_men_n579_), .Y(men_men_n581_));
  NO3        u0553(.A(men_men_n574_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n582_));
  NO4        u0554(.A(men_men_n578_), .B(men_men_n532_), .C(men_men_n143_), .D(men_men_n75_), .Y(men_men_n583_));
  OR2        u0555(.A(men_men_n583_), .B(men_men_n582_), .Y(men_men_n584_));
  NAi31      u0556(.An(men_men_n584_), .B(men_men_n581_), .C(men_men_n573_), .Y(men_men_n585_));
  NAi31      u0557(.An(f), .B(h), .C(g), .Y(men_men_n586_));
  NO4        u0558(.A(men_men_n299_), .B(men_men_n586_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n587_));
  NOi32      u0559(.An(b), .Bn(a), .C(c), .Y(men_men_n588_));
  NOi41      u0560(.An(men_men_n588_), .B(men_men_n342_), .C(men_men_n69_), .D(men_men_n115_), .Y(men_men_n589_));
  OR2        u0561(.A(men_men_n589_), .B(men_men_n587_), .Y(men_men_n590_));
  NOi32      u0562(.An(d), .Bn(a), .C(e), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n112_), .Y(men_men_n592_));
  NO2        u0564(.A(n), .B(c), .Y(men_men_n593_));
  NA3        u0565(.A(men_men_n593_), .B(men_men_n29_), .C(m), .Y(men_men_n594_));
  NA2        u0566(.A(men_men_n594_), .B(men_men_n592_), .Y(men_men_n595_));
  NOi32      u0567(.An(e), .Bn(a), .C(d), .Y(men_men_n596_));
  AOI210     u0568(.A0(men_men_n29_), .A1(d), .B0(men_men_n596_), .Y(men_men_n597_));
  AOI210     u0569(.A0(men_men_n597_), .A1(men_men_n201_), .B0(men_men_n540_), .Y(men_men_n598_));
  AOI210     u0570(.A0(men_men_n598_), .A1(men_men_n595_), .B0(men_men_n590_), .Y(men_men_n599_));
  OAI210     u0571(.A0(men_men_n236_), .A1(men_men_n89_), .B0(men_men_n599_), .Y(men_men_n600_));
  AOI210     u0572(.A0(men_men_n585_), .A1(men_men_n572_), .B0(men_men_n600_), .Y(men_men_n601_));
  NO3        u0573(.A(men_men_n306_), .B(men_men_n61_), .C(n), .Y(men_men_n602_));
  NA3        u0574(.A(men_men_n500_), .B(men_men_n165_), .C(men_men_n164_), .Y(men_men_n603_));
  NA2        u0575(.A(men_men_n449_), .B(men_men_n218_), .Y(men_men_n604_));
  OR2        u0576(.A(men_men_n604_), .B(men_men_n603_), .Y(men_men_n605_));
  NA2        u0577(.A(men_men_n76_), .B(men_men_n112_), .Y(men_men_n606_));
  NO2        u0578(.A(men_men_n606_), .B(men_men_n45_), .Y(men_men_n607_));
  AOI220     u0579(.A0(men_men_n607_), .A1(men_men_n527_), .B0(men_men_n605_), .B1(men_men_n602_), .Y(men_men_n608_));
  NO2        u0580(.A(men_men_n608_), .B(men_men_n89_), .Y(men_men_n609_));
  NA3        u0581(.A(men_men_n542_), .B(men_men_n330_), .C(men_men_n46_), .Y(men_men_n610_));
  NOi32      u0582(.An(e), .Bn(c), .C(f), .Y(men_men_n611_));
  NOi21      u0583(.An(f), .B(g), .Y(men_men_n612_));
  NO2        u0584(.A(men_men_n612_), .B(men_men_n200_), .Y(men_men_n613_));
  AOI220     u0585(.A0(men_men_n613_), .A1(men_men_n383_), .B0(men_men_n611_), .B1(men_men_n169_), .Y(men_men_n614_));
  NA3        u0586(.A(men_men_n614_), .B(men_men_n610_), .C(men_men_n172_), .Y(men_men_n615_));
  AOI210     u0587(.A0(men_men_n526_), .A1(men_men_n387_), .B0(men_men_n290_), .Y(men_men_n616_));
  NA2        u0588(.A(men_men_n616_), .B(men_men_n252_), .Y(men_men_n617_));
  NOi21      u0589(.An(j), .B(l), .Y(men_men_n618_));
  NAi21      u0590(.An(k), .B(h), .Y(men_men_n619_));
  NO2        u0591(.A(men_men_n619_), .B(men_men_n250_), .Y(men_men_n620_));
  NA2        u0592(.A(men_men_n620_), .B(men_men_n618_), .Y(men_men_n621_));
  OR2        u0593(.A(men_men_n621_), .B(men_men_n577_), .Y(men_men_n622_));
  NOi31      u0594(.An(m), .B(n), .C(k), .Y(men_men_n623_));
  NA2        u0595(.A(men_men_n618_), .B(men_men_n623_), .Y(men_men_n624_));
  AOI210     u0596(.A0(men_men_n387_), .A1(men_men_n361_), .B0(men_men_n290_), .Y(men_men_n625_));
  NAi21      u0597(.An(men_men_n624_), .B(men_men_n625_), .Y(men_men_n626_));
  NO2        u0598(.A(men_men_n265_), .B(men_men_n49_), .Y(men_men_n627_));
  NO2        u0599(.A(men_men_n299_), .B(men_men_n586_), .Y(men_men_n628_));
  NO2        u0600(.A(men_men_n523_), .B(men_men_n49_), .Y(men_men_n629_));
  NA2        u0601(.A(men_men_n629_), .B(men_men_n628_), .Y(men_men_n630_));
  NA4        u0602(.A(men_men_n630_), .B(men_men_n626_), .C(men_men_n622_), .D(men_men_n617_), .Y(men_men_n631_));
  NA2        u0603(.A(men_men_n108_), .B(men_men_n36_), .Y(men_men_n632_));
  NO2        u0604(.A(k), .B(men_men_n202_), .Y(men_men_n633_));
  INV        u0605(.A(men_men_n350_), .Y(men_men_n634_));
  NO2        u0606(.A(men_men_n634_), .B(n), .Y(men_men_n635_));
  NAi31      u0607(.An(men_men_n632_), .B(men_men_n635_), .C(men_men_n633_), .Y(men_men_n636_));
  NO2        u0608(.A(men_men_n522_), .B(men_men_n170_), .Y(men_men_n637_));
  NA3        u0609(.A(men_men_n543_), .B(men_men_n259_), .C(men_men_n139_), .Y(men_men_n638_));
  NA2        u0610(.A(men_men_n496_), .B(men_men_n153_), .Y(men_men_n639_));
  NO3        u0611(.A(men_men_n384_), .B(men_men_n639_), .C(men_men_n89_), .Y(men_men_n640_));
  AOI210     u0612(.A0(men_men_n638_), .A1(men_men_n637_), .B0(men_men_n640_), .Y(men_men_n641_));
  AN3        u0613(.A(f), .B(d), .C(b), .Y(men_men_n642_));
  OAI210     u0614(.A0(men_men_n642_), .A1(men_men_n126_), .B0(n), .Y(men_men_n643_));
  NA3        u0615(.A(men_men_n496_), .B(men_men_n153_), .C(men_men_n202_), .Y(men_men_n644_));
  AOI210     u0616(.A0(men_men_n643_), .A1(men_men_n220_), .B0(men_men_n644_), .Y(men_men_n645_));
  NAi31      u0617(.An(m), .B(n), .C(k), .Y(men_men_n646_));
  OR2        u0618(.A(men_men_n130_), .B(men_men_n61_), .Y(men_men_n647_));
  OAI210     u0619(.A0(men_men_n647_), .A1(men_men_n646_), .B0(men_men_n238_), .Y(men_men_n648_));
  OAI210     u0620(.A0(men_men_n648_), .A1(men_men_n645_), .B0(j), .Y(men_men_n649_));
  NA3        u0621(.A(men_men_n649_), .B(men_men_n641_), .C(men_men_n636_), .Y(men_men_n650_));
  NO4        u0622(.A(men_men_n650_), .B(men_men_n631_), .C(men_men_n615_), .D(men_men_n609_), .Y(men_men_n651_));
  NA2        u0623(.A(men_men_n371_), .B(men_men_n156_), .Y(men_men_n652_));
  NAi31      u0624(.An(g), .B(h), .C(f), .Y(men_men_n653_));
  OR3        u0625(.A(men_men_n653_), .B(men_men_n265_), .C(n), .Y(men_men_n654_));
  OA210      u0626(.A0(men_men_n523_), .A1(n), .B0(men_men_n575_), .Y(men_men_n655_));
  NA3        u0627(.A(men_men_n404_), .B(men_men_n119_), .C(men_men_n86_), .Y(men_men_n656_));
  OAI210     u0628(.A0(men_men_n655_), .A1(men_men_n93_), .B0(men_men_n656_), .Y(men_men_n657_));
  NOi21      u0629(.An(men_men_n654_), .B(men_men_n657_), .Y(men_men_n658_));
  AOI210     u0630(.A0(men_men_n658_), .A1(men_men_n652_), .B0(men_men_n517_), .Y(men_men_n659_));
  NO3        u0631(.A(g), .B(men_men_n201_), .C(men_men_n56_), .Y(men_men_n660_));
  NO2        u0632(.A(men_men_n503_), .B(men_men_n89_), .Y(men_men_n661_));
  OAI210     u0633(.A0(men_men_n661_), .A1(men_men_n383_), .B0(men_men_n660_), .Y(men_men_n662_));
  OR2        u0634(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n663_));
  NA2        u0635(.A(men_men_n588_), .B(men_men_n332_), .Y(men_men_n664_));
  OA220      u0636(.A0(men_men_n624_), .A1(men_men_n664_), .B0(men_men_n621_), .B1(men_men_n663_), .Y(men_men_n665_));
  NA3        u0637(.A(men_men_n514_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n666_));
  AN2        u0638(.A(h), .B(f), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n667_), .B(men_men_n37_), .Y(men_men_n668_));
  NA2        u0640(.A(men_men_n101_), .B(men_men_n46_), .Y(men_men_n669_));
  OAI220     u0641(.A0(men_men_n669_), .A1(men_men_n321_), .B0(men_men_n668_), .B1(men_men_n453_), .Y(men_men_n670_));
  AOI210     u0642(.A0(men_men_n556_), .A1(men_men_n415_), .B0(men_men_n49_), .Y(men_men_n671_));
  OAI220     u0643(.A0(men_men_n578_), .A1(men_men_n571_), .B0(men_men_n314_), .B1(men_men_n515_), .Y(men_men_n672_));
  AOI210     u0644(.A0(men_men_n672_), .A1(men_men_n671_), .B0(men_men_n670_), .Y(men_men_n673_));
  NA4        u0645(.A(men_men_n673_), .B(men_men_n666_), .C(men_men_n665_), .D(men_men_n662_), .Y(men_men_n674_));
  NO2        u0646(.A(men_men_n240_), .B(f), .Y(men_men_n675_));
  NO2        u0647(.A(men_men_n612_), .B(men_men_n61_), .Y(men_men_n676_));
  NO3        u0648(.A(men_men_n676_), .B(men_men_n675_), .C(men_men_n34_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n317_), .B(men_men_n135_), .Y(men_men_n678_));
  NA2        u0650(.A(men_men_n128_), .B(men_men_n49_), .Y(men_men_n679_));
  AOI220     u0651(.A0(men_men_n679_), .A1(men_men_n520_), .B0(men_men_n350_), .B1(men_men_n112_), .Y(men_men_n680_));
  OA220      u0652(.A0(men_men_n680_), .A1(men_men_n540_), .B0(men_men_n349_), .B1(men_men_n110_), .Y(men_men_n681_));
  OAI210     u0653(.A0(men_men_n678_), .A1(men_men_n677_), .B0(men_men_n681_), .Y(men_men_n682_));
  NO3        u0654(.A(men_men_n392_), .B(men_men_n182_), .C(men_men_n181_), .Y(men_men_n683_));
  NA2        u0655(.A(men_men_n683_), .B(men_men_n218_), .Y(men_men_n684_));
  NA3        u0656(.A(men_men_n684_), .B(men_men_n242_), .C(j), .Y(men_men_n685_));
  NA2        u0657(.A(men_men_n452_), .B(men_men_n86_), .Y(men_men_n686_));
  NO4        u0658(.A(men_men_n517_), .B(men_men_n686_), .C(men_men_n127_), .D(men_men_n201_), .Y(men_men_n687_));
  INV        u0659(.A(men_men_n687_), .Y(men_men_n688_));
  NA3        u0660(.A(men_men_n688_), .B(men_men_n685_), .C(men_men_n390_), .Y(men_men_n689_));
  NO4        u0661(.A(men_men_n689_), .B(men_men_n682_), .C(men_men_n674_), .D(men_men_n659_), .Y(men_men_n690_));
  NA4        u0662(.A(men_men_n690_), .B(men_men_n651_), .C(men_men_n601_), .D(men_men_n569_), .Y(men08));
  NO2        u0663(.A(k), .B(h), .Y(men_men_n692_));
  AO210      u0664(.A0(men_men_n240_), .A1(men_men_n439_), .B0(men_men_n692_), .Y(men_men_n693_));
  NO2        u0665(.A(men_men_n693_), .B(men_men_n288_), .Y(men_men_n694_));
  NA2        u0666(.A(men_men_n611_), .B(men_men_n86_), .Y(men_men_n695_));
  NA2        u0667(.A(men_men_n695_), .B(men_men_n449_), .Y(men_men_n696_));
  NA2        u0668(.A(men_men_n696_), .B(men_men_n694_), .Y(men_men_n697_));
  NA2        u0669(.A(men_men_n86_), .B(men_men_n109_), .Y(men_men_n698_));
  NO2        u0670(.A(men_men_n698_), .B(men_men_n57_), .Y(men_men_n699_));
  NA2        u0671(.A(men_men_n566_), .B(men_men_n220_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n700_), .B(men_men_n338_), .Y(men_men_n701_));
  AOI210     u0673(.A0(men_men_n566_), .A1(men_men_n149_), .B0(men_men_n86_), .Y(men_men_n702_));
  NA4        u0674(.A(men_men_n204_), .B(men_men_n135_), .C(men_men_n45_), .D(h), .Y(men_men_n703_));
  AN2        u0675(.A(l), .B(k), .Y(men_men_n704_));
  NA4        u0676(.A(men_men_n704_), .B(men_men_n108_), .C(men_men_n75_), .D(men_men_n202_), .Y(men_men_n705_));
  OAI210     u0677(.A0(men_men_n703_), .A1(g), .B0(men_men_n705_), .Y(men_men_n706_));
  NA2        u0678(.A(men_men_n706_), .B(men_men_n702_), .Y(men_men_n707_));
  NA4        u0679(.A(men_men_n707_), .B(men_men_n701_), .C(men_men_n697_), .D(men_men_n340_), .Y(men_men_n708_));
  AN2        u0680(.A(men_men_n524_), .B(men_men_n97_), .Y(men_men_n709_));
  NO4        u0681(.A(men_men_n167_), .B(men_men_n382_), .C(men_men_n111_), .D(g), .Y(men_men_n710_));
  AOI210     u0682(.A0(men_men_n710_), .A1(men_men_n700_), .B0(men_men_n509_), .Y(men_men_n711_));
  NAi21      u0683(.An(men_men_n709_), .B(men_men_n711_), .Y(men_men_n712_));
  NO2        u0684(.A(men_men_n526_), .B(men_men_n35_), .Y(men_men_n713_));
  OAI210     u0685(.A0(men_men_n543_), .A1(men_men_n47_), .B0(men_men_n647_), .Y(men_men_n714_));
  NO2        u0686(.A(men_men_n472_), .B(men_men_n128_), .Y(men_men_n715_));
  AOI210     u0687(.A0(men_men_n715_), .A1(men_men_n714_), .B0(men_men_n713_), .Y(men_men_n716_));
  INV        u0688(.A(men_men_n705_), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n693_), .B(men_men_n131_), .Y(men_men_n718_));
  AOI220     u0690(.A0(men_men_n718_), .A1(men_men_n391_), .B0(men_men_n717_), .B1(men_men_n78_), .Y(men_men_n719_));
  OAI210     u0691(.A0(men_men_n716_), .A1(men_men_n89_), .B0(men_men_n719_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n350_), .B(men_men_n43_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n684_), .B(men_men_n323_), .C(men_men_n374_), .Y(men_men_n722_));
  NA2        u0694(.A(men_men_n704_), .B(men_men_n208_), .Y(men_men_n723_));
  NO2        u0695(.A(men_men_n723_), .B(men_men_n316_), .Y(men_men_n724_));
  AOI210     u0696(.A0(men_men_n724_), .A1(men_men_n675_), .B0(men_men_n479_), .Y(men_men_n725_));
  NA3        u0697(.A(m), .B(l), .C(k), .Y(men_men_n726_));
  AOI210     u0698(.A0(men_men_n656_), .A1(men_men_n654_), .B0(men_men_n726_), .Y(men_men_n727_));
  NO2        u0699(.A(men_men_n525_), .B(men_men_n260_), .Y(men_men_n728_));
  NOi21      u0700(.An(men_men_n728_), .B(men_men_n521_), .Y(men_men_n729_));
  NA4        u0701(.A(men_men_n112_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n730_));
  NA3        u0702(.A(men_men_n119_), .B(men_men_n400_), .C(i), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n731_), .B(men_men_n730_), .Y(men_men_n732_));
  NO3        u0704(.A(men_men_n732_), .B(men_men_n729_), .C(men_men_n727_), .Y(men_men_n733_));
  NA4        u0705(.A(men_men_n733_), .B(men_men_n725_), .C(men_men_n722_), .D(men_men_n721_), .Y(men_men_n734_));
  NO4        u0706(.A(men_men_n734_), .B(men_men_n720_), .C(men_men_n712_), .D(men_men_n708_), .Y(men_men_n735_));
  INV        u0707(.A(men_men_n490_), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n736_), .B(men_men_n239_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n704_), .B(men_men_n75_), .Y(men_men_n738_));
  NO4        u0710(.A(men_men_n683_), .B(men_men_n167_), .C(n), .D(i), .Y(men_men_n739_));
  NOi21      u0711(.An(h), .B(j), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n740_), .B(f), .Y(men_men_n741_));
  NO2        u0713(.A(men_men_n741_), .B(men_men_n233_), .Y(men_men_n742_));
  NO2        u0714(.A(men_men_n742_), .B(men_men_n739_), .Y(men_men_n743_));
  OAI220     u0715(.A0(men_men_n743_), .A1(men_men_n738_), .B0(men_men_n581_), .B1(men_men_n62_), .Y(men_men_n744_));
  AOI210     u0716(.A0(men_men_n737_), .A1(l), .B0(men_men_n744_), .Y(men_men_n745_));
  NO2        u0717(.A(j), .B(i), .Y(men_men_n746_));
  NA2        u0718(.A(men_men_n746_), .B(men_men_n33_), .Y(men_men_n747_));
  NA2        u0719(.A(men_men_n409_), .B(men_men_n119_), .Y(men_men_n748_));
  OR2        u0720(.A(men_men_n748_), .B(men_men_n747_), .Y(men_men_n749_));
  NO3        u0721(.A(men_men_n144_), .B(men_men_n49_), .C(men_men_n109_), .Y(men_men_n750_));
  NO3        u0722(.A(men_men_n532_), .B(men_men_n143_), .C(men_men_n75_), .Y(men_men_n751_));
  NO3        u0723(.A(men_men_n472_), .B(men_men_n427_), .C(j), .Y(men_men_n752_));
  OAI210     u0724(.A0(men_men_n751_), .A1(men_men_n750_), .B0(men_men_n752_), .Y(men_men_n753_));
  INV        u0725(.A(men_men_n753_), .Y(men_men_n754_));
  NA2        u0726(.A(k), .B(j), .Y(men_men_n755_));
  AOI210     u0727(.A0(men_men_n520_), .A1(n), .B0(men_men_n542_), .Y(men_men_n756_));
  NA2        u0728(.A(men_men_n756_), .B(men_men_n545_), .Y(men_men_n757_));
  NO3        u0729(.A(men_men_n167_), .B(men_men_n382_), .C(men_men_n111_), .Y(men_men_n758_));
  AOI220     u0730(.A0(men_men_n758_), .A1(men_men_n234_), .B0(men_men_n604_), .B1(men_men_n297_), .Y(men_men_n759_));
  INV        u0731(.A(men_men_n759_), .Y(men_men_n760_));
  NO2        u0732(.A(men_men_n288_), .B(men_men_n131_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n761_), .B(men_men_n613_), .Y(men_men_n762_));
  NO2        u0734(.A(men_men_n726_), .B(men_men_n93_), .Y(men_men_n763_));
  NA2        u0735(.A(men_men_n763_), .B(men_men_n576_), .Y(men_men_n764_));
  NO2        u0736(.A(men_men_n578_), .B(men_men_n115_), .Y(men_men_n765_));
  OAI210     u0737(.A0(men_men_n765_), .A1(men_men_n752_), .B0(men_men_n671_), .Y(men_men_n766_));
  NA3        u0738(.A(men_men_n766_), .B(men_men_n764_), .C(men_men_n762_), .Y(men_men_n767_));
  OR3        u0739(.A(men_men_n767_), .B(men_men_n760_), .C(men_men_n754_), .Y(men_men_n768_));
  NA3        u0740(.A(men_men_n756_), .B(men_men_n545_), .C(men_men_n544_), .Y(men_men_n769_));
  NA4        u0741(.A(men_men_n769_), .B(men_men_n204_), .C(men_men_n439_), .D(men_men_n34_), .Y(men_men_n770_));
  OAI220     u0742(.A0(men_men_n703_), .A1(men_men_n695_), .B0(men_men_n321_), .B1(men_men_n38_), .Y(men_men_n771_));
  INV        u0743(.A(men_men_n771_), .Y(men_men_n772_));
  NA3        u0744(.A(men_men_n535_), .B(men_men_n281_), .C(h), .Y(men_men_n773_));
  NOi21      u0745(.An(men_men_n671_), .B(men_men_n773_), .Y(men_men_n774_));
  NO2        u0746(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n775_));
  NO2        u0747(.A(men_men_n773_), .B(men_men_n594_), .Y(men_men_n776_));
  AOI210     u0748(.A0(men_men_n775_), .A1(men_men_n635_), .B0(men_men_n776_), .Y(men_men_n777_));
  NAi41      u0749(.An(men_men_n774_), .B(men_men_n777_), .C(men_men_n772_), .D(men_men_n770_), .Y(men_men_n778_));
  OR2        u0750(.A(men_men_n763_), .B(men_men_n97_), .Y(men_men_n779_));
  AOI220     u0751(.A0(men_men_n779_), .A1(men_men_n226_), .B0(men_men_n752_), .B1(men_men_n627_), .Y(men_men_n780_));
  INV        u0752(.A(men_men_n325_), .Y(men_men_n781_));
  OAI210     u0753(.A0(men_men_n726_), .A1(men_men_n653_), .B0(men_men_n508_), .Y(men_men_n782_));
  NA3        u0754(.A(men_men_n237_), .B(men_men_n59_), .C(b), .Y(men_men_n783_));
  AOI220     u0755(.A0(men_men_n593_), .A1(men_men_n29_), .B0(men_men_n452_), .B1(men_men_n86_), .Y(men_men_n784_));
  NA2        u0756(.A(men_men_n784_), .B(men_men_n783_), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n773_), .B(men_men_n478_), .Y(men_men_n786_));
  AOI210     u0758(.A0(men_men_n785_), .A1(men_men_n782_), .B0(men_men_n786_), .Y(men_men_n787_));
  NA3        u0759(.A(men_men_n787_), .B(men_men_n781_), .C(men_men_n780_), .Y(men_men_n788_));
  NOi41      u0760(.An(men_men_n749_), .B(men_men_n788_), .C(men_men_n778_), .D(men_men_n768_), .Y(men_men_n789_));
  OR3        u0761(.A(men_men_n703_), .B(men_men_n220_), .C(g), .Y(men_men_n790_));
  NO3        u0762(.A(men_men_n331_), .B(men_men_n290_), .C(men_men_n111_), .Y(men_men_n791_));
  NA2        u0763(.A(men_men_n791_), .B(men_men_n757_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n793_), .B(men_men_n747_), .C(men_men_n265_), .Y(men_men_n794_));
  INV        u0766(.A(men_men_n794_), .Y(men_men_n795_));
  NA4        u0767(.A(men_men_n795_), .B(men_men_n792_), .C(men_men_n790_), .D(men_men_n393_), .Y(men_men_n796_));
  OR2        u0768(.A(men_men_n653_), .B(men_men_n94_), .Y(men_men_n797_));
  NOi31      u0769(.An(b), .B(d), .C(a), .Y(men_men_n798_));
  NO2        u0770(.A(men_men_n798_), .B(men_men_n591_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n799_), .B(n), .Y(men_men_n800_));
  NOi21      u0772(.An(men_men_n784_), .B(men_men_n800_), .Y(men_men_n801_));
  OAI220     u0773(.A0(men_men_n801_), .A1(men_men_n797_), .B0(men_men_n773_), .B1(men_men_n592_), .Y(men_men_n802_));
  NO2        u0774(.A(men_men_n543_), .B(men_men_n86_), .Y(men_men_n803_));
  NO3        u0775(.A(men_men_n612_), .B(men_men_n316_), .C(men_men_n115_), .Y(men_men_n804_));
  NOi21      u0776(.An(men_men_n804_), .B(men_men_n154_), .Y(men_men_n805_));
  AOI210     u0777(.A0(men_men_n791_), .A1(men_men_n803_), .B0(men_men_n805_), .Y(men_men_n806_));
  OAI210     u0778(.A0(men_men_n703_), .A1(men_men_n384_), .B0(men_men_n806_), .Y(men_men_n807_));
  NO2        u0779(.A(men_men_n683_), .B(n), .Y(men_men_n808_));
  AOI220     u0780(.A0(men_men_n761_), .A1(men_men_n660_), .B0(men_men_n808_), .B1(men_men_n694_), .Y(men_men_n809_));
  NA2        u0781(.A(men_men_n119_), .B(men_men_n86_), .Y(men_men_n810_));
  AOI210     u0782(.A0(men_men_n413_), .A1(men_men_n405_), .B0(men_men_n810_), .Y(men_men_n811_));
  NA2        u0783(.A(men_men_n724_), .B(men_men_n34_), .Y(men_men_n812_));
  NAi21      u0784(.An(men_men_n730_), .B(men_men_n423_), .Y(men_men_n813_));
  NO2        u0785(.A(men_men_n260_), .B(i), .Y(men_men_n814_));
  NA2        u0786(.A(men_men_n710_), .B(men_men_n339_), .Y(men_men_n815_));
  OAI210     u0787(.A0(men_men_n583_), .A1(men_men_n582_), .B0(men_men_n351_), .Y(men_men_n816_));
  AN3        u0788(.A(men_men_n816_), .B(men_men_n815_), .C(men_men_n813_), .Y(men_men_n817_));
  NAi41      u0789(.An(men_men_n811_), .B(men_men_n817_), .C(men_men_n812_), .D(men_men_n809_), .Y(men_men_n818_));
  NO4        u0790(.A(men_men_n818_), .B(men_men_n807_), .C(men_men_n802_), .D(men_men_n796_), .Y(men_men_n819_));
  NA4        u0791(.A(men_men_n819_), .B(men_men_n789_), .C(men_men_n745_), .D(men_men_n735_), .Y(men09));
  INV        u0792(.A(men_men_n120_), .Y(men_men_n821_));
  NA2        u0793(.A(f), .B(e), .Y(men_men_n822_));
  NO2        u0794(.A(men_men_n213_), .B(men_men_n111_), .Y(men_men_n823_));
  NA2        u0795(.A(men_men_n823_), .B(g), .Y(men_men_n824_));
  NA4        u0796(.A(men_men_n299_), .B(men_men_n461_), .C(men_men_n249_), .D(men_men_n117_), .Y(men_men_n825_));
  AOI210     u0797(.A0(men_men_n825_), .A1(g), .B0(men_men_n458_), .Y(men_men_n826_));
  AOI210     u0798(.A0(men_men_n826_), .A1(men_men_n824_), .B0(men_men_n822_), .Y(men_men_n827_));
  NA2        u0799(.A(men_men_n433_), .B(e), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n828_), .B(men_men_n500_), .Y(men_men_n829_));
  AOI210     u0801(.A0(men_men_n827_), .A1(men_men_n821_), .B0(men_men_n829_), .Y(men_men_n830_));
  NO2        u0802(.A(men_men_n194_), .B(men_men_n201_), .Y(men_men_n831_));
  NA3        u0803(.A(m), .B(l), .C(i), .Y(men_men_n832_));
  OAI220     u0804(.A0(men_men_n578_), .A1(men_men_n832_), .B0(men_men_n342_), .B1(men_men_n516_), .Y(men_men_n833_));
  NA4        u0805(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n834_));
  NAi31      u0806(.An(men_men_n833_), .B(men_men_n834_), .C(men_men_n428_), .Y(men_men_n835_));
  OR2        u0807(.A(men_men_n835_), .B(men_men_n831_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n797_), .B(men_men_n555_), .C(men_men_n508_), .Y(men_men_n837_));
  OA210      u0809(.A0(men_men_n837_), .A1(men_men_n836_), .B0(men_men_n800_), .Y(men_men_n838_));
  INV        u0810(.A(men_men_n328_), .Y(men_men_n839_));
  NO2        u0811(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n840_));
  NOi31      u0812(.An(k), .B(m), .C(l), .Y(men_men_n841_));
  NO2        u0813(.A(men_men_n330_), .B(men_men_n841_), .Y(men_men_n842_));
  AOI210     u0814(.A0(men_men_n842_), .A1(men_men_n840_), .B0(men_men_n586_), .Y(men_men_n843_));
  NA2        u0815(.A(men_men_n783_), .B(men_men_n321_), .Y(men_men_n844_));
  NA2        u0816(.A(men_men_n332_), .B(men_men_n334_), .Y(men_men_n845_));
  OAI210     u0817(.A0(men_men_n194_), .A1(men_men_n201_), .B0(men_men_n845_), .Y(men_men_n846_));
  AOI220     u0818(.A0(men_men_n846_), .A1(men_men_n844_), .B0(men_men_n843_), .B1(men_men_n839_), .Y(men_men_n847_));
  NA2        u0819(.A(men_men_n161_), .B(men_men_n113_), .Y(men_men_n848_));
  NA3        u0820(.A(men_men_n848_), .B(men_men_n693_), .C(men_men_n131_), .Y(men_men_n849_));
  NA3        u0821(.A(men_men_n849_), .B(men_men_n180_), .C(men_men_n31_), .Y(men_men_n850_));
  NA4        u0822(.A(men_men_n850_), .B(men_men_n847_), .C(men_men_n614_), .D(men_men_n84_), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n574_), .B(men_men_n486_), .Y(men_men_n852_));
  NA2        u0824(.A(men_men_n852_), .B(men_men_n180_), .Y(men_men_n853_));
  NOi21      u0825(.An(f), .B(d), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n854_), .B(m), .Y(men_men_n855_));
  NO2        u0827(.A(men_men_n855_), .B(men_men_n52_), .Y(men_men_n856_));
  NOi32      u0828(.An(g), .Bn(f), .C(d), .Y(men_men_n857_));
  NA4        u0829(.A(men_men_n857_), .B(men_men_n593_), .C(men_men_n29_), .D(m), .Y(men_men_n858_));
  NOi21      u0830(.An(men_men_n300_), .B(men_men_n858_), .Y(men_men_n859_));
  AOI210     u0831(.A0(men_men_n856_), .A1(men_men_n533_), .B0(men_men_n859_), .Y(men_men_n860_));
  NA3        u0832(.A(men_men_n299_), .B(men_men_n249_), .C(men_men_n117_), .Y(men_men_n861_));
  AN2        u0833(.A(f), .B(d), .Y(men_men_n862_));
  NA3        u0834(.A(men_men_n465_), .B(men_men_n862_), .C(men_men_n86_), .Y(men_men_n863_));
  NO3        u0835(.A(men_men_n863_), .B(men_men_n75_), .C(men_men_n202_), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n274_), .B(men_men_n56_), .Y(men_men_n865_));
  NA2        u0837(.A(men_men_n861_), .B(men_men_n864_), .Y(men_men_n866_));
  NAi41      u0838(.An(men_men_n477_), .B(men_men_n866_), .C(men_men_n860_), .D(men_men_n853_), .Y(men_men_n867_));
  NO4        u0839(.A(men_men_n612_), .B(men_men_n128_), .C(men_men_n316_), .D(men_men_n145_), .Y(men_men_n868_));
  NO2        u0840(.A(men_men_n646_), .B(men_men_n316_), .Y(men_men_n869_));
  AN2        u0841(.A(men_men_n869_), .B(men_men_n675_), .Y(men_men_n870_));
  NO3        u0842(.A(men_men_n870_), .B(men_men_n868_), .C(men_men_n222_), .Y(men_men_n871_));
  NA2        u0843(.A(men_men_n591_), .B(men_men_n86_), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n863_), .B(men_men_n417_), .Y(men_men_n873_));
  NOi31      u0845(.An(men_men_n211_), .B(men_men_n873_), .C(men_men_n295_), .Y(men_men_n874_));
  NA2        u0846(.A(c), .B(men_men_n114_), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n875_), .B(men_men_n397_), .Y(men_men_n876_));
  NA3        u0848(.A(men_men_n876_), .B(men_men_n498_), .C(f), .Y(men_men_n877_));
  OR2        u0849(.A(men_men_n653_), .B(men_men_n529_), .Y(men_men_n878_));
  INV        u0850(.A(men_men_n878_), .Y(men_men_n879_));
  NA2        u0851(.A(men_men_n799_), .B(men_men_n110_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n880_), .B(men_men_n879_), .Y(men_men_n881_));
  NA4        u0853(.A(men_men_n881_), .B(men_men_n877_), .C(men_men_n874_), .D(men_men_n871_), .Y(men_men_n882_));
  NO4        u0854(.A(men_men_n882_), .B(men_men_n867_), .C(men_men_n851_), .D(men_men_n838_), .Y(men_men_n883_));
  OR2        u0855(.A(men_men_n863_), .B(men_men_n75_), .Y(men_men_n884_));
  NA2        u0856(.A(men_men_n111_), .B(j), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n823_), .B(g), .Y(men_men_n886_));
  AOI210     u0858(.A0(men_men_n886_), .A1(men_men_n282_), .B0(men_men_n884_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n321_), .B(men_men_n834_), .Y(men_men_n888_));
  NO2        u0860(.A(men_men_n218_), .B(men_men_n212_), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n889_), .B(men_men_n215_), .Y(men_men_n890_));
  NO2        u0862(.A(men_men_n417_), .B(men_men_n822_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n891_), .B(men_men_n550_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n892_), .B(men_men_n890_), .Y(men_men_n893_));
  NA2        u0865(.A(e), .B(d), .Y(men_men_n894_));
  OAI220     u0866(.A0(men_men_n894_), .A1(c), .B0(men_men_n311_), .B1(d), .Y(men_men_n895_));
  NA3        u0867(.A(men_men_n895_), .B(men_men_n442_), .C(men_men_n496_), .Y(men_men_n896_));
  AOI210     u0868(.A0(men_men_n503_), .A1(men_men_n174_), .B0(men_men_n218_), .Y(men_men_n897_));
  INV        u0869(.A(men_men_n897_), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n274_), .B(men_men_n159_), .Y(men_men_n899_));
  NA2        u0871(.A(men_men_n864_), .B(men_men_n899_), .Y(men_men_n900_));
  NA3        u0872(.A(men_men_n160_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n901_));
  NA4        u0873(.A(men_men_n901_), .B(men_men_n900_), .C(men_men_n898_), .D(men_men_n896_), .Y(men_men_n902_));
  NO4        u0874(.A(men_men_n902_), .B(men_men_n893_), .C(men_men_n888_), .D(men_men_n887_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n839_), .B(men_men_n31_), .Y(men_men_n904_));
  AO210      u0876(.A0(men_men_n904_), .A1(men_men_n695_), .B0(men_men_n205_), .Y(men_men_n905_));
  OAI220     u0877(.A0(men_men_n612_), .A1(men_men_n61_), .B0(men_men_n290_), .B1(j), .Y(men_men_n906_));
  AOI220     u0878(.A0(men_men_n906_), .A1(men_men_n869_), .B0(men_men_n602_), .B1(men_men_n611_), .Y(men_men_n907_));
  OAI210     u0879(.A0(men_men_n828_), .A1(men_men_n164_), .B0(men_men_n907_), .Y(men_men_n908_));
  OAI210     u0880(.A0(men_men_n823_), .A1(men_men_n899_), .B0(men_men_n857_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n909_), .B(men_men_n594_), .Y(men_men_n910_));
  AOI210     u0882(.A0(men_men_n116_), .A1(men_men_n115_), .B0(men_men_n248_), .Y(men_men_n911_));
  NO2        u0883(.A(men_men_n911_), .B(men_men_n858_), .Y(men_men_n912_));
  BUFFER     u0884(.A(men_men_n912_), .Y(men_men_n913_));
  NOi31      u0885(.An(men_men_n533_), .B(men_men_n855_), .C(men_men_n282_), .Y(men_men_n914_));
  NO4        u0886(.A(men_men_n914_), .B(men_men_n913_), .C(men_men_n910_), .D(men_men_n908_), .Y(men_men_n915_));
  AO220      u0887(.A0(men_men_n442_), .A1(men_men_n740_), .B0(men_men_n169_), .B1(f), .Y(men_men_n916_));
  OAI210     u0888(.A0(men_men_n916_), .A1(men_men_n445_), .B0(men_men_n895_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n427_), .B(men_men_n71_), .Y(men_men_n918_));
  OAI210     u0890(.A0(men_men_n837_), .A1(men_men_n918_), .B0(men_men_n699_), .Y(men_men_n919_));
  AN4        u0891(.A(men_men_n919_), .B(men_men_n917_), .C(men_men_n915_), .D(men_men_n905_), .Y(men_men_n920_));
  NA4        u0892(.A(men_men_n920_), .B(men_men_n903_), .C(men_men_n883_), .D(men_men_n830_), .Y(men12));
  NO2        u0893(.A(men_men_n440_), .B(c), .Y(men_men_n922_));
  NO4        u0894(.A(men_men_n432_), .B(men_men_n240_), .C(men_men_n570_), .D(men_men_n202_), .Y(men_men_n923_));
  NA2        u0895(.A(men_men_n923_), .B(men_men_n922_), .Y(men_men_n924_));
  NA2        u0896(.A(men_men_n533_), .B(men_men_n918_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n440_), .B(men_men_n114_), .Y(men_men_n926_));
  NO2        u0898(.A(men_men_n840_), .B(men_men_n342_), .Y(men_men_n927_));
  NO2        u0899(.A(men_men_n653_), .B(men_men_n368_), .Y(men_men_n928_));
  AOI220     u0900(.A0(men_men_n928_), .A1(men_men_n531_), .B0(men_men_n927_), .B1(men_men_n926_), .Y(men_men_n929_));
  NA4        u0901(.A(men_men_n929_), .B(men_men_n925_), .C(men_men_n924_), .D(men_men_n431_), .Y(men_men_n930_));
  AOI210     u0902(.A0(men_men_n221_), .A1(men_men_n327_), .B0(men_men_n191_), .Y(men_men_n931_));
  OR2        u0903(.A(men_men_n931_), .B(men_men_n923_), .Y(men_men_n932_));
  AOI210     u0904(.A0(men_men_n324_), .A1(men_men_n380_), .B0(men_men_n202_), .Y(men_men_n933_));
  OAI210     u0905(.A0(men_men_n933_), .A1(men_men_n932_), .B0(men_men_n392_), .Y(men_men_n934_));
  NO2        u0906(.A(men_men_n632_), .B(men_men_n250_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n578_), .B(men_men_n832_), .Y(men_men_n936_));
  NO2        u0908(.A(men_men_n144_), .B(men_men_n225_), .Y(men_men_n937_));
  NA3        u0909(.A(men_men_n937_), .B(men_men_n228_), .C(i), .Y(men_men_n938_));
  NA2        u0910(.A(men_men_n938_), .B(men_men_n934_), .Y(men_men_n939_));
  OR2        u0911(.A(men_men_n312_), .B(men_men_n926_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n940_), .B(men_men_n343_), .Y(men_men_n941_));
  NA4        u0913(.A(men_men_n433_), .B(men_men_n425_), .C(men_men_n175_), .D(g), .Y(men_men_n942_));
  NA2        u0914(.A(men_men_n942_), .B(men_men_n941_), .Y(men_men_n943_));
  NO3        u0915(.A(men_men_n658_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n944_));
  NO4        u0916(.A(men_men_n944_), .B(men_men_n943_), .C(men_men_n939_), .D(men_men_n930_), .Y(men_men_n945_));
  NO2        u0917(.A(men_men_n358_), .B(men_men_n357_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n575_), .B(men_men_n73_), .Y(men_men_n947_));
  NA2        u0919(.A(men_men_n543_), .B(men_men_n139_), .Y(men_men_n948_));
  NOi21      u0920(.An(men_men_n34_), .B(men_men_n646_), .Y(men_men_n949_));
  AOI220     u0921(.A0(men_men_n949_), .A1(men_men_n948_), .B0(men_men_n947_), .B1(men_men_n946_), .Y(men_men_n950_));
  OAI210     u0922(.A0(men_men_n238_), .A1(men_men_n45_), .B0(men_men_n950_), .Y(men_men_n951_));
  NA2        u0923(.A(men_men_n423_), .B(men_men_n252_), .Y(men_men_n952_));
  NO3        u0924(.A(men_men_n810_), .B(men_men_n91_), .C(men_men_n397_), .Y(men_men_n953_));
  NAi21      u0925(.An(men_men_n953_), .B(men_men_n952_), .Y(men_men_n954_));
  NO2        u0926(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n955_));
  NO2        u0927(.A(men_men_n493_), .B(men_men_n290_), .Y(men_men_n956_));
  INV        u0928(.A(men_men_n956_), .Y(men_men_n957_));
  NO2        u0929(.A(men_men_n957_), .B(men_men_n139_), .Y(men_men_n958_));
  NA2        u0930(.A(men_men_n623_), .B(men_men_n351_), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n731_), .A1(men_men_n959_), .B0(men_men_n355_), .Y(men_men_n960_));
  NO4        u0932(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n954_), .D(men_men_n951_), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n337_), .B(g), .Y(men_men_n962_));
  NA2        u0934(.A(men_men_n156_), .B(i), .Y(men_men_n963_));
  NA2        u0935(.A(men_men_n46_), .B(i), .Y(men_men_n964_));
  OAI220     u0936(.A0(men_men_n964_), .A1(men_men_n190_), .B0(men_men_n963_), .B1(men_men_n94_), .Y(men_men_n965_));
  AOI210     u0937(.A0(men_men_n407_), .A1(men_men_n37_), .B0(men_men_n965_), .Y(men_men_n966_));
  NO2        u0938(.A(men_men_n139_), .B(men_men_n86_), .Y(men_men_n967_));
  OR2        u0939(.A(men_men_n967_), .B(men_men_n542_), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n543_), .B(men_men_n372_), .Y(men_men_n969_));
  AOI210     u0941(.A0(men_men_n969_), .A1(n), .B0(men_men_n968_), .Y(men_men_n970_));
  OAI220     u0942(.A0(men_men_n970_), .A1(men_men_n962_), .B0(men_men_n966_), .B1(men_men_n321_), .Y(men_men_n971_));
  NO2        u0943(.A(men_men_n653_), .B(men_men_n486_), .Y(men_men_n972_));
  NA3        u0944(.A(men_men_n332_), .B(men_men_n618_), .C(i), .Y(men_men_n973_));
  OAI210     u0945(.A0(men_men_n427_), .A1(men_men_n299_), .B0(men_men_n973_), .Y(men_men_n974_));
  OAI220     u0946(.A0(men_men_n974_), .A1(men_men_n972_), .B0(men_men_n671_), .B1(men_men_n751_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n596_), .B(men_men_n112_), .Y(men_men_n976_));
  OR3        u0948(.A(men_men_n299_), .B(men_men_n422_), .C(f), .Y(men_men_n977_));
  NA3        u0949(.A(men_men_n618_), .B(men_men_n82_), .C(i), .Y(men_men_n978_));
  OA220      u0950(.A0(men_men_n978_), .A1(men_men_n976_), .B0(men_men_n977_), .B1(men_men_n577_), .Y(men_men_n979_));
  NA3        u0951(.A(men_men_n313_), .B(men_men_n116_), .C(g), .Y(men_men_n980_));
  AOI210     u0952(.A0(men_men_n668_), .A1(men_men_n980_), .B0(m), .Y(men_men_n981_));
  OAI210     u0953(.A0(men_men_n981_), .A1(men_men_n927_), .B0(men_men_n312_), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n686_), .B(men_men_n872_), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n834_), .B(men_men_n428_), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n209_), .B(men_men_n79_), .Y(men_men_n985_));
  NA3        u0957(.A(men_men_n985_), .B(men_men_n978_), .C(men_men_n977_), .Y(men_men_n986_));
  AOI220     u0958(.A0(men_men_n986_), .A1(men_men_n246_), .B0(men_men_n984_), .B1(men_men_n983_), .Y(men_men_n987_));
  NA4        u0959(.A(men_men_n987_), .B(men_men_n982_), .C(men_men_n979_), .D(men_men_n975_), .Y(men_men_n988_));
  NO2        u0960(.A(men_men_n368_), .B(men_men_n93_), .Y(men_men_n989_));
  OAI210     u0961(.A0(men_men_n989_), .A1(men_men_n935_), .B0(men_men_n226_), .Y(men_men_n990_));
  NA2        u0962(.A(men_men_n657_), .B(men_men_n90_), .Y(men_men_n991_));
  NO2        u0963(.A(men_men_n448_), .B(men_men_n202_), .Y(men_men_n992_));
  AOI220     u0964(.A0(men_men_n992_), .A1(men_men_n373_), .B0(men_men_n940_), .B1(men_men_n206_), .Y(men_men_n993_));
  AOI220     u0965(.A0(men_men_n928_), .A1(men_men_n937_), .B0(men_men_n576_), .B1(men_men_n92_), .Y(men_men_n994_));
  NA4        u0966(.A(men_men_n994_), .B(men_men_n993_), .C(men_men_n991_), .D(men_men_n990_), .Y(men_men_n995_));
  OAI210     u0967(.A0(men_men_n984_), .A1(men_men_n936_), .B0(men_men_n531_), .Y(men_men_n996_));
  AOI210     u0968(.A0(men_men_n408_), .A1(men_men_n401_), .B0(men_men_n810_), .Y(men_men_n997_));
  INV        u0969(.A(men_men_n997_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n981_), .B(men_men_n926_), .Y(men_men_n999_));
  NO3        u0971(.A(men_men_n885_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1000_));
  AOI220     u0972(.A0(men_men_n1000_), .A1(men_men_n616_), .B0(men_men_n637_), .B1(men_men_n520_), .Y(men_men_n1001_));
  NA4        u0973(.A(men_men_n1001_), .B(men_men_n999_), .C(men_men_n998_), .D(men_men_n996_), .Y(men_men_n1002_));
  NO4        u0974(.A(men_men_n1002_), .B(men_men_n995_), .C(men_men_n988_), .D(men_men_n971_), .Y(men_men_n1003_));
  NAi31      u0975(.An(men_men_n136_), .B(men_men_n409_), .C(n), .Y(men_men_n1004_));
  NO3        u0976(.A(men_men_n124_), .B(men_men_n330_), .C(men_men_n841_), .Y(men_men_n1005_));
  NO2        u0977(.A(men_men_n1005_), .B(men_men_n1004_), .Y(men_men_n1006_));
  NA2        u0978(.A(men_men_n218_), .B(men_men_n165_), .Y(men_men_n1007_));
  NO3        u0979(.A(men_men_n297_), .B(men_men_n433_), .C(men_men_n169_), .Y(men_men_n1008_));
  NOi31      u0980(.An(men_men_n1007_), .B(men_men_n1008_), .C(men_men_n202_), .Y(men_men_n1009_));
  NAi21      u0981(.An(men_men_n543_), .B(men_men_n992_), .Y(men_men_n1010_));
  NA2        u0982(.A(men_men_n426_), .B(men_men_n872_), .Y(men_men_n1011_));
  NO3        u0983(.A(men_men_n427_), .B(men_men_n299_), .C(men_men_n75_), .Y(men_men_n1012_));
  AOI220     u0984(.A0(men_men_n1012_), .A1(men_men_n1011_), .B0(men_men_n469_), .B1(g), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n1013_), .B(men_men_n1010_), .Y(men_men_n1014_));
  NO2        u0986(.A(men_men_n654_), .B(men_men_n368_), .Y(men_men_n1015_));
  NA2        u0987(.A(men_men_n931_), .B(men_men_n922_), .Y(men_men_n1016_));
  NO3        u0988(.A(men_men_n532_), .B(men_men_n143_), .C(men_men_n201_), .Y(men_men_n1017_));
  OAI210     u0989(.A0(men_men_n1017_), .A1(men_men_n514_), .B0(men_men_n369_), .Y(men_men_n1018_));
  OAI220     u0990(.A0(men_men_n928_), .A1(men_men_n936_), .B0(men_men_n533_), .B1(men_men_n416_), .Y(men_men_n1019_));
  NA4        u0991(.A(men_men_n1019_), .B(men_men_n1018_), .C(men_men_n1016_), .D(men_men_n610_), .Y(men_men_n1020_));
  OAI210     u0992(.A0(men_men_n931_), .A1(men_men_n923_), .B0(men_men_n1007_), .Y(men_men_n1021_));
  NA3        u0993(.A(men_men_n969_), .B(men_men_n474_), .C(men_men_n46_), .Y(men_men_n1022_));
  AOI210     u0994(.A0(men_men_n371_), .A1(men_men_n369_), .B0(men_men_n320_), .Y(men_men_n1023_));
  NA4        u0995(.A(men_men_n1023_), .B(men_men_n1022_), .C(men_men_n1021_), .D(men_men_n261_), .Y(men_men_n1024_));
  OR3        u0996(.A(men_men_n1024_), .B(men_men_n1020_), .C(men_men_n1015_), .Y(men_men_n1025_));
  NO4        u0997(.A(men_men_n1025_), .B(men_men_n1014_), .C(men_men_n1009_), .D(men_men_n1006_), .Y(men_men_n1026_));
  NA4        u0998(.A(men_men_n1026_), .B(men_men_n1003_), .C(men_men_n961_), .D(men_men_n945_), .Y(men13));
  AN2        u0999(.A(c), .B(b), .Y(men_men_n1028_));
  NA3        u1000(.A(men_men_n237_), .B(men_men_n1028_), .C(m), .Y(men_men_n1029_));
  NA2        u1001(.A(men_men_n484_), .B(f), .Y(men_men_n1030_));
  NO4        u1002(.A(men_men_n1030_), .B(men_men_n1029_), .C(j), .D(men_men_n571_), .Y(men_men_n1031_));
  NA2        u1003(.A(men_men_n252_), .B(men_men_n1028_), .Y(men_men_n1032_));
  NO4        u1004(.A(men_men_n1032_), .B(men_men_n1030_), .C(men_men_n963_), .D(a), .Y(men_men_n1033_));
  NAi32      u1005(.An(d), .Bn(c), .C(e), .Y(men_men_n1034_));
  NA2        u1006(.A(men_men_n135_), .B(men_men_n45_), .Y(men_men_n1035_));
  NO4        u1007(.A(men_men_n1035_), .B(men_men_n1034_), .C(men_men_n578_), .D(men_men_n296_), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n400_), .B(men_men_n201_), .Y(men_men_n1037_));
  AN2        u1009(.A(d), .B(c), .Y(men_men_n1038_));
  NA2        u1010(.A(men_men_n1038_), .B(men_men_n114_), .Y(men_men_n1039_));
  NO4        u1011(.A(men_men_n1039_), .B(men_men_n1037_), .C(men_men_n170_), .D(men_men_n161_), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n484_), .B(c), .Y(men_men_n1041_));
  NO4        u1013(.A(men_men_n1035_), .B(men_men_n574_), .C(men_men_n1041_), .D(men_men_n296_), .Y(men_men_n1042_));
  OR2        u1014(.A(men_men_n1040_), .B(men_men_n1042_), .Y(men_men_n1043_));
  OR4        u1015(.A(men_men_n1043_), .B(men_men_n1036_), .C(men_men_n1033_), .D(men_men_n1031_), .Y(men_men_n1044_));
  NAi32      u1016(.An(f), .Bn(e), .C(c), .Y(men_men_n1045_));
  NO2        u1017(.A(men_men_n1045_), .B(men_men_n140_), .Y(men_men_n1046_));
  NA2        u1018(.A(men_men_n1046_), .B(g), .Y(men_men_n1047_));
  OR3        u1019(.A(men_men_n212_), .B(men_men_n170_), .C(men_men_n161_), .Y(men_men_n1048_));
  NO2        u1020(.A(men_men_n1048_), .B(men_men_n1047_), .Y(men_men_n1049_));
  NO2        u1021(.A(men_men_n1041_), .B(men_men_n296_), .Y(men_men_n1050_));
  NA2        u1022(.A(men_men_n620_), .B(men_men_n1512_), .Y(men_men_n1051_));
  NOi21      u1023(.An(men_men_n1050_), .B(men_men_n1051_), .Y(men_men_n1052_));
  NO2        u1024(.A(men_men_n755_), .B(men_men_n111_), .Y(men_men_n1053_));
  NOi41      u1025(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1054_));
  NA2        u1026(.A(men_men_n1054_), .B(men_men_n1053_), .Y(men_men_n1055_));
  NO2        u1027(.A(men_men_n1055_), .B(men_men_n1047_), .Y(men_men_n1056_));
  NA3        u1028(.A(k), .B(j), .C(i), .Y(men_men_n1057_));
  NO3        u1029(.A(men_men_n1057_), .B(men_men_n296_), .C(men_men_n93_), .Y(men_men_n1058_));
  OR3        u1030(.A(men_men_n1056_), .B(men_men_n1052_), .C(men_men_n1049_), .Y(men_men_n1059_));
  NO2        u1031(.A(f), .B(c), .Y(men_men_n1060_));
  NOi21      u1032(.An(men_men_n1060_), .B(men_men_n432_), .Y(men_men_n1061_));
  OR2        u1033(.A(men_men_n1059_), .B(men_men_n1044_), .Y(men02));
  OR3        u1034(.A(n), .B(m), .C(i), .Y(men_men_n1063_));
  NOi31      u1035(.An(e), .B(d), .C(c), .Y(men_men_n1064_));
  AOI210     u1036(.A0(men_men_n1058_), .A1(men_men_n1064_), .B0(men_men_n1036_), .Y(men_men_n1065_));
  AN3        u1037(.A(g), .B(f), .C(c), .Y(men_men_n1066_));
  NA3        u1038(.A(men_men_n1066_), .B(men_men_n455_), .C(h), .Y(men_men_n1067_));
  OR2        u1039(.A(men_men_n1057_), .B(men_men_n296_), .Y(men_men_n1068_));
  OR2        u1040(.A(men_men_n1068_), .B(men_men_n1067_), .Y(men_men_n1069_));
  INV        u1041(.A(men_men_n1049_), .Y(men_men_n1070_));
  NA3        u1042(.A(l), .B(k), .C(j), .Y(men_men_n1071_));
  NA2        u1043(.A(i), .B(h), .Y(men_men_n1072_));
  NO3        u1044(.A(men_men_n1072_), .B(men_men_n1071_), .C(men_men_n128_), .Y(men_men_n1073_));
  NO3        u1045(.A(men_men_n137_), .B(men_men_n272_), .C(men_men_n202_), .Y(men_men_n1074_));
  AOI210     u1046(.A0(men_men_n1074_), .A1(men_men_n1073_), .B0(men_men_n1052_), .Y(men_men_n1075_));
  NA3        u1047(.A(c), .B(b), .C(a), .Y(men_men_n1076_));
  NO3        u1048(.A(men_men_n1076_), .B(men_men_n894_), .C(men_men_n201_), .Y(men_men_n1077_));
  NO3        u1049(.A(men_men_n1057_), .B(men_men_n49_), .C(men_men_n111_), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n1078_), .B(men_men_n1077_), .Y(men_men_n1079_));
  AN4        u1051(.A(men_men_n1079_), .B(men_men_n1075_), .C(men_men_n1070_), .D(men_men_n1069_), .Y(men_men_n1080_));
  NO2        u1052(.A(men_men_n1039_), .B(men_men_n1037_), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n1055_), .B(men_men_n1048_), .Y(men_men_n1082_));
  AOI210     u1054(.A0(men_men_n1082_), .A1(men_men_n1081_), .B0(men_men_n1031_), .Y(men_men_n1083_));
  NA3        u1055(.A(men_men_n1083_), .B(men_men_n1080_), .C(men_men_n1065_), .Y(men03));
  NA4        u1056(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n201_), .Y(men_men_n1085_));
  NA4        u1057(.A(men_men_n563_), .B(m), .C(men_men_n111_), .D(men_men_n201_), .Y(men_men_n1086_));
  NA3        u1058(.A(men_men_n1086_), .B(men_men_n359_), .C(men_men_n1085_), .Y(men_men_n1087_));
  INV        u1059(.A(men_men_n1087_), .Y(men_men_n1088_));
  NOi31      u1060(.An(men_men_n797_), .B(men_men_n846_), .C(men_men_n835_), .Y(men_men_n1089_));
  OAI220     u1061(.A0(men_men_n1089_), .A1(men_men_n686_), .B0(men_men_n1088_), .B1(men_men_n575_), .Y(men_men_n1090_));
  NOi31      u1062(.An(i), .B(k), .C(j), .Y(men_men_n1091_));
  NA4        u1063(.A(men_men_n1091_), .B(men_men_n1064_), .C(men_men_n332_), .D(men_men_n323_), .Y(men_men_n1092_));
  OAI210     u1064(.A0(men_men_n810_), .A1(men_men_n410_), .B0(men_men_n1092_), .Y(men_men_n1093_));
  NOi31      u1065(.An(m), .B(n), .C(f), .Y(men_men_n1094_));
  NA2        u1066(.A(men_men_n1094_), .B(men_men_n51_), .Y(men_men_n1095_));
  AN2        u1067(.A(e), .B(c), .Y(men_men_n1096_));
  NA2        u1068(.A(men_men_n1096_), .B(a), .Y(men_men_n1097_));
  OAI220     u1069(.A0(men_men_n1097_), .A1(men_men_n1095_), .B0(men_men_n878_), .B1(men_men_n415_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n496_), .B(l), .Y(men_men_n1099_));
  NOi31      u1071(.An(men_men_n857_), .B(men_men_n1029_), .C(men_men_n1099_), .Y(men_men_n1100_));
  NO4        u1072(.A(men_men_n1100_), .B(men_men_n1098_), .C(men_men_n1093_), .D(men_men_n997_), .Y(men_men_n1101_));
  NO2        u1073(.A(men_men_n272_), .B(a), .Y(men_men_n1102_));
  INV        u1074(.A(men_men_n1036_), .Y(men_men_n1103_));
  NO2        u1075(.A(men_men_n89_), .B(g), .Y(men_men_n1104_));
  NA2        u1076(.A(men_men_n1103_), .B(men_men_n1101_), .Y(men_men_n1105_));
  NO4        u1077(.A(men_men_n1105_), .B(men_men_n1090_), .C(men_men_n811_), .D(men_men_n552_), .Y(men_men_n1106_));
  NA2        u1078(.A(c), .B(b), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n698_), .B(men_men_n1107_), .Y(men_men_n1108_));
  OAI210     u1080(.A0(men_men_n855_), .A1(men_men_n826_), .B0(men_men_n403_), .Y(men_men_n1109_));
  OAI210     u1081(.A0(men_men_n1109_), .A1(men_men_n856_), .B0(men_men_n1108_), .Y(men_men_n1110_));
  NAi21      u1082(.An(men_men_n411_), .B(men_men_n1108_), .Y(men_men_n1111_));
  NA3        u1083(.A(men_men_n416_), .B(men_men_n548_), .C(f), .Y(men_men_n1112_));
  OAI210     u1084(.A0(men_men_n537_), .A1(men_men_n39_), .B0(men_men_n1102_), .Y(men_men_n1113_));
  NA3        u1085(.A(men_men_n1113_), .B(men_men_n1112_), .C(men_men_n1111_), .Y(men_men_n1114_));
  NA2        u1086(.A(men_men_n249_), .B(men_men_n117_), .Y(men_men_n1115_));
  OAI210     u1087(.A0(men_men_n1115_), .A1(men_men_n276_), .B0(g), .Y(men_men_n1116_));
  NAi21      u1088(.An(f), .B(d), .Y(men_men_n1117_));
  NO2        u1089(.A(men_men_n1117_), .B(men_men_n1076_), .Y(men_men_n1118_));
  INV        u1090(.A(men_men_n1118_), .Y(men_men_n1119_));
  AOI210     u1091(.A0(men_men_n1116_), .A1(men_men_n282_), .B0(men_men_n1119_), .Y(men_men_n1120_));
  AOI210     u1092(.A0(men_men_n1120_), .A1(men_men_n112_), .B0(men_men_n1114_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n458_), .B(men_men_n457_), .Y(men_men_n1122_));
  NO2        u1094(.A(men_men_n176_), .B(men_men_n225_), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n1123_), .B(m), .Y(men_men_n1124_));
  NA3        u1096(.A(men_men_n911_), .B(men_men_n1099_), .C(men_men_n461_), .Y(men_men_n1125_));
  OAI210     u1097(.A0(men_men_n1125_), .A1(men_men_n300_), .B0(men_men_n459_), .Y(men_men_n1126_));
  AOI210     u1098(.A0(men_men_n1126_), .A1(men_men_n1122_), .B0(men_men_n1124_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n550_), .B(men_men_n399_), .Y(men_men_n1128_));
  NA2        u1100(.A(men_men_n152_), .B(men_men_n33_), .Y(men_men_n1129_));
  AOI210     u1101(.A0(men_men_n959_), .A1(men_men_n1129_), .B0(men_men_n202_), .Y(men_men_n1130_));
  OAI210     u1102(.A0(men_men_n1130_), .A1(men_men_n436_), .B0(men_men_n1118_), .Y(men_men_n1131_));
  NO2        u1103(.A(men_men_n362_), .B(men_men_n361_), .Y(men_men_n1132_));
  AOI210     u1104(.A0(men_men_n1123_), .A1(men_men_n418_), .B0(men_men_n953_), .Y(men_men_n1133_));
  NAi41      u1105(.An(men_men_n1132_), .B(men_men_n1133_), .C(men_men_n1131_), .D(men_men_n1128_), .Y(men_men_n1134_));
  NO2        u1106(.A(men_men_n1134_), .B(men_men_n1127_), .Y(men_men_n1135_));
  NA4        u1107(.A(men_men_n1135_), .B(men_men_n1121_), .C(men_men_n1110_), .D(men_men_n1106_), .Y(men00));
  AOI210     u1108(.A0(men_men_n289_), .A1(men_men_n202_), .B0(men_men_n264_), .Y(men_men_n1137_));
  NO2        u1109(.A(men_men_n1137_), .B(men_men_n566_), .Y(men_men_n1138_));
  AOI210     u1110(.A0(men_men_n891_), .A1(men_men_n937_), .B0(men_men_n1093_), .Y(men_men_n1139_));
  NO2        u1111(.A(men_men_n953_), .B(men_men_n709_), .Y(men_men_n1140_));
  NA3        u1112(.A(men_men_n1140_), .B(men_men_n1139_), .C(men_men_n998_), .Y(men_men_n1141_));
  NA2        u1113(.A(men_men_n498_), .B(f), .Y(men_men_n1142_));
  OAI210     u1114(.A0(men_men_n1005_), .A1(men_men_n40_), .B0(men_men_n639_), .Y(men_men_n1143_));
  NA3        u1115(.A(men_men_n1143_), .B(men_men_n245_), .C(n), .Y(men_men_n1144_));
  AOI210     u1116(.A0(men_men_n1144_), .A1(men_men_n1142_), .B0(men_men_n1039_), .Y(men_men_n1145_));
  NO4        u1117(.A(men_men_n1145_), .B(men_men_n1141_), .C(men_men_n1138_), .D(men_men_n1059_), .Y(men_men_n1146_));
  NA3        u1118(.A(men_men_n160_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1147_));
  NA3        u1119(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1148_));
  NOi31      u1120(.An(n), .B(m), .C(i), .Y(men_men_n1149_));
  NA3        u1121(.A(men_men_n1149_), .B(men_men_n642_), .C(men_men_n51_), .Y(men_men_n1150_));
  OAI210     u1122(.A0(men_men_n1148_), .A1(men_men_n1147_), .B0(men_men_n1150_), .Y(men_men_n1151_));
  INV        u1123(.A(men_men_n565_), .Y(men_men_n1152_));
  NO4        u1124(.A(men_men_n1152_), .B(men_men_n1151_), .C(men_men_n1132_), .D(men_men_n914_), .Y(men_men_n1153_));
  NO4        u1125(.A(men_men_n475_), .B(men_men_n345_), .C(men_men_n1107_), .D(men_men_n59_), .Y(men_men_n1154_));
  NA3        u1126(.A(men_men_n374_), .B(men_men_n208_), .C(g), .Y(men_men_n1155_));
  OA220      u1127(.A0(men_men_n1155_), .A1(men_men_n1148_), .B0(men_men_n375_), .B1(men_men_n130_), .Y(men_men_n1156_));
  NO2        u1128(.A(h), .B(g), .Y(men_men_n1157_));
  NA4        u1129(.A(men_men_n487_), .B(men_men_n455_), .C(men_men_n1157_), .D(men_men_n1028_), .Y(men_men_n1158_));
  AOI220     u1130(.A0(men_men_n307_), .A1(men_men_n234_), .B0(men_men_n171_), .B1(men_men_n142_), .Y(men_men_n1159_));
  NA3        u1131(.A(men_men_n1159_), .B(men_men_n1158_), .C(men_men_n1156_), .Y(men_men_n1160_));
  NO3        u1132(.A(men_men_n1160_), .B(men_men_n1154_), .C(men_men_n254_), .Y(men_men_n1161_));
  INV        u1133(.A(men_men_n310_), .Y(men_men_n1162_));
  NA2        u1134(.A(men_men_n234_), .B(men_men_n337_), .Y(men_men_n1163_));
  NA3        u1135(.A(men_men_n1163_), .B(men_men_n1162_), .C(men_men_n147_), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n227_), .B(men_men_n175_), .Y(men_men_n1165_));
  NA2        u1137(.A(men_men_n1165_), .B(men_men_n416_), .Y(men_men_n1166_));
  NA3        u1138(.A(men_men_n173_), .B(men_men_n111_), .C(g), .Y(men_men_n1167_));
  NA2        u1139(.A(men_men_n455_), .B(f), .Y(men_men_n1168_));
  NOi31      u1140(.An(men_men_n865_), .B(men_men_n1168_), .C(men_men_n1167_), .Y(men_men_n1169_));
  NAi31      u1141(.An(men_men_n178_), .B(men_men_n852_), .C(men_men_n455_), .Y(men_men_n1170_));
  NAi31      u1142(.An(men_men_n1169_), .B(men_men_n1170_), .C(men_men_n1166_), .Y(men_men_n1171_));
  NO2        u1143(.A(men_men_n263_), .B(men_men_n75_), .Y(men_men_n1172_));
  NO3        u1144(.A(men_men_n415_), .B(men_men_n822_), .C(n), .Y(men_men_n1173_));
  NA2        u1145(.A(men_men_n1173_), .B(men_men_n1172_), .Y(men_men_n1174_));
  NAi31      u1146(.An(men_men_n1042_), .B(men_men_n1174_), .C(men_men_n74_), .Y(men_men_n1175_));
  NO4        u1147(.A(men_men_n1175_), .B(men_men_n1171_), .C(men_men_n1164_), .D(men_men_n507_), .Y(men_men_n1176_));
  AN3        u1148(.A(men_men_n1176_), .B(men_men_n1161_), .C(men_men_n1153_), .Y(men_men_n1177_));
  NA3        u1149(.A(men_men_n1094_), .B(men_men_n596_), .C(men_men_n454_), .Y(men_men_n1178_));
  NA3        u1150(.A(men_men_n1178_), .B(men_men_n551_), .C(men_men_n230_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n1087_), .B(men_men_n524_), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n1180_), .B(men_men_n286_), .Y(men_men_n1181_));
  OAI210     u1153(.A0(men_men_n453_), .A1(men_men_n118_), .B0(men_men_n858_), .Y(men_men_n1182_));
  AOI220     u1154(.A0(men_men_n1182_), .A1(men_men_n1125_), .B0(men_men_n550_), .B1(men_men_n399_), .Y(men_men_n1183_));
  OR4        u1155(.A(men_men_n1039_), .B(men_men_n260_), .C(men_men_n210_), .D(e), .Y(men_men_n1184_));
  NO2        u1156(.A(men_men_n205_), .B(men_men_n202_), .Y(men_men_n1185_));
  NA2        u1157(.A(n), .B(e), .Y(men_men_n1186_));
  NO2        u1158(.A(men_men_n1186_), .B(men_men_n140_), .Y(men_men_n1187_));
  AOI220     u1159(.A0(men_men_n1187_), .A1(men_men_n262_), .B0(men_men_n839_), .B1(men_men_n1185_), .Y(men_men_n1188_));
  OAI210     u1160(.A0(men_men_n346_), .A1(men_men_n301_), .B0(men_men_n438_), .Y(men_men_n1189_));
  NA4        u1161(.A(men_men_n1189_), .B(men_men_n1188_), .C(men_men_n1184_), .D(men_men_n1183_), .Y(men_men_n1190_));
  AOI210     u1162(.A0(men_men_n1187_), .A1(men_men_n843_), .B0(men_men_n811_), .Y(men_men_n1191_));
  NO2        u1163(.A(men_men_n68_), .B(h), .Y(men_men_n1192_));
  NO3        u1164(.A(men_men_n1039_), .B(men_men_n1037_), .C(men_men_n723_), .Y(men_men_n1193_));
  INV        u1165(.A(men_men_n128_), .Y(men_men_n1194_));
  AN2        u1166(.A(men_men_n1194_), .B(men_men_n1074_), .Y(men_men_n1195_));
  OAI210     u1167(.A0(men_men_n1195_), .A1(men_men_n1193_), .B0(men_men_n1192_), .Y(men_men_n1196_));
  NA3        u1168(.A(men_men_n1196_), .B(men_men_n1191_), .C(men_men_n860_), .Y(men_men_n1197_));
  NO4        u1169(.A(men_men_n1197_), .B(men_men_n1190_), .C(men_men_n1181_), .D(men_men_n1179_), .Y(men_men_n1198_));
  NA2        u1170(.A(men_men_n827_), .B(men_men_n750_), .Y(men_men_n1199_));
  NA4        u1171(.A(men_men_n1199_), .B(men_men_n1198_), .C(men_men_n1177_), .D(men_men_n1146_), .Y(men01));
  AN2        u1172(.A(men_men_n1018_), .B(men_men_n1016_), .Y(men_men_n1201_));
  NO3        u1173(.A(men_men_n794_), .B(men_men_n786_), .C(men_men_n270_), .Y(men_men_n1202_));
  NA2        u1174(.A(men_men_n385_), .B(i), .Y(men_men_n1203_));
  NA3        u1175(.A(men_men_n1203_), .B(men_men_n1202_), .C(men_men_n1201_), .Y(men_men_n1204_));
  NA2        u1176(.A(men_men_n576_), .B(men_men_n92_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n543_), .B(men_men_n259_), .Y(men_men_n1206_));
  NA2        u1178(.A(men_men_n956_), .B(men_men_n1206_), .Y(men_men_n1207_));
  NA4        u1179(.A(men_men_n1207_), .B(men_men_n1205_), .C(men_men_n907_), .D(men_men_n322_), .Y(men_men_n1208_));
  NA2        u1180(.A(men_men_n45_), .B(f), .Y(men_men_n1209_));
  NA2        u1181(.A(men_men_n704_), .B(men_men_n98_), .Y(men_men_n1210_));
  NO2        u1182(.A(men_men_n1210_), .B(men_men_n1209_), .Y(men_men_n1211_));
  NO2        u1183(.A(men_men_n773_), .B(men_men_n592_), .Y(men_men_n1212_));
  AOI210     u1184(.A0(men_men_n1211_), .A1(men_men_n627_), .B0(men_men_n1212_), .Y(men_men_n1213_));
  INV        u1185(.A(men_men_n116_), .Y(men_men_n1214_));
  OA220      u1186(.A0(men_men_n1214_), .A1(men_men_n573_), .B0(men_men_n655_), .B1(men_men_n359_), .Y(men_men_n1215_));
  NAi41      u1187(.An(men_men_n155_), .B(men_men_n1215_), .C(men_men_n1213_), .D(men_men_n890_), .Y(men_men_n1216_));
  NO3        u1188(.A(men_men_n774_), .B(men_men_n670_), .C(men_men_n501_), .Y(men_men_n1217_));
  NA4        u1189(.A(men_men_n704_), .B(men_men_n98_), .C(men_men_n45_), .D(men_men_n201_), .Y(men_men_n1218_));
  OA220      u1190(.A0(men_men_n1218_), .A1(men_men_n663_), .B0(men_men_n185_), .B1(men_men_n183_), .Y(men_men_n1219_));
  NA3        u1191(.A(men_men_n1219_), .B(men_men_n1217_), .C(men_men_n133_), .Y(men_men_n1220_));
  NO4        u1192(.A(men_men_n1220_), .B(men_men_n1216_), .C(men_men_n1208_), .D(men_men_n1204_), .Y(men_men_n1221_));
  INV        u1193(.A(men_men_n1155_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n1222_), .B(men_men_n520_), .Y(men_men_n1223_));
  AOI210     u1195(.A0(men_men_n194_), .A1(men_men_n91_), .B0(men_men_n201_), .Y(men_men_n1224_));
  OAI210     u1196(.A0(men_men_n800_), .A1(men_men_n416_), .B0(men_men_n1224_), .Y(men_men_n1225_));
  NA2        u1197(.A(men_men_n193_), .B(men_men_n34_), .Y(men_men_n1226_));
  OR2        u1198(.A(men_men_n1226_), .B(men_men_n321_), .Y(men_men_n1227_));
  NA3        u1199(.A(men_men_n1227_), .B(men_men_n1225_), .C(men_men_n1223_), .Y(men_men_n1228_));
  AOI210     u1200(.A0(men_men_n584_), .A1(men_men_n116_), .B0(men_men_n590_), .Y(men_men_n1229_));
  OAI210     u1201(.A0(men_men_n1214_), .A1(men_men_n581_), .B0(men_men_n1229_), .Y(men_men_n1230_));
  NA2        u1202(.A(men_men_n269_), .B(men_men_n185_), .Y(men_men_n1231_));
  NA2        u1203(.A(men_men_n1231_), .B(men_men_n660_), .Y(men_men_n1232_));
  NO3        u1204(.A(men_men_n810_), .B(men_men_n194_), .C(men_men_n397_), .Y(men_men_n1233_));
  NO2        u1205(.A(men_men_n1233_), .B(men_men_n953_), .Y(men_men_n1234_));
  OAI210     u1206(.A0(men_men_n1211_), .A1(men_men_n315_), .B0(men_men_n671_), .Y(men_men_n1235_));
  NA4        u1207(.A(men_men_n1235_), .B(men_men_n1234_), .C(men_men_n1232_), .D(men_men_n777_), .Y(men_men_n1236_));
  NO3        u1208(.A(men_men_n1236_), .B(men_men_n1230_), .C(men_men_n1228_), .Y(men_men_n1237_));
  NA3        u1209(.A(men_men_n593_), .B(men_men_n29_), .C(f), .Y(men_men_n1238_));
  NO2        u1210(.A(men_men_n1238_), .B(men_men_n194_), .Y(men_men_n1239_));
  AOI210     u1211(.A0(men_men_n494_), .A1(men_men_n58_), .B0(men_men_n1239_), .Y(men_men_n1240_));
  OR3        u1212(.A(men_men_n1210_), .B(men_men_n594_), .C(men_men_n1209_), .Y(men_men_n1241_));
  NO2        u1213(.A(men_men_n1218_), .B(men_men_n976_), .Y(men_men_n1242_));
  NO2        u1214(.A(men_men_n1242_), .B(men_men_n1151_), .Y(men_men_n1243_));
  NA4        u1215(.A(men_men_n1243_), .B(men_men_n1241_), .C(men_men_n1240_), .D(men_men_n749_), .Y(men_men_n1244_));
  NO2        u1216(.A(men_men_n963_), .B(men_men_n220_), .Y(men_men_n1245_));
  NO2        u1217(.A(men_men_n964_), .B(men_men_n545_), .Y(men_men_n1246_));
  OAI210     u1218(.A0(men_men_n1246_), .A1(men_men_n1245_), .B0(men_men_n330_), .Y(men_men_n1247_));
  NA2        u1219(.A(men_men_n559_), .B(men_men_n557_), .Y(men_men_n1248_));
  NO3        u1220(.A(men_men_n81_), .B(men_men_n290_), .C(men_men_n45_), .Y(men_men_n1249_));
  NA2        u1221(.A(men_men_n1249_), .B(men_men_n542_), .Y(men_men_n1250_));
  NA3        u1222(.A(men_men_n1250_), .B(men_men_n1248_), .C(men_men_n665_), .Y(men_men_n1251_));
  OR2        u1223(.A(men_men_n1155_), .B(men_men_n1148_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n359_), .B(men_men_n73_), .Y(men_men_n1253_));
  INV        u1225(.A(men_men_n1253_), .Y(men_men_n1254_));
  NA2        u1226(.A(men_men_n1249_), .B(men_men_n803_), .Y(men_men_n1255_));
  NA4        u1227(.A(men_men_n1255_), .B(men_men_n1254_), .C(men_men_n1252_), .D(men_men_n377_), .Y(men_men_n1256_));
  NOi41      u1228(.An(men_men_n1247_), .B(men_men_n1256_), .C(men_men_n1251_), .D(men_men_n1244_), .Y(men_men_n1257_));
  INV        u1229(.A(men_men_n130_), .Y(men_men_n1258_));
  NO3        u1230(.A(men_men_n1072_), .B(men_men_n170_), .C(men_men_n89_), .Y(men_men_n1259_));
  AOI220     u1231(.A0(men_men_n1259_), .A1(men_men_n1258_), .B0(men_men_n1249_), .B1(men_men_n967_), .Y(men_men_n1260_));
  INV        u1232(.A(men_men_n1260_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n604_), .B(men_men_n603_), .Y(men_men_n1262_));
  NO4        u1234(.A(men_men_n1072_), .B(men_men_n1262_), .C(men_men_n168_), .D(men_men_n89_), .Y(men_men_n1263_));
  NO3        u1235(.A(men_men_n1263_), .B(men_men_n1261_), .C(men_men_n631_), .Y(men_men_n1264_));
  NA4        u1236(.A(men_men_n1264_), .B(men_men_n1257_), .C(men_men_n1237_), .D(men_men_n1221_), .Y(men06));
  NO2        u1237(.A(men_men_n398_), .B(men_men_n549_), .Y(men_men_n1266_));
  INV        u1238(.A(men_men_n730_), .Y(men_men_n1267_));
  OAI210     u1239(.A0(men_men_n1267_), .A1(men_men_n255_), .B0(men_men_n1266_), .Y(men_men_n1268_));
  NO2        u1240(.A(men_men_n212_), .B(men_men_n103_), .Y(men_men_n1269_));
  OAI210     u1241(.A0(men_men_n1269_), .A1(men_men_n1259_), .B0(men_men_n373_), .Y(men_men_n1270_));
  NO3        u1242(.A(men_men_n588_), .B(men_men_n798_), .C(men_men_n591_), .Y(men_men_n1271_));
  OR2        u1243(.A(men_men_n1271_), .B(men_men_n878_), .Y(men_men_n1272_));
  NA4        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n1268_), .D(men_men_n1247_), .Y(men_men_n1273_));
  NO3        u1245(.A(men_men_n1273_), .B(men_men_n1251_), .C(men_men_n244_), .Y(men_men_n1274_));
  NO2        u1246(.A(men_men_n290_), .B(men_men_n45_), .Y(men_men_n1275_));
  AOI210     u1247(.A0(men_men_n1275_), .A1(men_men_n968_), .B0(men_men_n1245_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n1275_), .B(men_men_n546_), .Y(men_men_n1277_));
  AOI210     u1249(.A0(men_men_n1277_), .A1(men_men_n1276_), .B0(men_men_n327_), .Y(men_men_n1278_));
  INV        u1250(.A(men_men_n669_), .Y(men_men_n1279_));
  NA2        u1251(.A(men_men_n1279_), .B(men_men_n635_), .Y(men_men_n1280_));
  NO2        u1252(.A(men_men_n503_), .B(men_men_n165_), .Y(men_men_n1281_));
  NOi21      u1253(.An(men_men_n132_), .B(men_men_n45_), .Y(men_men_n1282_));
  NO2        u1254(.A(men_men_n597_), .B(men_men_n1095_), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n449_), .B(men_men_n235_), .Y(men_men_n1284_));
  NO4        u1256(.A(men_men_n1284_), .B(men_men_n1283_), .C(men_men_n1282_), .D(men_men_n1281_), .Y(men_men_n1285_));
  OR2        u1257(.A(men_men_n589_), .B(men_men_n587_), .Y(men_men_n1286_));
  NO2        u1258(.A(men_men_n358_), .B(men_men_n131_), .Y(men_men_n1287_));
  AOI210     u1259(.A0(men_men_n1287_), .A1(men_men_n576_), .B0(men_men_n1286_), .Y(men_men_n1288_));
  NA3        u1260(.A(men_men_n1288_), .B(men_men_n1285_), .C(men_men_n1280_), .Y(men_men_n1289_));
  NO2        u1261(.A(men_men_n741_), .B(men_men_n357_), .Y(men_men_n1290_));
  NO3        u1262(.A(men_men_n671_), .B(men_men_n751_), .C(men_men_n627_), .Y(men_men_n1291_));
  NOi21      u1263(.An(men_men_n1290_), .B(men_men_n1291_), .Y(men_men_n1292_));
  AN2        u1264(.A(men_men_n949_), .B(men_men_n638_), .Y(men_men_n1293_));
  NO4        u1265(.A(men_men_n1293_), .B(men_men_n1292_), .C(men_men_n1289_), .D(men_men_n1278_), .Y(men_men_n1294_));
  NO2        u1266(.A(men_men_n793_), .B(men_men_n265_), .Y(men_men_n1295_));
  OAI220     u1267(.A0(men_men_n730_), .A1(men_men_n47_), .B0(men_men_n212_), .B1(men_men_n606_), .Y(men_men_n1296_));
  OAI210     u1268(.A0(men_men_n265_), .A1(c), .B0(men_men_n634_), .Y(men_men_n1297_));
  AOI220     u1269(.A0(men_men_n1297_), .A1(men_men_n1296_), .B0(men_men_n1295_), .B1(men_men_n255_), .Y(men_men_n1298_));
  NO3        u1270(.A(men_men_n232_), .B(men_men_n103_), .C(men_men_n272_), .Y(men_men_n1299_));
  OAI220     u1271(.A0(men_men_n695_), .A1(men_men_n235_), .B0(men_men_n500_), .B1(men_men_n503_), .Y(men_men_n1300_));
  NO3        u1272(.A(men_men_n1300_), .B(men_men_n1299_), .C(men_men_n1098_), .Y(men_men_n1301_));
  NA4        u1273(.A(men_men_n784_), .B(men_men_n783_), .C(men_men_n426_), .D(men_men_n872_), .Y(men_men_n1302_));
  NAi31      u1274(.An(men_men_n741_), .B(men_men_n1302_), .C(men_men_n193_), .Y(men_men_n1303_));
  NA3        u1275(.A(men_men_n1303_), .B(men_men_n1301_), .C(men_men_n1298_), .Y(men_men_n1304_));
  NOi31      u1276(.An(men_men_n1271_), .B(men_men_n452_), .C(men_men_n386_), .Y(men_men_n1305_));
  OR3        u1277(.A(men_men_n1305_), .B(men_men_n773_), .C(men_men_n529_), .Y(men_men_n1306_));
  OR3        u1278(.A(men_men_n361_), .B(men_men_n212_), .C(men_men_n606_), .Y(men_men_n1307_));
  AOI210     u1279(.A0(men_men_n559_), .A1(men_men_n438_), .B0(men_men_n363_), .Y(men_men_n1308_));
  NA3        u1280(.A(men_men_n1308_), .B(men_men_n1307_), .C(men_men_n1306_), .Y(men_men_n1309_));
  AOI220     u1281(.A0(men_men_n1290_), .A1(men_men_n750_), .B0(men_men_n1287_), .B1(men_men_n226_), .Y(men_men_n1310_));
  AN2        u1282(.A(men_men_n923_), .B(men_men_n922_), .Y(men_men_n1311_));
  NO4        u1283(.A(men_men_n1311_), .B(men_men_n870_), .C(men_men_n490_), .D(men_men_n469_), .Y(men_men_n1312_));
  NA3        u1284(.A(men_men_n1312_), .B(men_men_n1310_), .C(men_men_n1255_), .Y(men_men_n1313_));
  NAi21      u1285(.An(j), .B(i), .Y(men_men_n1314_));
  NO4        u1286(.A(men_men_n1262_), .B(men_men_n1314_), .C(men_men_n432_), .D(men_men_n223_), .Y(men_men_n1315_));
  NO4        u1287(.A(men_men_n1315_), .B(men_men_n1313_), .C(men_men_n1309_), .D(men_men_n1304_), .Y(men_men_n1316_));
  NA4        u1288(.A(men_men_n1316_), .B(men_men_n1294_), .C(men_men_n1274_), .D(men_men_n1264_), .Y(men07));
  NAi32      u1289(.An(m), .Bn(b), .C(n), .Y(men_men_n1318_));
  NO3        u1290(.A(men_men_n1318_), .B(g), .C(f), .Y(men_men_n1319_));
  OAI210     u1291(.A0(men_men_n309_), .A1(men_men_n471_), .B0(men_men_n1319_), .Y(men_men_n1320_));
  NAi21      u1292(.An(f), .B(c), .Y(men_men_n1321_));
  OR2        u1293(.A(e), .B(d), .Y(men_men_n1322_));
  OAI220     u1294(.A0(men_men_n1322_), .A1(men_men_n1321_), .B0(men_men_n619_), .B1(men_men_n311_), .Y(men_men_n1323_));
  NA3        u1295(.A(men_men_n1323_), .B(men_men_n1512_), .C(men_men_n173_), .Y(men_men_n1324_));
  NOi31      u1296(.An(n), .B(m), .C(b), .Y(men_men_n1325_));
  NO3        u1297(.A(men_men_n128_), .B(men_men_n439_), .C(h), .Y(men_men_n1326_));
  NA2        u1298(.A(men_men_n1324_), .B(men_men_n1320_), .Y(men_men_n1327_));
  NOi41      u1299(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1328_));
  NA3        u1300(.A(men_men_n1328_), .B(men_men_n862_), .C(men_men_n400_), .Y(men_men_n1329_));
  NO2        u1301(.A(men_men_n1329_), .B(men_men_n56_), .Y(men_men_n1330_));
  NA2        u1302(.A(men_men_n1074_), .B(men_men_n208_), .Y(men_men_n1331_));
  NO2        u1303(.A(men_men_n1331_), .B(men_men_n61_), .Y(men_men_n1332_));
  NO2        u1304(.A(k), .B(i), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n1045_), .B(men_men_n432_), .Y(men_men_n1335_));
  NA3        u1307(.A(men_men_n1335_), .B(men_men_n1334_), .C(men_men_n202_), .Y(men_men_n1336_));
  NO2        u1308(.A(men_men_n1057_), .B(men_men_n296_), .Y(men_men_n1337_));
  NA2        u1309(.A(men_men_n1192_), .B(men_men_n280_), .Y(men_men_n1338_));
  NA2        u1310(.A(men_men_n1338_), .B(men_men_n1336_), .Y(men_men_n1339_));
  NO4        u1311(.A(men_men_n1339_), .B(men_men_n1332_), .C(men_men_n1330_), .D(men_men_n1327_), .Y(men_men_n1340_));
  NO3        u1312(.A(e), .B(d), .C(c), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n128_), .B(men_men_n202_), .Y(men_men_n1342_));
  NA2        u1314(.A(men_men_n1342_), .B(men_men_n1341_), .Y(men_men_n1343_));
  NO2        u1315(.A(men_men_n1343_), .B(c), .Y(men_men_n1344_));
  OR2        u1316(.A(h), .B(f), .Y(men_men_n1345_));
  NO3        u1317(.A(n), .B(m), .C(i), .Y(men_men_n1346_));
  OAI210     u1318(.A0(men_men_n1096_), .A1(men_men_n150_), .B0(men_men_n1346_), .Y(men_men_n1347_));
  NO2        u1319(.A(i), .B(g), .Y(men_men_n1348_));
  OR3        u1320(.A(men_men_n1348_), .B(men_men_n1318_), .C(men_men_n72_), .Y(men_men_n1349_));
  OAI220     u1321(.A0(men_men_n1349_), .A1(men_men_n471_), .B0(men_men_n1347_), .B1(men_men_n1345_), .Y(men_men_n1350_));
  NA3        u1322(.A(men_men_n692_), .B(men_men_n679_), .C(men_men_n111_), .Y(men_men_n1351_));
  NA3        u1323(.A(men_men_n1325_), .B(men_men_n1053_), .C(men_men_n667_), .Y(men_men_n1352_));
  AOI210     u1324(.A0(men_men_n1352_), .A1(men_men_n1351_), .B0(men_men_n45_), .Y(men_men_n1353_));
  NO2        u1325(.A(l), .B(k), .Y(men_men_n1354_));
  NOi41      u1326(.An(men_men_n535_), .B(men_men_n1354_), .C(men_men_n466_), .D(men_men_n432_), .Y(men_men_n1355_));
  NO3        u1327(.A(men_men_n432_), .B(d), .C(c), .Y(men_men_n1356_));
  NO4        u1328(.A(men_men_n1355_), .B(men_men_n1353_), .C(men_men_n1350_), .D(men_men_n1344_), .Y(men_men_n1357_));
  NO2        u1329(.A(men_men_n141_), .B(h), .Y(men_men_n1358_));
  NO2        u1330(.A(g), .B(c), .Y(men_men_n1359_));
  NO2        u1331(.A(men_men_n440_), .B(a), .Y(men_men_n1360_));
  NA3        u1332(.A(men_men_n1360_), .B(k), .C(men_men_n112_), .Y(men_men_n1361_));
  NO2        u1333(.A(i), .B(h), .Y(men_men_n1362_));
  NA2        u1334(.A(men_men_n1362_), .B(men_men_n208_), .Y(men_men_n1363_));
  AOI210     u1335(.A0(men_men_n1117_), .A1(h), .B0(men_men_n404_), .Y(men_men_n1364_));
  NA2        u1336(.A(men_men_n134_), .B(men_men_n208_), .Y(men_men_n1365_));
  AOI210     u1337(.A0(men_men_n245_), .A1(men_men_n114_), .B0(men_men_n520_), .Y(men_men_n1366_));
  OAI220     u1338(.A0(men_men_n1366_), .A1(men_men_n1363_), .B0(men_men_n1365_), .B1(men_men_n1364_), .Y(men_men_n1367_));
  NO2        u1339(.A(men_men_n747_), .B(men_men_n179_), .Y(men_men_n1368_));
  NOi31      u1340(.An(m), .B(n), .C(b), .Y(men_men_n1369_));
  NOi31      u1341(.An(f), .B(d), .C(c), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n1370_), .B(men_men_n1369_), .Y(men_men_n1371_));
  INV        u1343(.A(men_men_n1371_), .Y(men_men_n1372_));
  NO3        u1344(.A(men_men_n1372_), .B(men_men_n1368_), .C(men_men_n1367_), .Y(men_men_n1373_));
  NA2        u1345(.A(men_men_n1066_), .B(men_men_n455_), .Y(men_men_n1374_));
  NO4        u1346(.A(men_men_n1374_), .B(men_men_n1053_), .C(men_men_n432_), .D(men_men_n45_), .Y(men_men_n1375_));
  OAI210     u1347(.A0(men_men_n176_), .A1(men_men_n515_), .B0(men_men_n1054_), .Y(men_men_n1376_));
  NO3        u1348(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1377_));
  INV        u1349(.A(men_men_n1376_), .Y(men_men_n1378_));
  NO2        u1350(.A(men_men_n1378_), .B(men_men_n1375_), .Y(men_men_n1379_));
  AN3        u1351(.A(men_men_n1379_), .B(men_men_n1373_), .C(men_men_n1361_), .Y(men_men_n1380_));
  NA2        u1352(.A(men_men_n1325_), .B(men_men_n370_), .Y(men_men_n1381_));
  NA2        u1353(.A(men_men_n1356_), .B(men_men_n203_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n179_), .B(b), .Y(men_men_n1383_));
  AOI220     u1355(.A0(men_men_n1149_), .A1(men_men_n1383_), .B0(men_men_n1073_), .B1(men_men_n1374_), .Y(men_men_n1384_));
  NO2        u1356(.A(i), .B(men_men_n201_), .Y(men_men_n1385_));
  NA4        u1357(.A(men_men_n1123_), .B(men_men_n1385_), .C(men_men_n104_), .D(m), .Y(men_men_n1386_));
  NA3        u1358(.A(men_men_n1386_), .B(men_men_n1384_), .C(men_men_n1382_), .Y(men_men_n1387_));
  NO4        u1359(.A(men_men_n128_), .B(g), .C(f), .D(e), .Y(men_men_n1388_));
  NA3        u1360(.A(men_men_n1333_), .B(men_men_n281_), .C(h), .Y(men_men_n1389_));
  NA2        u1361(.A(men_men_n30_), .B(h), .Y(men_men_n1390_));
  NO2        u1362(.A(men_men_n1390_), .B(men_men_n1063_), .Y(men_men_n1391_));
  NOi41      u1363(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1392_));
  NA2        u1364(.A(men_men_n1392_), .B(men_men_n112_), .Y(men_men_n1393_));
  NA2        u1365(.A(men_men_n1328_), .B(men_men_n1354_), .Y(men_men_n1394_));
  NA2        u1366(.A(men_men_n1394_), .B(men_men_n1393_), .Y(men_men_n1395_));
  OR3        u1367(.A(men_men_n529_), .B(men_men_n528_), .C(men_men_n111_), .Y(men_men_n1396_));
  NA2        u1368(.A(men_men_n1094_), .B(men_men_n397_), .Y(men_men_n1397_));
  OAI220     u1369(.A0(men_men_n1397_), .A1(men_men_n425_), .B0(men_men_n1396_), .B1(men_men_n290_), .Y(men_men_n1398_));
  AO210      u1370(.A0(men_men_n1398_), .A1(men_men_n114_), .B0(men_men_n1395_), .Y(men_men_n1399_));
  NO3        u1371(.A(men_men_n1399_), .B(men_men_n1391_), .C(men_men_n1387_), .Y(men_men_n1400_));
  NA4        u1372(.A(men_men_n1400_), .B(men_men_n1380_), .C(men_men_n1357_), .D(men_men_n1340_), .Y(men_men_n1401_));
  NO2        u1373(.A(men_men_n382_), .B(j), .Y(men_men_n1402_));
  NA3        u1374(.A(men_men_n1377_), .B(men_men_n1322_), .C(men_men_n1094_), .Y(men_men_n1403_));
  NA2        u1375(.A(men_men_n1061_), .B(e), .Y(men_men_n1404_));
  NA2        u1376(.A(men_men_n1404_), .B(men_men_n1403_), .Y(men_men_n1405_));
  NA3        u1377(.A(g), .B(men_men_n1402_), .C(men_men_n152_), .Y(men_men_n1406_));
  INV        u1378(.A(men_men_n1406_), .Y(men_men_n1407_));
  NO3        u1379(.A(men_men_n741_), .B(men_men_n168_), .C(men_men_n400_), .Y(men_men_n1408_));
  NO3        u1380(.A(men_men_n1408_), .B(men_men_n1407_), .C(men_men_n1405_), .Y(men_men_n1409_));
  NO3        u1381(.A(men_men_n1063_), .B(men_men_n570_), .C(g), .Y(men_men_n1410_));
  INV        u1382(.A(men_men_n1410_), .Y(men_men_n1411_));
  NO2        u1383(.A(men_men_n1411_), .B(men_men_n1045_), .Y(men_men_n1412_));
  OR2        u1384(.A(n), .B(i), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n1413_), .B(men_men_n49_), .Y(men_men_n1414_));
  AOI220     u1386(.A0(men_men_n1414_), .A1(men_men_n1157_), .B0(men_men_n814_), .B1(men_men_n184_), .Y(men_men_n1415_));
  INV        u1387(.A(men_men_n1415_), .Y(men_men_n1416_));
  NO2        u1388(.A(men_men_n212_), .B(k), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n1416_), .B(men_men_n1412_), .Y(men_men_n1418_));
  INV        u1390(.A(men_men_n49_), .Y(men_men_n1419_));
  NO3        u1391(.A(men_men_n1076_), .B(men_men_n1322_), .C(men_men_n49_), .Y(men_men_n1420_));
  NA2        u1392(.A(men_men_n1077_), .B(men_men_n1419_), .Y(men_men_n1421_));
  NO2        u1393(.A(men_men_n1063_), .B(h), .Y(men_men_n1422_));
  NA2        u1394(.A(men_men_n1422_), .B(d), .Y(men_men_n1423_));
  OAI220     u1395(.A0(men_men_n1423_), .A1(c), .B0(men_men_n1421_), .B1(j), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n173_), .B(men_men_n111_), .Y(men_men_n1425_));
  AOI210     u1397(.A0(men_men_n515_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1426_));
  NA2        u1398(.A(men_men_n1426_), .B(men_men_n1360_), .Y(men_men_n1427_));
  NO2        u1399(.A(men_men_n1314_), .B(men_men_n168_), .Y(men_men_n1428_));
  NOi21      u1400(.An(d), .B(f), .Y(men_men_n1429_));
  NO2        u1401(.A(men_men_n1322_), .B(f), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n290_), .B(c), .Y(men_men_n1431_));
  NA2        u1403(.A(men_men_n1431_), .B(men_men_n530_), .Y(men_men_n1432_));
  NA2        u1404(.A(men_men_n1432_), .B(men_men_n1427_), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n1433_), .B(men_men_n1424_), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1434_), .B(men_men_n1418_), .C(men_men_n1409_), .Y(men_men_n1435_));
  NO2        u1407(.A(men_men_n1066_), .B(men_men_n40_), .Y(men_men_n1436_));
  NO2        u1408(.A(men_men_n455_), .B(men_men_n290_), .Y(men_men_n1437_));
  OAI210     u1409(.A0(men_men_n1437_), .A1(men_men_n1436_), .B0(men_men_n1337_), .Y(men_men_n1438_));
  OAI210     u1410(.A0(men_men_n1388_), .A1(men_men_n1325_), .B0(men_men_n875_), .Y(men_men_n1439_));
  NO2        u1411(.A(men_men_n1034_), .B(men_men_n128_), .Y(men_men_n1440_));
  NA2        u1412(.A(men_men_n1440_), .B(men_men_n612_), .Y(men_men_n1441_));
  NA3        u1413(.A(men_men_n1441_), .B(men_men_n1439_), .C(men_men_n1438_), .Y(men_men_n1442_));
  NA2        u1414(.A(men_men_n1359_), .B(men_men_n1429_), .Y(men_men_n1443_));
  NO2        u1415(.A(men_men_n1443_), .B(m), .Y(men_men_n1444_));
  NA3        u1416(.A(men_men_n1074_), .B(men_men_n108_), .C(men_men_n208_), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n144_), .B(men_men_n175_), .Y(men_men_n1446_));
  OAI210     u1418(.A0(men_men_n1446_), .A1(men_men_n109_), .B0(men_men_n1369_), .Y(men_men_n1447_));
  NA2        u1419(.A(men_men_n1447_), .B(men_men_n1445_), .Y(men_men_n1448_));
  NO3        u1420(.A(men_men_n1448_), .B(men_men_n1444_), .C(men_men_n1442_), .Y(men_men_n1449_));
  NO2        u1421(.A(men_men_n1321_), .B(e), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1450_), .B(men_men_n395_), .Y(men_men_n1451_));
  OAI210     u1423(.A0(men_men_n1430_), .A1(men_men_n1104_), .B0(men_men_n623_), .Y(men_men_n1452_));
  OR3        u1424(.A(men_men_n1417_), .B(men_men_n1192_), .C(men_men_n128_), .Y(men_men_n1453_));
  OAI220     u1425(.A0(men_men_n1453_), .A1(men_men_n1451_), .B0(men_men_n1452_), .B1(men_men_n434_), .Y(men_men_n1454_));
  NO3        u1426(.A(men_men_n1396_), .B(men_men_n342_), .C(a), .Y(men_men_n1455_));
  NO2        u1427(.A(men_men_n1455_), .B(men_men_n1454_), .Y(men_men_n1456_));
  NA2        u1428(.A(men_men_n1450_), .B(men_men_n173_), .Y(men_men_n1457_));
  AOI210     u1429(.A0(men_men_n522_), .A1(men_men_n357_), .B0(men_men_n1457_), .Y(men_men_n1458_));
  NA2        u1430(.A(men_men_n528_), .B(g), .Y(men_men_n1459_));
  AOI210     u1431(.A0(men_men_n1459_), .A1(men_men_n1356_), .B0(men_men_n1420_), .Y(men_men_n1460_));
  NA2        u1432(.A(men_men_n1104_), .B(a), .Y(men_men_n1461_));
  OAI210     u1433(.A0(men_men_n1461_), .A1(men_men_n69_), .B0(men_men_n1460_), .Y(men_men_n1462_));
  OR2        u1434(.A(h), .B(men_men_n528_), .Y(men_men_n1463_));
  NO2        u1435(.A(men_men_n1463_), .B(men_men_n168_), .Y(men_men_n1464_));
  NA4        u1436(.A(men_men_n1074_), .B(men_men_n1071_), .C(men_men_n208_), .D(men_men_n68_), .Y(men_men_n1465_));
  NA2        u1437(.A(men_men_n1326_), .B(men_men_n176_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n49_), .B(l), .Y(men_men_n1467_));
  INV        u1439(.A(men_men_n471_), .Y(men_men_n1468_));
  OAI210     u1440(.A0(men_men_n1468_), .A1(men_men_n1077_), .B0(men_men_n1467_), .Y(men_men_n1469_));
  NO2        u1441(.A(m), .B(i), .Y(men_men_n1470_));
  BUFFER     u1442(.A(men_men_n1470_), .Y(men_men_n1471_));
  NA2        u1443(.A(men_men_n1471_), .B(men_men_n1358_), .Y(men_men_n1472_));
  NA4        u1444(.A(men_men_n1472_), .B(men_men_n1469_), .C(men_men_n1466_), .D(men_men_n1465_), .Y(men_men_n1473_));
  NO4        u1445(.A(men_men_n1473_), .B(men_men_n1464_), .C(men_men_n1462_), .D(men_men_n1458_), .Y(men_men_n1474_));
  NA3        u1446(.A(men_men_n1474_), .B(men_men_n1456_), .C(men_men_n1449_), .Y(men_men_n1475_));
  NA3        u1447(.A(men_men_n955_), .B(men_men_n134_), .C(men_men_n46_), .Y(men_men_n1476_));
  AOI210     u1448(.A0(men_men_n142_), .A1(c), .B0(men_men_n1476_), .Y(men_men_n1477_));
  INV        u1449(.A(men_men_n177_), .Y(men_men_n1478_));
  NA2        u1450(.A(men_men_n1478_), .B(men_men_n1422_), .Y(men_men_n1479_));
  AO210      u1451(.A0(men_men_n129_), .A1(l), .B0(men_men_n1381_), .Y(men_men_n1480_));
  NO2        u1452(.A(men_men_n72_), .B(c), .Y(men_men_n1481_));
  NO4        u1453(.A(men_men_n1345_), .B(men_men_n178_), .C(men_men_n439_), .D(men_men_n45_), .Y(men_men_n1482_));
  AOI210     u1454(.A0(men_men_n1428_), .A1(men_men_n1481_), .B0(men_men_n1482_), .Y(men_men_n1483_));
  NA3        u1455(.A(men_men_n1483_), .B(men_men_n1480_), .C(men_men_n1479_), .Y(men_men_n1484_));
  NO2        u1456(.A(men_men_n1484_), .B(men_men_n1477_), .Y(men_men_n1485_));
  NO4        u1457(.A(men_men_n212_), .B(men_men_n178_), .C(men_men_n245_), .D(k), .Y(men_men_n1486_));
  AOI210     u1458(.A0(men_men_n150_), .A1(men_men_n56_), .B0(men_men_n1450_), .Y(men_men_n1487_));
  NO2        u1459(.A(men_men_n1487_), .B(men_men_n1425_), .Y(men_men_n1488_));
  NO2        u1460(.A(men_men_n1476_), .B(men_men_n109_), .Y(men_men_n1489_));
  NOi21      u1461(.An(men_men_n1326_), .B(e), .Y(men_men_n1490_));
  NO4        u1462(.A(men_men_n1490_), .B(men_men_n1489_), .C(men_men_n1488_), .D(men_men_n1486_), .Y(men_men_n1491_));
  AOI220     u1463(.A0(men_men_n1470_), .A1(men_men_n633_), .B0(men_men_n1512_), .B1(men_men_n153_), .Y(men_men_n1492_));
  NOi31      u1464(.An(men_men_n30_), .B(men_men_n1492_), .C(n), .Y(men_men_n1493_));
  INV        u1465(.A(men_men_n1493_), .Y(men_men_n1494_));
  NA2        u1466(.A(men_men_n59_), .B(a), .Y(men_men_n1495_));
  NO2        u1467(.A(men_men_n1333_), .B(men_men_n116_), .Y(men_men_n1496_));
  OAI220     u1468(.A0(men_men_n1496_), .A1(men_men_n1381_), .B0(men_men_n1397_), .B1(men_men_n1495_), .Y(men_men_n1497_));
  NA4        u1469(.A(men_men_n1511_), .B(men_men_n1494_), .C(men_men_n1491_), .D(men_men_n1485_), .Y(men_men_n1498_));
  OR4        u1470(.A(men_men_n1498_), .B(men_men_n1475_), .C(men_men_n1435_), .D(men_men_n1401_), .Y(men04));
  NOi31      u1471(.An(men_men_n1388_), .B(men_men_n1389_), .C(men_men_n1039_), .Y(men_men_n1500_));
  NA2        u1472(.A(men_men_n1430_), .B(men_men_n814_), .Y(men_men_n1501_));
  NO4        u1473(.A(men_men_n1501_), .B(men_men_n1029_), .C(men_men_n472_), .D(j), .Y(men_men_n1502_));
  OR3        u1474(.A(men_men_n1502_), .B(men_men_n1500_), .C(men_men_n1056_), .Y(men_men_n1503_));
  NO3        u1475(.A(men_men_n1334_), .B(men_men_n93_), .C(k), .Y(men_men_n1504_));
  AOI210     u1476(.A0(men_men_n1504_), .A1(men_men_n1050_), .B0(men_men_n1169_), .Y(men_men_n1505_));
  NA2        u1477(.A(men_men_n1505_), .B(men_men_n1196_), .Y(men_men_n1506_));
  NO3        u1478(.A(men_men_n1506_), .B(men_men_n1503_), .C(men_men_n1044_), .Y(men_men_n1507_));
  NA3        u1479(.A(men_men_n1507_), .B(men_men_n1092_), .C(men_men_n1080_), .Y(men05));
  INV        u1480(.A(men_men_n1497_), .Y(men_men_n1511_));
  INV        u1481(.A(j), .Y(men_men_n1512_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule