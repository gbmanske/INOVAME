library verilog;
use verilog.vl_types.all;
entity tb_maquinaVenda is
end tb_maquinaVenda;
