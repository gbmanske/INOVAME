// Benchmark "top" written by ABC on Fri Jun 21 17:49:20 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n142_, new_new_n143_,
    new_new_n144_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n827_, new_new_n828_, new_new_n829_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1107_, new_new_n1111_,
    new_new_n1112_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  OAI210     g0034(.A0(new_new_n56_), .A1(new_new_n53_), .B0(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  OAI210     g0068(.A0(new_new_n86_), .A1(new_new_n83_), .B0(i_2_), .Y(new_new_n91_));
  NAi21      g0069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g0070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n64_), .Y(new_new_n94_));
  NA2        g0072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g0073(.A(new_new_n95_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g0074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g0075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n81_), .Y(new_new_n98_));
  AN3        g0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g0077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g0078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g0079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g0080(.A0(new_new_n102_), .A1(new_new_n63_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g0081(.A(i_7_), .Y(new_new_n104_));
  NA2        g0082(.A(new_new_n47_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g0083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g0084(.A(new_new_n106_), .B(new_new_n87_), .Y(new_new_n107_));
  NA2        g0085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g0086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g0087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g0088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  NO3        g0089(.A(new_new_n111_), .B(new_new_n92_), .C(new_new_n54_), .Y(new_new_n112_));
  AN2        g0090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g0092(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n115_));
  NO2        g0093(.A(i_8_), .B(new_new_n104_), .Y(new_new_n116_));
  NO3        g0094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g0095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g0097(.A(new_new_n119_), .B(i_0_), .Y(new_new_n120_));
  NA2        g0098(.A(i_11_), .B(i_12_), .Y(new_new_n121_));
  OAI210     g0099(.A0(new_new_n120_), .A1(new_new_n118_), .B0(new_new_n121_), .Y(new_new_n122_));
  NO2        g0100(.A(new_new_n122_), .B(new_new_n117_), .Y(new_new_n123_));
  NAi41      g0101(.An(new_new_n112_), .B(new_new_n123_), .C(new_new_n110_), .D(new_new_n103_), .Y(new_new_n124_));
  NOi21      g0102(.An(i_1_), .B(i_5_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(i_11_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g0105(.A(i_7_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NO2        g0107(.A(new_new_n129_), .B(new_new_n47_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n131_));
  NAi21      g0109(.An(i_3_), .B(i_8_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(new_new_n63_), .Y(new_new_n133_));
  NOi31      g0111(.An(new_new_n133_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n134_));
  NO2        g0112(.A(i_1_), .B(new_new_n87_), .Y(new_new_n135_));
  NO2        g0113(.A(i_6_), .B(i_5_), .Y(new_new_n136_));
  NA2        g0114(.A(new_new_n136_), .B(i_3_), .Y(new_new_n137_));
  AO210      g0115(.A0(new_new_n137_), .A1(new_new_n48_), .B0(new_new_n135_), .Y(new_new_n138_));
  OAI220     g0116(.A0(new_new_n138_), .A1(new_new_n111_), .B0(new_new_n134_), .B1(new_new_n126_), .Y(new_new_n139_));
  NO3        g0117(.A(new_new_n139_), .B(new_new_n124_), .C(new_new_n98_), .Y(new_new_n140_));
  NA3        g0118(.A(new_new_n140_), .B(new_new_n80_), .C(new_new_n57_), .Y(men2));
  NO2        g0119(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n142_));
  NA2        g0120(.A(i_6_), .B(new_new_n25_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NA4        g0122(.A(new_new_n144_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(men0));
  AN2        g0123(.A(i_8_), .B(i_7_), .Y(new_new_n146_));
  NA2        g0124(.A(new_new_n146_), .B(i_6_), .Y(new_new_n147_));
  NO2        g0125(.A(i_12_), .B(i_13_), .Y(new_new_n148_));
  NAi21      g0126(.An(i_5_), .B(i_11_), .Y(new_new_n149_));
  NOi21      g0127(.An(new_new_n148_), .B(new_new_n149_), .Y(new_new_n150_));
  NO2        g0128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NA2        g0129(.A(i_2_), .B(i_3_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(i_4_), .Y(new_new_n153_));
  NA3        g0131(.A(new_new_n153_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n154_));
  OR2        g0132(.A(new_new_n154_), .B(new_new_n25_), .Y(new_new_n155_));
  AN2        g0133(.A(new_new_n148_), .B(new_new_n84_), .Y(new_new_n156_));
  NO2        g0134(.A(new_new_n156_), .B(new_new_n27_), .Y(new_new_n157_));
  NA2        g0135(.A(i_1_), .B(i_5_), .Y(new_new_n158_));
  NO2        g0136(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n159_));
  NA2        g0137(.A(new_new_n159_), .B(new_new_n36_), .Y(new_new_n160_));
  NO3        g0138(.A(new_new_n160_), .B(new_new_n158_), .C(new_new_n157_), .Y(new_new_n161_));
  OR2        g0139(.A(i_0_), .B(i_1_), .Y(new_new_n162_));
  NO3        g0140(.A(new_new_n162_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n163_));
  NAi32      g0141(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n164_));
  NAi21      g0142(.An(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  NOi21      g0143(.An(i_4_), .B(i_10_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n40_), .Y(new_new_n167_));
  NO2        g0145(.A(i_3_), .B(i_5_), .Y(new_new_n168_));
  NO3        g0146(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n169_));
  NA2        g0147(.A(new_new_n169_), .B(new_new_n168_), .Y(new_new_n170_));
  OAI210     g0148(.A0(new_new_n170_), .A1(new_new_n167_), .B0(new_new_n165_), .Y(new_new_n171_));
  NO2        g0149(.A(new_new_n171_), .B(new_new_n161_), .Y(new_new_n172_));
  AOI210     g0150(.A0(new_new_n172_), .A1(new_new_n155_), .B0(new_new_n147_), .Y(new_new_n173_));
  NA3        g0151(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n174_));
  NA2        g0152(.A(i_3_), .B(new_new_n49_), .Y(new_new_n175_));
  NOi21      g0153(.An(i_4_), .B(i_9_), .Y(new_new_n176_));
  NOi21      g0154(.An(i_11_), .B(i_13_), .Y(new_new_n177_));
  NA2        g0155(.A(new_new_n177_), .B(new_new_n176_), .Y(new_new_n178_));
  OR2        g0156(.A(new_new_n178_), .B(new_new_n175_), .Y(new_new_n179_));
  NO2        g0157(.A(i_4_), .B(i_5_), .Y(new_new_n180_));
  NAi21      g0158(.An(i_12_), .B(i_11_), .Y(new_new_n181_));
  NO2        g0159(.A(new_new_n181_), .B(i_13_), .Y(new_new_n182_));
  NA3        g0160(.A(new_new_n182_), .B(new_new_n180_), .C(new_new_n84_), .Y(new_new_n183_));
  AOI210     g0161(.A0(new_new_n183_), .A1(new_new_n179_), .B0(new_new_n174_), .Y(new_new_n184_));
  NO2        g0162(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n185_));
  NA2        g0163(.A(new_new_n185_), .B(new_new_n47_), .Y(new_new_n186_));
  NA2        g0164(.A(new_new_n36_), .B(i_5_), .Y(new_new_n187_));
  NAi31      g0165(.An(new_new_n187_), .B(new_new_n156_), .C(i_11_), .Y(new_new_n188_));
  NA2        g0166(.A(i_3_), .B(i_5_), .Y(new_new_n189_));
  OR2        g0167(.A(new_new_n189_), .B(new_new_n178_), .Y(new_new_n190_));
  AOI210     g0168(.A0(new_new_n190_), .A1(new_new_n188_), .B0(new_new_n186_), .Y(new_new_n191_));
  NO2        g0169(.A(new_new_n74_), .B(i_5_), .Y(new_new_n192_));
  NO2        g0170(.A(i_13_), .B(i_10_), .Y(new_new_n193_));
  NA3        g0171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n45_), .Y(new_new_n194_));
  NO2        g0172(.A(i_2_), .B(i_1_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(i_3_), .Y(new_new_n196_));
  NAi21      g0174(.An(i_4_), .B(i_12_), .Y(new_new_n197_));
  NO4        g0175(.A(new_new_n197_), .B(new_new_n196_), .C(new_new_n194_), .D(new_new_n25_), .Y(new_new_n198_));
  NO3        g0176(.A(new_new_n198_), .B(new_new_n191_), .C(new_new_n184_), .Y(new_new_n199_));
  INV        g0177(.A(i_8_), .Y(new_new_n200_));
  NO2        g0178(.A(new_new_n200_), .B(i_7_), .Y(new_new_n201_));
  NA2        g0179(.A(new_new_n201_), .B(i_6_), .Y(new_new_n202_));
  NO3        g0180(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n203_));
  NA2        g0181(.A(new_new_n203_), .B(new_new_n116_), .Y(new_new_n204_));
  NO3        g0182(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n205_));
  NA3        g0183(.A(new_new_n205_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n206_));
  NO3        g0184(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n207_));
  OAI210     g0185(.A0(new_new_n99_), .A1(i_12_), .B0(new_new_n207_), .Y(new_new_n208_));
  AOI210     g0186(.A0(new_new_n208_), .A1(new_new_n206_), .B0(new_new_n204_), .Y(new_new_n209_));
  NO2        g0187(.A(i_3_), .B(i_8_), .Y(new_new_n210_));
  NO3        g0188(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n211_));
  NA3        g0189(.A(new_new_n211_), .B(new_new_n210_), .C(new_new_n40_), .Y(new_new_n212_));
  NO2        g0190(.A(new_new_n106_), .B(new_new_n59_), .Y(new_new_n213_));
  NO2        g0191(.A(i_13_), .B(i_9_), .Y(new_new_n214_));
  NA3        g0192(.A(new_new_n214_), .B(i_6_), .C(new_new_n200_), .Y(new_new_n215_));
  NAi21      g0193(.An(i_12_), .B(i_3_), .Y(new_new_n216_));
  OR2        g0194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n45_), .B(i_5_), .Y(new_new_n218_));
  NO3        g0196(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n219_));
  NA2        g0197(.A(new_new_n219_), .B(i_10_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n220_), .A1(new_new_n217_), .B0(new_new_n106_), .B1(new_new_n212_), .Y(new_new_n221_));
  AOI210     g0199(.A0(new_new_n221_), .A1(i_7_), .B0(new_new_n209_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(i_4_), .B0(new_new_n202_), .B1(new_new_n199_), .Y(new_new_n223_));
  NAi21      g0201(.An(i_12_), .B(i_7_), .Y(new_new_n224_));
  NA3        g0202(.A(i_13_), .B(new_new_n200_), .C(i_10_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  NA2        g0204(.A(i_0_), .B(i_5_), .Y(new_new_n227_));
  OAI220     g0205(.A0(new_new_n87_), .A1(new_new_n196_), .B0(new_new_n186_), .B1(new_new_n137_), .Y(new_new_n228_));
  NAi31      g0206(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n36_), .B(i_13_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n231_));
  NA3        g0209(.A(new_new_n231_), .B(i_0_), .C(new_new_n230_), .Y(new_new_n232_));
  INV        g0210(.A(i_13_), .Y(new_new_n233_));
  NO2        g0211(.A(i_12_), .B(new_new_n233_), .Y(new_new_n234_));
  NA3        g0212(.A(new_new_n234_), .B(new_new_n205_), .C(new_new_n203_), .Y(new_new_n235_));
  OAI210     g0213(.A0(new_new_n232_), .A1(new_new_n229_), .B0(new_new_n235_), .Y(new_new_n236_));
  AOI220     g0214(.A0(new_new_n236_), .A1(new_new_n146_), .B0(new_new_n228_), .B1(new_new_n226_), .Y(new_new_n237_));
  NO2        g0215(.A(i_12_), .B(new_new_n37_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n189_), .B(i_4_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  OR2        g0218(.A(i_8_), .B(i_7_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n241_), .B(new_new_n87_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n54_), .B(i_1_), .Y(new_new_n243_));
  NA2        g0221(.A(new_new_n243_), .B(new_new_n242_), .Y(new_new_n244_));
  INV        g0222(.A(i_12_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n45_), .B(new_new_n245_), .Y(new_new_n246_));
  NO3        g0224(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(i_2_), .B(i_1_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n244_), .B(new_new_n240_), .Y(new_new_n249_));
  NO3        g0227(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n250_));
  NAi21      g0228(.An(i_4_), .B(i_3_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n251_), .B(new_new_n76_), .Y(new_new_n252_));
  NO2        g0230(.A(i_0_), .B(i_6_), .Y(new_new_n253_));
  NOi41      g0231(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n254_));
  NA2        g0232(.A(new_new_n254_), .B(new_new_n253_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n248_), .B(new_new_n189_), .Y(new_new_n256_));
  NAi21      g0234(.An(new_new_n255_), .B(new_new_n256_), .Y(new_new_n257_));
  INV        g0235(.A(new_new_n257_), .Y(new_new_n258_));
  AOI220     g0236(.A0(new_new_n258_), .A1(new_new_n40_), .B0(new_new_n249_), .B1(new_new_n214_), .Y(new_new_n259_));
  NO2        g0237(.A(i_11_), .B(new_new_n233_), .Y(new_new_n260_));
  NOi21      g0238(.An(i_1_), .B(i_6_), .Y(new_new_n261_));
  NAi21      g0239(.An(i_3_), .B(i_7_), .Y(new_new_n262_));
  NO2        g0240(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n263_));
  NO2        g0241(.A(i_12_), .B(i_3_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n74_), .B(i_5_), .Y(new_new_n265_));
  NA2        g0243(.A(i_3_), .B(i_9_), .Y(new_new_n266_));
  NAi21      g0244(.An(i_7_), .B(i_10_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n267_), .B(new_new_n266_), .Y(new_new_n268_));
  NA3        g0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n269_));
  INV        g0247(.A(new_new_n147_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n245_), .B(i_13_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n76_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n272_), .B(new_new_n270_), .Y(new_new_n273_));
  NO2        g0251(.A(new_new_n241_), .B(new_new_n37_), .Y(new_new_n274_));
  NA2        g0252(.A(i_12_), .B(i_6_), .Y(new_new_n275_));
  OR2        g0253(.A(i_13_), .B(i_9_), .Y(new_new_n276_));
  NO3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n49_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n251_), .B(i_2_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n277_), .C(new_new_n45_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n260_), .B(i_9_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n265_), .B(new_new_n162_), .C(new_new_n65_), .Y(new_new_n281_));
  OAI210     g0259(.A0(new_new_n281_), .A1(new_new_n280_), .B0(new_new_n279_), .Y(new_new_n282_));
  NA2        g0260(.A(new_new_n159_), .B(new_new_n64_), .Y(new_new_n283_));
  NO3        g0261(.A(i_11_), .B(new_new_n233_), .C(new_new_n25_), .Y(new_new_n284_));
  NO2        g0262(.A(new_new_n262_), .B(i_8_), .Y(new_new_n285_));
  NO2        g0263(.A(i_6_), .B(new_new_n49_), .Y(new_new_n286_));
  NA3        g0264(.A(new_new_n286_), .B(new_new_n285_), .C(new_new_n284_), .Y(new_new_n287_));
  NO3        g0265(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n288_));
  NA3        g0266(.A(new_new_n288_), .B(new_new_n274_), .C(new_new_n234_), .Y(new_new_n289_));
  AOI210     g0267(.A0(new_new_n289_), .A1(new_new_n287_), .B0(new_new_n283_), .Y(new_new_n290_));
  AOI210     g0268(.A0(new_new_n282_), .A1(new_new_n274_), .B0(new_new_n290_), .Y(new_new_n291_));
  NA4        g0269(.A(new_new_n291_), .B(new_new_n273_), .C(new_new_n259_), .D(new_new_n237_), .Y(new_new_n292_));
  NO3        g0270(.A(i_12_), .B(new_new_n233_), .C(new_new_n37_), .Y(new_new_n293_));
  INV        g0271(.A(new_new_n293_), .Y(new_new_n294_));
  NA2        g0272(.A(i_8_), .B(new_new_n104_), .Y(new_new_n295_));
  NO3        g0273(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n296_));
  AOI220     g0274(.A0(new_new_n296_), .A1(new_new_n203_), .B0(new_new_n168_), .B1(new_new_n243_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(new_new_n295_), .Y(new_new_n298_));
  NO3        g0276(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n248_), .B(i_0_), .Y(new_new_n300_));
  AOI220     g0278(.A0(new_new_n300_), .A1(new_new_n201_), .B0(new_new_n299_), .B1(new_new_n146_), .Y(new_new_n301_));
  NA2        g0279(.A(new_new_n286_), .B(new_new_n26_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n302_), .B(new_new_n301_), .Y(new_new_n303_));
  NA2        g0281(.A(i_0_), .B(i_1_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n304_), .B(i_2_), .Y(new_new_n305_));
  NO2        g0283(.A(new_new_n60_), .B(i_6_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(new_new_n305_), .C(new_new_n168_), .Y(new_new_n307_));
  OAI210     g0285(.A0(new_new_n170_), .A1(new_new_n147_), .B0(new_new_n307_), .Y(new_new_n308_));
  NO3        g0286(.A(new_new_n308_), .B(new_new_n303_), .C(new_new_n298_), .Y(new_new_n309_));
  NO2        g0287(.A(i_3_), .B(i_10_), .Y(new_new_n310_));
  NA3        g0288(.A(new_new_n310_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n311_));
  NO2        g0289(.A(i_2_), .B(new_new_n104_), .Y(new_new_n312_));
  NA2        g0290(.A(i_1_), .B(new_new_n36_), .Y(new_new_n313_));
  NOi21      g0291(.An(new_new_n227_), .B(new_new_n106_), .Y(new_new_n314_));
  NA3        g0292(.A(new_new_n314_), .B(i_1_), .C(new_new_n312_), .Y(new_new_n315_));
  AN2        g0293(.A(i_3_), .B(i_10_), .Y(new_new_n316_));
  NA4        g0294(.A(new_new_n316_), .B(new_new_n205_), .C(new_new_n182_), .D(new_new_n180_), .Y(new_new_n317_));
  NO2        g0295(.A(i_5_), .B(new_new_n37_), .Y(new_new_n318_));
  NO2        g0296(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n319_));
  OR2        g0297(.A(new_new_n315_), .B(new_new_n311_), .Y(new_new_n320_));
  OAI220     g0298(.A0(new_new_n320_), .A1(i_6_), .B0(new_new_n309_), .B1(new_new_n294_), .Y(new_new_n321_));
  NO4        g0299(.A(new_new_n321_), .B(new_new_n292_), .C(new_new_n223_), .D(new_new_n173_), .Y(new_new_n322_));
  NO3        g0300(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n323_));
  NO2        g0301(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n324_));
  NA2        g0302(.A(new_new_n300_), .B(new_new_n324_), .Y(new_new_n325_));
  NO3        g0303(.A(i_6_), .B(new_new_n200_), .C(i_7_), .Y(new_new_n326_));
  NA2        g0304(.A(new_new_n326_), .B(new_new_n205_), .Y(new_new_n327_));
  AOI210     g0305(.A0(new_new_n327_), .A1(new_new_n325_), .B0(new_new_n175_), .Y(new_new_n328_));
  NO2        g0306(.A(i_2_), .B(i_3_), .Y(new_new_n329_));
  OR2        g0307(.A(i_0_), .B(i_5_), .Y(new_new_n330_));
  NA2        g0308(.A(new_new_n227_), .B(new_new_n330_), .Y(new_new_n331_));
  NA4        g0309(.A(new_new_n331_), .B(new_new_n242_), .C(new_new_n329_), .D(i_1_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n300_), .B(new_new_n168_), .C(new_new_n116_), .Y(new_new_n333_));
  NAi21      g0311(.An(i_8_), .B(i_7_), .Y(new_new_n334_));
  NO2        g0312(.A(new_new_n334_), .B(i_6_), .Y(new_new_n335_));
  NO2        g0313(.A(new_new_n162_), .B(new_new_n47_), .Y(new_new_n336_));
  NA3        g0314(.A(new_new_n336_), .B(new_new_n335_), .C(new_new_n168_), .Y(new_new_n337_));
  NA3        g0315(.A(new_new_n337_), .B(new_new_n333_), .C(new_new_n332_), .Y(new_new_n338_));
  OAI210     g0316(.A0(new_new_n338_), .A1(new_new_n328_), .B0(i_4_), .Y(new_new_n339_));
  NO2        g0317(.A(i_12_), .B(i_10_), .Y(new_new_n340_));
  NOi21      g0318(.An(i_5_), .B(i_0_), .Y(new_new_n341_));
  AOI210     g0319(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n104_), .Y(new_new_n342_));
  NO4        g0320(.A(new_new_n342_), .B(new_new_n313_), .C(new_new_n341_), .D(new_new_n132_), .Y(new_new_n343_));
  NA4        g0321(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n344_));
  NA2        g0322(.A(new_new_n343_), .B(new_new_n340_), .Y(new_new_n345_));
  NO2        g0323(.A(i_6_), .B(i_8_), .Y(new_new_n346_));
  NOi21      g0324(.An(i_0_), .B(i_2_), .Y(new_new_n347_));
  AN2        g0325(.A(new_new_n347_), .B(new_new_n346_), .Y(new_new_n348_));
  NO2        g0326(.A(i_1_), .B(i_7_), .Y(new_new_n349_));
  AO220      g0327(.A0(new_new_n349_), .A1(new_new_n348_), .B0(new_new_n335_), .B1(new_new_n243_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n350_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n351_));
  NA3        g0329(.A(new_new_n351_), .B(new_new_n345_), .C(new_new_n339_), .Y(new_new_n352_));
  NO3        g0330(.A(new_new_n241_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n353_));
  NO3        g0331(.A(new_new_n334_), .B(i_2_), .C(i_1_), .Y(new_new_n354_));
  OAI210     g0332(.A0(new_new_n354_), .A1(new_new_n353_), .B0(i_6_), .Y(new_new_n355_));
  NA3        g0333(.A(new_new_n261_), .B(new_new_n312_), .C(new_new_n200_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n356_), .A1(new_new_n355_), .B0(new_new_n331_), .Y(new_new_n357_));
  NOi21      g0335(.An(new_new_n158_), .B(new_new_n107_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n358_), .B(new_new_n128_), .Y(new_new_n359_));
  OAI210     g0337(.A0(new_new_n359_), .A1(new_new_n357_), .B0(i_3_), .Y(new_new_n360_));
  INV        g0338(.A(new_new_n85_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n304_), .B(new_new_n82_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n136_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n95_), .B(new_new_n200_), .Y(new_new_n364_));
  NA3        g0342(.A(new_new_n314_), .B(new_new_n364_), .C(new_new_n64_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n365_), .A1(new_new_n363_), .B0(new_new_n361_), .Y(new_new_n366_));
  NO2        g0344(.A(new_new_n200_), .B(i_9_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n213_), .C(new_new_n162_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n368_), .B(new_new_n47_), .Y(new_new_n369_));
  NO3        g0347(.A(new_new_n369_), .B(new_new_n366_), .C(new_new_n303_), .Y(new_new_n370_));
  AOI210     g0348(.A0(new_new_n370_), .A1(new_new_n360_), .B0(new_new_n167_), .Y(new_new_n371_));
  AOI210     g0349(.A0(new_new_n352_), .A1(new_new_n323_), .B0(new_new_n371_), .Y(new_new_n372_));
  NOi32      g0350(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n373_));
  INV        g0351(.A(new_new_n373_), .Y(new_new_n374_));
  NAi21      g0352(.An(i_0_), .B(i_6_), .Y(new_new_n375_));
  NAi21      g0353(.An(i_1_), .B(i_5_), .Y(new_new_n376_));
  NA2        g0354(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n377_));
  NA2        g0355(.A(new_new_n377_), .B(new_new_n25_), .Y(new_new_n378_));
  OAI210     g0356(.A0(new_new_n378_), .A1(new_new_n164_), .B0(new_new_n255_), .Y(new_new_n379_));
  NAi41      g0357(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n380_));
  OAI220     g0358(.A0(new_new_n380_), .A1(new_new_n376_), .B0(new_new_n229_), .B1(new_new_n164_), .Y(new_new_n381_));
  AOI210     g0359(.A0(new_new_n380_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n382_));
  NOi32      g0360(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n383_));
  NAi21      g0361(.An(i_6_), .B(i_1_), .Y(new_new_n384_));
  NA3        g0362(.A(new_new_n384_), .B(new_new_n383_), .C(new_new_n47_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(i_0_), .Y(new_new_n386_));
  OR3        g0364(.A(new_new_n386_), .B(new_new_n382_), .C(new_new_n381_), .Y(new_new_n387_));
  NO2        g0365(.A(i_1_), .B(new_new_n104_), .Y(new_new_n388_));
  NAi21      g0366(.An(i_3_), .B(i_4_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n389_), .B(i_9_), .Y(new_new_n390_));
  AN2        g0368(.A(i_6_), .B(i_7_), .Y(new_new_n391_));
  OAI210     g0369(.A0(new_new_n391_), .A1(new_new_n388_), .B0(new_new_n390_), .Y(new_new_n392_));
  NA2        g0370(.A(i_2_), .B(i_7_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n389_), .B(i_10_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n392_), .B(new_new_n192_), .Y(new_new_n395_));
  AOI210     g0373(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n396_));
  OAI210     g0374(.A0(new_new_n396_), .A1(new_new_n195_), .B0(new_new_n394_), .Y(new_new_n397_));
  AOI220     g0375(.A0(new_new_n394_), .A1(new_new_n349_), .B0(new_new_n247_), .B1(new_new_n195_), .Y(new_new_n398_));
  AOI210     g0376(.A0(new_new_n398_), .A1(new_new_n397_), .B0(i_5_), .Y(new_new_n399_));
  NO4        g0377(.A(new_new_n399_), .B(new_new_n395_), .C(new_new_n387_), .D(new_new_n379_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n400_), .B(new_new_n374_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n402_));
  AN2        g0380(.A(i_12_), .B(i_5_), .Y(new_new_n403_));
  NO2        g0381(.A(i_4_), .B(new_new_n26_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n404_), .B(new_new_n403_), .Y(new_new_n405_));
  NO2        g0383(.A(i_11_), .B(i_6_), .Y(new_new_n406_));
  NA3        g0384(.A(new_new_n406_), .B(new_new_n336_), .C(new_new_n233_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n405_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n251_), .B(i_5_), .Y(new_new_n409_));
  NO2        g0387(.A(i_5_), .B(i_10_), .Y(new_new_n410_));
  AOI220     g0388(.A0(new_new_n410_), .A1(new_new_n278_), .B0(new_new_n409_), .B1(new_new_n205_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n148_), .B(new_new_n46_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n412_), .B(new_new_n411_), .Y(new_new_n413_));
  OAI210     g0391(.A0(new_new_n413_), .A1(new_new_n408_), .B0(new_new_n402_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n154_), .B(new_new_n87_), .Y(new_new_n416_));
  OAI210     g0394(.A0(new_new_n416_), .A1(new_new_n408_), .B0(new_new_n415_), .Y(new_new_n417_));
  NO3        g0395(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n418_));
  NO2        g0396(.A(i_3_), .B(new_new_n104_), .Y(new_new_n419_));
  NO2        g0397(.A(i_11_), .B(i_12_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n410_), .B(new_new_n245_), .Y(new_new_n421_));
  NA3        g0399(.A(new_new_n116_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n422_));
  OAI220     g0400(.A0(new_new_n422_), .A1(new_new_n229_), .B0(new_new_n421_), .B1(new_new_n344_), .Y(new_new_n423_));
  NAi21      g0401(.An(i_13_), .B(i_0_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(new_new_n248_), .Y(new_new_n425_));
  NA2        g0403(.A(new_new_n423_), .B(new_new_n425_), .Y(new_new_n426_));
  NA3        g0404(.A(new_new_n426_), .B(new_new_n417_), .C(new_new_n414_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n45_), .B(new_new_n233_), .Y(new_new_n428_));
  NO3        g0406(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n429_));
  NO2        g0407(.A(i_0_), .B(i_11_), .Y(new_new_n430_));
  INV        g0408(.A(i_5_), .Y(new_new_n431_));
  AN2        g0409(.A(i_1_), .B(i_6_), .Y(new_new_n432_));
  NOi21      g0410(.An(i_2_), .B(i_12_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n433_), .B(new_new_n432_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n434_), .B(new_new_n431_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n146_), .B(i_9_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(i_4_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n435_), .B(new_new_n437_), .Y(new_new_n438_));
  OR2        g0416(.A(i_13_), .B(i_10_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n178_), .B(new_new_n127_), .Y(new_new_n440_));
  OR2        g0418(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n293_), .B(new_new_n442_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n286_), .B(new_new_n219_), .Y(new_new_n444_));
  OAI220     g0422(.A0(new_new_n444_), .A1(new_new_n441_), .B0(new_new_n443_), .B1(new_new_n358_), .Y(new_new_n445_));
  INV        g0423(.A(new_new_n445_), .Y(new_new_n446_));
  AOI210     g0424(.A0(new_new_n446_), .A1(new_new_n438_), .B0(new_new_n26_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n333_), .B(new_new_n332_), .Y(new_new_n448_));
  AOI220     g0426(.A0(new_new_n306_), .A1(new_new_n296_), .B0(new_new_n300_), .B1(new_new_n324_), .Y(new_new_n449_));
  NO2        g0427(.A(new_new_n449_), .B(new_new_n175_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n189_), .B(new_new_n87_), .Y(new_new_n451_));
  AOI220     g0429(.A0(new_new_n451_), .A1(new_new_n305_), .B0(new_new_n288_), .B1(new_new_n219_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n452_), .B(new_new_n295_), .Y(new_new_n453_));
  NO3        g0431(.A(new_new_n453_), .B(new_new_n450_), .C(new_new_n448_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n203_), .B(new_new_n99_), .Y(new_new_n455_));
  NA3        g0433(.A(new_new_n336_), .B(new_new_n168_), .C(new_new_n87_), .Y(new_new_n456_));
  AOI210     g0434(.A0(new_new_n456_), .A1(new_new_n455_), .B0(new_new_n334_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n306_), .B(new_new_n243_), .Y(new_new_n458_));
  NO2        g0436(.A(new_new_n458_), .B(new_new_n189_), .Y(new_new_n459_));
  NO2        g0437(.A(i_3_), .B(new_new_n49_), .Y(new_new_n460_));
  NA3        g0438(.A(new_new_n349_), .B(new_new_n348_), .C(new_new_n460_), .Y(new_new_n461_));
  NA2        g0439(.A(new_new_n326_), .B(new_new_n331_), .Y(new_new_n462_));
  OAI210     g0440(.A0(new_new_n462_), .A1(new_new_n196_), .B0(new_new_n461_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n463_), .B(new_new_n459_), .C(new_new_n457_), .Y(new_new_n464_));
  AOI210     g0442(.A0(new_new_n464_), .A1(new_new_n454_), .B0(new_new_n280_), .Y(new_new_n465_));
  NO4        g0443(.A(new_new_n465_), .B(new_new_n447_), .C(new_new_n427_), .D(new_new_n401_), .Y(new_new_n466_));
  NO2        g0444(.A(new_new_n64_), .B(i_4_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n74_), .B(i_13_), .Y(new_new_n468_));
  NA3        g0446(.A(new_new_n468_), .B(new_new_n467_), .C(i_2_), .Y(new_new_n469_));
  NO2        g0447(.A(i_10_), .B(i_9_), .Y(new_new_n470_));
  NAi21      g0448(.An(i_12_), .B(i_8_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n471_), .B(i_3_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n472_), .B(new_new_n470_), .Y(new_new_n473_));
  NO2        g0451(.A(new_new_n47_), .B(i_4_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n474_), .B(new_new_n107_), .Y(new_new_n475_));
  OAI220     g0453(.A0(new_new_n475_), .A1(new_new_n212_), .B0(new_new_n473_), .B1(new_new_n469_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n319_), .B(i_0_), .Y(new_new_n477_));
  NO3        g0455(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n275_), .B(new_new_n100_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n479_), .B(new_new_n478_), .Y(new_new_n480_));
  NA2        g0458(.A(i_8_), .B(i_9_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n480_), .B(new_new_n477_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n260_), .B(new_new_n318_), .Y(new_new_n483_));
  NO3        g0461(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n484_));
  AOI210     g0462(.A0(new_new_n264_), .A1(new_new_n195_), .B0(new_new_n484_), .Y(new_new_n485_));
  NA3        g0463(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n486_));
  NA4        g0464(.A(new_new_n149_), .B(new_new_n119_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n487_));
  OAI220     g0465(.A0(new_new_n487_), .A1(new_new_n486_), .B0(new_new_n485_), .B1(new_new_n483_), .Y(new_new_n488_));
  NO3        g0466(.A(new_new_n488_), .B(new_new_n482_), .C(new_new_n476_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n305_), .B(new_new_n111_), .Y(new_new_n490_));
  OR2        g0468(.A(new_new_n490_), .B(new_new_n215_), .Y(new_new_n491_));
  OA210      g0469(.A0(new_new_n368_), .A1(new_new_n104_), .B0(new_new_n307_), .Y(new_new_n492_));
  OA220      g0470(.A0(new_new_n492_), .A1(new_new_n167_), .B0(new_new_n491_), .B1(new_new_n240_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n99_), .B(i_13_), .Y(new_new_n494_));
  NA2        g0472(.A(new_new_n451_), .B(new_new_n402_), .Y(new_new_n495_));
  NO2        g0473(.A(i_2_), .B(i_13_), .Y(new_new_n496_));
  NA3        g0474(.A(new_new_n496_), .B(new_new_n166_), .C(new_new_n102_), .Y(new_new_n497_));
  OAI220     g0475(.A0(new_new_n497_), .A1(new_new_n245_), .B0(new_new_n495_), .B1(new_new_n494_), .Y(new_new_n498_));
  NO3        g0476(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n499_));
  NO2        g0477(.A(i_6_), .B(i_7_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n500_), .B(new_new_n499_), .Y(new_new_n501_));
  NO2        g0479(.A(i_11_), .B(i_1_), .Y(new_new_n502_));
  OR2        g0480(.A(i_11_), .B(i_8_), .Y(new_new_n503_));
  NOi21      g0481(.An(i_2_), .B(i_7_), .Y(new_new_n504_));
  NAi31      g0482(.An(new_new_n503_), .B(new_new_n504_), .C(i_0_), .Y(new_new_n505_));
  NO2        g0483(.A(new_new_n439_), .B(i_6_), .Y(new_new_n506_));
  NA3        g0484(.A(new_new_n506_), .B(new_new_n467_), .C(new_new_n76_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n507_), .B(new_new_n505_), .Y(new_new_n508_));
  NO2        g0486(.A(i_3_), .B(new_new_n200_), .Y(new_new_n509_));
  NO2        g0487(.A(i_6_), .B(i_10_), .Y(new_new_n510_));
  NA4        g0488(.A(new_new_n510_), .B(new_new_n323_), .C(new_new_n509_), .D(new_new_n245_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n511_), .B(new_new_n160_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n162_), .B(i_3_), .Y(new_new_n514_));
  NAi31      g0492(.An(new_new_n513_), .B(new_new_n514_), .C(new_new_n234_), .Y(new_new_n515_));
  NA3        g0493(.A(new_new_n415_), .B(new_new_n185_), .C(new_new_n153_), .Y(new_new_n516_));
  NA2        g0494(.A(new_new_n516_), .B(new_new_n515_), .Y(new_new_n517_));
  NO4        g0495(.A(new_new_n517_), .B(new_new_n512_), .C(new_new_n508_), .D(new_new_n498_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n478_), .B(new_new_n403_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n484_), .B(new_new_n410_), .Y(new_new_n520_));
  NO2        g0498(.A(new_new_n520_), .B(new_new_n232_), .Y(new_new_n521_));
  NAi21      g0499(.An(new_new_n225_), .B(new_new_n420_), .Y(new_new_n522_));
  NA2        g0500(.A(new_new_n349_), .B(new_new_n227_), .Y(new_new_n523_));
  NO2        g0501(.A(new_new_n26_), .B(i_5_), .Y(new_new_n524_));
  NO2        g0502(.A(i_0_), .B(new_new_n87_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n525_), .B(new_new_n524_), .C(new_new_n146_), .Y(new_new_n526_));
  OR3        g0504(.A(new_new_n313_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n527_));
  OAI220     g0505(.A0(new_new_n527_), .A1(new_new_n526_), .B0(new_new_n523_), .B1(new_new_n522_), .Y(new_new_n528_));
  NA4        g0506(.A(new_new_n316_), .B(new_new_n231_), .C(new_new_n74_), .D(new_new_n245_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n529_), .B(new_new_n501_), .Y(new_new_n530_));
  NO3        g0508(.A(new_new_n530_), .B(new_new_n528_), .C(new_new_n521_), .Y(new_new_n531_));
  NA4        g0509(.A(new_new_n531_), .B(new_new_n518_), .C(new_new_n493_), .D(new_new_n489_), .Y(new_new_n532_));
  NA3        g0510(.A(new_new_n316_), .B(new_new_n182_), .C(new_new_n180_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n311_), .A1(new_new_n187_), .B0(new_new_n533_), .Y(new_new_n534_));
  AN2        g0512(.A(new_new_n296_), .B(new_new_n242_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n535_), .B(new_new_n534_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n126_), .B(new_new_n115_), .Y(new_new_n537_));
  AN2        g0515(.A(new_new_n537_), .B(new_new_n478_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n323_), .B(new_new_n169_), .Y(new_new_n539_));
  OAI210     g0517(.A0(new_new_n539_), .A1(new_new_n240_), .B0(new_new_n317_), .Y(new_new_n540_));
  AOI220     g0518(.A0(new_new_n540_), .A1(new_new_n335_), .B0(new_new_n538_), .B1(new_new_n319_), .Y(new_new_n541_));
  NA4        g0519(.A(new_new_n468_), .B(new_new_n467_), .C(new_new_n210_), .D(i_2_), .Y(new_new_n542_));
  INV        g0520(.A(new_new_n542_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n373_), .B(new_new_n74_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n391_), .B(new_new_n383_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n36_), .B(i_8_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n39_), .B(i_13_), .Y(new_new_n547_));
  INV        g0525(.A(new_new_n547_), .Y(new_new_n548_));
  AOI210     g0526(.A0(new_new_n543_), .A1(new_new_n211_), .B0(new_new_n548_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n265_), .B(new_new_n65_), .Y(new_new_n550_));
  OAI210     g0528(.A0(i_8_), .A1(new_new_n550_), .B0(new_new_n138_), .Y(new_new_n551_));
  AOI210     g0529(.A0(new_new_n201_), .A1(i_9_), .B0(new_new_n274_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n552_), .B(new_new_n206_), .Y(new_new_n553_));
  NO2        g0531(.A(new_new_n189_), .B(new_new_n87_), .Y(new_new_n554_));
  AOI220     g0532(.A0(new_new_n554_), .A1(new_new_n553_), .B0(new_new_n551_), .B1(new_new_n440_), .Y(new_new_n555_));
  NA4        g0533(.A(new_new_n555_), .B(new_new_n549_), .C(new_new_n541_), .D(new_new_n536_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n409_), .B(new_new_n305_), .Y(new_new_n557_));
  OAI210     g0535(.A0(new_new_n405_), .A1(new_new_n174_), .B0(new_new_n557_), .Y(new_new_n558_));
  NO2        g0536(.A(i_12_), .B(new_new_n200_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n559_), .B(new_new_n233_), .Y(new_new_n560_));
  NA2        g0538(.A(new_new_n510_), .B(new_new_n27_), .Y(new_new_n561_));
  NO3        g0539(.A(new_new_n561_), .B(new_new_n560_), .C(new_new_n490_), .Y(new_new_n562_));
  NOi31      g0540(.An(new_new_n326_), .B(new_new_n439_), .C(new_new_n38_), .Y(new_new_n563_));
  OAI210     g0541(.A0(new_new_n563_), .A1(new_new_n562_), .B0(new_new_n558_), .Y(new_new_n564_));
  NO2        g0542(.A(i_8_), .B(i_7_), .Y(new_new_n565_));
  OAI210     g0543(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n566_), .B(new_new_n231_), .Y(new_new_n567_));
  AOI220     g0545(.A0(new_new_n336_), .A1(new_new_n40_), .B0(new_new_n243_), .B1(new_new_n214_), .Y(new_new_n568_));
  OAI220     g0546(.A0(new_new_n568_), .A1(new_new_n189_), .B0(new_new_n567_), .B1(new_new_n251_), .Y(new_new_n569_));
  NA2        g0547(.A(new_new_n45_), .B(i_10_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n570_), .B(i_6_), .Y(new_new_n571_));
  NA3        g0549(.A(new_new_n571_), .B(new_new_n569_), .C(new_new_n565_), .Y(new_new_n572_));
  AOI220     g0550(.A0(new_new_n451_), .A1(new_new_n336_), .B0(new_new_n256_), .B1(new_new_n253_), .Y(new_new_n573_));
  OAI220     g0551(.A0(new_new_n573_), .A1(new_new_n271_), .B0(new_new_n494_), .B1(new_new_n137_), .Y(new_new_n574_));
  NA2        g0552(.A(new_new_n574_), .B(new_new_n274_), .Y(new_new_n575_));
  NOi31      g0553(.An(new_new_n300_), .B(new_new_n311_), .C(new_new_n187_), .Y(new_new_n576_));
  NA3        g0554(.A(new_new_n316_), .B(new_new_n180_), .C(new_new_n99_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n230_), .B(new_new_n45_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n162_), .B(i_5_), .Y(new_new_n579_));
  NA3        g0557(.A(new_new_n579_), .B(new_new_n428_), .C(new_new_n329_), .Y(new_new_n580_));
  OAI210     g0558(.A0(new_new_n580_), .A1(new_new_n578_), .B0(new_new_n577_), .Y(new_new_n581_));
  OAI210     g0559(.A0(new_new_n581_), .A1(new_new_n576_), .B0(new_new_n484_), .Y(new_new_n582_));
  NA4        g0560(.A(new_new_n582_), .B(new_new_n575_), .C(new_new_n572_), .D(new_new_n564_), .Y(new_new_n583_));
  NA2        g0561(.A(new_new_n293_), .B(new_new_n85_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n363_), .B(new_new_n584_), .Y(new_new_n585_));
  NA2        g0563(.A(new_new_n306_), .B(new_new_n296_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n586_), .B(new_new_n179_), .Y(new_new_n587_));
  AOI210     g0565(.A0(new_new_n384_), .A1(new_new_n47_), .B0(new_new_n388_), .Y(new_new_n588_));
  NA2        g0566(.A(i_0_), .B(new_new_n49_), .Y(new_new_n589_));
  NA3        g0567(.A(new_new_n559_), .B(new_new_n284_), .C(new_new_n589_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n588_), .B(new_new_n590_), .Y(new_new_n591_));
  NO3        g0569(.A(new_new_n591_), .B(new_new_n587_), .C(new_new_n585_), .Y(new_new_n592_));
  NO4        g0570(.A(new_new_n261_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n593_));
  NO3        g0571(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n594_));
  NO2        g0572(.A(new_new_n241_), .B(new_new_n36_), .Y(new_new_n595_));
  AN2        g0573(.A(new_new_n595_), .B(new_new_n594_), .Y(new_new_n596_));
  OA210      g0574(.A0(new_new_n596_), .A1(new_new_n593_), .B0(new_new_n373_), .Y(new_new_n597_));
  NO2        g0575(.A(new_new_n439_), .B(i_1_), .Y(new_new_n598_));
  NOi31      g0576(.An(new_new_n598_), .B(new_new_n479_), .C(new_new_n74_), .Y(new_new_n599_));
  AN4        g0577(.A(new_new_n599_), .B(new_new_n437_), .C(new_new_n524_), .D(i_2_), .Y(new_new_n600_));
  NO2        g0578(.A(new_new_n449_), .B(new_new_n183_), .Y(new_new_n601_));
  NO3        g0579(.A(new_new_n601_), .B(new_new_n600_), .C(new_new_n597_), .Y(new_new_n602_));
  NOi21      g0580(.An(i_10_), .B(i_6_), .Y(new_new_n603_));
  NO2        g0581(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n604_));
  AOI220     g0582(.A0(new_new_n293_), .A1(new_new_n604_), .B0(new_new_n284_), .B1(new_new_n603_), .Y(new_new_n605_));
  NO2        g0583(.A(new_new_n605_), .B(new_new_n477_), .Y(new_new_n606_));
  NO2        g0584(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n607_));
  NA2        g0585(.A(new_new_n326_), .B(new_new_n169_), .Y(new_new_n608_));
  AOI220     g0586(.A0(new_new_n608_), .A1(new_new_n458_), .B0(new_new_n190_), .B1(new_new_n188_), .Y(new_new_n609_));
  NO2        g0587(.A(new_new_n205_), .B(new_new_n37_), .Y(new_new_n610_));
  NOi31      g0588(.An(new_new_n150_), .B(new_new_n610_), .C(new_new_n344_), .Y(new_new_n611_));
  NO3        g0589(.A(new_new_n611_), .B(new_new_n609_), .C(new_new_n606_), .Y(new_new_n612_));
  NO2        g0590(.A(new_new_n544_), .B(new_new_n398_), .Y(new_new_n613_));
  INV        g0591(.A(new_new_n329_), .Y(new_new_n614_));
  NO2        g0592(.A(i_12_), .B(new_new_n87_), .Y(new_new_n615_));
  NA3        g0593(.A(new_new_n615_), .B(new_new_n284_), .C(new_new_n589_), .Y(new_new_n616_));
  NA3        g0594(.A(new_new_n406_), .B(new_new_n293_), .C(new_new_n227_), .Y(new_new_n617_));
  AOI210     g0595(.A0(new_new_n617_), .A1(new_new_n616_), .B0(new_new_n614_), .Y(new_new_n618_));
  NO3        g0596(.A(i_4_), .B(new_new_n355_), .C(new_new_n311_), .Y(new_new_n619_));
  OR2        g0597(.A(i_2_), .B(i_5_), .Y(new_new_n620_));
  NO3        g0598(.A(new_new_n619_), .B(new_new_n618_), .C(new_new_n613_), .Y(new_new_n621_));
  NA4        g0599(.A(new_new_n621_), .B(new_new_n612_), .C(new_new_n602_), .D(new_new_n592_), .Y(new_new_n622_));
  NO4        g0600(.A(new_new_n622_), .B(new_new_n583_), .C(new_new_n556_), .D(new_new_n532_), .Y(new_new_n623_));
  NA4        g0601(.A(new_new_n623_), .B(new_new_n466_), .C(new_new_n372_), .D(new_new_n322_), .Y(men7));
  NO2        g0602(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n625_));
  NO2        g0603(.A(new_new_n111_), .B(new_new_n92_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n404_), .B(new_new_n626_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n510_), .B(new_new_n85_), .Y(new_new_n628_));
  NA2        g0606(.A(i_11_), .B(new_new_n200_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n148_), .B(new_new_n629_), .Y(new_new_n630_));
  OAI210     g0608(.A0(new_new_n630_), .A1(new_new_n628_), .B0(new_new_n627_), .Y(new_new_n631_));
  NA3        g0609(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n245_), .B(i_4_), .Y(new_new_n633_));
  NA2        g0611(.A(new_new_n633_), .B(i_8_), .Y(new_new_n634_));
  NO2        g0612(.A(new_new_n108_), .B(new_new_n632_), .Y(new_new_n635_));
  NA2        g0613(.A(i_2_), .B(new_new_n87_), .Y(new_new_n636_));
  OAI210     g0614(.A0(new_new_n90_), .A1(new_new_n210_), .B0(new_new_n211_), .Y(new_new_n637_));
  NO2        g0615(.A(i_7_), .B(new_new_n37_), .Y(new_new_n638_));
  NA2        g0616(.A(i_4_), .B(i_8_), .Y(new_new_n639_));
  AOI210     g0617(.A0(new_new_n639_), .A1(new_new_n316_), .B0(new_new_n638_), .Y(new_new_n640_));
  OAI220     g0618(.A0(new_new_n640_), .A1(new_new_n636_), .B0(new_new_n637_), .B1(i_13_), .Y(new_new_n641_));
  NO4        g0619(.A(new_new_n641_), .B(new_new_n635_), .C(new_new_n631_), .D(new_new_n625_), .Y(new_new_n642_));
  AOI210     g0620(.A0(new_new_n132_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n643_));
  AOI210     g0621(.A0(new_new_n643_), .A1(new_new_n245_), .B0(new_new_n166_), .Y(new_new_n644_));
  OR2        g0622(.A(i_6_), .B(i_10_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n645_), .B(new_new_n23_), .Y(new_new_n646_));
  OR3        g0624(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n647_));
  NO3        g0625(.A(new_new_n647_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n648_));
  INV        g0626(.A(new_new_n207_), .Y(new_new_n649_));
  NO2        g0627(.A(new_new_n648_), .B(new_new_n646_), .Y(new_new_n650_));
  OA220      g0628(.A0(new_new_n650_), .A1(new_new_n614_), .B0(new_new_n644_), .B1(new_new_n276_), .Y(new_new_n651_));
  AOI210     g0629(.A0(new_new_n651_), .A1(new_new_n642_), .B0(new_new_n64_), .Y(new_new_n652_));
  NOi21      g0630(.An(i_11_), .B(i_7_), .Y(new_new_n653_));
  AO210      g0631(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n654_), .B(new_new_n653_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n655_), .B(new_new_n214_), .Y(new_new_n656_));
  NA3        g0634(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n657_));
  NAi31      g0635(.An(new_new_n657_), .B(new_new_n224_), .C(i_11_), .Y(new_new_n658_));
  AOI210     g0636(.A0(new_new_n658_), .A1(new_new_n656_), .B0(new_new_n64_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n660_));
  AO210      g0638(.A0(new_new_n660_), .A1(new_new_n398_), .B0(new_new_n41_), .Y(new_new_n661_));
  NO3        g0639(.A(new_new_n267_), .B(new_new_n216_), .C(new_new_n629_), .Y(new_new_n662_));
  OAI210     g0640(.A0(new_new_n662_), .A1(new_new_n234_), .B0(new_new_n64_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n433_), .B(new_new_n31_), .Y(new_new_n664_));
  OR2        g0642(.A(new_new_n216_), .B(new_new_n111_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n665_), .B(new_new_n664_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n64_), .B(i_9_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n667_), .B(i_4_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n668_), .B(new_new_n666_), .Y(new_new_n669_));
  NO2        g0647(.A(i_1_), .B(i_12_), .Y(new_new_n670_));
  NA3        g0648(.A(new_new_n670_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n671_));
  NA4        g0649(.A(new_new_n671_), .B(new_new_n669_), .C(new_new_n663_), .D(new_new_n661_), .Y(new_new_n672_));
  OAI210     g0650(.A0(new_new_n672_), .A1(new_new_n659_), .B0(i_6_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n245_), .B(new_new_n87_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(i_11_), .Y(new_new_n675_));
  INV        g0653(.A(new_new_n480_), .Y(new_new_n676_));
  NO4        g0654(.A(new_new_n224_), .B(new_new_n132_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n677_));
  NA2        g0655(.A(new_new_n677_), .B(new_new_n667_), .Y(new_new_n678_));
  NA2        g0656(.A(new_new_n245_), .B(i_6_), .Y(new_new_n679_));
  NO3        g0657(.A(new_new_n645_), .B(new_new_n241_), .C(new_new_n23_), .Y(new_new_n680_));
  AOI210     g0658(.A0(i_1_), .A1(new_new_n268_), .B0(new_new_n680_), .Y(new_new_n681_));
  OAI210     g0659(.A0(new_new_n681_), .A1(new_new_n45_), .B0(new_new_n678_), .Y(new_new_n682_));
  NA3        g0660(.A(new_new_n565_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n142_), .B(i_9_), .Y(new_new_n684_));
  NA3        g0662(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n47_), .B(i_1_), .Y(new_new_n686_));
  NA3        g0664(.A(new_new_n686_), .B(new_new_n275_), .C(new_new_n45_), .Y(new_new_n687_));
  OAI220     g0665(.A0(new_new_n687_), .A1(new_new_n685_), .B0(new_new_n684_), .B1(new_new_n1112_), .Y(new_new_n688_));
  NA3        g0666(.A(new_new_n667_), .B(new_new_n329_), .C(i_6_), .Y(new_new_n689_));
  NO2        g0667(.A(new_new_n689_), .B(new_new_n23_), .Y(new_new_n690_));
  AOI210     g0668(.A0(new_new_n502_), .A1(new_new_n442_), .B0(new_new_n250_), .Y(new_new_n691_));
  NO2        g0669(.A(new_new_n691_), .B(new_new_n636_), .Y(new_new_n692_));
  NAi21      g0670(.An(new_new_n683_), .B(new_new_n94_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n686_), .B(new_new_n275_), .Y(new_new_n694_));
  NO2        g0672(.A(i_11_), .B(new_new_n37_), .Y(new_new_n695_));
  NA2        g0673(.A(new_new_n695_), .B(new_new_n24_), .Y(new_new_n696_));
  OAI210     g0674(.A0(new_new_n696_), .A1(new_new_n694_), .B0(new_new_n693_), .Y(new_new_n697_));
  OR4        g0675(.A(new_new_n697_), .B(new_new_n692_), .C(new_new_n690_), .D(new_new_n688_), .Y(new_new_n698_));
  NO3        g0676(.A(new_new_n698_), .B(new_new_n682_), .C(new_new_n676_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n245_), .B(new_new_n104_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n700_), .B(new_new_n653_), .Y(new_new_n701_));
  NA2        g0679(.A(new_new_n701_), .B(i_1_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n702_), .B(new_new_n647_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n703_), .B(new_new_n47_), .Y(new_new_n704_));
  NA2        g0682(.A(i_3_), .B(new_new_n200_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n118_), .Y(new_new_n706_));
  AN2        g0684(.A(new_new_n706_), .B(new_new_n571_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n241_), .B(new_new_n45_), .Y(new_new_n708_));
  NO3        g0686(.A(new_new_n708_), .B(new_new_n319_), .C(new_new_n246_), .Y(new_new_n709_));
  NO2        g0687(.A(new_new_n121_), .B(new_new_n37_), .Y(new_new_n710_));
  NO2        g0688(.A(new_new_n710_), .B(i_6_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n87_), .B(i_9_), .Y(new_new_n712_));
  NO2        g0690(.A(new_new_n712_), .B(new_new_n64_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n713_), .B(new_new_n670_), .Y(new_new_n714_));
  NO4        g0692(.A(new_new_n714_), .B(new_new_n711_), .C(new_new_n709_), .D(i_4_), .Y(new_new_n715_));
  NA2        g0693(.A(i_1_), .B(i_3_), .Y(new_new_n716_));
  NO2        g0694(.A(new_new_n481_), .B(new_new_n95_), .Y(new_new_n717_));
  AOI210     g0695(.A0(new_new_n708_), .A1(new_new_n603_), .B0(new_new_n717_), .Y(new_new_n718_));
  NO2        g0696(.A(new_new_n718_), .B(new_new_n716_), .Y(new_new_n719_));
  NO3        g0697(.A(new_new_n719_), .B(new_new_n715_), .C(new_new_n707_), .Y(new_new_n720_));
  NA4        g0698(.A(new_new_n720_), .B(new_new_n704_), .C(new_new_n699_), .D(new_new_n673_), .Y(new_new_n721_));
  NO3        g0699(.A(new_new_n503_), .B(i_3_), .C(i_7_), .Y(new_new_n722_));
  NOi21      g0700(.An(new_new_n722_), .B(i_10_), .Y(new_new_n723_));
  OA210      g0701(.A0(new_new_n723_), .A1(new_new_n254_), .B0(new_new_n87_), .Y(new_new_n724_));
  NA2        g0702(.A(new_new_n391_), .B(new_new_n390_), .Y(new_new_n725_));
  NA3        g0703(.A(new_new_n510_), .B(new_new_n546_), .C(new_new_n47_), .Y(new_new_n726_));
  NO3        g0704(.A(new_new_n504_), .B(new_new_n639_), .C(new_new_n87_), .Y(new_new_n727_));
  NA2        g0705(.A(new_new_n727_), .B(new_new_n25_), .Y(new_new_n728_));
  NA3        g0706(.A(new_new_n166_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n729_));
  NA4        g0707(.A(new_new_n729_), .B(new_new_n728_), .C(new_new_n726_), .D(new_new_n725_), .Y(new_new_n730_));
  OAI210     g0708(.A0(new_new_n730_), .A1(new_new_n724_), .B0(i_1_), .Y(new_new_n731_));
  AOI210     g0709(.A0(new_new_n275_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n732_));
  NO2        g0710(.A(new_new_n389_), .B(i_2_), .Y(new_new_n733_));
  NA2        g0711(.A(new_new_n733_), .B(new_new_n732_), .Y(new_new_n734_));
  OAI210     g0712(.A0(new_new_n689_), .A1(new_new_n471_), .B0(new_new_n734_), .Y(new_new_n735_));
  INV        g0713(.A(new_new_n735_), .Y(new_new_n736_));
  AOI210     g0714(.A0(new_new_n736_), .A1(new_new_n731_), .B0(i_13_), .Y(new_new_n737_));
  OR2        g0715(.A(i_11_), .B(i_7_), .Y(new_new_n738_));
  NA3        g0716(.A(new_new_n738_), .B(new_new_n109_), .C(new_new_n142_), .Y(new_new_n739_));
  AOI220     g0717(.A0(new_new_n496_), .A1(new_new_n166_), .B0(new_new_n474_), .B1(new_new_n142_), .Y(new_new_n740_));
  OAI210     g0718(.A0(new_new_n740_), .A1(new_new_n45_), .B0(new_new_n739_), .Y(new_new_n741_));
  AOI210     g0719(.A0(new_new_n685_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n1111_), .B(new_new_n95_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n741_), .A1(new_new_n346_), .B0(new_new_n743_), .Y(new_new_n744_));
  NA2        g0722(.A(new_new_n118_), .B(new_new_n111_), .Y(new_new_n745_));
  AOI220     g0723(.A0(new_new_n745_), .A1(new_new_n73_), .B0(new_new_n406_), .B1(new_new_n686_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n746_), .B(new_new_n251_), .Y(new_new_n747_));
  AOI210     g0725(.A0(new_new_n471_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n131_), .B(i_13_), .Y(new_new_n749_));
  NO2        g0727(.A(new_new_n685_), .B(new_new_n118_), .Y(new_new_n750_));
  NO2        g0728(.A(new_new_n749_), .B(new_new_n732_), .Y(new_new_n751_));
  NO3        g0729(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n26_), .B(new_new_n200_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n753_), .B(i_7_), .Y(new_new_n754_));
  NO3        g0732(.A(new_new_n504_), .B(new_new_n245_), .C(new_new_n87_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n755_), .A1(new_new_n754_), .B0(new_new_n752_), .Y(new_new_n756_));
  AOI220     g0734(.A0(new_new_n406_), .A1(new_new_n686_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n757_));
  OAI220     g0735(.A0(new_new_n757_), .A1(new_new_n634_), .B0(new_new_n756_), .B1(new_new_n649_), .Y(new_new_n758_));
  NO3        g0736(.A(new_new_n758_), .B(new_new_n751_), .C(new_new_n747_), .Y(new_new_n759_));
  OR2        g0737(.A(i_11_), .B(i_6_), .Y(new_new_n760_));
  NA3        g0738(.A(new_new_n633_), .B(new_new_n753_), .C(i_7_), .Y(new_new_n761_));
  NO2        g0739(.A(new_new_n761_), .B(new_new_n760_), .Y(new_new_n762_));
  NA3        g0740(.A(new_new_n433_), .B(new_new_n638_), .C(new_new_n100_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n675_), .B(i_13_), .Y(new_new_n764_));
  NAi21      g0742(.An(i_11_), .B(i_12_), .Y(new_new_n765_));
  NOi41      g0743(.An(new_new_n114_), .B(new_new_n765_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n766_));
  NO3        g0744(.A(new_new_n504_), .B(new_new_n615_), .C(new_new_n639_), .Y(new_new_n767_));
  AOI220     g0745(.A0(new_new_n767_), .A1(new_new_n323_), .B0(new_new_n766_), .B1(new_new_n47_), .Y(new_new_n768_));
  NA3        g0746(.A(new_new_n768_), .B(new_new_n764_), .C(new_new_n763_), .Y(new_new_n769_));
  OAI210     g0747(.A0(new_new_n769_), .A1(new_new_n762_), .B0(new_new_n64_), .Y(new_new_n770_));
  NO2        g0748(.A(i_2_), .B(i_12_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n388_), .B(new_new_n771_), .Y(new_new_n772_));
  NA2        g0750(.A(i_8_), .B(new_new_n25_), .Y(new_new_n773_));
  NO3        g0751(.A(new_new_n773_), .B(new_new_n404_), .C(new_new_n633_), .Y(new_new_n774_));
  OAI210     g0752(.A0(new_new_n774_), .A1(new_new_n390_), .B0(new_new_n388_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n132_), .B(i_2_), .Y(new_new_n776_));
  NA2        g0754(.A(new_new_n776_), .B(new_new_n670_), .Y(new_new_n777_));
  NA3        g0755(.A(new_new_n777_), .B(new_new_n775_), .C(new_new_n772_), .Y(new_new_n778_));
  NA3        g0756(.A(new_new_n778_), .B(new_new_n46_), .C(new_new_n233_), .Y(new_new_n779_));
  NA4        g0757(.A(new_new_n779_), .B(new_new_n770_), .C(new_new_n759_), .D(new_new_n744_), .Y(new_new_n780_));
  OR4        g0758(.A(new_new_n780_), .B(new_new_n737_), .C(new_new_n721_), .D(new_new_n652_), .Y(men5));
  AOI210     g0759(.A0(new_new_n701_), .A1(new_new_n278_), .B0(new_new_n440_), .Y(new_new_n782_));
  AN2        g0760(.A(new_new_n24_), .B(i_10_), .Y(new_new_n783_));
  NA3        g0761(.A(new_new_n783_), .B(new_new_n771_), .C(new_new_n111_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n634_), .B(i_11_), .Y(new_new_n785_));
  OAI210     g0763(.A0(new_new_n638_), .A1(new_new_n90_), .B0(new_new_n785_), .Y(new_new_n786_));
  NA3        g0764(.A(new_new_n786_), .B(new_new_n784_), .C(new_new_n782_), .Y(new_new_n787_));
  NO3        g0765(.A(i_11_), .B(new_new_n245_), .C(i_13_), .Y(new_new_n788_));
  NO2        g0766(.A(new_new_n128_), .B(new_new_n23_), .Y(new_new_n789_));
  NA2        g0767(.A(i_12_), .B(i_8_), .Y(new_new_n790_));
  OAI210     g0768(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n790_), .Y(new_new_n791_));
  INV        g0769(.A(new_new_n470_), .Y(new_new_n792_));
  AOI220     g0770(.A0(new_new_n329_), .A1(new_new_n607_), .B0(new_new_n791_), .B1(new_new_n789_), .Y(new_new_n793_));
  INV        g0771(.A(new_new_n793_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n794_), .B(new_new_n787_), .Y(new_new_n795_));
  INV        g0773(.A(new_new_n177_), .Y(new_new_n796_));
  INV        g0774(.A(new_new_n254_), .Y(new_new_n797_));
  OAI210     g0775(.A0(new_new_n733_), .A1(new_new_n472_), .B0(new_new_n114_), .Y(new_new_n798_));
  AOI210     g0776(.A0(new_new_n798_), .A1(new_new_n797_), .B0(new_new_n796_), .Y(new_new_n799_));
  NO2        g0777(.A(new_new_n481_), .B(new_new_n26_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n800_), .B(new_new_n442_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n801_), .B(i_2_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n802_), .Y(new_new_n803_));
  AOI210     g0781(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n439_), .Y(new_new_n804_));
  AOI210     g0782(.A0(new_new_n804_), .A1(new_new_n803_), .B0(new_new_n799_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n197_), .B(new_new_n129_), .Y(new_new_n806_));
  OAI210     g0784(.A0(new_new_n806_), .A1(new_new_n789_), .B0(i_2_), .Y(new_new_n807_));
  INV        g0785(.A(new_new_n178_), .Y(new_new_n808_));
  NO3        g0786(.A(new_new_n654_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n809_));
  AOI210     g0787(.A0(new_new_n808_), .A1(new_new_n90_), .B0(new_new_n809_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n810_), .A1(new_new_n807_), .B0(new_new_n200_), .Y(new_new_n811_));
  OA210      g0789(.A0(new_new_n655_), .A1(new_new_n130_), .B0(i_13_), .Y(new_new_n812_));
  NA2        g0790(.A(new_new_n207_), .B(new_new_n210_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n156_), .B(new_new_n629_), .Y(new_new_n814_));
  AOI210     g0792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n393_), .Y(new_new_n815_));
  AOI210     g0793(.A0(new_new_n216_), .A1(new_new_n152_), .B0(new_new_n546_), .Y(new_new_n816_));
  OAI210     g0794(.A0(new_new_n816_), .A1(new_new_n234_), .B0(new_new_n442_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n105_), .B(new_new_n45_), .Y(new_new_n818_));
  INV        g0796(.A(new_new_n312_), .Y(new_new_n819_));
  NA4        g0797(.A(new_new_n819_), .B(new_new_n316_), .C(new_new_n128_), .D(new_new_n43_), .Y(new_new_n820_));
  OAI210     g0798(.A0(new_new_n820_), .A1(new_new_n818_), .B0(new_new_n817_), .Y(new_new_n821_));
  NO4        g0799(.A(new_new_n821_), .B(new_new_n815_), .C(new_new_n812_), .D(new_new_n811_), .Y(new_new_n822_));
  NA2        g0800(.A(new_new_n607_), .B(new_new_n28_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n788_), .B(new_new_n285_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n824_), .B(new_new_n823_), .Y(new_new_n825_));
  NO2        g0803(.A(new_new_n63_), .B(i_12_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n826_), .B(new_new_n130_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n827_), .B(new_new_n629_), .Y(new_new_n828_));
  AOI220     g0806(.A0(new_new_n828_), .A1(new_new_n36_), .B0(new_new_n825_), .B1(new_new_n47_), .Y(new_new_n829_));
  NA4        g0807(.A(new_new_n829_), .B(new_new_n822_), .C(new_new_n805_), .D(new_new_n795_), .Y(men6));
  NO3        g0808(.A(new_new_n263_), .B(new_new_n318_), .C(i_1_), .Y(new_new_n831_));
  NO2        g0809(.A(new_new_n192_), .B(new_new_n143_), .Y(new_new_n832_));
  OAI210     g0810(.A0(new_new_n832_), .A1(new_new_n831_), .B0(new_new_n776_), .Y(new_new_n833_));
  NA4        g0811(.A(new_new_n410_), .B(new_new_n509_), .C(new_new_n72_), .D(new_new_n104_), .Y(new_new_n834_));
  INV        g0812(.A(new_new_n834_), .Y(new_new_n835_));
  NO2        g0813(.A(i_11_), .B(i_9_), .Y(new_new_n836_));
  NO2        g0814(.A(new_new_n835_), .B(new_new_n341_), .Y(new_new_n837_));
  AO210      g0815(.A0(new_new_n837_), .A1(new_new_n833_), .B0(i_12_), .Y(new_new_n838_));
  NA2        g0816(.A(new_new_n394_), .B(new_new_n349_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n615_), .B(new_new_n64_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n723_), .B(new_new_n72_), .Y(new_new_n841_));
  NA4        g0819(.A(new_new_n660_), .B(new_new_n841_), .C(new_new_n840_), .D(new_new_n839_), .Y(new_new_n842_));
  INV        g0820(.A(new_new_n204_), .Y(new_new_n843_));
  AOI220     g0821(.A0(new_new_n843_), .A1(new_new_n836_), .B0(new_new_n842_), .B1(new_new_n74_), .Y(new_new_n844_));
  INV        g0822(.A(new_new_n340_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n76_), .B(new_new_n135_), .Y(new_new_n846_));
  INV        g0824(.A(new_new_n128_), .Y(new_new_n847_));
  NA2        g0825(.A(new_new_n847_), .B(new_new_n47_), .Y(new_new_n848_));
  AOI210     g0826(.A0(new_new_n848_), .A1(new_new_n846_), .B0(new_new_n845_), .Y(new_new_n849_));
  NO2        g0827(.A(new_new_n545_), .B(new_new_n192_), .Y(new_new_n850_));
  NO2        g0828(.A(new_new_n32_), .B(i_11_), .Y(new_new_n851_));
  NA3        g0829(.A(new_new_n851_), .B(new_new_n500_), .C(new_new_n410_), .Y(new_new_n852_));
  NAi32      g0830(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n853_));
  AOI210     g0831(.A0(new_new_n760_), .A1(new_new_n88_), .B0(new_new_n853_), .Y(new_new_n854_));
  OAI210     g0832(.A0(new_new_n722_), .A1(new_new_n595_), .B0(new_new_n594_), .Y(new_new_n855_));
  NAi31      g0833(.An(new_new_n854_), .B(new_new_n855_), .C(new_new_n852_), .Y(new_new_n856_));
  OR3        g0834(.A(new_new_n856_), .B(new_new_n850_), .C(new_new_n849_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n738_), .B(i_2_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n859_));
  OAI210     g0837(.A0(new_new_n859_), .A1(new_new_n432_), .B0(new_new_n378_), .Y(new_new_n860_));
  NA2        g0838(.A(new_new_n860_), .B(new_new_n858_), .Y(new_new_n861_));
  AO220      g0839(.A0(new_new_n377_), .A1(new_new_n367_), .B0(new_new_n418_), .B1(new_new_n629_), .Y(new_new_n862_));
  NA3        g0840(.A(new_new_n862_), .B(new_new_n264_), .C(i_7_), .Y(new_new_n863_));
  OR2        g0841(.A(new_new_n655_), .B(new_new_n472_), .Y(new_new_n864_));
  NA3        g0842(.A(new_new_n864_), .B(new_new_n151_), .C(new_new_n70_), .Y(new_new_n865_));
  AO210      g0843(.A0(new_new_n520_), .A1(new_new_n792_), .B0(new_new_n36_), .Y(new_new_n866_));
  NA4        g0844(.A(new_new_n866_), .B(new_new_n865_), .C(new_new_n863_), .D(new_new_n861_), .Y(new_new_n867_));
  OAI210     g0845(.A0(new_new_n674_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n868_), .B(new_new_n594_), .Y(new_new_n869_));
  NA3        g0847(.A(new_new_n393_), .B(new_new_n247_), .C(new_new_n151_), .Y(new_new_n870_));
  OAI210     g0848(.A0(new_new_n418_), .A1(new_new_n211_), .B0(new_new_n71_), .Y(new_new_n871_));
  NA4        g0849(.A(new_new_n871_), .B(new_new_n870_), .C(new_new_n869_), .D(new_new_n637_), .Y(new_new_n872_));
  AO210      g0850(.A0(new_new_n546_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n873_));
  NA3        g0851(.A(new_new_n873_), .B(new_new_n510_), .C(new_new_n227_), .Y(new_new_n874_));
  AOI210     g0852(.A0(new_new_n472_), .A1(new_new_n470_), .B0(new_new_n593_), .Y(new_new_n875_));
  NO2        g0853(.A(new_new_n645_), .B(new_new_n105_), .Y(new_new_n876_));
  OAI210     g0854(.A0(new_new_n876_), .A1(new_new_n115_), .B0(new_new_n430_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n253_), .B(new_new_n47_), .Y(new_new_n878_));
  NA3        g0856(.A(new_new_n877_), .B(new_new_n875_), .C(new_new_n874_), .Y(new_new_n879_));
  NO4        g0857(.A(new_new_n879_), .B(new_new_n872_), .C(new_new_n867_), .D(new_new_n857_), .Y(new_new_n880_));
  NA4        g0858(.A(new_new_n880_), .B(new_new_n844_), .C(new_new_n838_), .D(new_new_n400_), .Y(men3));
  NA2        g0859(.A(i_6_), .B(i_7_), .Y(new_new_n882_));
  NO2        g0860(.A(new_new_n882_), .B(i_0_), .Y(new_new_n883_));
  NO2        g0861(.A(i_11_), .B(new_new_n245_), .Y(new_new_n884_));
  OAI210     g0862(.A0(new_new_n883_), .A1(new_new_n300_), .B0(new_new_n884_), .Y(new_new_n885_));
  NO2        g0863(.A(new_new_n885_), .B(new_new_n200_), .Y(new_new_n886_));
  NO3        g0864(.A(new_new_n477_), .B(new_new_n92_), .C(new_new_n45_), .Y(new_new_n887_));
  OA210      g0865(.A0(new_new_n887_), .A1(new_new_n886_), .B0(new_new_n180_), .Y(new_new_n888_));
  NA3        g0866(.A(new_new_n870_), .B(new_new_n637_), .C(new_new_n392_), .Y(new_new_n889_));
  NA2        g0867(.A(new_new_n889_), .B(new_new_n40_), .Y(new_new_n890_));
  NOi21      g0868(.An(new_new_n99_), .B(new_new_n801_), .Y(new_new_n891_));
  NO3        g0869(.A(new_new_n665_), .B(new_new_n481_), .C(new_new_n135_), .Y(new_new_n892_));
  NA2        g0870(.A(new_new_n433_), .B(new_new_n46_), .Y(new_new_n893_));
  AN2        g0871(.A(new_new_n479_), .B(new_new_n56_), .Y(new_new_n894_));
  NO3        g0872(.A(new_new_n894_), .B(new_new_n892_), .C(new_new_n891_), .Y(new_new_n895_));
  AOI210     g0873(.A0(new_new_n895_), .A1(new_new_n890_), .B0(new_new_n49_), .Y(new_new_n896_));
  NO4        g0874(.A(new_new_n396_), .B(new_new_n403_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n192_), .B(new_new_n603_), .Y(new_new_n898_));
  NOi31      g0876(.An(new_new_n898_), .B(new_new_n897_), .C(new_new_n39_), .Y(new_new_n899_));
  NA2        g0877(.A(new_new_n748_), .B(new_new_n712_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n347_), .B(new_new_n460_), .Y(new_new_n901_));
  OAI220     g0879(.A0(new_new_n901_), .A1(new_new_n900_), .B0(new_new_n899_), .B1(new_new_n64_), .Y(new_new_n902_));
  NOi21      g0880(.An(i_5_), .B(i_9_), .Y(new_new_n903_));
  NA2        g0881(.A(new_new_n903_), .B(new_new_n468_), .Y(new_new_n904_));
  AOI210     g0882(.A0(new_new_n275_), .A1(new_new_n502_), .B0(new_new_n727_), .Y(new_new_n905_));
  NO3        g0883(.A(new_new_n436_), .B(new_new_n275_), .C(new_new_n74_), .Y(new_new_n906_));
  NO2        g0884(.A(new_new_n181_), .B(new_new_n152_), .Y(new_new_n907_));
  AOI210     g0885(.A0(new_new_n907_), .A1(new_new_n253_), .B0(new_new_n906_), .Y(new_new_n908_));
  OAI220     g0886(.A0(new_new_n908_), .A1(new_new_n187_), .B0(new_new_n905_), .B1(new_new_n904_), .Y(new_new_n909_));
  NO4        g0887(.A(new_new_n909_), .B(new_new_n902_), .C(new_new_n896_), .D(new_new_n888_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n192_), .B(new_new_n24_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n710_), .B(new_new_n626_), .Y(new_new_n912_));
  NO2        g0890(.A(new_new_n912_), .B(new_new_n911_), .Y(new_new_n913_));
  NA2        g0891(.A(new_new_n323_), .B(new_new_n133_), .Y(new_new_n914_));
  NAi21      g0892(.An(new_new_n167_), .B(new_new_n460_), .Y(new_new_n915_));
  OAI220     g0893(.A0(new_new_n915_), .A1(new_new_n878_), .B0(new_new_n914_), .B1(new_new_n421_), .Y(new_new_n916_));
  NO2        g0894(.A(new_new_n916_), .B(new_new_n913_), .Y(new_new_n917_));
  NO2        g0895(.A(new_new_n410_), .B(new_new_n304_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n918_), .B(new_new_n750_), .Y(new_new_n919_));
  NA2        g0897(.A(new_new_n604_), .B(i_0_), .Y(new_new_n920_));
  NO3        g0898(.A(new_new_n920_), .B(new_new_n405_), .C(new_new_n90_), .Y(new_new_n921_));
  NO4        g0899(.A(new_new_n620_), .B(new_new_n224_), .C(new_new_n439_), .D(new_new_n432_), .Y(new_new_n922_));
  AOI210     g0900(.A0(new_new_n922_), .A1(i_11_), .B0(new_new_n921_), .Y(new_new_n923_));
  INV        g0901(.A(new_new_n500_), .Y(new_new_n924_));
  AN2        g0902(.A(new_new_n99_), .B(new_new_n252_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n788_), .B(new_new_n341_), .Y(new_new_n926_));
  AOI210     g0904(.A0(new_new_n510_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n927_));
  OAI220     g0905(.A0(new_new_n927_), .A1(new_new_n926_), .B0(new_new_n696_), .B1(new_new_n567_), .Y(new_new_n928_));
  NA2        g0906(.A(i_0_), .B(i_10_), .Y(new_new_n929_));
  OAI210     g0907(.A0(new_new_n929_), .A1(new_new_n87_), .B0(new_new_n570_), .Y(new_new_n930_));
  NO4        g0908(.A(new_new_n118_), .B(new_new_n59_), .C(new_new_n705_), .D(i_5_), .Y(new_new_n931_));
  AN2        g0909(.A(new_new_n931_), .B(new_new_n930_), .Y(new_new_n932_));
  AOI220     g0910(.A0(new_new_n347_), .A1(new_new_n101_), .B0(new_new_n192_), .B1(new_new_n85_), .Y(new_new_n933_));
  NA2        g0911(.A(new_new_n598_), .B(i_4_), .Y(new_new_n934_));
  NA2        g0912(.A(new_new_n195_), .B(new_new_n210_), .Y(new_new_n935_));
  OAI220     g0913(.A0(new_new_n935_), .A1(new_new_n926_), .B0(new_new_n934_), .B1(new_new_n933_), .Y(new_new_n936_));
  NO4        g0914(.A(new_new_n936_), .B(new_new_n932_), .C(new_new_n928_), .D(new_new_n925_), .Y(new_new_n937_));
  NA4        g0915(.A(new_new_n937_), .B(new_new_n923_), .C(new_new_n919_), .D(new_new_n917_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n939_));
  NA2        g0917(.A(i_11_), .B(i_9_), .Y(new_new_n940_));
  NO3        g0918(.A(i_12_), .B(new_new_n940_), .C(new_new_n636_), .Y(new_new_n941_));
  AO220      g0919(.A0(new_new_n941_), .A1(new_new_n939_), .B0(new_new_n277_), .B1(new_new_n89_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n49_), .B(i_7_), .Y(new_new_n943_));
  NA2        g0921(.A(new_new_n415_), .B(new_new_n185_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n944_), .B(new_new_n165_), .Y(new_new_n945_));
  NO2        g0923(.A(new_new_n940_), .B(new_new_n74_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n181_), .B(i_0_), .Y(new_new_n947_));
  INV        g0925(.A(new_new_n947_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n500_), .B(new_new_n239_), .Y(new_new_n949_));
  AOI210     g0927(.A0(new_new_n391_), .A1(new_new_n42_), .B0(new_new_n429_), .Y(new_new_n950_));
  OAI220     g0928(.A0(new_new_n950_), .A1(new_new_n904_), .B0(new_new_n949_), .B1(new_new_n948_), .Y(new_new_n951_));
  NO3        g0929(.A(new_new_n951_), .B(new_new_n945_), .C(new_new_n942_), .Y(new_new_n952_));
  NA2        g0930(.A(new_new_n695_), .B(new_new_n125_), .Y(new_new_n953_));
  NO2        g0931(.A(i_6_), .B(new_new_n953_), .Y(new_new_n954_));
  AOI210     g0932(.A0(new_new_n471_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n177_), .B(new_new_n106_), .Y(new_new_n956_));
  NOi32      g0934(.An(new_new_n955_), .Bn(new_new_n195_), .C(new_new_n956_), .Y(new_new_n957_));
  AOI210     g0935(.A0(new_new_n638_), .A1(new_new_n341_), .B0(new_new_n252_), .Y(new_new_n958_));
  NO2        g0936(.A(new_new_n958_), .B(new_new_n893_), .Y(new_new_n959_));
  NO3        g0937(.A(new_new_n959_), .B(new_new_n957_), .C(new_new_n954_), .Y(new_new_n960_));
  NOi21      g0938(.An(i_7_), .B(i_5_), .Y(new_new_n961_));
  NOi31      g0939(.An(new_new_n961_), .B(i_0_), .C(new_new_n765_), .Y(new_new_n962_));
  NA3        g0940(.A(new_new_n962_), .B(new_new_n404_), .C(i_6_), .Y(new_new_n963_));
  OA210      g0941(.A0(new_new_n956_), .A1(new_new_n545_), .B0(new_new_n963_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n424_), .B(new_new_n380_), .C(new_new_n376_), .Y(new_new_n965_));
  NO2        g0943(.A(new_new_n269_), .B(new_new_n330_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n765_), .B(new_new_n266_), .Y(new_new_n967_));
  AOI210     g0945(.A0(new_new_n967_), .A1(new_new_n966_), .B0(new_new_n965_), .Y(new_new_n968_));
  NA4        g0946(.A(new_new_n968_), .B(new_new_n964_), .C(new_new_n960_), .D(new_new_n952_), .Y(new_new_n969_));
  NO2        g0947(.A(new_new_n911_), .B(new_new_n248_), .Y(new_new_n970_));
  AN2        g0948(.A(new_new_n346_), .B(new_new_n341_), .Y(new_new_n971_));
  AO220      g0949(.A0(new_new_n971_), .A1(new_new_n907_), .B0(new_new_n362_), .B1(new_new_n27_), .Y(new_new_n972_));
  OAI210     g0950(.A0(new_new_n972_), .A1(new_new_n970_), .B0(i_10_), .Y(new_new_n973_));
  OA210      g0951(.A0(new_new_n500_), .A1(new_new_n231_), .B0(new_new_n499_), .Y(new_new_n974_));
  NA3        g0952(.A(new_new_n499_), .B(new_new_n433_), .C(new_new_n46_), .Y(new_new_n975_));
  OAI210     g0953(.A0(new_new_n915_), .A1(new_new_n924_), .B0(new_new_n975_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n946_), .B(new_new_n316_), .Y(new_new_n977_));
  NA2        g0955(.A(new_new_n194_), .B(new_new_n977_), .Y(new_new_n978_));
  AOI220     g0956(.A0(new_new_n978_), .A1(new_new_n500_), .B0(new_new_n976_), .B1(new_new_n74_), .Y(new_new_n979_));
  NA3        g0957(.A(new_new_n859_), .B(new_new_n402_), .C(new_new_n674_), .Y(new_new_n980_));
  NA2        g0958(.A(new_new_n95_), .B(new_new_n45_), .Y(new_new_n981_));
  NO2        g0959(.A(new_new_n76_), .B(new_new_n790_), .Y(new_new_n982_));
  AOI220     g0960(.A0(new_new_n982_), .A1(new_new_n981_), .B0(new_new_n180_), .B1(new_new_n626_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n983_), .A1(new_new_n980_), .B0(new_new_n48_), .Y(new_new_n984_));
  NO3        g0962(.A(new_new_n620_), .B(new_new_n375_), .C(new_new_n24_), .Y(new_new_n985_));
  INV        g0963(.A(new_new_n985_), .Y(new_new_n986_));
  NAi21      g0964(.An(i_9_), .B(i_5_), .Y(new_new_n987_));
  NO2        g0965(.A(new_new_n632_), .B(new_new_n108_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n988_), .B(i_0_), .Y(new_new_n989_));
  OAI220     g0967(.A0(new_new_n989_), .A1(new_new_n87_), .B0(new_new_n986_), .B1(new_new_n178_), .Y(new_new_n990_));
  NO2        g0968(.A(new_new_n990_), .B(new_new_n984_), .Y(new_new_n991_));
  NA3        g0969(.A(new_new_n991_), .B(new_new_n979_), .C(new_new_n973_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n992_), .B(new_new_n969_), .C(new_new_n938_), .Y(new_new_n993_));
  NO2        g0971(.A(i_0_), .B(new_new_n765_), .Y(new_new_n994_));
  NA2        g0972(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n929_), .B(new_new_n995_), .Y(new_new_n996_));
  NO3        g0974(.A(new_new_n108_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n997_));
  AO220      g0975(.A0(new_new_n997_), .A1(new_new_n996_), .B0(new_new_n994_), .B1(new_new_n180_), .Y(new_new_n998_));
  AOI210     g0976(.A0(new_new_n840_), .A1(new_new_n725_), .B0(new_new_n956_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n998_), .A1(new_new_n364_), .B0(new_new_n999_), .Y(new_new_n1000_));
  NA2        g0978(.A(new_new_n776_), .B(new_new_n150_), .Y(new_new_n1001_));
  INV        g0979(.A(new_new_n1001_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n1002_), .B(new_new_n712_), .C(new_new_n74_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n855_), .B(new_new_n424_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n883_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n884_), .B(i_9_), .Y(new_new_n1006_));
  AOI210     g0984(.A0(new_new_n1005_), .A1(new_new_n526_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n253_), .A1(i_9_), .B0(new_new_n238_), .Y(new_new_n1008_));
  AOI210     g0986(.A0(new_new_n1008_), .A1(new_new_n920_), .B0(new_new_n158_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n1009_), .B(new_new_n1007_), .C(new_new_n1004_), .Y(new_new_n1010_));
  NA3        g0988(.A(new_new_n1010_), .B(new_new_n1003_), .C(new_new_n1000_), .Y(new_new_n1011_));
  NA2        g0989(.A(new_new_n971_), .B(new_new_n393_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n311_), .A1(new_new_n167_), .B0(new_new_n1012_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n1014_));
  NA2        g0992(.A(new_new_n943_), .B(new_new_n514_), .Y(new_new_n1015_));
  AOI210     g0993(.A0(new_new_n1014_), .A1(new_new_n167_), .B0(new_new_n1015_), .Y(new_new_n1016_));
  NO2        g0994(.A(new_new_n1016_), .B(new_new_n1013_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n929_), .B(new_new_n903_), .C(new_new_n197_), .Y(new_new_n1018_));
  AOI220     g0996(.A0(new_new_n1018_), .A1(i_11_), .B0(new_new_n599_), .B1(new_new_n76_), .Y(new_new_n1019_));
  NO3        g0997(.A(new_new_n218_), .B(new_new_n403_), .C(i_0_), .Y(new_new_n1020_));
  OAI210     g0998(.A0(new_new_n1020_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n1021_));
  INV        g0999(.A(new_new_n227_), .Y(new_new_n1022_));
  OAI220     g1000(.A0(new_new_n560_), .A1(new_new_n143_), .B0(new_new_n679_), .B1(new_new_n649_), .Y(new_new_n1023_));
  NA3        g1001(.A(new_new_n1023_), .B(new_new_n419_), .C(new_new_n1022_), .Y(new_new_n1024_));
  NA4        g1002(.A(new_new_n1024_), .B(new_new_n1021_), .C(new_new_n1019_), .D(new_new_n1017_), .Y(new_new_n1025_));
  NO2        g1003(.A(new_new_n251_), .B(new_new_n95_), .Y(new_new_n1026_));
  AOI210     g1004(.A0(new_new_n1026_), .A1(new_new_n994_), .B0(new_new_n112_), .Y(new_new_n1027_));
  AOI220     g1005(.A0(new_new_n961_), .A1(new_new_n514_), .B0(new_new_n883_), .B1(new_new_n168_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n367_), .B(new_new_n182_), .Y(new_new_n1029_));
  OA220      g1007(.A0(new_new_n1029_), .A1(new_new_n1028_), .B0(new_new_n1027_), .B1(i_5_), .Y(new_new_n1030_));
  AOI210     g1008(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n181_), .Y(new_new_n1031_));
  NA2        g1009(.A(new_new_n1031_), .B(new_new_n974_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n646_), .B(new_new_n192_), .C(new_new_n85_), .Y(new_new_n1033_));
  NA2        g1011(.A(new_new_n1033_), .B(new_new_n577_), .Y(new_new_n1034_));
  NA2        g1012(.A(new_new_n519_), .B(new_new_n497_), .Y(new_new_n1035_));
  NO2        g1013(.A(new_new_n1035_), .B(new_new_n1034_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n410_), .B(new_new_n177_), .C(new_new_n176_), .Y(new_new_n1037_));
  NA3        g1015(.A(new_new_n943_), .B(new_new_n300_), .C(new_new_n238_), .Y(new_new_n1038_));
  NA2        g1016(.A(new_new_n1038_), .B(new_new_n1037_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n410_), .B(new_new_n348_), .C(new_new_n230_), .Y(new_new_n1040_));
  OAI210     g1018(.A0(new_new_n898_), .A1(new_new_n683_), .B0(new_new_n1040_), .Y(new_new_n1041_));
  NOi31      g1019(.An(new_new_n409_), .B(new_new_n995_), .C(new_new_n248_), .Y(new_new_n1042_));
  NO3        g1020(.A(new_new_n940_), .B(new_new_n227_), .C(new_new_n197_), .Y(new_new_n1043_));
  NO4        g1021(.A(new_new_n1043_), .B(new_new_n1042_), .C(new_new_n1041_), .D(new_new_n1039_), .Y(new_new_n1044_));
  NA4        g1022(.A(new_new_n1044_), .B(new_new_n1036_), .C(new_new_n1032_), .D(new_new_n1030_), .Y(new_new_n1045_));
  INV        g1023(.A(new_new_n648_), .Y(new_new_n1046_));
  NO3        g1024(.A(new_new_n1046_), .B(new_new_n589_), .C(new_new_n361_), .Y(new_new_n1047_));
  INV        g1025(.A(new_new_n1047_), .Y(new_new_n1048_));
  NA3        g1026(.A(new_new_n316_), .B(i_5_), .C(new_new_n200_), .Y(new_new_n1049_));
  NAi31      g1027(.An(new_new_n250_), .B(new_new_n1049_), .C(new_new_n251_), .Y(new_new_n1050_));
  NO4        g1028(.A(new_new_n248_), .B(new_new_n218_), .C(i_0_), .D(i_12_), .Y(new_new_n1051_));
  AOI220     g1029(.A0(new_new_n1051_), .A1(new_new_n1050_), .B0(new_new_n835_), .B1(new_new_n182_), .Y(new_new_n1052_));
  AN2        g1030(.A(new_new_n929_), .B(new_new_n158_), .Y(new_new_n1053_));
  NO4        g1031(.A(new_new_n1053_), .B(i_12_), .C(new_new_n683_), .D(new_new_n135_), .Y(new_new_n1054_));
  NA2        g1032(.A(new_new_n1054_), .B(new_new_n227_), .Y(new_new_n1055_));
  NA3        g1033(.A(new_new_n101_), .B(new_new_n603_), .C(i_11_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n1056_), .B(new_new_n160_), .Y(new_new_n1057_));
  NA2        g1035(.A(new_new_n65_), .B(new_new_n104_), .Y(new_new_n1058_));
  NO2        g1036(.A(new_new_n1058_), .B(new_new_n1049_), .Y(new_new_n1059_));
  AOI210     g1037(.A0(new_new_n1059_), .A1(new_new_n947_), .B0(new_new_n1057_), .Y(new_new_n1060_));
  NA4        g1038(.A(new_new_n1060_), .B(new_new_n1055_), .C(new_new_n1052_), .D(new_new_n1048_), .Y(new_new_n1061_));
  NO4        g1039(.A(new_new_n1061_), .B(new_new_n1045_), .C(new_new_n1025_), .D(new_new_n1011_), .Y(new_new_n1062_));
  OAI210     g1040(.A0(new_new_n858_), .A1(new_new_n851_), .B0(new_new_n37_), .Y(new_new_n1063_));
  NA3        g1041(.A(new_new_n955_), .B(new_new_n388_), .C(i_5_), .Y(new_new_n1064_));
  NA3        g1042(.A(new_new_n1064_), .B(new_new_n1063_), .C(new_new_n644_), .Y(new_new_n1065_));
  NA2        g1043(.A(new_new_n1065_), .B(new_new_n214_), .Y(new_new_n1066_));
  NA2        g1044(.A(new_new_n193_), .B(new_new_n195_), .Y(new_new_n1067_));
  AO210      g1045(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1067_), .Y(new_new_n1068_));
  OAI210     g1046(.A0(new_new_n648_), .A1(new_new_n646_), .B0(new_new_n329_), .Y(new_new_n1069_));
  NAi31      g1047(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1070_));
  AOI210     g1048(.A0(new_new_n121_), .A1(new_new_n71_), .B0(new_new_n1070_), .Y(new_new_n1071_));
  NO2        g1049(.A(new_new_n1071_), .B(new_new_n680_), .Y(new_new_n1072_));
  NA3        g1050(.A(new_new_n1072_), .B(new_new_n1069_), .C(new_new_n1068_), .Y(new_new_n1073_));
  NO2        g1051(.A(new_new_n486_), .B(new_new_n275_), .Y(new_new_n1074_));
  NO4        g1052(.A(new_new_n241_), .B(new_new_n149_), .C(new_new_n716_), .D(new_new_n37_), .Y(new_new_n1075_));
  NO3        g1053(.A(new_new_n1075_), .B(new_new_n1074_), .C(new_new_n922_), .Y(new_new_n1076_));
  OAI210     g1054(.A0(new_new_n1056_), .A1(new_new_n152_), .B0(new_new_n1076_), .Y(new_new_n1077_));
  AOI210     g1055(.A0(new_new_n1073_), .A1(new_new_n49_), .B0(new_new_n1077_), .Y(new_new_n1078_));
  AOI210     g1056(.A0(new_new_n1078_), .A1(new_new_n1066_), .B0(new_new_n74_), .Y(new_new_n1079_));
  NO2        g1057(.A(new_new_n596_), .B(new_new_n399_), .Y(new_new_n1080_));
  NO2        g1058(.A(new_new_n1080_), .B(new_new_n796_), .Y(new_new_n1081_));
  INV        g1059(.A(new_new_n77_), .Y(new_new_n1082_));
  AOI210     g1060(.A0(new_new_n1031_), .A1(new_new_n943_), .B0(new_new_n962_), .Y(new_new_n1083_));
  AOI210     g1061(.A0(new_new_n1083_), .A1(new_new_n1082_), .B0(new_new_n716_), .Y(new_new_n1084_));
  NA2        g1062(.A(new_new_n269_), .B(new_new_n58_), .Y(new_new_n1085_));
  AOI220     g1063(.A0(new_new_n1085_), .A1(new_new_n77_), .B0(new_new_n362_), .B1(new_new_n263_), .Y(new_new_n1086_));
  NO2        g1064(.A(new_new_n1086_), .B(new_new_n245_), .Y(new_new_n1087_));
  NA3        g1065(.A(new_new_n99_), .B(new_new_n318_), .C(new_new_n31_), .Y(new_new_n1088_));
  INV        g1066(.A(new_new_n1088_), .Y(new_new_n1089_));
  NO3        g1067(.A(new_new_n1089_), .B(new_new_n1087_), .C(new_new_n1084_), .Y(new_new_n1090_));
  OAI210     g1068(.A0(new_new_n277_), .A1(new_new_n163_), .B0(new_new_n90_), .Y(new_new_n1091_));
  NA3        g1069(.A(new_new_n800_), .B(new_new_n300_), .C(new_new_n81_), .Y(new_new_n1092_));
  AOI210     g1070(.A0(new_new_n1092_), .A1(new_new_n1091_), .B0(i_11_), .Y(new_new_n1093_));
  NA2        g1071(.A(new_new_n639_), .B(new_new_n224_), .Y(new_new_n1094_));
  OAI210     g1072(.A0(new_new_n1094_), .A1(new_new_n955_), .B0(new_new_n214_), .Y(new_new_n1095_));
  NA2        g1073(.A(new_new_n169_), .B(i_5_), .Y(new_new_n1096_));
  AOI210     g1074(.A0(new_new_n1095_), .A1(new_new_n813_), .B0(new_new_n1096_), .Y(new_new_n1097_));
  NO3        g1075(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1098_));
  OAI210     g1076(.A0(new_new_n966_), .A1(new_new_n318_), .B0(new_new_n1098_), .Y(new_new_n1099_));
  NO2        g1077(.A(new_new_n1099_), .B(new_new_n765_), .Y(new_new_n1100_));
  NO4        g1078(.A(new_new_n987_), .B(new_new_n503_), .C(new_new_n262_), .D(new_new_n261_), .Y(new_new_n1101_));
  NO2        g1079(.A(new_new_n1101_), .B(new_new_n593_), .Y(new_new_n1102_));
  NO2        g1080(.A(new_new_n854_), .B(new_new_n381_), .Y(new_new_n1103_));
  AOI210     g1081(.A0(new_new_n1103_), .A1(new_new_n1102_), .B0(new_new_n41_), .Y(new_new_n1104_));
  NO4        g1082(.A(new_new_n1104_), .B(new_new_n1100_), .C(new_new_n1097_), .D(new_new_n1093_), .Y(new_new_n1105_));
  OAI210     g1083(.A0(new_new_n1090_), .A1(i_4_), .B0(new_new_n1105_), .Y(new_new_n1106_));
  NO3        g1084(.A(new_new_n1106_), .B(new_new_n1081_), .C(new_new_n1079_), .Y(new_new_n1107_));
  NA4        g1085(.A(new_new_n1107_), .B(new_new_n1062_), .C(new_new_n993_), .D(new_new_n910_), .Y(men4));
  INV        g1086(.A(new_new_n742_), .Y(new_new_n1111_));
  INV        g1087(.A(i_2_), .Y(new_new_n1112_));
endmodule


