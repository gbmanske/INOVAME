//Benchmark atmr_misex3_1774_0.0313

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1218_, ori_ori_n1219_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1522_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1595_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  AN2        o0001(.A(f), .B(e), .Y(ori_ori_n30_));
  NOi32      o0002(.An(m), .Bn(l), .C(n), .Y(ori_ori_n31_));
  NOi32      o0003(.An(i), .Bn(g), .C(h), .Y(ori_ori_n32_));
  NA2        o0004(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  AN2        o0005(.A(m), .B(l), .Y(ori_ori_n34_));
  NOi32      o0006(.An(j), .Bn(g), .C(k), .Y(ori_ori_n35_));
  NA2        o0007(.A(ori_ori_n35_), .B(ori_ori_n34_), .Y(ori_ori_n36_));
  NO2        o0008(.A(ori_ori_n36_), .B(n), .Y(ori_ori_n37_));
  INV        o0009(.A(h), .Y(ori_ori_n38_));
  NAi21      o0010(.An(j), .B(l), .Y(ori_ori_n39_));
  NAi32      o0011(.An(n), .Bn(g), .C(m), .Y(ori_ori_n40_));
  NO3        o0012(.A(ori_ori_n40_), .B(ori_ori_n39_), .C(ori_ori_n38_), .Y(ori_ori_n41_));
  NAi31      o0013(.An(n), .B(m), .C(l), .Y(ori_ori_n42_));
  INV        o0014(.A(i), .Y(ori_ori_n43_));
  AN2        o0015(.A(h), .B(g), .Y(ori_ori_n44_));
  NA2        o0016(.A(ori_ori_n44_), .B(ori_ori_n43_), .Y(ori_ori_n45_));
  NO2        o0017(.A(ori_ori_n45_), .B(ori_ori_n42_), .Y(ori_ori_n46_));
  NAi21      o0018(.An(n), .B(m), .Y(ori_ori_n47_));
  NOi32      o0019(.An(k), .Bn(h), .C(l), .Y(ori_ori_n48_));
  NOi32      o0020(.An(k), .Bn(h), .C(g), .Y(ori_ori_n49_));
  INV        o0021(.A(ori_ori_n49_), .Y(ori_ori_n50_));
  NO2        o0022(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n51_));
  INV        o0023(.A(c), .Y(ori_ori_n52_));
  NA2        o0024(.A(e), .B(b), .Y(ori_ori_n53_));
  NO2        o0025(.A(ori_ori_n53_), .B(ori_ori_n52_), .Y(ori_ori_n54_));
  INV        o0026(.A(d), .Y(ori_ori_n55_));
  NAi21      o0027(.An(i), .B(h), .Y(ori_ori_n56_));
  NAi41      o0028(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n57_));
  NA2        o0029(.A(g), .B(f), .Y(ori_ori_n58_));
  NAi21      o0030(.An(i), .B(j), .Y(ori_ori_n59_));
  NAi32      o0031(.An(n), .Bn(k), .C(m), .Y(ori_ori_n60_));
  NAi31      o0032(.An(l), .B(m), .C(k), .Y(ori_ori_n61_));
  NAi21      o0033(.An(e), .B(h), .Y(ori_ori_n62_));
  NAi41      o0034(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n63_));
  INV        o0035(.A(m), .Y(ori_ori_n64_));
  NOi21      o0036(.An(k), .B(l), .Y(ori_ori_n65_));
  NA2        o0037(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  AN4        o0038(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n67_));
  NOi31      o0039(.An(h), .B(g), .C(f), .Y(ori_ori_n68_));
  NA2        o0040(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  NAi32      o0041(.An(m), .Bn(k), .C(j), .Y(ori_ori_n70_));
  NOi32      o0042(.An(h), .Bn(g), .C(f), .Y(ori_ori_n71_));
  NA2        o0043(.A(ori_ori_n71_), .B(ori_ori_n67_), .Y(ori_ori_n72_));
  OA220      o0044(.A0(ori_ori_n72_), .A1(ori_ori_n70_), .B0(ori_ori_n69_), .B1(ori_ori_n66_), .Y(ori_ori_n73_));
  INV        o0045(.A(ori_ori_n73_), .Y(ori_ori_n74_));
  INV        o0046(.A(n), .Y(ori_ori_n75_));
  NOi32      o0047(.An(e), .Bn(b), .C(d), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  INV        o0049(.A(j), .Y(ori_ori_n78_));
  AN3        o0050(.A(m), .B(k), .C(i), .Y(ori_ori_n79_));
  NA3        o0051(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .Y(ori_ori_n80_));
  NO2        o0052(.A(ori_ori_n80_), .B(f), .Y(ori_ori_n81_));
  NAi32      o0053(.An(g), .Bn(f), .C(h), .Y(ori_ori_n82_));
  NAi31      o0054(.An(j), .B(m), .C(l), .Y(ori_ori_n83_));
  NO2        o0055(.A(ori_ori_n83_), .B(ori_ori_n82_), .Y(ori_ori_n84_));
  NA2        o0056(.A(m), .B(l), .Y(ori_ori_n85_));
  NAi31      o0057(.An(k), .B(j), .C(g), .Y(ori_ori_n86_));
  NO3        o0058(.A(ori_ori_n86_), .B(ori_ori_n85_), .C(f), .Y(ori_ori_n87_));
  AN2        o0059(.A(j), .B(g), .Y(ori_ori_n88_));
  NOi32      o0060(.An(m), .Bn(l), .C(i), .Y(ori_ori_n89_));
  NOi21      o0061(.An(g), .B(i), .Y(ori_ori_n90_));
  NOi32      o0062(.An(m), .Bn(j), .C(k), .Y(ori_ori_n91_));
  AOI220     o0063(.A0(ori_ori_n91_), .A1(ori_ori_n90_), .B0(ori_ori_n89_), .B1(ori_ori_n88_), .Y(ori_ori_n92_));
  NO2        o0064(.A(ori_ori_n92_), .B(f), .Y(ori_ori_n93_));
  NO3        o0065(.A(ori_ori_n87_), .B(ori_ori_n84_), .C(ori_ori_n81_), .Y(ori_ori_n94_));
  NAi41      o0066(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n95_));
  AN2        o0067(.A(e), .B(b), .Y(ori_ori_n96_));
  NOi31      o0068(.An(c), .B(h), .C(f), .Y(ori_ori_n97_));
  NA2        o0069(.A(ori_ori_n97_), .B(ori_ori_n96_), .Y(ori_ori_n98_));
  NO2        o0070(.A(ori_ori_n98_), .B(ori_ori_n95_), .Y(ori_ori_n99_));
  NOi21      o0071(.An(g), .B(f), .Y(ori_ori_n100_));
  NOi21      o0072(.An(i), .B(h), .Y(ori_ori_n101_));
  INV        o0073(.A(a), .Y(ori_ori_n102_));
  NA2        o0074(.A(ori_ori_n96_), .B(ori_ori_n102_), .Y(ori_ori_n103_));
  INV        o0075(.A(l), .Y(ori_ori_n104_));
  NOi21      o0076(.An(m), .B(n), .Y(ori_ori_n105_));
  AN2        o0077(.A(k), .B(h), .Y(ori_ori_n106_));
  INV        o0078(.A(b), .Y(ori_ori_n107_));
  NA2        o0079(.A(l), .B(j), .Y(ori_ori_n108_));
  AN2        o0080(.A(k), .B(i), .Y(ori_ori_n109_));
  NA2        o0081(.A(ori_ori_n109_), .B(ori_ori_n108_), .Y(ori_ori_n110_));
  NA2        o0082(.A(g), .B(e), .Y(ori_ori_n111_));
  NOi32      o0083(.An(c), .Bn(a), .C(d), .Y(ori_ori_n112_));
  NA2        o0084(.A(ori_ori_n112_), .B(ori_ori_n105_), .Y(ori_ori_n113_));
  INV        o0085(.A(ori_ori_n99_), .Y(ori_ori_n114_));
  OAI210     o0086(.A0(ori_ori_n94_), .A1(ori_ori_n77_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  NOi31      o0087(.An(k), .B(m), .C(j), .Y(ori_ori_n116_));
  NA3        o0088(.A(ori_ori_n116_), .B(ori_ori_n68_), .C(ori_ori_n67_), .Y(ori_ori_n117_));
  NOi31      o0089(.An(k), .B(m), .C(i), .Y(ori_ori_n118_));
  INV        o0090(.A(ori_ori_n117_), .Y(ori_ori_n119_));
  NOi32      o0091(.An(f), .Bn(b), .C(e), .Y(ori_ori_n120_));
  NAi21      o0092(.An(g), .B(h), .Y(ori_ori_n121_));
  NAi21      o0093(.An(m), .B(n), .Y(ori_ori_n122_));
  NAi21      o0094(.An(j), .B(k), .Y(ori_ori_n123_));
  NO3        o0095(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(ori_ori_n121_), .Y(ori_ori_n124_));
  NAi41      o0096(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n125_));
  NAi31      o0097(.An(j), .B(k), .C(h), .Y(ori_ori_n126_));
  NA2        o0098(.A(ori_ori_n124_), .B(ori_ori_n120_), .Y(ori_ori_n127_));
  NO2        o0099(.A(k), .B(j), .Y(ori_ori_n128_));
  NO2        o0100(.A(ori_ori_n128_), .B(ori_ori_n122_), .Y(ori_ori_n129_));
  AN2        o0101(.A(k), .B(j), .Y(ori_ori_n130_));
  NAi21      o0102(.An(c), .B(b), .Y(ori_ori_n131_));
  NA2        o0103(.A(f), .B(d), .Y(ori_ori_n132_));
  NO4        o0104(.A(ori_ori_n132_), .B(ori_ori_n131_), .C(ori_ori_n130_), .D(ori_ori_n121_), .Y(ori_ori_n133_));
  NA2        o0105(.A(h), .B(c), .Y(ori_ori_n134_));
  NAi31      o0106(.An(f), .B(e), .C(b), .Y(ori_ori_n135_));
  NA2        o0107(.A(ori_ori_n133_), .B(ori_ori_n129_), .Y(ori_ori_n136_));
  NA2        o0108(.A(d), .B(b), .Y(ori_ori_n137_));
  NAi21      o0109(.An(e), .B(f), .Y(ori_ori_n138_));
  NO2        o0110(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n139_));
  NA2        o0111(.A(b), .B(a), .Y(ori_ori_n140_));
  NAi21      o0112(.An(e), .B(g), .Y(ori_ori_n141_));
  NAi21      o0113(.An(c), .B(d), .Y(ori_ori_n142_));
  NAi31      o0114(.An(l), .B(k), .C(h), .Y(ori_ori_n143_));
  NO2        o0115(.A(ori_ori_n122_), .B(ori_ori_n143_), .Y(ori_ori_n144_));
  NA2        o0116(.A(ori_ori_n144_), .B(ori_ori_n139_), .Y(ori_ori_n145_));
  NAi41      o0117(.An(ori_ori_n119_), .B(ori_ori_n145_), .C(ori_ori_n136_), .D(ori_ori_n127_), .Y(ori_ori_n146_));
  NAi31      o0118(.An(e), .B(f), .C(b), .Y(ori_ori_n147_));
  NOi21      o0119(.An(g), .B(d), .Y(ori_ori_n148_));
  NO2        o0120(.A(ori_ori_n148_), .B(ori_ori_n147_), .Y(ori_ori_n149_));
  NOi21      o0121(.An(h), .B(i), .Y(ori_ori_n150_));
  NOi21      o0122(.An(k), .B(m), .Y(ori_ori_n151_));
  NA3        o0123(.A(ori_ori_n151_), .B(ori_ori_n150_), .C(n), .Y(ori_ori_n152_));
  NOi21      o0124(.An(ori_ori_n149_), .B(ori_ori_n152_), .Y(ori_ori_n153_));
  NOi21      o0125(.An(h), .B(g), .Y(ori_ori_n154_));
  NAi31      o0126(.An(l), .B(j), .C(h), .Y(ori_ori_n155_));
  NOi32      o0127(.An(n), .Bn(k), .C(m), .Y(ori_ori_n156_));
  INV        o0128(.A(l), .Y(ori_ori_n157_));
  NAi31      o0129(.An(d), .B(f), .C(c), .Y(ori_ori_n158_));
  NAi31      o0130(.An(e), .B(f), .C(c), .Y(ori_ori_n159_));
  NA2        o0131(.A(ori_ori_n159_), .B(ori_ori_n158_), .Y(ori_ori_n160_));
  NA2        o0132(.A(j), .B(h), .Y(ori_ori_n161_));
  OR3        o0133(.A(n), .B(m), .C(k), .Y(ori_ori_n162_));
  NO2        o0134(.A(ori_ori_n162_), .B(ori_ori_n161_), .Y(ori_ori_n163_));
  NAi32      o0135(.An(m), .Bn(k), .C(n), .Y(ori_ori_n164_));
  NO2        o0136(.A(ori_ori_n164_), .B(ori_ori_n161_), .Y(ori_ori_n165_));
  AOI220     o0137(.A0(ori_ori_n165_), .A1(ori_ori_n149_), .B0(ori_ori_n163_), .B1(ori_ori_n160_), .Y(ori_ori_n166_));
  NO2        o0138(.A(n), .B(m), .Y(ori_ori_n167_));
  NA2        o0139(.A(ori_ori_n167_), .B(ori_ori_n48_), .Y(ori_ori_n168_));
  NAi21      o0140(.An(f), .B(e), .Y(ori_ori_n169_));
  NA2        o0141(.A(d), .B(c), .Y(ori_ori_n170_));
  NO2        o0142(.A(ori_ori_n170_), .B(ori_ori_n169_), .Y(ori_ori_n171_));
  NOi21      o0143(.An(ori_ori_n171_), .B(ori_ori_n168_), .Y(ori_ori_n172_));
  NAi31      o0144(.An(m), .B(n), .C(b), .Y(ori_ori_n173_));
  NA2        o0145(.A(k), .B(i), .Y(ori_ori_n174_));
  NAi21      o0146(.An(h), .B(f), .Y(ori_ori_n175_));
  NO2        o0147(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  NO2        o0148(.A(ori_ori_n173_), .B(ori_ori_n142_), .Y(ori_ori_n177_));
  NA2        o0149(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  NOi32      o0150(.An(f), .Bn(c), .C(d), .Y(ori_ori_n179_));
  NOi32      o0151(.An(f), .Bn(c), .C(e), .Y(ori_ori_n180_));
  NO2        o0152(.A(ori_ori_n180_), .B(ori_ori_n179_), .Y(ori_ori_n181_));
  NO3        o0153(.A(n), .B(m), .C(j), .Y(ori_ori_n182_));
  NA2        o0154(.A(ori_ori_n182_), .B(ori_ori_n106_), .Y(ori_ori_n183_));
  AO210      o0155(.A0(ori_ori_n183_), .A1(ori_ori_n168_), .B0(ori_ori_n181_), .Y(ori_ori_n184_));
  NAi41      o0156(.An(ori_ori_n172_), .B(ori_ori_n184_), .C(ori_ori_n178_), .D(ori_ori_n166_), .Y(ori_ori_n185_));
  OR3        o0157(.A(ori_ori_n185_), .B(ori_ori_n153_), .C(ori_ori_n146_), .Y(ori_ori_n186_));
  NO3        o0158(.A(ori_ori_n186_), .B(ori_ori_n115_), .C(ori_ori_n74_), .Y(ori_ori_n187_));
  NA3        o0159(.A(m), .B(ori_ori_n104_), .C(j), .Y(ori_ori_n188_));
  NAi31      o0160(.An(n), .B(h), .C(g), .Y(ori_ori_n189_));
  NO2        o0161(.A(ori_ori_n189_), .B(ori_ori_n188_), .Y(ori_ori_n190_));
  NOi32      o0162(.An(m), .Bn(k), .C(l), .Y(ori_ori_n191_));
  NA3        o0163(.A(ori_ori_n191_), .B(ori_ori_n78_), .C(g), .Y(ori_ori_n192_));
  NO2        o0164(.A(ori_ori_n192_), .B(n), .Y(ori_ori_n193_));
  NOi21      o0165(.An(k), .B(j), .Y(ori_ori_n194_));
  NA4        o0166(.A(ori_ori_n194_), .B(ori_ori_n105_), .C(i), .D(g), .Y(ori_ori_n195_));
  NAi41      o0167(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n196_));
  INV        o0168(.A(ori_ori_n196_), .Y(ori_ori_n197_));
  INV        o0169(.A(f), .Y(ori_ori_n198_));
  INV        o0170(.A(g), .Y(ori_ori_n199_));
  NOi31      o0171(.An(i), .B(j), .C(h), .Y(ori_ori_n200_));
  NOi21      o0172(.An(l), .B(m), .Y(ori_ori_n201_));
  NA2        o0173(.A(ori_ori_n201_), .B(ori_ori_n200_), .Y(ori_ori_n202_));
  NO3        o0174(.A(ori_ori_n202_), .B(ori_ori_n199_), .C(ori_ori_n198_), .Y(ori_ori_n203_));
  NA2        o0175(.A(ori_ori_n203_), .B(ori_ori_n197_), .Y(ori_ori_n204_));
  INV        o0176(.A(ori_ori_n204_), .Y(ori_ori_n205_));
  NOi21      o0177(.An(n), .B(m), .Y(ori_ori_n206_));
  OR2        o0178(.A(ori_ori_n70_), .B(ori_ori_n69_), .Y(ori_ori_n207_));
  NAi21      o0179(.An(j), .B(h), .Y(ori_ori_n208_));
  XN2        o0180(.A(i), .B(h), .Y(ori_ori_n209_));
  NA2        o0181(.A(ori_ori_n209_), .B(ori_ori_n208_), .Y(ori_ori_n210_));
  NOi31      o0182(.An(k), .B(n), .C(m), .Y(ori_ori_n211_));
  NOi31      o0183(.An(ori_ori_n211_), .B(ori_ori_n170_), .C(ori_ori_n169_), .Y(ori_ori_n212_));
  NA2        o0184(.A(ori_ori_n212_), .B(ori_ori_n210_), .Y(ori_ori_n213_));
  NAi31      o0185(.An(f), .B(e), .C(c), .Y(ori_ori_n214_));
  NO4        o0186(.A(ori_ori_n214_), .B(ori_ori_n162_), .C(ori_ori_n161_), .D(ori_ori_n55_), .Y(ori_ori_n215_));
  NA3        o0187(.A(e), .B(c), .C(b), .Y(ori_ori_n216_));
  NAi32      o0188(.An(m), .Bn(i), .C(k), .Y(ori_ori_n217_));
  INV        o0189(.A(k), .Y(ori_ori_n218_));
  INV        o0190(.A(ori_ori_n215_), .Y(ori_ori_n219_));
  NAi21      o0191(.An(n), .B(a), .Y(ori_ori_n220_));
  NO2        o0192(.A(ori_ori_n220_), .B(ori_ori_n137_), .Y(ori_ori_n221_));
  NAi41      o0193(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n222_));
  NO2        o0194(.A(ori_ori_n222_), .B(e), .Y(ori_ori_n223_));
  NA2        o0195(.A(ori_ori_n223_), .B(ori_ori_n221_), .Y(ori_ori_n224_));
  AN4        o0196(.A(ori_ori_n224_), .B(ori_ori_n219_), .C(ori_ori_n213_), .D(ori_ori_n207_), .Y(ori_ori_n225_));
  OR2        o0197(.A(h), .B(g), .Y(ori_ori_n226_));
  NO2        o0198(.A(ori_ori_n226_), .B(ori_ori_n95_), .Y(ori_ori_n227_));
  NA2        o0199(.A(ori_ori_n227_), .B(ori_ori_n120_), .Y(ori_ori_n228_));
  NAi41      o0200(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n229_));
  NO2        o0201(.A(ori_ori_n229_), .B(ori_ori_n198_), .Y(ori_ori_n230_));
  NA2        o0202(.A(ori_ori_n151_), .B(ori_ori_n101_), .Y(ori_ori_n231_));
  NAi21      o0203(.An(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NO2        o0204(.A(n), .B(a), .Y(ori_ori_n233_));
  NAi31      o0205(.An(ori_ori_n222_), .B(ori_ori_n233_), .C(ori_ori_n96_), .Y(ori_ori_n234_));
  AN2        o0206(.A(ori_ori_n234_), .B(ori_ori_n232_), .Y(ori_ori_n235_));
  NAi21      o0207(.An(h), .B(i), .Y(ori_ori_n236_));
  NA2        o0208(.A(ori_ori_n167_), .B(k), .Y(ori_ori_n237_));
  NO2        o0209(.A(ori_ori_n237_), .B(ori_ori_n236_), .Y(ori_ori_n238_));
  NA2        o0210(.A(ori_ori_n238_), .B(ori_ori_n179_), .Y(ori_ori_n239_));
  NA3        o0211(.A(ori_ori_n239_), .B(ori_ori_n235_), .C(ori_ori_n228_), .Y(ori_ori_n240_));
  NOi21      o0212(.An(g), .B(e), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n63_), .B(ori_ori_n64_), .Y(ori_ori_n242_));
  NA2        o0214(.A(ori_ori_n242_), .B(ori_ori_n241_), .Y(ori_ori_n243_));
  NOi32      o0215(.An(l), .Bn(j), .C(i), .Y(ori_ori_n244_));
  AOI210     o0216(.A0(ori_ori_n65_), .A1(ori_ori_n78_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NAi21      o0217(.An(f), .B(g), .Y(ori_ori_n246_));
  NO2        o0218(.A(ori_ori_n246_), .B(ori_ori_n57_), .Y(ori_ori_n247_));
  NO2        o0219(.A(ori_ori_n245_), .B(ori_ori_n243_), .Y(ori_ori_n248_));
  NOi41      o0220(.An(ori_ori_n225_), .B(ori_ori_n248_), .C(ori_ori_n240_), .D(ori_ori_n205_), .Y(ori_ori_n249_));
  NO4        o0221(.A(ori_ori_n190_), .B(ori_ori_n46_), .C(ori_ori_n41_), .D(ori_ori_n37_), .Y(ori_ori_n250_));
  NO2        o0222(.A(ori_ori_n250_), .B(ori_ori_n103_), .Y(ori_ori_n251_));
  NA3        o0223(.A(ori_ori_n55_), .B(c), .C(b), .Y(ori_ori_n252_));
  NAi21      o0224(.An(h), .B(g), .Y(ori_ori_n253_));
  NO2        o0225(.A(ori_ori_n231_), .B(ori_ori_n246_), .Y(ori_ori_n254_));
  NAi31      o0226(.An(g), .B(k), .C(h), .Y(ori_ori_n255_));
  NA4        o0227(.A(ori_ori_n151_), .B(ori_ori_n71_), .C(ori_ori_n67_), .D(ori_ori_n108_), .Y(ori_ori_n256_));
  NA3        o0228(.A(ori_ori_n151_), .B(ori_ori_n150_), .C(ori_ori_n75_), .Y(ori_ori_n257_));
  NO2        o0229(.A(ori_ori_n257_), .B(ori_ori_n181_), .Y(ori_ori_n258_));
  NOi21      o0230(.An(ori_ori_n256_), .B(ori_ori_n258_), .Y(ori_ori_n259_));
  NA3        o0231(.A(e), .B(c), .C(b), .Y(ori_ori_n260_));
  NAi31      o0232(.An(h), .B(l), .C(i), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n261_), .B(ori_ori_n155_), .Y(ori_ori_n262_));
  NOi21      o0234(.An(ori_ori_n262_), .B(ori_ori_n47_), .Y(ori_ori_n263_));
  NA2        o0235(.A(ori_ori_n247_), .B(ori_ori_n263_), .Y(ori_ori_n264_));
  NAi21      o0236(.An(l), .B(k), .Y(ori_ori_n265_));
  NO2        o0237(.A(ori_ori_n265_), .B(ori_ori_n47_), .Y(ori_ori_n266_));
  NOi21      o0238(.An(l), .B(j), .Y(ori_ori_n267_));
  NAi32      o0239(.An(j), .Bn(h), .C(i), .Y(ori_ori_n268_));
  NAi21      o0240(.An(m), .B(l), .Y(ori_ori_n269_));
  NO3        o0241(.A(ori_ori_n269_), .B(ori_ori_n268_), .C(ori_ori_n75_), .Y(ori_ori_n270_));
  NA2        o0242(.A(h), .B(g), .Y(ori_ori_n271_));
  NA2        o0243(.A(ori_ori_n264_), .B(ori_ori_n259_), .Y(ori_ori_n272_));
  NO2        o0244(.A(ori_ori_n135_), .B(d), .Y(ori_ori_n273_));
  NA2        o0245(.A(ori_ori_n273_), .B(ori_ori_n51_), .Y(ori_ori_n274_));
  NO2        o0246(.A(ori_ori_n98_), .B(ori_ori_n95_), .Y(ori_ori_n275_));
  NAi32      o0247(.An(n), .Bn(m), .C(l), .Y(ori_ori_n276_));
  NO2        o0248(.A(ori_ori_n276_), .B(ori_ori_n268_), .Y(ori_ori_n277_));
  NA2        o0249(.A(ori_ori_n277_), .B(ori_ori_n171_), .Y(ori_ori_n278_));
  NAi31      o0250(.An(k), .B(l), .C(j), .Y(ori_ori_n279_));
  OAI210     o0251(.A0(ori_ori_n265_), .A1(j), .B0(ori_ori_n279_), .Y(ori_ori_n280_));
  NOi21      o0252(.An(ori_ori_n280_), .B(ori_ori_n111_), .Y(ori_ori_n281_));
  NA2        o0253(.A(ori_ori_n278_), .B(ori_ori_n274_), .Y(ori_ori_n282_));
  NO3        o0254(.A(ori_ori_n282_), .B(ori_ori_n272_), .C(ori_ori_n251_), .Y(ori_ori_n283_));
  NA2        o0255(.A(ori_ori_n238_), .B(ori_ori_n180_), .Y(ori_ori_n284_));
  NAi21      o0256(.An(m), .B(k), .Y(ori_ori_n285_));
  NO2        o0257(.A(ori_ori_n209_), .B(ori_ori_n285_), .Y(ori_ori_n286_));
  NAi41      o0258(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n287_));
  NO2        o0259(.A(ori_ori_n287_), .B(ori_ori_n141_), .Y(ori_ori_n288_));
  NA2        o0260(.A(ori_ori_n288_), .B(ori_ori_n286_), .Y(ori_ori_n289_));
  NA2        o0261(.A(e), .B(c), .Y(ori_ori_n290_));
  NO3        o0262(.A(ori_ori_n290_), .B(n), .C(d), .Y(ori_ori_n291_));
  NOi21      o0263(.An(f), .B(h), .Y(ori_ori_n292_));
  NA2        o0264(.A(ori_ori_n292_), .B(ori_ori_n109_), .Y(ori_ori_n293_));
  NO2        o0265(.A(ori_ori_n293_), .B(ori_ori_n199_), .Y(ori_ori_n294_));
  NAi31      o0266(.An(d), .B(e), .C(b), .Y(ori_ori_n295_));
  NO2        o0267(.A(ori_ori_n122_), .B(ori_ori_n295_), .Y(ori_ori_n296_));
  NA2        o0268(.A(ori_ori_n296_), .B(ori_ori_n294_), .Y(ori_ori_n297_));
  NA3        o0269(.A(ori_ori_n297_), .B(ori_ori_n289_), .C(ori_ori_n284_), .Y(ori_ori_n298_));
  NO4        o0270(.A(ori_ori_n287_), .B(ori_ori_n70_), .C(ori_ori_n62_), .D(ori_ori_n199_), .Y(ori_ori_n299_));
  NA2        o0271(.A(ori_ori_n233_), .B(ori_ori_n96_), .Y(ori_ori_n300_));
  OR2        o0272(.A(ori_ori_n300_), .B(ori_ori_n192_), .Y(ori_ori_n301_));
  NOi31      o0273(.An(l), .B(n), .C(m), .Y(ori_ori_n302_));
  NA2        o0274(.A(ori_ori_n302_), .B(ori_ori_n200_), .Y(ori_ori_n303_));
  NO2        o0275(.A(ori_ori_n303_), .B(ori_ori_n181_), .Y(ori_ori_n304_));
  NAi32      o0276(.An(ori_ori_n304_), .Bn(ori_ori_n299_), .C(ori_ori_n301_), .Y(ori_ori_n305_));
  NAi32      o0277(.An(m), .Bn(j), .C(k), .Y(ori_ori_n306_));
  NAi41      o0278(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n307_));
  OAI210     o0279(.A0(ori_ori_n196_), .A1(ori_ori_n306_), .B0(ori_ori_n307_), .Y(ori_ori_n308_));
  NOi31      o0280(.An(j), .B(m), .C(k), .Y(ori_ori_n309_));
  NO2        o0281(.A(ori_ori_n116_), .B(ori_ori_n309_), .Y(ori_ori_n310_));
  AN3        o0282(.A(h), .B(g), .C(f), .Y(ori_ori_n311_));
  NAi31      o0283(.An(ori_ori_n310_), .B(ori_ori_n311_), .C(ori_ori_n308_), .Y(ori_ori_n312_));
  NOi32      o0284(.An(m), .Bn(j), .C(l), .Y(ori_ori_n313_));
  NO2        o0285(.A(ori_ori_n313_), .B(ori_ori_n89_), .Y(ori_ori_n314_));
  NAi32      o0286(.An(ori_ori_n314_), .Bn(ori_ori_n189_), .C(ori_ori_n273_), .Y(ori_ori_n315_));
  NO2        o0287(.A(ori_ori_n269_), .B(ori_ori_n268_), .Y(ori_ori_n316_));
  NO2        o0288(.A(ori_ori_n202_), .B(g), .Y(ori_ori_n317_));
  NO2        o0289(.A(ori_ori_n147_), .B(ori_ori_n75_), .Y(ori_ori_n318_));
  AOI220     o0290(.A0(ori_ori_n318_), .A1(ori_ori_n317_), .B0(ori_ori_n230_), .B1(ori_ori_n316_), .Y(ori_ori_n319_));
  NA2        o0291(.A(ori_ori_n217_), .B(ori_ori_n70_), .Y(ori_ori_n320_));
  NA3        o0292(.A(ori_ori_n320_), .B(ori_ori_n311_), .C(ori_ori_n197_), .Y(ori_ori_n321_));
  NA4        o0293(.A(ori_ori_n321_), .B(ori_ori_n319_), .C(ori_ori_n315_), .D(ori_ori_n312_), .Y(ori_ori_n322_));
  NA3        o0294(.A(h), .B(g), .C(f), .Y(ori_ori_n323_));
  NO2        o0295(.A(ori_ori_n323_), .B(ori_ori_n66_), .Y(ori_ori_n324_));
  NA2        o0296(.A(ori_ori_n307_), .B(ori_ori_n196_), .Y(ori_ori_n325_));
  NA2        o0297(.A(ori_ori_n154_), .B(e), .Y(ori_ori_n326_));
  NO2        o0298(.A(ori_ori_n326_), .B(ori_ori_n39_), .Y(ori_ori_n327_));
  NA2        o0299(.A(ori_ori_n325_), .B(ori_ori_n324_), .Y(ori_ori_n328_));
  NOi32      o0300(.An(j), .Bn(g), .C(i), .Y(ori_ori_n329_));
  NA3        o0301(.A(ori_ori_n329_), .B(ori_ori_n265_), .C(ori_ori_n105_), .Y(ori_ori_n330_));
  OR2        o0302(.A(ori_ori_n103_), .B(ori_ori_n330_), .Y(ori_ori_n331_));
  NOi32      o0303(.An(e), .Bn(b), .C(a), .Y(ori_ori_n332_));
  AN2        o0304(.A(l), .B(j), .Y(ori_ori_n333_));
  NO2        o0305(.A(ori_ori_n285_), .B(ori_ori_n333_), .Y(ori_ori_n334_));
  NO3        o0306(.A(ori_ori_n287_), .B(ori_ori_n62_), .C(ori_ori_n199_), .Y(ori_ori_n335_));
  NA2        o0307(.A(ori_ori_n195_), .B(ori_ori_n33_), .Y(ori_ori_n336_));
  AOI220     o0308(.A0(ori_ori_n336_), .A1(ori_ori_n332_), .B0(ori_ori_n335_), .B1(ori_ori_n334_), .Y(ori_ori_n337_));
  NA4        o0309(.A(ori_ori_n191_), .B(ori_ori_n78_), .C(g), .D(ori_ori_n198_), .Y(ori_ori_n338_));
  NA2        o0310(.A(ori_ori_n49_), .B(ori_ori_n105_), .Y(ori_ori_n339_));
  NA3        o0311(.A(ori_ori_n337_), .B(ori_ori_n331_), .C(ori_ori_n328_), .Y(ori_ori_n340_));
  NO4        o0312(.A(ori_ori_n340_), .B(ori_ori_n322_), .C(ori_ori_n305_), .D(ori_ori_n298_), .Y(ori_ori_n341_));
  NA4        o0313(.A(ori_ori_n341_), .B(ori_ori_n283_), .C(ori_ori_n249_), .D(ori_ori_n187_), .Y(ori10));
  NA3        o0314(.A(m), .B(k), .C(i), .Y(ori_ori_n343_));
  NOi21      o0315(.An(e), .B(f), .Y(ori_ori_n344_));
  NO4        o0316(.A(ori_ori_n142_), .B(ori_ori_n344_), .C(n), .D(ori_ori_n102_), .Y(ori_ori_n345_));
  NAi31      o0317(.An(b), .B(f), .C(c), .Y(ori_ori_n346_));
  INV        o0318(.A(ori_ori_n346_), .Y(ori_ori_n347_));
  NOi32      o0319(.An(k), .Bn(h), .C(j), .Y(ori_ori_n348_));
  NA2        o0320(.A(ori_ori_n348_), .B(ori_ori_n206_), .Y(ori_ori_n349_));
  NA2        o0321(.A(ori_ori_n152_), .B(ori_ori_n349_), .Y(ori_ori_n350_));
  NA2        o0322(.A(ori_ori_n350_), .B(ori_ori_n347_), .Y(ori_ori_n351_));
  AN2        o0323(.A(j), .B(h), .Y(ori_ori_n352_));
  NO3        o0324(.A(n), .B(m), .C(k), .Y(ori_ori_n353_));
  NA2        o0325(.A(ori_ori_n353_), .B(ori_ori_n352_), .Y(ori_ori_n354_));
  NO3        o0326(.A(ori_ori_n354_), .B(ori_ori_n142_), .C(ori_ori_n198_), .Y(ori_ori_n355_));
  OR2        o0327(.A(m), .B(k), .Y(ori_ori_n356_));
  NO2        o0328(.A(ori_ori_n161_), .B(ori_ori_n356_), .Y(ori_ori_n357_));
  NA4        o0329(.A(n), .B(f), .C(c), .D(ori_ori_n107_), .Y(ori_ori_n358_));
  NOi21      o0330(.An(ori_ori_n357_), .B(ori_ori_n358_), .Y(ori_ori_n359_));
  NOi32      o0331(.An(d), .Bn(a), .C(c), .Y(ori_ori_n360_));
  NA2        o0332(.A(ori_ori_n360_), .B(ori_ori_n169_), .Y(ori_ori_n361_));
  NO2        o0333(.A(ori_ori_n359_), .B(ori_ori_n355_), .Y(ori_ori_n362_));
  NO2        o0334(.A(ori_ori_n358_), .B(ori_ori_n269_), .Y(ori_ori_n363_));
  NOi32      o0335(.An(f), .Bn(d), .C(c), .Y(ori_ori_n364_));
  AOI220     o0336(.A0(ori_ori_n364_), .A1(ori_ori_n277_), .B0(ori_ori_n363_), .B1(ori_ori_n200_), .Y(ori_ori_n365_));
  NA3        o0337(.A(ori_ori_n365_), .B(ori_ori_n362_), .C(ori_ori_n351_), .Y(ori_ori_n366_));
  NO2        o0338(.A(ori_ori_n55_), .B(ori_ori_n107_), .Y(ori_ori_n367_));
  NA2        o0339(.A(ori_ori_n233_), .B(ori_ori_n367_), .Y(ori_ori_n368_));
  INV        o0340(.A(e), .Y(ori_ori_n369_));
  NA2        o0341(.A(ori_ori_n44_), .B(e), .Y(ori_ori_n370_));
  OAI220     o0342(.A0(ori_ori_n370_), .A1(ori_ori_n188_), .B0(ori_ori_n192_), .B1(ori_ori_n369_), .Y(ori_ori_n371_));
  NO2        o0343(.A(ori_ori_n80_), .B(ori_ori_n369_), .Y(ori_ori_n372_));
  NO2        o0344(.A(ori_ori_n92_), .B(ori_ori_n369_), .Y(ori_ori_n373_));
  NO3        o0345(.A(ori_ori_n373_), .B(ori_ori_n372_), .C(ori_ori_n371_), .Y(ori_ori_n374_));
  NOi32      o0346(.An(h), .Bn(e), .C(g), .Y(ori_ori_n375_));
  NA3        o0347(.A(ori_ori_n375_), .B(ori_ori_n267_), .C(m), .Y(ori_ori_n376_));
  NOi21      o0348(.An(g), .B(h), .Y(ori_ori_n377_));
  AN3        o0349(.A(m), .B(l), .C(i), .Y(ori_ori_n378_));
  NA3        o0350(.A(ori_ori_n378_), .B(ori_ori_n377_), .C(e), .Y(ori_ori_n379_));
  AN3        o0351(.A(h), .B(g), .C(e), .Y(ori_ori_n380_));
  NA2        o0352(.A(ori_ori_n380_), .B(ori_ori_n89_), .Y(ori_ori_n381_));
  AN3        o0353(.A(ori_ori_n381_), .B(ori_ori_n379_), .C(ori_ori_n376_), .Y(ori_ori_n382_));
  AOI210     o0354(.A0(ori_ori_n382_), .A1(ori_ori_n374_), .B0(ori_ori_n368_), .Y(ori_ori_n383_));
  NA3        o0355(.A(ori_ori_n360_), .B(ori_ori_n169_), .C(ori_ori_n75_), .Y(ori_ori_n384_));
  NAi31      o0356(.An(b), .B(c), .C(a), .Y(ori_ori_n385_));
  NO2        o0357(.A(ori_ori_n385_), .B(n), .Y(ori_ori_n386_));
  NA2        o0358(.A(ori_ori_n49_), .B(m), .Y(ori_ori_n387_));
  NO2        o0359(.A(ori_ori_n387_), .B(ori_ori_n138_), .Y(ori_ori_n388_));
  NA2        o0360(.A(ori_ori_n388_), .B(ori_ori_n386_), .Y(ori_ori_n389_));
  INV        o0361(.A(ori_ori_n389_), .Y(ori_ori_n390_));
  NO3        o0362(.A(ori_ori_n390_), .B(ori_ori_n383_), .C(ori_ori_n366_), .Y(ori_ori_n391_));
  NA2        o0363(.A(i), .B(g), .Y(ori_ori_n392_));
  NOi21      o0364(.An(a), .B(n), .Y(ori_ori_n393_));
  NOi21      o0365(.An(d), .B(c), .Y(ori_ori_n394_));
  NA2        o0366(.A(ori_ori_n394_), .B(ori_ori_n393_), .Y(ori_ori_n395_));
  NA3        o0367(.A(i), .B(g), .C(f), .Y(ori_ori_n396_));
  OR2        o0368(.A(ori_ori_n396_), .B(ori_ori_n61_), .Y(ori_ori_n397_));
  NO2        o0369(.A(ori_ori_n397_), .B(ori_ori_n395_), .Y(ori_ori_n398_));
  INV        o0370(.A(ori_ori_n398_), .Y(ori_ori_n399_));
  OR2        o0371(.A(n), .B(m), .Y(ori_ori_n400_));
  NO2        o0372(.A(ori_ori_n400_), .B(ori_ori_n143_), .Y(ori_ori_n401_));
  NO2        o0373(.A(ori_ori_n170_), .B(ori_ori_n138_), .Y(ori_ori_n402_));
  OAI210     o0374(.A0(ori_ori_n401_), .A1(ori_ori_n163_), .B0(ori_ori_n402_), .Y(ori_ori_n403_));
  INV        o0375(.A(ori_ori_n339_), .Y(ori_ori_n404_));
  NA3        o0376(.A(ori_ori_n404_), .B(ori_ori_n332_), .C(d), .Y(ori_ori_n405_));
  NO2        o0377(.A(ori_ori_n385_), .B(ori_ori_n47_), .Y(ori_ori_n406_));
  NO3        o0378(.A(ori_ori_n58_), .B(ori_ori_n104_), .C(e), .Y(ori_ori_n407_));
  NAi21      o0379(.An(k), .B(j), .Y(ori_ori_n408_));
  NA2        o0380(.A(ori_ori_n236_), .B(ori_ori_n408_), .Y(ori_ori_n409_));
  NA3        o0381(.A(ori_ori_n409_), .B(ori_ori_n407_), .C(ori_ori_n406_), .Y(ori_ori_n410_));
  NAi21      o0382(.An(e), .B(d), .Y(ori_ori_n411_));
  INV        o0383(.A(ori_ori_n411_), .Y(ori_ori_n412_));
  NO2        o0384(.A(ori_ori_n237_), .B(ori_ori_n198_), .Y(ori_ori_n413_));
  NA3        o0385(.A(ori_ori_n413_), .B(ori_ori_n412_), .C(ori_ori_n210_), .Y(ori_ori_n414_));
  NA4        o0386(.A(ori_ori_n414_), .B(ori_ori_n410_), .C(ori_ori_n405_), .D(ori_ori_n403_), .Y(ori_ori_n415_));
  NO2        o0387(.A(ori_ori_n303_), .B(ori_ori_n198_), .Y(ori_ori_n416_));
  NA2        o0388(.A(ori_ori_n416_), .B(ori_ori_n412_), .Y(ori_ori_n417_));
  NOi31      o0389(.An(n), .B(m), .C(k), .Y(ori_ori_n418_));
  AOI220     o0390(.A0(ori_ori_n418_), .A1(ori_ori_n352_), .B0(ori_ori_n206_), .B1(ori_ori_n48_), .Y(ori_ori_n419_));
  NAi31      o0391(.An(g), .B(f), .C(c), .Y(ori_ori_n420_));
  OR3        o0392(.A(ori_ori_n420_), .B(ori_ori_n419_), .C(e), .Y(ori_ori_n421_));
  NA3        o0393(.A(ori_ori_n421_), .B(ori_ori_n417_), .C(ori_ori_n278_), .Y(ori_ori_n422_));
  NO3        o0394(.A(ori_ori_n422_), .B(ori_ori_n415_), .C(ori_ori_n248_), .Y(ori_ori_n423_));
  NOi32      o0395(.An(c), .Bn(a), .C(b), .Y(ori_ori_n424_));
  NA2        o0396(.A(ori_ori_n424_), .B(ori_ori_n105_), .Y(ori_ori_n425_));
  INV        o0397(.A(ori_ori_n255_), .Y(ori_ori_n426_));
  AN2        o0398(.A(e), .B(d), .Y(ori_ori_n427_));
  NA2        o0399(.A(ori_ori_n427_), .B(ori_ori_n426_), .Y(ori_ori_n428_));
  INV        o0400(.A(ori_ori_n138_), .Y(ori_ori_n429_));
  NO2        o0401(.A(ori_ori_n121_), .B(ori_ori_n39_), .Y(ori_ori_n430_));
  NO2        o0402(.A(ori_ori_n58_), .B(e), .Y(ori_ori_n431_));
  NA3        o0403(.A(ori_ori_n155_), .B(ori_ori_n245_), .C(ori_ori_n110_), .Y(ori_ori_n432_));
  AOI220     o0404(.A0(ori_ori_n432_), .A1(ori_ori_n431_), .B0(ori_ori_n430_), .B1(ori_ori_n429_), .Y(ori_ori_n433_));
  AOI210     o0405(.A0(ori_ori_n433_), .A1(ori_ori_n428_), .B0(ori_ori_n425_), .Y(ori_ori_n434_));
  INV        o0406(.A(ori_ori_n193_), .Y(ori_ori_n435_));
  NOi21      o0407(.An(a), .B(b), .Y(ori_ori_n436_));
  NA3        o0408(.A(e), .B(d), .C(c), .Y(ori_ori_n437_));
  NAi21      o0409(.An(ori_ori_n437_), .B(ori_ori_n436_), .Y(ori_ori_n438_));
  NO2        o0410(.A(ori_ori_n384_), .B(ori_ori_n192_), .Y(ori_ori_n439_));
  NOi21      o0411(.An(ori_ori_n438_), .B(ori_ori_n439_), .Y(ori_ori_n440_));
  AOI210     o0412(.A0(ori_ori_n250_), .A1(ori_ori_n435_), .B0(ori_ori_n440_), .Y(ori_ori_n441_));
  NO4        o0413(.A(ori_ori_n175_), .B(ori_ori_n95_), .C(ori_ori_n52_), .D(b), .Y(ori_ori_n442_));
  NA2        o0414(.A(ori_ori_n347_), .B(ori_ori_n144_), .Y(ori_ori_n443_));
  OR2        o0415(.A(k), .B(j), .Y(ori_ori_n444_));
  NA2        o0416(.A(l), .B(k), .Y(ori_ori_n445_));
  NA3        o0417(.A(ori_ori_n445_), .B(ori_ori_n444_), .C(ori_ori_n206_), .Y(ori_ori_n446_));
  AOI210     o0418(.A0(ori_ori_n217_), .A1(ori_ori_n306_), .B0(ori_ori_n75_), .Y(ori_ori_n447_));
  NOi21      o0419(.An(ori_ori_n446_), .B(ori_ori_n447_), .Y(ori_ori_n448_));
  OR3        o0420(.A(ori_ori_n448_), .B(ori_ori_n134_), .C(ori_ori_n125_), .Y(ori_ori_n449_));
  NA2        o0421(.A(ori_ori_n256_), .B(ori_ori_n117_), .Y(ori_ori_n450_));
  INV        o0422(.A(ori_ori_n450_), .Y(ori_ori_n451_));
  NA3        o0423(.A(ori_ori_n451_), .B(ori_ori_n449_), .C(ori_ori_n443_), .Y(ori_ori_n452_));
  NO4        o0424(.A(ori_ori_n452_), .B(ori_ori_n442_), .C(ori_ori_n441_), .D(ori_ori_n434_), .Y(ori_ori_n453_));
  INV        o0425(.A(e), .Y(ori_ori_n454_));
  NO2        o0426(.A(ori_ori_n175_), .B(ori_ori_n52_), .Y(ori_ori_n455_));
  NAi31      o0427(.An(j), .B(l), .C(i), .Y(ori_ori_n456_));
  OAI210     o0428(.A0(ori_ori_n456_), .A1(ori_ori_n122_), .B0(ori_ori_n95_), .Y(ori_ori_n457_));
  NA3        o0429(.A(ori_ori_n457_), .B(ori_ori_n455_), .C(ori_ori_n454_), .Y(ori_ori_n458_));
  NO3        o0430(.A(ori_ori_n361_), .B(ori_ori_n314_), .C(ori_ori_n189_), .Y(ori_ori_n459_));
  NO2        o0431(.A(ori_ori_n361_), .B(ori_ori_n339_), .Y(ori_ori_n460_));
  NO4        o0432(.A(ori_ori_n460_), .B(ori_ori_n459_), .C(ori_ori_n172_), .D(ori_ori_n275_), .Y(ori_ori_n461_));
  NA3        o0433(.A(ori_ori_n461_), .B(ori_ori_n458_), .C(ori_ori_n225_), .Y(ori_ori_n462_));
  OAI210     o0434(.A0(ori_ori_n118_), .A1(ori_ori_n116_), .B0(n), .Y(ori_ori_n463_));
  NO2        o0435(.A(ori_ori_n463_), .B(ori_ori_n121_), .Y(ori_ori_n464_));
  AN2        o0436(.A(ori_ori_n464_), .B(ori_ori_n180_), .Y(ori_ori_n465_));
  XO2        o0437(.A(i), .B(h), .Y(ori_ori_n466_));
  NA3        o0438(.A(ori_ori_n466_), .B(ori_ori_n151_), .C(n), .Y(ori_ori_n467_));
  NAi41      o0439(.An(ori_ori_n270_), .B(ori_ori_n467_), .C(ori_ori_n419_), .D(ori_ori_n349_), .Y(ori_ori_n468_));
  NOi32      o0440(.An(ori_ori_n468_), .Bn(ori_ori_n431_), .C(ori_ori_n252_), .Y(ori_ori_n469_));
  NAi31      o0441(.An(c), .B(f), .C(d), .Y(ori_ori_n470_));
  AOI210     o0442(.A0(ori_ori_n257_), .A1(ori_ori_n183_), .B0(ori_ori_n470_), .Y(ori_ori_n471_));
  NOi21      o0443(.An(ori_ori_n73_), .B(ori_ori_n471_), .Y(ori_ori_n472_));
  NA2        o0444(.A(ori_ori_n211_), .B(ori_ori_n101_), .Y(ori_ori_n473_));
  AOI210     o0445(.A0(ori_ori_n473_), .A1(ori_ori_n168_), .B0(ori_ori_n470_), .Y(ori_ori_n474_));
  INV        o0446(.A(ori_ori_n474_), .Y(ori_ori_n475_));
  AN2        o0447(.A(ori_ori_n263_), .B(ori_ori_n247_), .Y(ori_ori_n476_));
  NA3        o0448(.A(ori_ori_n35_), .B(ori_ori_n34_), .C(f), .Y(ori_ori_n477_));
  NAi31      o0449(.An(ori_ori_n476_), .B(ori_ori_n475_), .C(ori_ori_n472_), .Y(ori_ori_n478_));
  NO4        o0450(.A(ori_ori_n478_), .B(ori_ori_n469_), .C(ori_ori_n465_), .D(ori_ori_n462_), .Y(ori_ori_n479_));
  NA4        o0451(.A(ori_ori_n479_), .B(ori_ori_n453_), .C(ori_ori_n423_), .D(ori_ori_n391_), .Y(ori11));
  NO2        o0452(.A(ori_ori_n63_), .B(f), .Y(ori_ori_n481_));
  NA2        o0453(.A(j), .B(g), .Y(ori_ori_n482_));
  NAi31      o0454(.An(i), .B(m), .C(l), .Y(ori_ori_n483_));
  NA3        o0455(.A(m), .B(k), .C(j), .Y(ori_ori_n484_));
  OAI220     o0456(.A0(ori_ori_n484_), .A1(ori_ori_n121_), .B0(ori_ori_n483_), .B1(ori_ori_n482_), .Y(ori_ori_n485_));
  NA2        o0457(.A(ori_ori_n485_), .B(ori_ori_n481_), .Y(ori_ori_n486_));
  NOi32      o0458(.An(e), .Bn(b), .C(f), .Y(ori_ori_n487_));
  NA2        o0459(.A(ori_ori_n44_), .B(j), .Y(ori_ori_n488_));
  NAi31      o0460(.An(d), .B(e), .C(a), .Y(ori_ori_n489_));
  NO2        o0461(.A(ori_ori_n489_), .B(n), .Y(ori_ori_n490_));
  NA2        o0462(.A(ori_ori_n490_), .B(ori_ori_n93_), .Y(ori_ori_n491_));
  NA2        o0463(.A(j), .B(i), .Y(ori_ori_n492_));
  NAi31      o0464(.An(n), .B(m), .C(k), .Y(ori_ori_n493_));
  NO3        o0465(.A(ori_ori_n493_), .B(ori_ori_n492_), .C(ori_ori_n104_), .Y(ori_ori_n494_));
  NO4        o0466(.A(n), .B(d), .C(ori_ori_n107_), .D(a), .Y(ori_ori_n495_));
  OR2        o0467(.A(n), .B(c), .Y(ori_ori_n496_));
  NO2        o0468(.A(ori_ori_n496_), .B(ori_ori_n140_), .Y(ori_ori_n497_));
  NO2        o0469(.A(ori_ori_n497_), .B(ori_ori_n495_), .Y(ori_ori_n498_));
  NA2        o0470(.A(ori_ori_n485_), .B(f), .Y(ori_ori_n499_));
  NO2        o0471(.A(ori_ori_n255_), .B(ori_ori_n47_), .Y(ori_ori_n500_));
  NO2        o0472(.A(ori_ori_n499_), .B(ori_ori_n498_), .Y(ori_ori_n501_));
  INV        o0473(.A(ori_ori_n501_), .Y(ori_ori_n502_));
  NA2        o0474(.A(ori_ori_n130_), .B(ori_ori_n32_), .Y(ori_ori_n503_));
  OAI220     o0475(.A0(ori_ori_n503_), .A1(m), .B0(ori_ori_n488_), .B1(ori_ori_n217_), .Y(ori_ori_n504_));
  NOi41      o0476(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n505_));
  NAi32      o0477(.An(e), .Bn(b), .C(c), .Y(ori_ori_n506_));
  OR2        o0478(.A(ori_ori_n506_), .B(ori_ori_n75_), .Y(ori_ori_n507_));
  AN2        o0479(.A(ori_ori_n307_), .B(ori_ori_n287_), .Y(ori_ori_n508_));
  NA2        o0480(.A(ori_ori_n508_), .B(ori_ori_n507_), .Y(ori_ori_n509_));
  OA210      o0481(.A0(ori_ori_n509_), .A1(ori_ori_n505_), .B0(ori_ori_n504_), .Y(ori_ori_n510_));
  NO2        o0482(.A(ori_ori_n483_), .B(ori_ori_n482_), .Y(ori_ori_n511_));
  INV        o0483(.A(ori_ori_n386_), .Y(ori_ori_n512_));
  NA2        o0484(.A(ori_ori_n511_), .B(f), .Y(ori_ori_n513_));
  NAi32      o0485(.An(d), .Bn(a), .C(b), .Y(ori_ori_n514_));
  NO2        o0486(.A(ori_ori_n514_), .B(ori_ori_n47_), .Y(ori_ori_n515_));
  NA2        o0487(.A(h), .B(f), .Y(ori_ori_n516_));
  NO2        o0488(.A(ori_ori_n516_), .B(ori_ori_n86_), .Y(ori_ori_n517_));
  NO3        o0489(.A(ori_ori_n164_), .B(ori_ori_n161_), .C(g), .Y(ori_ori_n518_));
  AOI220     o0490(.A0(ori_ori_n518_), .A1(ori_ori_n54_), .B0(ori_ori_n517_), .B1(ori_ori_n515_), .Y(ori_ori_n519_));
  OAI210     o0491(.A0(ori_ori_n513_), .A1(ori_ori_n512_), .B0(ori_ori_n519_), .Y(ori_ori_n520_));
  AN3        o0492(.A(j), .B(h), .C(g), .Y(ori_ori_n521_));
  NO2        o0493(.A(ori_ori_n137_), .B(c), .Y(ori_ori_n522_));
  NA3        o0494(.A(ori_ori_n522_), .B(ori_ori_n521_), .C(ori_ori_n418_), .Y(ori_ori_n523_));
  NA3        o0495(.A(f), .B(d), .C(b), .Y(ori_ori_n524_));
  NO4        o0496(.A(ori_ori_n524_), .B(ori_ori_n164_), .C(ori_ori_n161_), .D(g), .Y(ori_ori_n525_));
  NAi21      o0497(.An(ori_ori_n525_), .B(ori_ori_n523_), .Y(ori_ori_n526_));
  NO3        o0498(.A(ori_ori_n526_), .B(ori_ori_n520_), .C(ori_ori_n510_), .Y(ori_ori_n527_));
  AN4        o0499(.A(ori_ori_n527_), .B(ori_ori_n502_), .C(ori_ori_n491_), .D(ori_ori_n486_), .Y(ori_ori_n528_));
  INV        o0500(.A(k), .Y(ori_ori_n529_));
  NA3        o0501(.A(l), .B(ori_ori_n529_), .C(i), .Y(ori_ori_n530_));
  INV        o0502(.A(ori_ori_n530_), .Y(ori_ori_n531_));
  NAi32      o0503(.An(h), .Bn(f), .C(g), .Y(ori_ori_n532_));
  NAi41      o0504(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n533_));
  OAI210     o0505(.A0(ori_ori_n489_), .A1(n), .B0(ori_ori_n533_), .Y(ori_ori_n534_));
  NA2        o0506(.A(ori_ori_n534_), .B(m), .Y(ori_ori_n535_));
  NAi31      o0507(.An(h), .B(g), .C(f), .Y(ori_ori_n536_));
  OR2        o0508(.A(ori_ori_n535_), .B(ori_ori_n532_), .Y(ori_ori_n537_));
  NO3        o0509(.A(ori_ori_n532_), .B(ori_ori_n63_), .C(ori_ori_n64_), .Y(ori_ori_n538_));
  NAi21      o0510(.An(ori_ori_n538_), .B(ori_ori_n537_), .Y(ori_ori_n539_));
  NAi31      o0511(.An(f), .B(h), .C(g), .Y(ori_ori_n540_));
  NOi32      o0512(.An(b), .Bn(a), .C(c), .Y(ori_ori_n541_));
  NOi32      o0513(.An(d), .Bn(a), .C(e), .Y(ori_ori_n542_));
  NO2        o0514(.A(n), .B(c), .Y(ori_ori_n543_));
  NOi32      o0515(.An(e), .Bn(a), .C(d), .Y(ori_ori_n544_));
  AOI210     o0516(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n544_), .Y(ori_ori_n545_));
  NO2        o0517(.A(ori_ori_n232_), .B(ori_ori_n78_), .Y(ori_ori_n546_));
  AOI210     o0518(.A0(ori_ori_n539_), .A1(ori_ori_n531_), .B0(ori_ori_n546_), .Y(ori_ori_n547_));
  NO3        o0519(.A(ori_ori_n285_), .B(ori_ori_n56_), .C(n), .Y(ori_ori_n548_));
  NA3        o0520(.A(ori_ori_n470_), .B(ori_ori_n159_), .C(ori_ori_n158_), .Y(ori_ori_n549_));
  NA2        o0521(.A(ori_ori_n420_), .B(ori_ori_n214_), .Y(ori_ori_n550_));
  OR2        o0522(.A(ori_ori_n550_), .B(ori_ori_n549_), .Y(ori_ori_n551_));
  NA2        o0523(.A(ori_ori_n551_), .B(ori_ori_n548_), .Y(ori_ori_n552_));
  NO2        o0524(.A(ori_ori_n552_), .B(ori_ori_n78_), .Y(ori_ori_n553_));
  NA3        o0525(.A(ori_ori_n505_), .B(ori_ori_n309_), .C(ori_ori_n44_), .Y(ori_ori_n554_));
  NOi32      o0526(.An(e), .Bn(c), .C(f), .Y(ori_ori_n555_));
  NOi21      o0527(.An(f), .B(g), .Y(ori_ori_n556_));
  NO2        o0528(.A(ori_ori_n556_), .B(ori_ori_n196_), .Y(ori_ori_n557_));
  AOI220     o0529(.A0(ori_ori_n557_), .A1(ori_ori_n357_), .B0(ori_ori_n555_), .B1(ori_ori_n163_), .Y(ori_ori_n558_));
  NA3        o0530(.A(ori_ori_n558_), .B(ori_ori_n554_), .C(ori_ori_n166_), .Y(ori_ori_n559_));
  NOi21      o0531(.An(j), .B(l), .Y(ori_ori_n560_));
  NAi21      o0532(.An(k), .B(h), .Y(ori_ori_n561_));
  NO2        o0533(.A(ori_ori_n561_), .B(ori_ori_n246_), .Y(ori_ori_n562_));
  NA2        o0534(.A(ori_ori_n562_), .B(ori_ori_n560_), .Y(ori_ori_n563_));
  OR2        o0535(.A(ori_ori_n563_), .B(ori_ori_n535_), .Y(ori_ori_n564_));
  NO2        o0536(.A(ori_ori_n279_), .B(ori_ori_n540_), .Y(ori_ori_n565_));
  NO2        o0537(.A(ori_ori_n489_), .B(ori_ori_n47_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n565_), .Y(ori_ori_n567_));
  NA2        o0539(.A(ori_ori_n567_), .B(ori_ori_n564_), .Y(ori_ori_n568_));
  NA2        o0540(.A(ori_ori_n101_), .B(ori_ori_n34_), .Y(ori_ori_n569_));
  NO2        o0541(.A(k), .B(ori_ori_n199_), .Y(ori_ori_n570_));
  INV        o0542(.A(ori_ori_n332_), .Y(ori_ori_n571_));
  NO2        o0543(.A(ori_ori_n571_), .B(n), .Y(ori_ori_n572_));
  NAi31      o0544(.An(ori_ori_n569_), .B(ori_ori_n572_), .C(ori_ori_n570_), .Y(ori_ori_n573_));
  NO2        o0545(.A(ori_ori_n488_), .B(ori_ori_n164_), .Y(ori_ori_n574_));
  NA3        o0546(.A(ori_ori_n506_), .B(ori_ori_n252_), .C(ori_ori_n135_), .Y(ori_ori_n575_));
  NA2        o0547(.A(ori_ori_n466_), .B(ori_ori_n151_), .Y(ori_ori_n576_));
  NO3        o0548(.A(ori_ori_n358_), .B(ori_ori_n576_), .C(ori_ori_n78_), .Y(ori_ori_n577_));
  AOI210     o0549(.A0(ori_ori_n575_), .A1(ori_ori_n574_), .B0(ori_ori_n577_), .Y(ori_ori_n578_));
  AN3        o0550(.A(f), .B(d), .C(b), .Y(ori_ori_n579_));
  OAI210     o0551(.A0(ori_ori_n579_), .A1(ori_ori_n120_), .B0(n), .Y(ori_ori_n580_));
  NA3        o0552(.A(ori_ori_n466_), .B(ori_ori_n151_), .C(ori_ori_n199_), .Y(ori_ori_n581_));
  AOI210     o0553(.A0(ori_ori_n580_), .A1(ori_ori_n216_), .B0(ori_ori_n581_), .Y(ori_ori_n582_));
  NAi31      o0554(.An(m), .B(n), .C(k), .Y(ori_ori_n583_));
  OR2        o0555(.A(ori_ori_n125_), .B(ori_ori_n56_), .Y(ori_ori_n584_));
  OAI210     o0556(.A0(ori_ori_n584_), .A1(ori_ori_n583_), .B0(ori_ori_n234_), .Y(ori_ori_n585_));
  OAI210     o0557(.A0(ori_ori_n585_), .A1(ori_ori_n582_), .B0(j), .Y(ori_ori_n586_));
  NA3        o0558(.A(ori_ori_n586_), .B(ori_ori_n578_), .C(ori_ori_n573_), .Y(ori_ori_n587_));
  NO4        o0559(.A(ori_ori_n587_), .B(ori_ori_n568_), .C(ori_ori_n559_), .D(ori_ori_n553_), .Y(ori_ori_n588_));
  NA2        o0560(.A(ori_ori_n345_), .B(ori_ori_n154_), .Y(ori_ori_n589_));
  NAi31      o0561(.An(g), .B(h), .C(f), .Y(ori_ori_n590_));
  OA210      o0562(.A0(ori_ori_n489_), .A1(n), .B0(ori_ori_n533_), .Y(ori_ori_n591_));
  NO2        o0563(.A(ori_ori_n591_), .B(ori_ori_n82_), .Y(ori_ori_n592_));
  INV        o0564(.A(ori_ori_n592_), .Y(ori_ori_n593_));
  AOI210     o0565(.A0(ori_ori_n593_), .A1(ori_ori_n589_), .B0(ori_ori_n484_), .Y(ori_ori_n594_));
  NO3        o0566(.A(g), .B(ori_ori_n198_), .C(ori_ori_n52_), .Y(ori_ori_n595_));
  NAi21      o0567(.An(h), .B(j), .Y(ori_ori_n596_));
  NO2        o0568(.A(ori_ori_n473_), .B(ori_ori_n78_), .Y(ori_ori_n597_));
  OAI210     o0569(.A0(ori_ori_n597_), .A1(ori_ori_n357_), .B0(ori_ori_n595_), .Y(ori_ori_n598_));
  OR2        o0570(.A(ori_ori_n63_), .B(ori_ori_n64_), .Y(ori_ori_n599_));
  OR2        o0571(.A(ori_ori_n563_), .B(ori_ori_n599_), .Y(ori_ori_n600_));
  AN2        o0572(.A(h), .B(f), .Y(ori_ori_n601_));
  NA2        o0573(.A(ori_ori_n601_), .B(ori_ori_n35_), .Y(ori_ori_n602_));
  NA2        o0574(.A(ori_ori_n91_), .B(ori_ori_n44_), .Y(ori_ori_n603_));
  OAI220     o0575(.A0(ori_ori_n603_), .A1(ori_ori_n300_), .B0(ori_ori_n602_), .B1(ori_ori_n425_), .Y(ori_ori_n604_));
  AOI210     o0576(.A0(ori_ori_n514_), .A1(ori_ori_n385_), .B0(ori_ori_n47_), .Y(ori_ori_n605_));
  OAI220     o0577(.A0(ori_ori_n536_), .A1(ori_ori_n530_), .B0(ori_ori_n293_), .B1(ori_ori_n482_), .Y(ori_ori_n606_));
  AOI210     o0578(.A0(ori_ori_n606_), .A1(ori_ori_n605_), .B0(ori_ori_n604_), .Y(ori_ori_n607_));
  NA3        o0579(.A(ori_ori_n607_), .B(ori_ori_n600_), .C(ori_ori_n598_), .Y(ori_ori_n608_));
  NO2        o0580(.A(ori_ori_n556_), .B(ori_ori_n56_), .Y(ori_ori_n609_));
  NO2        o0581(.A(ori_ori_n609_), .B(ori_ori_n32_), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n296_), .B(ori_ori_n130_), .Y(ori_ori_n611_));
  NA2        o0583(.A(ori_ori_n122_), .B(ori_ori_n47_), .Y(ori_ori_n612_));
  AOI220     o0584(.A0(ori_ori_n612_), .A1(ori_ori_n487_), .B0(ori_ori_n332_), .B1(ori_ori_n105_), .Y(ori_ori_n613_));
  OA220      o0585(.A0(ori_ori_n613_), .A1(ori_ori_n503_), .B0(ori_ori_n330_), .B1(ori_ori_n103_), .Y(ori_ori_n614_));
  OAI210     o0586(.A0(ori_ori_n611_), .A1(ori_ori_n610_), .B0(ori_ori_n614_), .Y(ori_ori_n615_));
  NO3        o0587(.A(ori_ori_n364_), .B(ori_ori_n180_), .C(ori_ori_n179_), .Y(ori_ori_n616_));
  NA2        o0588(.A(ori_ori_n616_), .B(ori_ori_n214_), .Y(ori_ori_n617_));
  NA3        o0589(.A(ori_ori_n617_), .B(ori_ori_n238_), .C(j), .Y(ori_ori_n618_));
  NO3        o0590(.A(ori_ori_n420_), .B(ori_ori_n161_), .C(i), .Y(ori_ori_n619_));
  NA2        o0591(.A(ori_ori_n424_), .B(ori_ori_n75_), .Y(ori_ori_n620_));
  NO4        o0592(.A(ori_ori_n484_), .B(ori_ori_n620_), .C(ori_ori_n121_), .D(ori_ori_n198_), .Y(ori_ori_n621_));
  INV        o0593(.A(ori_ori_n621_), .Y(ori_ori_n622_));
  NA3        o0594(.A(ori_ori_n622_), .B(ori_ori_n618_), .C(ori_ori_n362_), .Y(ori_ori_n623_));
  NO4        o0595(.A(ori_ori_n623_), .B(ori_ori_n615_), .C(ori_ori_n608_), .D(ori_ori_n594_), .Y(ori_ori_n624_));
  NA4        o0596(.A(ori_ori_n624_), .B(ori_ori_n588_), .C(ori_ori_n547_), .D(ori_ori_n528_), .Y(ori08));
  NO2        o0597(.A(k), .B(h), .Y(ori_ori_n626_));
  AO210      o0598(.A0(ori_ori_n236_), .A1(ori_ori_n408_), .B0(ori_ori_n626_), .Y(ori_ori_n627_));
  NO2        o0599(.A(ori_ori_n627_), .B(ori_ori_n269_), .Y(ori_ori_n628_));
  NA2        o0600(.A(ori_ori_n555_), .B(ori_ori_n75_), .Y(ori_ori_n629_));
  NA2        o0601(.A(ori_ori_n629_), .B(ori_ori_n420_), .Y(ori_ori_n630_));
  NA2        o0602(.A(ori_ori_n630_), .B(ori_ori_n628_), .Y(ori_ori_n631_));
  NA2        o0603(.A(ori_ori_n75_), .B(ori_ori_n102_), .Y(ori_ori_n632_));
  NO2        o0604(.A(ori_ori_n632_), .B(ori_ori_n53_), .Y(ori_ori_n633_));
  NO4        o0605(.A(ori_ori_n343_), .B(ori_ori_n104_), .C(j), .D(ori_ori_n199_), .Y(ori_ori_n634_));
  NA2        o0606(.A(ori_ori_n524_), .B(ori_ori_n216_), .Y(ori_ori_n635_));
  AOI220     o0607(.A0(ori_ori_n635_), .A1(ori_ori_n317_), .B0(ori_ori_n634_), .B1(ori_ori_n633_), .Y(ori_ori_n636_));
  AOI210     o0608(.A0(ori_ori_n524_), .A1(ori_ori_n147_), .B0(ori_ori_n75_), .Y(ori_ori_n637_));
  NA4        o0609(.A(ori_ori_n201_), .B(ori_ori_n130_), .C(ori_ori_n43_), .D(h), .Y(ori_ori_n638_));
  AN2        o0610(.A(l), .B(k), .Y(ori_ori_n639_));
  NA4        o0611(.A(ori_ori_n639_), .B(ori_ori_n101_), .C(ori_ori_n64_), .D(ori_ori_n199_), .Y(ori_ori_n640_));
  OAI210     o0612(.A0(ori_ori_n638_), .A1(g), .B0(ori_ori_n640_), .Y(ori_ori_n641_));
  NA2        o0613(.A(ori_ori_n641_), .B(ori_ori_n637_), .Y(ori_ori_n642_));
  NA4        o0614(.A(ori_ori_n642_), .B(ori_ori_n636_), .C(ori_ori_n631_), .D(ori_ori_n319_), .Y(ori_ori_n643_));
  AN2        o0615(.A(ori_ori_n490_), .B(ori_ori_n87_), .Y(ori_ori_n644_));
  NO4        o0616(.A(ori_ori_n161_), .B(ori_ori_n356_), .C(ori_ori_n104_), .D(g), .Y(ori_ori_n645_));
  NA2        o0617(.A(ori_ori_n645_), .B(ori_ori_n635_), .Y(ori_ori_n646_));
  NO2        o0618(.A(ori_ori_n36_), .B(ori_ori_n198_), .Y(ori_ori_n647_));
  NA2        o0619(.A(ori_ori_n557_), .B(ori_ori_n316_), .Y(ori_ori_n648_));
  NAi31      o0620(.An(ori_ori_n644_), .B(ori_ori_n648_), .C(ori_ori_n646_), .Y(ori_ori_n649_));
  OAI210     o0621(.A0(ori_ori_n506_), .A1(ori_ori_n45_), .B0(ori_ori_n584_), .Y(ori_ori_n650_));
  NO2        o0622(.A(ori_ori_n445_), .B(ori_ori_n122_), .Y(ori_ori_n651_));
  NA2        o0623(.A(ori_ori_n651_), .B(ori_ori_n650_), .Y(ori_ori_n652_));
  NO3        o0624(.A(ori_ori_n285_), .B(ori_ori_n121_), .C(ori_ori_n39_), .Y(ori_ori_n653_));
  NAi21      o0625(.An(ori_ori_n653_), .B(ori_ori_n640_), .Y(ori_ori_n654_));
  NA2        o0626(.A(ori_ori_n627_), .B(ori_ori_n126_), .Y(ori_ori_n655_));
  AOI220     o0627(.A0(ori_ori_n655_), .A1(ori_ori_n363_), .B0(ori_ori_n654_), .B1(ori_ori_n67_), .Y(ori_ori_n656_));
  NA2        o0628(.A(ori_ori_n652_), .B(ori_ori_n656_), .Y(ori_ori_n657_));
  NA2        o0629(.A(ori_ori_n332_), .B(ori_ori_n41_), .Y(ori_ori_n658_));
  NA3        o0630(.A(ori_ori_n617_), .B(ori_ori_n302_), .C(ori_ori_n348_), .Y(ori_ori_n659_));
  NA3        o0631(.A(m), .B(l), .C(k), .Y(ori_ori_n660_));
  NA3        o0632(.A(ori_ori_n105_), .B(k), .C(ori_ori_n78_), .Y(ori_ori_n661_));
  NA2        o0633(.A(ori_ori_n659_), .B(ori_ori_n658_), .Y(ori_ori_n662_));
  NO4        o0634(.A(ori_ori_n662_), .B(ori_ori_n657_), .C(ori_ori_n649_), .D(ori_ori_n643_), .Y(ori_ori_n663_));
  NA2        o0635(.A(ori_ori_n557_), .B(ori_ori_n357_), .Y(ori_ori_n664_));
  INV        o0636(.A(ori_ori_n460_), .Y(ori_ori_n665_));
  NA3        o0637(.A(ori_ori_n665_), .B(ori_ori_n664_), .C(ori_ori_n235_), .Y(ori_ori_n666_));
  NA2        o0638(.A(ori_ori_n639_), .B(ori_ori_n64_), .Y(ori_ori_n667_));
  NO4        o0639(.A(ori_ori_n616_), .B(ori_ori_n161_), .C(n), .D(i), .Y(ori_ori_n668_));
  NOi21      o0640(.An(h), .B(j), .Y(ori_ori_n669_));
  NA2        o0641(.A(ori_ori_n669_), .B(f), .Y(ori_ori_n670_));
  NO2        o0642(.A(ori_ori_n668_), .B(ori_ori_n619_), .Y(ori_ori_n671_));
  NO2        o0643(.A(ori_ori_n671_), .B(ori_ori_n667_), .Y(ori_ori_n672_));
  AOI210     o0644(.A0(ori_ori_n666_), .A1(l), .B0(ori_ori_n672_), .Y(ori_ori_n673_));
  NO2        o0645(.A(j), .B(i), .Y(ori_ori_n674_));
  NA3        o0646(.A(ori_ori_n674_), .B(ori_ori_n71_), .C(l), .Y(ori_ori_n675_));
  NA2        o0647(.A(ori_ori_n674_), .B(ori_ori_n31_), .Y(ori_ori_n676_));
  OR2        o0648(.A(ori_ori_n675_), .B(ori_ori_n535_), .Y(ori_ori_n677_));
  NO3        o0649(.A(ori_ori_n142_), .B(ori_ori_n47_), .C(ori_ori_n102_), .Y(ori_ori_n678_));
  NO3        o0650(.A(ori_ori_n445_), .B(ori_ori_n396_), .C(j), .Y(ori_ori_n679_));
  INV        o0651(.A(j), .Y(ori_ori_n680_));
  NO3        o0652(.A(ori_ori_n269_), .B(ori_ori_n680_), .C(ori_ori_n38_), .Y(ori_ori_n681_));
  AOI210     o0653(.A0(ori_ori_n487_), .A1(n), .B0(ori_ori_n505_), .Y(ori_ori_n682_));
  NA2        o0654(.A(ori_ori_n682_), .B(ori_ori_n508_), .Y(ori_ori_n683_));
  AN3        o0655(.A(ori_ori_n683_), .B(ori_ori_n681_), .C(ori_ori_n90_), .Y(ori_ori_n684_));
  NO3        o0656(.A(ori_ori_n161_), .B(ori_ori_n356_), .C(ori_ori_n104_), .Y(ori_ori_n685_));
  AOI220     o0657(.A0(ori_ori_n685_), .A1(ori_ori_n230_), .B0(ori_ori_n550_), .B1(ori_ori_n277_), .Y(ori_ori_n686_));
  NAi31      o0658(.An(ori_ori_n545_), .B(ori_ori_n84_), .C(ori_ori_n75_), .Y(ori_ori_n687_));
  NA2        o0659(.A(ori_ori_n687_), .B(ori_ori_n686_), .Y(ori_ori_n688_));
  NO2        o0660(.A(ori_ori_n269_), .B(ori_ori_n126_), .Y(ori_ori_n689_));
  AOI220     o0661(.A0(ori_ori_n689_), .A1(ori_ori_n557_), .B0(ori_ori_n653_), .B1(ori_ori_n637_), .Y(ori_ori_n690_));
  NO2        o0662(.A(ori_ori_n660_), .B(ori_ori_n82_), .Y(ori_ori_n691_));
  NA2        o0663(.A(ori_ori_n691_), .B(ori_ori_n534_), .Y(ori_ori_n692_));
  NO2        o0664(.A(ori_ori_n536_), .B(ori_ori_n108_), .Y(ori_ori_n693_));
  OAI210     o0665(.A0(ori_ori_n693_), .A1(ori_ori_n679_), .B0(ori_ori_n605_), .Y(ori_ori_n694_));
  NA3        o0666(.A(ori_ori_n694_), .B(ori_ori_n692_), .C(ori_ori_n690_), .Y(ori_ori_n695_));
  OR3        o0667(.A(ori_ori_n695_), .B(ori_ori_n688_), .C(ori_ori_n684_), .Y(ori_ori_n696_));
  NA3        o0668(.A(ori_ori_n682_), .B(ori_ori_n508_), .C(ori_ori_n507_), .Y(ori_ori_n697_));
  NA4        o0669(.A(ori_ori_n697_), .B(ori_ori_n201_), .C(ori_ori_n408_), .D(ori_ori_n32_), .Y(ori_ori_n698_));
  NO4        o0670(.A(ori_ori_n445_), .B(ori_ori_n392_), .C(j), .D(f), .Y(ori_ori_n699_));
  OAI220     o0671(.A0(ori_ori_n638_), .A1(ori_ori_n629_), .B0(ori_ori_n300_), .B1(ori_ori_n36_), .Y(ori_ori_n700_));
  AOI210     o0672(.A0(ori_ori_n699_), .A1(ori_ori_n242_), .B0(ori_ori_n700_), .Y(ori_ori_n701_));
  NO2        o0673(.A(ori_ori_n83_), .B(ori_ori_n45_), .Y(ori_ori_n702_));
  NA2        o0674(.A(ori_ori_n702_), .B(ori_ori_n572_), .Y(ori_ori_n703_));
  NA3        o0675(.A(ori_ori_n703_), .B(ori_ori_n701_), .C(ori_ori_n698_), .Y(ori_ori_n704_));
  BUFFER     o0676(.A(ori_ori_n691_), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n705_), .B(ori_ori_n221_), .Y(ori_ori_n706_));
  NO2        o0678(.A(ori_ori_n591_), .B(ori_ori_n64_), .Y(ori_ori_n707_));
  AOI210     o0679(.A0(ori_ori_n699_), .A1(ori_ori_n707_), .B0(ori_ori_n304_), .Y(ori_ori_n708_));
  OAI210     o0680(.A0(ori_ori_n660_), .A1(ori_ori_n590_), .B0(ori_ori_n477_), .Y(ori_ori_n709_));
  NA3        o0681(.A(ori_ori_n233_), .B(ori_ori_n55_), .C(b), .Y(ori_ori_n710_));
  AOI220     o0682(.A0(ori_ori_n543_), .A1(ori_ori_n29_), .B0(ori_ori_n424_), .B1(ori_ori_n75_), .Y(ori_ori_n711_));
  NA2        o0683(.A(ori_ori_n711_), .B(ori_ori_n710_), .Y(ori_ori_n712_));
  NA2        o0684(.A(ori_ori_n712_), .B(ori_ori_n709_), .Y(ori_ori_n713_));
  NA3        o0685(.A(ori_ori_n713_), .B(ori_ori_n708_), .C(ori_ori_n706_), .Y(ori_ori_n714_));
  NOi41      o0686(.An(ori_ori_n677_), .B(ori_ori_n714_), .C(ori_ori_n704_), .D(ori_ori_n696_), .Y(ori_ori_n715_));
  NO3        o0687(.A(ori_ori_n310_), .B(ori_ori_n271_), .C(ori_ori_n104_), .Y(ori_ori_n716_));
  NA2        o0688(.A(ori_ori_n716_), .B(ori_ori_n683_), .Y(ori_ori_n717_));
  NO3        o0689(.A(ori_ori_n482_), .B(ori_ori_n85_), .C(h), .Y(ori_ori_n718_));
  NA2        o0690(.A(ori_ori_n718_), .B(ori_ori_n633_), .Y(ori_ori_n719_));
  NA3        o0691(.A(ori_ori_n719_), .B(ori_ori_n717_), .C(ori_ori_n365_), .Y(ori_ori_n720_));
  OR2        o0692(.A(ori_ori_n590_), .B(ori_ori_n83_), .Y(ori_ori_n721_));
  NOi31      o0693(.An(b), .B(d), .C(a), .Y(ori_ori_n722_));
  NO2        o0694(.A(ori_ori_n722_), .B(ori_ori_n542_), .Y(ori_ori_n723_));
  NO2        o0695(.A(ori_ori_n723_), .B(n), .Y(ori_ori_n724_));
  NOi21      o0696(.An(ori_ori_n711_), .B(ori_ori_n724_), .Y(ori_ori_n725_));
  NO2        o0697(.A(ori_ori_n725_), .B(ori_ori_n721_), .Y(ori_ori_n726_));
  NO2        o0698(.A(ori_ori_n506_), .B(ori_ori_n75_), .Y(ori_ori_n727_));
  NA2        o0699(.A(ori_ori_n716_), .B(ori_ori_n727_), .Y(ori_ori_n728_));
  OAI210     o0700(.A0(ori_ori_n638_), .A1(ori_ori_n358_), .B0(ori_ori_n728_), .Y(ori_ori_n729_));
  NO2        o0701(.A(ori_ori_n616_), .B(n), .Y(ori_ori_n730_));
  AOI220     o0702(.A0(ori_ori_n689_), .A1(ori_ori_n595_), .B0(ori_ori_n730_), .B1(ori_ori_n628_), .Y(ori_ori_n731_));
  NO2        o0703(.A(ori_ori_n290_), .B(ori_ori_n220_), .Y(ori_ori_n732_));
  OAI210     o0704(.A0(ori_ori_n87_), .A1(ori_ori_n84_), .B0(ori_ori_n732_), .Y(ori_ori_n733_));
  INV        o0705(.A(ori_ori_n733_), .Y(ori_ori_n734_));
  NA2        o0706(.A(ori_ori_n645_), .B(ori_ori_n318_), .Y(ori_ori_n735_));
  NA2        o0707(.A(ori_ori_n538_), .B(ori_ori_n333_), .Y(ori_ori_n736_));
  AN2        o0708(.A(ori_ori_n736_), .B(ori_ori_n735_), .Y(ori_ori_n737_));
  NAi31      o0709(.An(ori_ori_n734_), .B(ori_ori_n737_), .C(ori_ori_n731_), .Y(ori_ori_n738_));
  NO4        o0710(.A(ori_ori_n738_), .B(ori_ori_n729_), .C(ori_ori_n726_), .D(ori_ori_n720_), .Y(ori_ori_n739_));
  NA4        o0711(.A(ori_ori_n739_), .B(ori_ori_n715_), .C(ori_ori_n673_), .D(ori_ori_n663_), .Y(ori09));
  INV        o0712(.A(ori_ori_n113_), .Y(ori_ori_n741_));
  NA2        o0713(.A(f), .B(e), .Y(ori_ori_n742_));
  NA4        o0714(.A(ori_ori_n279_), .B(ori_ori_n155_), .C(ori_ori_n245_), .D(ori_ori_n110_), .Y(ori_ori_n743_));
  AOI210     o0715(.A0(ori_ori_n743_), .A1(g), .B0(ori_ori_n430_), .Y(ori_ori_n744_));
  NO2        o0716(.A(ori_ori_n744_), .B(ori_ori_n742_), .Y(ori_ori_n745_));
  NA2        o0717(.A(ori_ori_n401_), .B(e), .Y(ori_ori_n746_));
  NO2        o0718(.A(ori_ori_n746_), .B(ori_ori_n470_), .Y(ori_ori_n747_));
  AOI210     o0719(.A0(ori_ori_n745_), .A1(ori_ori_n741_), .B0(ori_ori_n747_), .Y(ori_ori_n748_));
  NA3        o0720(.A(m), .B(l), .C(i), .Y(ori_ori_n749_));
  OAI220     o0721(.A0(ori_ori_n536_), .A1(ori_ori_n749_), .B0(ori_ori_n323_), .B1(ori_ori_n483_), .Y(ori_ori_n750_));
  NAi21      o0722(.An(ori_ori_n750_), .B(ori_ori_n397_), .Y(ori_ori_n751_));
  NA3        o0723(.A(ori_ori_n721_), .B(ori_ori_n513_), .C(ori_ori_n477_), .Y(ori_ori_n752_));
  OA210      o0724(.A0(ori_ori_n752_), .A1(ori_ori_n751_), .B0(ori_ori_n724_), .Y(ori_ori_n753_));
  INV        o0725(.A(ori_ori_n307_), .Y(ori_ori_n754_));
  NO2        o0726(.A(ori_ori_n118_), .B(ori_ori_n116_), .Y(ori_ori_n755_));
  NOi31      o0727(.An(k), .B(m), .C(l), .Y(ori_ori_n756_));
  NO2        o0728(.A(ori_ori_n309_), .B(ori_ori_n756_), .Y(ori_ori_n757_));
  AOI210     o0729(.A0(ori_ori_n757_), .A1(ori_ori_n755_), .B0(ori_ori_n540_), .Y(ori_ori_n758_));
  NA2        o0730(.A(ori_ori_n710_), .B(ori_ori_n300_), .Y(ori_ori_n759_));
  NA2        o0731(.A(ori_ori_n311_), .B(ori_ori_n313_), .Y(ori_ori_n760_));
  OAI210     o0732(.A0(ori_ori_n192_), .A1(ori_ori_n198_), .B0(ori_ori_n760_), .Y(ori_ori_n761_));
  AOI220     o0733(.A0(ori_ori_n761_), .A1(ori_ori_n759_), .B0(ori_ori_n758_), .B1(ori_ori_n754_), .Y(ori_ori_n762_));
  NA2        o0734(.A(ori_ori_n157_), .B(ori_ori_n106_), .Y(ori_ori_n763_));
  NA3        o0735(.A(ori_ori_n763_), .B(ori_ori_n627_), .C(ori_ori_n126_), .Y(ori_ori_n764_));
  NA3        o0736(.A(ori_ori_n764_), .B(ori_ori_n177_), .C(ori_ori_n30_), .Y(ori_ori_n765_));
  NA4        o0737(.A(ori_ori_n765_), .B(ori_ori_n762_), .C(ori_ori_n558_), .D(ori_ori_n73_), .Y(ori_ori_n766_));
  NO2        o0738(.A(ori_ori_n532_), .B(ori_ori_n456_), .Y(ori_ori_n767_));
  NA2        o0739(.A(ori_ori_n767_), .B(ori_ori_n177_), .Y(ori_ori_n768_));
  NOi21      o0740(.An(f), .B(d), .Y(ori_ori_n769_));
  NA2        o0741(.A(ori_ori_n769_), .B(m), .Y(ori_ori_n770_));
  NO2        o0742(.A(ori_ori_n770_), .B(ori_ori_n50_), .Y(ori_ori_n771_));
  NA2        o0743(.A(ori_ori_n771_), .B(ori_ori_n497_), .Y(ori_ori_n772_));
  NA3        o0744(.A(ori_ori_n279_), .B(ori_ori_n245_), .C(ori_ori_n110_), .Y(ori_ori_n773_));
  AN2        o0745(.A(f), .B(d), .Y(ori_ori_n774_));
  NA3        o0746(.A(ori_ori_n436_), .B(ori_ori_n774_), .C(ori_ori_n75_), .Y(ori_ori_n775_));
  NO3        o0747(.A(ori_ori_n775_), .B(ori_ori_n64_), .C(ori_ori_n199_), .Y(ori_ori_n776_));
  NA2        o0748(.A(ori_ori_n773_), .B(ori_ori_n776_), .Y(ori_ori_n777_));
  NAi41      o0749(.An(ori_ori_n450_), .B(ori_ori_n777_), .C(ori_ori_n772_), .D(ori_ori_n768_), .Y(ori_ori_n778_));
  NO4        o0750(.A(ori_ori_n556_), .B(ori_ori_n122_), .C(ori_ori_n295_), .D(ori_ori_n143_), .Y(ori_ori_n779_));
  NO2        o0751(.A(ori_ori_n583_), .B(ori_ori_n295_), .Y(ori_ori_n780_));
  INV        o0752(.A(ori_ori_n779_), .Y(ori_ori_n781_));
  NA3        o0753(.A(ori_ori_n151_), .B(ori_ori_n101_), .C(ori_ori_n100_), .Y(ori_ori_n782_));
  OAI220     o0754(.A0(ori_ori_n775_), .A1(ori_ori_n387_), .B0(ori_ori_n307_), .B1(ori_ori_n782_), .Y(ori_ori_n783_));
  NOi31      o0755(.An(ori_ori_n207_), .B(ori_ori_n783_), .C(ori_ori_n275_), .Y(ori_ori_n784_));
  NA2        o0756(.A(c), .B(ori_ori_n107_), .Y(ori_ori_n785_));
  NO2        o0757(.A(ori_ori_n785_), .B(ori_ori_n369_), .Y(ori_ori_n786_));
  NA3        o0758(.A(ori_ori_n786_), .B(ori_ori_n468_), .C(f), .Y(ori_ori_n787_));
  OR2        o0759(.A(ori_ori_n590_), .B(ori_ori_n493_), .Y(ori_ori_n788_));
  INV        o0760(.A(ori_ori_n788_), .Y(ori_ori_n789_));
  NA2        o0761(.A(ori_ori_n723_), .B(ori_ori_n103_), .Y(ori_ori_n790_));
  NA2        o0762(.A(ori_ori_n790_), .B(ori_ori_n789_), .Y(ori_ori_n791_));
  NA4        o0763(.A(ori_ori_n791_), .B(ori_ori_n787_), .C(ori_ori_n784_), .D(ori_ori_n781_), .Y(ori_ori_n792_));
  NO4        o0764(.A(ori_ori_n792_), .B(ori_ori_n778_), .C(ori_ori_n766_), .D(ori_ori_n753_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n126_), .B(ori_ori_n122_), .Y(ori_ori_n794_));
  NO2        o0766(.A(ori_ori_n214_), .B(ori_ori_n208_), .Y(ori_ori_n795_));
  AOI220     o0767(.A0(ori_ori_n795_), .A1(ori_ori_n211_), .B0(ori_ori_n273_), .B1(ori_ori_n794_), .Y(ori_ori_n796_));
  NO2        o0768(.A(ori_ori_n387_), .B(ori_ori_n742_), .Y(ori_ori_n797_));
  INV        o0769(.A(ori_ori_n796_), .Y(ori_ori_n798_));
  NA2        o0770(.A(e), .B(d), .Y(ori_ori_n799_));
  OAI220     o0771(.A0(ori_ori_n799_), .A1(c), .B0(ori_ori_n290_), .B1(d), .Y(ori_ori_n800_));
  NA3        o0772(.A(ori_ori_n800_), .B(ori_ori_n413_), .C(ori_ori_n466_), .Y(ori_ori_n801_));
  AOI210     o0773(.A0(ori_ori_n473_), .A1(ori_ori_n168_), .B0(ori_ori_n214_), .Y(ori_ori_n802_));
  AOI210     o0774(.A0(ori_ori_n557_), .A1(ori_ori_n316_), .B0(ori_ori_n802_), .Y(ori_ori_n803_));
  INV        o0775(.A(ori_ori_n155_), .Y(ori_ori_n804_));
  NA2        o0776(.A(ori_ori_n776_), .B(ori_ori_n804_), .Y(ori_ori_n805_));
  NA3        o0777(.A(ori_ori_n156_), .B(ori_ori_n76_), .C(ori_ori_n32_), .Y(ori_ori_n806_));
  NA4        o0778(.A(ori_ori_n806_), .B(ori_ori_n805_), .C(ori_ori_n803_), .D(ori_ori_n801_), .Y(ori_ori_n807_));
  NO2        o0779(.A(ori_ori_n807_), .B(ori_ori_n798_), .Y(ori_ori_n808_));
  OR2        o0780(.A(ori_ori_n629_), .B(ori_ori_n202_), .Y(ori_ori_n809_));
  OAI220     o0781(.A0(ori_ori_n556_), .A1(ori_ori_n56_), .B0(ori_ori_n271_), .B1(j), .Y(ori_ori_n810_));
  AOI220     o0782(.A0(ori_ori_n810_), .A1(ori_ori_n780_), .B0(ori_ori_n548_), .B1(ori_ori_n555_), .Y(ori_ori_n811_));
  OAI210     o0783(.A0(ori_ori_n746_), .A1(ori_ori_n158_), .B0(ori_ori_n811_), .Y(ori_ori_n812_));
  AN2        o0784(.A(ori_ori_n759_), .B(ori_ori_n750_), .Y(ori_ori_n813_));
  NO2        o0785(.A(ori_ori_n813_), .B(ori_ori_n812_), .Y(ori_ori_n814_));
  AO220      o0786(.A0(ori_ori_n413_), .A1(ori_ori_n669_), .B0(ori_ori_n163_), .B1(f), .Y(ori_ori_n815_));
  OAI210     o0787(.A0(ori_ori_n815_), .A1(ori_ori_n416_), .B0(ori_ori_n800_), .Y(ori_ori_n816_));
  NA2        o0788(.A(ori_ori_n752_), .B(ori_ori_n633_), .Y(ori_ori_n817_));
  AN4        o0789(.A(ori_ori_n817_), .B(ori_ori_n816_), .C(ori_ori_n814_), .D(ori_ori_n809_), .Y(ori_ori_n818_));
  NA4        o0790(.A(ori_ori_n818_), .B(ori_ori_n808_), .C(ori_ori_n793_), .D(ori_ori_n748_), .Y(ori12));
  NO2        o0791(.A(ori_ori_n411_), .B(c), .Y(ori_ori_n820_));
  NO4        o0792(.A(ori_ori_n400_), .B(ori_ori_n236_), .C(ori_ori_n529_), .D(ori_ori_n199_), .Y(ori_ori_n821_));
  NA2        o0793(.A(ori_ori_n821_), .B(ori_ori_n820_), .Y(ori_ori_n822_));
  NO2        o0794(.A(ori_ori_n411_), .B(ori_ori_n107_), .Y(ori_ori_n823_));
  NO2        o0795(.A(ori_ori_n755_), .B(ori_ori_n323_), .Y(ori_ori_n824_));
  NO2        o0796(.A(ori_ori_n590_), .B(ori_ori_n343_), .Y(ori_ori_n825_));
  AOI220     o0797(.A0(ori_ori_n825_), .A1(ori_ori_n495_), .B0(ori_ori_n824_), .B1(ori_ori_n823_), .Y(ori_ori_n826_));
  NA3        o0798(.A(ori_ori_n826_), .B(ori_ori_n822_), .C(ori_ori_n399_), .Y(ori_ori_n827_));
  AOI210     o0799(.A0(ori_ori_n217_), .A1(ori_ori_n306_), .B0(ori_ori_n189_), .Y(ori_ori_n828_));
  OR2        o0800(.A(ori_ori_n828_), .B(ori_ori_n821_), .Y(ori_ori_n829_));
  AOI210     o0801(.A0(ori_ori_n303_), .A1(ori_ori_n354_), .B0(ori_ori_n199_), .Y(ori_ori_n830_));
  OAI210     o0802(.A0(ori_ori_n830_), .A1(ori_ori_n829_), .B0(ori_ori_n364_), .Y(ori_ori_n831_));
  NO2        o0803(.A(ori_ori_n569_), .B(ori_ori_n246_), .Y(ori_ori_n832_));
  NO2        o0804(.A(ori_ori_n536_), .B(ori_ori_n749_), .Y(ori_ori_n833_));
  NO2        o0805(.A(ori_ori_n142_), .B(ori_ori_n220_), .Y(ori_ori_n834_));
  NA3        o0806(.A(ori_ori_n834_), .B(ori_ori_n223_), .C(i), .Y(ori_ori_n835_));
  NA2        o0807(.A(ori_ori_n835_), .B(ori_ori_n831_), .Y(ori_ori_n836_));
  OR2        o0808(.A(ori_ori_n291_), .B(ori_ori_n823_), .Y(ori_ori_n837_));
  NA2        o0809(.A(ori_ori_n837_), .B(ori_ori_n324_), .Y(ori_ori_n838_));
  NO3        o0810(.A(ori_ori_n122_), .B(ori_ori_n143_), .C(ori_ori_n199_), .Y(ori_ori_n839_));
  NA2        o0811(.A(ori_ori_n839_), .B(ori_ori_n487_), .Y(ori_ori_n840_));
  NA4        o0812(.A(ori_ori_n401_), .B(ori_ori_n394_), .C(ori_ori_n169_), .D(g), .Y(ori_ori_n841_));
  NA3        o0813(.A(ori_ori_n841_), .B(ori_ori_n840_), .C(ori_ori_n838_), .Y(ori_ori_n842_));
  NO3        o0814(.A(ori_ori_n593_), .B(ori_ori_n83_), .C(ori_ori_n43_), .Y(ori_ori_n843_));
  NO4        o0815(.A(ori_ori_n843_), .B(ori_ori_n842_), .C(ori_ori_n836_), .D(ori_ori_n827_), .Y(ori_ori_n844_));
  NA2        o0816(.A(ori_ori_n506_), .B(ori_ori_n135_), .Y(ori_ori_n845_));
  NOi21      o0817(.An(ori_ori_n32_), .B(ori_ori_n583_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n846_), .B(ori_ori_n845_), .Y(ori_ori_n847_));
  OAI210     o0819(.A0(ori_ori_n234_), .A1(ori_ori_n43_), .B0(ori_ori_n847_), .Y(ori_ori_n848_));
  INV        o0820(.A(ori_ori_n289_), .Y(ori_ori_n849_));
  NO2        o0821(.A(ori_ori_n47_), .B(ori_ori_n43_), .Y(ori_ori_n850_));
  NO2        o0822(.A(ori_ori_n463_), .B(ori_ori_n271_), .Y(ori_ori_n851_));
  INV        o0823(.A(ori_ori_n851_), .Y(ori_ori_n852_));
  NO2        o0824(.A(ori_ori_n852_), .B(ori_ori_n135_), .Y(ori_ori_n853_));
  INV        o0825(.A(ori_ori_n337_), .Y(ori_ori_n854_));
  NO4        o0826(.A(ori_ori_n854_), .B(ori_ori_n853_), .C(ori_ori_n849_), .D(ori_ori_n848_), .Y(ori_ori_n855_));
  NA2        o0827(.A(ori_ori_n316_), .B(g), .Y(ori_ori_n856_));
  NA2        o0828(.A(ori_ori_n154_), .B(i), .Y(ori_ori_n857_));
  NA2        o0829(.A(ori_ori_n44_), .B(i), .Y(ori_ori_n858_));
  OAI220     o0830(.A0(ori_ori_n858_), .A1(ori_ori_n188_), .B0(ori_ori_n857_), .B1(ori_ori_n83_), .Y(ori_ori_n859_));
  AOI210     o0831(.A0(ori_ori_n378_), .A1(ori_ori_n35_), .B0(ori_ori_n859_), .Y(ori_ori_n860_));
  NO2        o0832(.A(ori_ori_n135_), .B(ori_ori_n75_), .Y(ori_ori_n861_));
  OR2        o0833(.A(ori_ori_n861_), .B(ori_ori_n505_), .Y(ori_ori_n862_));
  NA2        o0834(.A(ori_ori_n506_), .B(ori_ori_n346_), .Y(ori_ori_n863_));
  AOI210     o0835(.A0(ori_ori_n863_), .A1(n), .B0(ori_ori_n862_), .Y(ori_ori_n864_));
  OAI220     o0836(.A0(ori_ori_n864_), .A1(ori_ori_n856_), .B0(ori_ori_n860_), .B1(ori_ori_n300_), .Y(ori_ori_n865_));
  NO2        o0837(.A(ori_ori_n590_), .B(ori_ori_n456_), .Y(ori_ori_n866_));
  NA3        o0838(.A(ori_ori_n311_), .B(ori_ori_n560_), .C(i), .Y(ori_ori_n867_));
  OAI210     o0839(.A0(ori_ori_n396_), .A1(ori_ori_n279_), .B0(ori_ori_n867_), .Y(ori_ori_n868_));
  OAI210     o0840(.A0(ori_ori_n868_), .A1(ori_ori_n866_), .B0(ori_ori_n605_), .Y(ori_ori_n869_));
  NA2        o0841(.A(ori_ori_n544_), .B(ori_ori_n105_), .Y(ori_ori_n870_));
  OR3        o0842(.A(ori_ori_n279_), .B(ori_ori_n392_), .C(f), .Y(ori_ori_n871_));
  NA3        o0843(.A(ori_ori_n560_), .B(ori_ori_n71_), .C(i), .Y(ori_ori_n872_));
  OA220      o0844(.A0(ori_ori_n872_), .A1(ori_ori_n870_), .B0(ori_ori_n871_), .B1(ori_ori_n535_), .Y(ori_ori_n873_));
  NA3        o0845(.A(ori_ori_n292_), .B(ori_ori_n109_), .C(g), .Y(ori_ori_n874_));
  AOI210     o0846(.A0(ori_ori_n602_), .A1(ori_ori_n874_), .B0(m), .Y(ori_ori_n875_));
  OAI210     o0847(.A0(ori_ori_n875_), .A1(ori_ori_n824_), .B0(ori_ori_n291_), .Y(ori_ori_n876_));
  INV        o0848(.A(ori_ori_n620_), .Y(ori_ori_n877_));
  INV        o0849(.A(ori_ori_n397_), .Y(ori_ori_n878_));
  INV        o0850(.A(ori_ori_n872_), .Y(ori_ori_n879_));
  AOI220     o0851(.A0(ori_ori_n879_), .A1(ori_ori_n242_), .B0(ori_ori_n878_), .B1(ori_ori_n877_), .Y(ori_ori_n880_));
  NA4        o0852(.A(ori_ori_n880_), .B(ori_ori_n876_), .C(ori_ori_n873_), .D(ori_ori_n869_), .Y(ori_ori_n881_));
  NO2        o0853(.A(ori_ori_n343_), .B(ori_ori_n82_), .Y(ori_ori_n882_));
  OAI210     o0854(.A0(ori_ori_n882_), .A1(ori_ori_n832_), .B0(ori_ori_n221_), .Y(ori_ori_n883_));
  NA2        o0855(.A(ori_ori_n592_), .B(ori_ori_n79_), .Y(ori_ori_n884_));
  NO2        o0856(.A(ori_ori_n419_), .B(ori_ori_n199_), .Y(ori_ori_n885_));
  AOI220     o0857(.A0(ori_ori_n885_), .A1(ori_ori_n347_), .B0(ori_ori_n837_), .B1(ori_ori_n203_), .Y(ori_ori_n886_));
  AOI220     o0858(.A0(ori_ori_n825_), .A1(ori_ori_n834_), .B0(ori_ori_n534_), .B1(ori_ori_n81_), .Y(ori_ori_n887_));
  NA4        o0859(.A(ori_ori_n887_), .B(ori_ori_n886_), .C(ori_ori_n884_), .D(ori_ori_n883_), .Y(ori_ori_n888_));
  OAI210     o0860(.A0(ori_ori_n878_), .A1(ori_ori_n833_), .B0(ori_ori_n495_), .Y(ori_ori_n889_));
  NA2        o0861(.A(ori_ori_n875_), .B(ori_ori_n823_), .Y(ori_ori_n890_));
  NA2        o0862(.A(ori_ori_n574_), .B(ori_ori_n487_), .Y(ori_ori_n891_));
  NA3        o0863(.A(ori_ori_n891_), .B(ori_ori_n890_), .C(ori_ori_n889_), .Y(ori_ori_n892_));
  NO4        o0864(.A(ori_ori_n892_), .B(ori_ori_n888_), .C(ori_ori_n881_), .D(ori_ori_n865_), .Y(ori_ori_n893_));
  NAi31      o0865(.An(ori_ori_n131_), .B(ori_ori_n380_), .C(n), .Y(ori_ori_n894_));
  NO3        o0866(.A(ori_ori_n116_), .B(ori_ori_n309_), .C(ori_ori_n756_), .Y(ori_ori_n895_));
  NO2        o0867(.A(ori_ori_n895_), .B(ori_ori_n894_), .Y(ori_ori_n896_));
  NO3        o0868(.A(ori_ori_n253_), .B(ori_ori_n131_), .C(ori_ori_n369_), .Y(ori_ori_n897_));
  AOI210     o0869(.A0(ori_ori_n897_), .A1(ori_ori_n457_), .B0(ori_ori_n896_), .Y(ori_ori_n898_));
  INV        o0870(.A(ori_ori_n898_), .Y(ori_ori_n899_));
  NA2        o0871(.A(ori_ori_n214_), .B(ori_ori_n159_), .Y(ori_ori_n900_));
  NO3        o0872(.A(ori_ori_n277_), .B(ori_ori_n401_), .C(ori_ori_n163_), .Y(ori_ori_n901_));
  NOi31      o0873(.An(ori_ori_n900_), .B(ori_ori_n901_), .C(ori_ori_n199_), .Y(ori_ori_n902_));
  NAi21      o0874(.An(ori_ori_n506_), .B(ori_ori_n885_), .Y(ori_ori_n903_));
  NA2        o0875(.A(ori_ori_n442_), .B(g), .Y(ori_ori_n904_));
  NA2        o0876(.A(ori_ori_n904_), .B(ori_ori_n903_), .Y(ori_ori_n905_));
  NA2        o0877(.A(ori_ori_n828_), .B(ori_ori_n820_), .Y(ori_ori_n906_));
  OAI220     o0878(.A0(ori_ori_n825_), .A1(ori_ori_n833_), .B0(ori_ori_n497_), .B1(ori_ori_n386_), .Y(ori_ori_n907_));
  NA3        o0879(.A(ori_ori_n907_), .B(ori_ori_n906_), .C(ori_ori_n554_), .Y(ori_ori_n908_));
  OAI210     o0880(.A0(ori_ori_n828_), .A1(ori_ori_n821_), .B0(ori_ori_n900_), .Y(ori_ori_n909_));
  NA3        o0881(.A(ori_ori_n863_), .B(ori_ori_n447_), .C(ori_ori_n44_), .Y(ori_ori_n910_));
  INV        o0882(.A(ori_ori_n299_), .Y(ori_ori_n911_));
  NA3        o0883(.A(ori_ori_n911_), .B(ori_ori_n910_), .C(ori_ori_n909_), .Y(ori_ori_n912_));
  OR2        o0884(.A(ori_ori_n912_), .B(ori_ori_n908_), .Y(ori_ori_n913_));
  NO4        o0885(.A(ori_ori_n913_), .B(ori_ori_n905_), .C(ori_ori_n902_), .D(ori_ori_n899_), .Y(ori_ori_n914_));
  NA4        o0886(.A(ori_ori_n914_), .B(ori_ori_n893_), .C(ori_ori_n855_), .D(ori_ori_n844_), .Y(ori13));
  AN2        o0887(.A(c), .B(b), .Y(ori_ori_n916_));
  NAi32      o0888(.An(d), .Bn(c), .C(e), .Y(ori_ori_n917_));
  AN2        o0889(.A(d), .B(c), .Y(ori_ori_n918_));
  NA2        o0890(.A(ori_ori_n918_), .B(ori_ori_n107_), .Y(ori_ori_n919_));
  NO3        o0891(.A(m), .B(i), .C(h), .Y(ori_ori_n920_));
  NA3        o0892(.A(k), .B(j), .C(i), .Y(ori_ori_n921_));
  NO2        o0893(.A(f), .B(c), .Y(ori_ori_n922_));
  NOi21      o0894(.An(ori_ori_n922_), .B(ori_ori_n400_), .Y(ori_ori_n923_));
  AN3        o0895(.A(g), .B(f), .C(c), .Y(ori_ori_n924_));
  NA3        o0896(.A(l), .B(k), .C(j), .Y(ori_ori_n925_));
  NA2        o0897(.A(i), .B(h), .Y(ori_ori_n926_));
  NO3        o0898(.A(ori_ori_n926_), .B(ori_ori_n925_), .C(ori_ori_n122_), .Y(ori_ori_n927_));
  NO3        o0899(.A(ori_ori_n132_), .B(ori_ori_n260_), .C(ori_ori_n199_), .Y(ori_ori_n928_));
  NA3        o0900(.A(c), .B(b), .C(a), .Y(ori_ori_n929_));
  NO2        o0901(.A(ori_ori_n483_), .B(ori_ori_n540_), .Y(ori_ori_n930_));
  NA4        o0902(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .D(ori_ori_n198_), .Y(ori_ori_n931_));
  NA4        o0903(.A(ori_ori_n521_), .B(m), .C(ori_ori_n104_), .D(ori_ori_n198_), .Y(ori_ori_n932_));
  NA3        o0904(.A(ori_ori_n932_), .B(ori_ori_n338_), .C(ori_ori_n931_), .Y(ori_ori_n933_));
  NO2        o0905(.A(ori_ori_n933_), .B(ori_ori_n930_), .Y(ori_ori_n934_));
  NOi41      o0906(.An(ori_ori_n721_), .B(ori_ori_n761_), .C(ori_ori_n751_), .D(ori_ori_n647_), .Y(ori_ori_n935_));
  OAI220     o0907(.A0(ori_ori_n935_), .A1(ori_ori_n620_), .B0(ori_ori_n934_), .B1(ori_ori_n533_), .Y(ori_ori_n936_));
  NOi31      o0908(.An(m), .B(n), .C(f), .Y(ori_ori_n937_));
  NA2        o0909(.A(ori_ori_n937_), .B(ori_ori_n49_), .Y(ori_ori_n938_));
  AN2        o0910(.A(e), .B(c), .Y(ori_ori_n939_));
  NA2        o0911(.A(ori_ori_n939_), .B(a), .Y(ori_ori_n940_));
  OAI220     o0912(.A0(ori_ori_n940_), .A1(ori_ori_n938_), .B0(ori_ori_n788_), .B1(ori_ori_n385_), .Y(ori_ori_n941_));
  NA2        o0913(.A(ori_ori_n466_), .B(l), .Y(ori_ori_n942_));
  NO2        o0914(.A(ori_ori_n260_), .B(a), .Y(ori_ori_n943_));
  NO2        o0915(.A(ori_ori_n78_), .B(g), .Y(ori_ori_n944_));
  NO3        o0916(.A(ori_ori_n941_), .B(ori_ori_n936_), .C(ori_ori_n734_), .Y(ori_ori_n945_));
  NA2        o0917(.A(c), .B(b), .Y(ori_ori_n946_));
  NO2        o0918(.A(ori_ori_n632_), .B(ori_ori_n946_), .Y(ori_ori_n947_));
  OAI210     o0919(.A0(ori_ori_n770_), .A1(ori_ori_n744_), .B0(ori_ori_n374_), .Y(ori_ori_n948_));
  OAI210     o0920(.A0(ori_ori_n948_), .A1(ori_ori_n771_), .B0(ori_ori_n947_), .Y(ori_ori_n949_));
  NAi21      o0921(.An(ori_ori_n382_), .B(ori_ori_n947_), .Y(ori_ori_n950_));
  OAI210     o0922(.A0(ori_ori_n500_), .A1(ori_ori_n37_), .B0(ori_ori_n943_), .Y(ori_ori_n951_));
  NA2        o0923(.A(ori_ori_n951_), .B(ori_ori_n950_), .Y(ori_ori_n952_));
  OAI210     o0924(.A0(ori_ori_n244_), .A1(ori_ori_n262_), .B0(g), .Y(ori_ori_n953_));
  NAi21      o0925(.An(f), .B(d), .Y(ori_ori_n954_));
  NO2        o0926(.A(ori_ori_n954_), .B(ori_ori_n929_), .Y(ori_ori_n955_));
  INV        o0927(.A(ori_ori_n955_), .Y(ori_ori_n956_));
  NO2        o0928(.A(ori_ori_n953_), .B(ori_ori_n956_), .Y(ori_ori_n957_));
  AOI210     o0929(.A0(ori_ori_n957_), .A1(ori_ori_n105_), .B0(ori_ori_n952_), .Y(ori_ori_n958_));
  NA2        o0930(.A(ori_ori_n942_), .B(ori_ori_n155_), .Y(ori_ori_n959_));
  NA2        o0931(.A(ori_ori_n404_), .B(ori_ori_n955_), .Y(ori_ori_n960_));
  NA4        o0932(.A(ori_ori_n960_), .B(ori_ori_n958_), .C(ori_ori_n949_), .D(ori_ori_n945_), .Y(ori00));
  NA2        o0933(.A(ori_ori_n797_), .B(ori_ori_n834_), .Y(ori_ori_n962_));
  INV        o0934(.A(ori_ori_n644_), .Y(ori_ori_n963_));
  NA2        o0935(.A(ori_ori_n963_), .B(ori_ori_n962_), .Y(ori_ori_n964_));
  NA2        o0936(.A(ori_ori_n468_), .B(f), .Y(ori_ori_n965_));
  OAI210     o0937(.A0(ori_ori_n895_), .A1(ori_ori_n38_), .B0(ori_ori_n576_), .Y(ori_ori_n966_));
  NA3        o0938(.A(ori_ori_n966_), .B(ori_ori_n241_), .C(n), .Y(ori_ori_n967_));
  AOI210     o0939(.A0(ori_ori_n967_), .A1(ori_ori_n965_), .B0(ori_ori_n919_), .Y(ori_ori_n968_));
  NO2        o0940(.A(ori_ori_n968_), .B(ori_ori_n964_), .Y(ori_ori_n969_));
  NA3        o0941(.A(ori_ori_n156_), .B(ori_ori_n44_), .C(ori_ori_n43_), .Y(ori_ori_n970_));
  NA3        o0942(.A(d), .B(ori_ori_n52_), .C(b), .Y(ori_ori_n971_));
  NO2        o0943(.A(ori_ori_n971_), .B(ori_ori_n970_), .Y(ori_ori_n972_));
  NO4        o0944(.A(ori_ori_n448_), .B(ori_ori_n326_), .C(ori_ori_n946_), .D(ori_ori_n55_), .Y(ori_ori_n973_));
  NA3        o0945(.A(ori_ori_n348_), .B(ori_ori_n206_), .C(g), .Y(ori_ori_n974_));
  OR2        o0946(.A(ori_ori_n974_), .B(ori_ori_n971_), .Y(ori_ori_n975_));
  NO2        o0947(.A(h), .B(g), .Y(ori_ori_n976_));
  NA4        o0948(.A(ori_ori_n457_), .B(ori_ori_n427_), .C(ori_ori_n976_), .D(ori_ori_n916_), .Y(ori_ori_n977_));
  OAI220     o0949(.A0(ori_ori_n483_), .A1(ori_ori_n540_), .B0(ori_ori_n83_), .B1(ori_ori_n82_), .Y(ori_ori_n978_));
  AOI220     o0950(.A0(ori_ori_n978_), .A1(ori_ori_n490_), .B0(ori_ori_n839_), .B1(ori_ori_n522_), .Y(ori_ori_n979_));
  AOI220     o0951(.A0(ori_ori_n286_), .A1(ori_ori_n230_), .B0(ori_ori_n165_), .B1(ori_ori_n139_), .Y(ori_ori_n980_));
  NA4        o0952(.A(ori_ori_n980_), .B(ori_ori_n979_), .C(ori_ori_n977_), .D(ori_ori_n975_), .Y(ori_ori_n981_));
  NO3        o0953(.A(ori_ori_n981_), .B(ori_ori_n973_), .C(ori_ori_n248_), .Y(ori_ori_n982_));
  AOI210     o0954(.A0(ori_ori_n230_), .A1(ori_ori_n316_), .B0(ori_ori_n525_), .Y(ori_ori_n983_));
  NA2        o0955(.A(ori_ori_n983_), .B(ori_ori_n145_), .Y(ori_ori_n984_));
  NO2        o0956(.A(ori_ori_n222_), .B(ori_ori_n169_), .Y(ori_ori_n985_));
  NA2        o0957(.A(ori_ori_n985_), .B(ori_ori_n386_), .Y(ori_ori_n986_));
  INV        o0958(.A(ori_ori_n986_), .Y(ori_ori_n987_));
  NO3        o0959(.A(ori_ori_n987_), .B(ori_ori_n984_), .C(ori_ori_n476_), .Y(ori_ori_n988_));
  AN3        o0960(.A(ori_ori_n988_), .B(ori_ori_n982_), .C(ori_ori_n523_), .Y(ori_ori_n989_));
  NA3        o0961(.A(ori_ori_n937_), .B(ori_ori_n544_), .C(ori_ori_n426_), .Y(ori_ori_n990_));
  NA2        o0962(.A(ori_ori_n990_), .B(ori_ori_n224_), .Y(ori_ori_n991_));
  NA2        o0963(.A(ori_ori_n933_), .B(ori_ori_n490_), .Y(ori_ori_n992_));
  NA4        o0964(.A(ori_ori_n579_), .B(ori_ori_n194_), .C(ori_ori_n206_), .D(ori_ori_n154_), .Y(ori_ori_n993_));
  NA2        o0965(.A(ori_ori_n993_), .B(ori_ori_n992_), .Y(ori_ori_n994_));
  NO2        o0966(.A(ori_ori_n425_), .B(ori_ori_n111_), .Y(ori_ori_n995_));
  NA2        o0967(.A(ori_ori_n995_), .B(ori_ori_n959_), .Y(ori_ori_n996_));
  NO2        o0968(.A(ori_ori_n202_), .B(ori_ori_n199_), .Y(ori_ori_n997_));
  NA2        o0969(.A(n), .B(e), .Y(ori_ori_n998_));
  NO2        o0970(.A(ori_ori_n998_), .B(ori_ori_n137_), .Y(ori_ori_n999_));
  AOI220     o0971(.A0(ori_ori_n999_), .A1(ori_ori_n254_), .B0(ori_ori_n754_), .B1(ori_ori_n997_), .Y(ori_ori_n1000_));
  OAI210     o0972(.A0(ori_ori_n327_), .A1(ori_ori_n281_), .B0(ori_ori_n406_), .Y(ori_ori_n1001_));
  NA3        o0973(.A(ori_ori_n1001_), .B(ori_ori_n1000_), .C(ori_ori_n996_), .Y(ori_ori_n1002_));
  NA2        o0974(.A(ori_ori_n999_), .B(ori_ori_n758_), .Y(ori_ori_n1003_));
  AOI220     o0975(.A0(ori_ori_n846_), .A1(ori_ori_n522_), .B0(ori_ori_n579_), .B1(ori_ori_n227_), .Y(ori_ori_n1004_));
  NO2        o0976(.A(ori_ori_n59_), .B(h), .Y(ori_ori_n1005_));
  NA3        o0977(.A(ori_ori_n1004_), .B(ori_ori_n1003_), .C(ori_ori_n772_), .Y(ori_ori_n1006_));
  NO4        o0978(.A(ori_ori_n1006_), .B(ori_ori_n1002_), .C(ori_ori_n994_), .D(ori_ori_n991_), .Y(ori_ori_n1007_));
  NA2        o0979(.A(ori_ori_n745_), .B(ori_ori_n678_), .Y(ori_ori_n1008_));
  NA4        o0980(.A(ori_ori_n1008_), .B(ori_ori_n1007_), .C(ori_ori_n989_), .D(ori_ori_n969_), .Y(ori01));
  NO2        o0981(.A(ori_ori_n439_), .B(ori_ori_n258_), .Y(ori_ori_n1010_));
  NA2        o0982(.A(ori_ori_n359_), .B(i), .Y(ori_ori_n1011_));
  NA3        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1010_), .C(ori_ori_n906_), .Y(ori_ori_n1012_));
  NA2        o0984(.A(ori_ori_n534_), .B(ori_ori_n81_), .Y(ori_ori_n1013_));
  NA2        o0985(.A(ori_ori_n506_), .B(ori_ori_n252_), .Y(ori_ori_n1014_));
  NA2        o0986(.A(ori_ori_n851_), .B(ori_ori_n1014_), .Y(ori_ori_n1015_));
  NA4        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1013_), .C(ori_ori_n811_), .D(ori_ori_n301_), .Y(ori_ori_n1016_));
  NA2        o0988(.A(ori_ori_n43_), .B(f), .Y(ori_ori_n1017_));
  NA2        o0989(.A(ori_ori_n639_), .B(ori_ori_n88_), .Y(ori_ori_n1018_));
  NO2        o0990(.A(ori_ori_n1018_), .B(ori_ori_n1017_), .Y(ori_ori_n1019_));
  OR2        o0991(.A(ori_ori_n591_), .B(ori_ori_n338_), .Y(ori_ori_n1020_));
  NAi41      o0992(.An(ori_ori_n153_), .B(ori_ori_n1020_), .C(ori_ori_n993_), .D(ori_ori_n796_), .Y(ori_ori_n1021_));
  NO2        o0993(.A(ori_ori_n604_), .B(ori_ori_n471_), .Y(ori_ori_n1022_));
  NA4        o0994(.A(ori_ori_n639_), .B(ori_ori_n88_), .C(ori_ori_n43_), .D(ori_ori_n198_), .Y(ori_ori_n1023_));
  OA220      o0995(.A0(ori_ori_n1023_), .A1(ori_ori_n599_), .B0(ori_ori_n183_), .B1(ori_ori_n181_), .Y(ori_ori_n1024_));
  NA3        o0996(.A(ori_ori_n1024_), .B(ori_ori_n1022_), .C(ori_ori_n127_), .Y(ori_ori_n1025_));
  NO4        o0997(.A(ori_ori_n1025_), .B(ori_ori_n1021_), .C(ori_ori_n1016_), .D(ori_ori_n1012_), .Y(ori_ori_n1026_));
  INV        o0998(.A(ori_ori_n974_), .Y(ori_ori_n1027_));
  NA2        o0999(.A(ori_ori_n1027_), .B(ori_ori_n487_), .Y(ori_ori_n1028_));
  AOI210     o1000(.A0(ori_ori_n192_), .A1(ori_ori_n80_), .B0(ori_ori_n198_), .Y(ori_ori_n1029_));
  OAI210     o1001(.A0(ori_ori_n724_), .A1(ori_ori_n386_), .B0(ori_ori_n1029_), .Y(ori_ori_n1030_));
  AN3        o1002(.A(m), .B(l), .C(k), .Y(ori_ori_n1031_));
  OAI210     o1003(.A0(ori_ori_n329_), .A1(ori_ori_n32_), .B0(ori_ori_n1031_), .Y(ori_ori_n1032_));
  OR2        o1004(.A(ori_ori_n1032_), .B(ori_ori_n300_), .Y(ori_ori_n1033_));
  NA3        o1005(.A(ori_ori_n1033_), .B(ori_ori_n1030_), .C(ori_ori_n1028_), .Y(ori_ori_n1034_));
  NA2        o1006(.A(ori_ori_n538_), .B(ori_ori_n109_), .Y(ori_ori_n1035_));
  INV        o1007(.A(ori_ori_n1035_), .Y(ori_ori_n1036_));
  NA2        o1008(.A(ori_ori_n257_), .B(ori_ori_n183_), .Y(ori_ori_n1037_));
  NA2        o1009(.A(ori_ori_n1037_), .B(ori_ori_n595_), .Y(ori_ori_n1038_));
  OAI210     o1010(.A0(ori_ori_n1019_), .A1(ori_ori_n294_), .B0(ori_ori_n605_), .Y(ori_ori_n1039_));
  NA3        o1011(.A(ori_ori_n1039_), .B(ori_ori_n1038_), .C(ori_ori_n703_), .Y(ori_ori_n1040_));
  NO3        o1012(.A(ori_ori_n1040_), .B(ori_ori_n1036_), .C(ori_ori_n1034_), .Y(ori_ori_n1041_));
  NA2        o1013(.A(ori_ori_n464_), .B(ori_ori_n54_), .Y(ori_ori_n1042_));
  NO2        o1014(.A(ori_ori_n1023_), .B(ori_ori_n870_), .Y(ori_ori_n1043_));
  NO2        o1015(.A(ori_ori_n195_), .B(ori_ori_n103_), .Y(ori_ori_n1044_));
  NO3        o1016(.A(ori_ori_n1044_), .B(ori_ori_n1043_), .C(ori_ori_n972_), .Y(ori_ori_n1045_));
  NA3        o1017(.A(ori_ori_n1045_), .B(ori_ori_n1042_), .C(ori_ori_n677_), .Y(ori_ori_n1046_));
  NO2        o1018(.A(ori_ori_n857_), .B(ori_ori_n216_), .Y(ori_ori_n1047_));
  NO2        o1019(.A(ori_ori_n858_), .B(ori_ori_n508_), .Y(ori_ori_n1048_));
  OAI210     o1020(.A0(ori_ori_n1048_), .A1(ori_ori_n1047_), .B0(ori_ori_n309_), .Y(ori_ori_n1049_));
  NA2        o1021(.A(ori_ori_n517_), .B(ori_ori_n515_), .Y(ori_ori_n1050_));
  NO3        o1022(.A(ori_ori_n70_), .B(ori_ori_n271_), .C(ori_ori_n43_), .Y(ori_ori_n1051_));
  NA2        o1023(.A(ori_ori_n1051_), .B(ori_ori_n505_), .Y(ori_ori_n1052_));
  NA3        o1024(.A(ori_ori_n1052_), .B(ori_ori_n1050_), .C(ori_ori_n600_), .Y(ori_ori_n1053_));
  OR2        o1025(.A(ori_ori_n974_), .B(ori_ori_n971_), .Y(ori_ori_n1054_));
  NA2        o1026(.A(ori_ori_n1051_), .B(ori_ori_n727_), .Y(ori_ori_n1055_));
  NA3        o1027(.A(ori_ori_n1055_), .B(ori_ori_n1054_), .C(ori_ori_n351_), .Y(ori_ori_n1056_));
  NOi41      o1028(.An(ori_ori_n1049_), .B(ori_ori_n1056_), .C(ori_ori_n1053_), .D(ori_ori_n1046_), .Y(ori_ori_n1057_));
  NO2        o1029(.A(ori_ori_n121_), .B(ori_ori_n43_), .Y(ori_ori_n1058_));
  NO2        o1030(.A(ori_ori_n43_), .B(ori_ori_n38_), .Y(ori_ori_n1059_));
  AO220      o1031(.A0(ori_ori_n1059_), .A1(ori_ori_n557_), .B0(ori_ori_n1058_), .B1(ori_ori_n637_), .Y(ori_ori_n1060_));
  NA2        o1032(.A(ori_ori_n1060_), .B(ori_ori_n309_), .Y(ori_ori_n1061_));
  INV        o1033(.A(ori_ori_n125_), .Y(ori_ori_n1062_));
  NO3        o1034(.A(ori_ori_n926_), .B(ori_ori_n164_), .C(ori_ori_n78_), .Y(ori_ori_n1063_));
  AOI220     o1035(.A0(ori_ori_n1063_), .A1(ori_ori_n1062_), .B0(ori_ori_n1051_), .B1(ori_ori_n861_), .Y(ori_ori_n1064_));
  NA2        o1036(.A(ori_ori_n1064_), .B(ori_ori_n1061_), .Y(ori_ori_n1065_));
  NO2        o1037(.A(ori_ori_n550_), .B(ori_ori_n549_), .Y(ori_ori_n1066_));
  NO4        o1038(.A(ori_ori_n926_), .B(ori_ori_n1066_), .C(ori_ori_n162_), .D(ori_ori_n78_), .Y(ori_ori_n1067_));
  NO3        o1039(.A(ori_ori_n1067_), .B(ori_ori_n1065_), .C(ori_ori_n568_), .Y(ori_ori_n1068_));
  NA4        o1040(.A(ori_ori_n1068_), .B(ori_ori_n1057_), .C(ori_ori_n1041_), .D(ori_ori_n1026_), .Y(ori06));
  NO2        o1041(.A(ori_ori_n208_), .B(ori_ori_n95_), .Y(ori_ori_n1070_));
  OAI210     o1042(.A0(ori_ori_n1070_), .A1(ori_ori_n1063_), .B0(ori_ori_n347_), .Y(ori_ori_n1071_));
  NO2        o1043(.A(ori_ori_n541_), .B(ori_ori_n722_), .Y(ori_ori_n1072_));
  OR2        o1044(.A(ori_ori_n1072_), .B(ori_ori_n788_), .Y(ori_ori_n1073_));
  NA3        o1045(.A(ori_ori_n1073_), .B(ori_ori_n1071_), .C(ori_ori_n1049_), .Y(ori_ori_n1074_));
  NO3        o1046(.A(ori_ori_n1074_), .B(ori_ori_n1053_), .C(ori_ori_n240_), .Y(ori_ori_n1075_));
  NO2        o1047(.A(ori_ori_n271_), .B(ori_ori_n43_), .Y(ori_ori_n1076_));
  AOI210     o1048(.A0(ori_ori_n1076_), .A1(ori_ori_n862_), .B0(ori_ori_n1047_), .Y(ori_ori_n1077_));
  AOI210     o1049(.A0(ori_ori_n1076_), .A1(ori_ori_n509_), .B0(ori_ori_n1060_), .Y(ori_ori_n1078_));
  AOI210     o1050(.A0(ori_ori_n1078_), .A1(ori_ori_n1077_), .B0(ori_ori_n306_), .Y(ori_ori_n1079_));
  OAI210     o1051(.A0(ori_ori_n80_), .A1(ori_ori_n38_), .B0(ori_ori_n603_), .Y(ori_ori_n1080_));
  NA2        o1052(.A(ori_ori_n1080_), .B(ori_ori_n572_), .Y(ori_ori_n1081_));
  NO2        o1053(.A(ori_ori_n473_), .B(ori_ori_n159_), .Y(ori_ori_n1082_));
  NO2        o1054(.A(ori_ori_n545_), .B(ori_ori_n938_), .Y(ori_ori_n1083_));
  OAI210     o1055(.A0(ori_ori_n420_), .A1(ori_ori_n231_), .B0(ori_ori_n806_), .Y(ori_ori_n1084_));
  NO3        o1056(.A(ori_ori_n1084_), .B(ori_ori_n1083_), .C(ori_ori_n1082_), .Y(ori_ori_n1085_));
  NA2        o1057(.A(ori_ori_n1085_), .B(ori_ori_n1081_), .Y(ori_ori_n1086_));
  AN2        o1058(.A(ori_ori_n846_), .B(ori_ori_n575_), .Y(ori_ori_n1087_));
  NO3        o1059(.A(ori_ori_n1087_), .B(ori_ori_n1086_), .C(ori_ori_n1079_), .Y(ori_ori_n1088_));
  NO2        o1060(.A(ori_ori_n661_), .B(ori_ori_n45_), .Y(ori_ori_n1089_));
  NA2        o1061(.A(ori_ori_n332_), .B(ori_ori_n1089_), .Y(ori_ori_n1090_));
  NO3        o1062(.A(ori_ori_n226_), .B(ori_ori_n95_), .C(ori_ori_n260_), .Y(ori_ori_n1091_));
  OAI220     o1063(.A0(ori_ori_n629_), .A1(ori_ori_n231_), .B0(ori_ori_n470_), .B1(ori_ori_n473_), .Y(ori_ori_n1092_));
  INV        o1064(.A(k), .Y(ori_ori_n1093_));
  NO3        o1065(.A(ori_ori_n1093_), .B(ori_ori_n540_), .C(j), .Y(ori_ori_n1094_));
  NO3        o1066(.A(ori_ori_n1092_), .B(ori_ori_n1091_), .C(ori_ori_n941_), .Y(ori_ori_n1095_));
  NA3        o1067(.A(ori_ori_n711_), .B(ori_ori_n710_), .C(ori_ori_n395_), .Y(ori_ori_n1096_));
  NAi31      o1068(.An(ori_ori_n670_), .B(ori_ori_n1096_), .C(ori_ori_n191_), .Y(ori_ori_n1097_));
  NA4        o1069(.A(ori_ori_n1097_), .B(ori_ori_n1095_), .C(ori_ori_n1090_), .D(ori_ori_n1004_), .Y(ori_ori_n1098_));
  NA2        o1070(.A(ori_ori_n517_), .B(ori_ori_n406_), .Y(ori_ori_n1099_));
  NA2        o1071(.A(ori_ori_n1094_), .B(ori_ori_n707_), .Y(ori_ori_n1100_));
  NA2        o1072(.A(ori_ori_n1100_), .B(ori_ori_n1099_), .Y(ori_ori_n1101_));
  AN2        o1073(.A(ori_ori_n821_), .B(ori_ori_n820_), .Y(ori_ori_n1102_));
  NO3        o1074(.A(ori_ori_n1102_), .B(ori_ori_n460_), .C(ori_ori_n442_), .Y(ori_ori_n1103_));
  NA2        o1075(.A(ori_ori_n1103_), .B(ori_ori_n1055_), .Y(ori_ori_n1104_));
  NAi21      o1076(.An(j), .B(i), .Y(ori_ori_n1105_));
  NO4        o1077(.A(ori_ori_n1066_), .B(ori_ori_n1105_), .C(ori_ori_n400_), .D(ori_ori_n218_), .Y(ori_ori_n1106_));
  NO4        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1104_), .C(ori_ori_n1101_), .D(ori_ori_n1098_), .Y(ori_ori_n1107_));
  NA4        o1079(.A(ori_ori_n1107_), .B(ori_ori_n1088_), .C(ori_ori_n1075_), .D(ori_ori_n1068_), .Y(ori07));
  NAi32      o1080(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1109_));
  NO3        o1081(.A(ori_ori_n1109_), .B(g), .C(f), .Y(ori_ori_n1110_));
  NAi21      o1082(.An(f), .B(c), .Y(ori_ori_n1111_));
  NOi31      o1083(.An(n), .B(m), .C(b), .Y(ori_ori_n1112_));
  NOi41      o1084(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1113_));
  NO2        o1085(.A(ori_ori_n921_), .B(ori_ori_n276_), .Y(ori_ori_n1114_));
  NA2        o1086(.A(ori_ori_n494_), .B(ori_ori_n71_), .Y(ori_ori_n1115_));
  NA2        o1087(.A(ori_ori_n1005_), .B(ori_ori_n266_), .Y(ori_ori_n1116_));
  NA2        o1088(.A(ori_ori_n1116_), .B(ori_ori_n1115_), .Y(ori_ori_n1117_));
  NO2        o1089(.A(ori_ori_n1117_), .B(ori_ori_n1110_), .Y(ori_ori_n1118_));
  NO3        o1090(.A(e), .B(d), .C(c), .Y(ori_ori_n1119_));
  NO2        o1091(.A(ori_ori_n122_), .B(ori_ori_n199_), .Y(ori_ori_n1120_));
  NA2        o1092(.A(ori_ori_n1120_), .B(ori_ori_n1119_), .Y(ori_ori_n1121_));
  INV        o1093(.A(ori_ori_n1121_), .Y(ori_ori_n1122_));
  NA3        o1094(.A(ori_ori_n626_), .B(ori_ori_n612_), .C(ori_ori_n104_), .Y(ori_ori_n1123_));
  NO2        o1095(.A(ori_ori_n1123_), .B(ori_ori_n43_), .Y(ori_ori_n1124_));
  NO2        o1096(.A(l), .B(k), .Y(ori_ori_n1125_));
  NO3        o1097(.A(ori_ori_n400_), .B(d), .C(c), .Y(ori_ori_n1126_));
  NO2        o1098(.A(ori_ori_n1124_), .B(ori_ori_n1122_), .Y(ori_ori_n1127_));
  NO2        o1099(.A(g), .B(c), .Y(ori_ori_n1128_));
  NO2        o1100(.A(ori_ori_n411_), .B(a), .Y(ori_ori_n1129_));
  NA2        o1101(.A(ori_ori_n1129_), .B(ori_ori_n105_), .Y(ori_ori_n1130_));
  NA2        o1102(.A(ori_ori_n128_), .B(ori_ori_n206_), .Y(ori_ori_n1131_));
  NO2        o1103(.A(ori_ori_n1131_), .B(ori_ori_n1219_), .Y(ori_ori_n1132_));
  NO2        o1104(.A(ori_ori_n676_), .B(ori_ori_n175_), .Y(ori_ori_n1133_));
  NOi31      o1105(.An(m), .B(n), .C(b), .Y(ori_ori_n1134_));
  NOi31      o1106(.An(f), .B(d), .C(c), .Y(ori_ori_n1135_));
  NA2        o1107(.A(ori_ori_n1135_), .B(ori_ori_n1134_), .Y(ori_ori_n1136_));
  INV        o1108(.A(ori_ori_n1136_), .Y(ori_ori_n1137_));
  NO3        o1109(.A(ori_ori_n1137_), .B(ori_ori_n1133_), .C(ori_ori_n1132_), .Y(ori_ori_n1138_));
  NA2        o1110(.A(ori_ori_n924_), .B(ori_ori_n427_), .Y(ori_ori_n1139_));
  NO2        o1111(.A(ori_ori_n1139_), .B(ori_ori_n400_), .Y(ori_ori_n1140_));
  NO3        o1112(.A(ori_ori_n39_), .B(i), .C(h), .Y(ori_ori_n1141_));
  NO2        o1113(.A(ori_ori_n920_), .B(ori_ori_n1140_), .Y(ori_ori_n1142_));
  AN3        o1114(.A(ori_ori_n1142_), .B(ori_ori_n1138_), .C(ori_ori_n1130_), .Y(ori_ori_n1143_));
  NA2        o1115(.A(ori_ori_n1112_), .B(ori_ori_n344_), .Y(ori_ori_n1144_));
  INV        o1116(.A(ori_ori_n1144_), .Y(ori_ori_n1145_));
  INV        o1117(.A(ori_ori_n927_), .Y(ori_ori_n1146_));
  NAi21      o1118(.An(ori_ori_n1145_), .B(ori_ori_n1146_), .Y(ori_ori_n1147_));
  NO4        o1119(.A(ori_ori_n122_), .B(g), .C(f), .D(e), .Y(ori_ori_n1148_));
  NA2        o1120(.A(ori_ori_n1113_), .B(ori_ori_n1125_), .Y(ori_ori_n1149_));
  INV        o1121(.A(ori_ori_n1149_), .Y(ori_ori_n1150_));
  OR3        o1122(.A(ori_ori_n493_), .B(ori_ori_n492_), .C(ori_ori_n104_), .Y(ori_ori_n1151_));
  NA2        o1123(.A(ori_ori_n937_), .B(ori_ori_n369_), .Y(ori_ori_n1152_));
  NO2        o1124(.A(ori_ori_n1152_), .B(ori_ori_n394_), .Y(ori_ori_n1153_));
  AO210      o1125(.A0(ori_ori_n1153_), .A1(ori_ori_n107_), .B0(ori_ori_n1150_), .Y(ori_ori_n1154_));
  NO2        o1126(.A(ori_ori_n1154_), .B(ori_ori_n1147_), .Y(ori_ori_n1155_));
  NA4        o1127(.A(ori_ori_n1155_), .B(ori_ori_n1143_), .C(ori_ori_n1127_), .D(ori_ori_n1118_), .Y(ori_ori_n1156_));
  NO2        o1128(.A(ori_ori_n946_), .B(ori_ori_n102_), .Y(ori_ori_n1157_));
  NO2        o1129(.A(ori_ori_n356_), .B(j), .Y(ori_ori_n1158_));
  NA2        o1130(.A(ori_ori_n1141_), .B(ori_ori_n937_), .Y(ori_ori_n1159_));
  NA2        o1131(.A(ori_ori_n923_), .B(ori_ori_n141_), .Y(ori_ori_n1160_));
  NA2        o1132(.A(ori_ori_n1160_), .B(ori_ori_n1159_), .Y(ori_ori_n1161_));
  NA2        o1133(.A(ori_ori_n1158_), .B(ori_ori_n150_), .Y(ori_ori_n1162_));
  INV        o1134(.A(ori_ori_n1162_), .Y(ori_ori_n1163_));
  NO2        o1135(.A(ori_ori_n1163_), .B(ori_ori_n1161_), .Y(ori_ori_n1164_));
  INV        o1136(.A(ori_ori_n47_), .Y(ori_ori_n1165_));
  NA2        o1137(.A(ori_ori_n1165_), .B(ori_ori_n976_), .Y(ori_ori_n1166_));
  INV        o1138(.A(ori_ori_n1166_), .Y(ori_ori_n1167_));
  NO2        o1139(.A(ori_ori_n596_), .B(ori_ori_n164_), .Y(ori_ori_n1168_));
  NO2        o1140(.A(ori_ori_n1168_), .B(ori_ori_n1167_), .Y(ori_ori_n1169_));
  NA2        o1141(.A(ori_ori_n1157_), .B(f), .Y(ori_ori_n1170_));
  INV        o1142(.A(ori_ori_n167_), .Y(ori_ori_n1171_));
  NO2        o1143(.A(ori_ori_n1218_), .B(ori_ori_n1170_), .Y(ori_ori_n1172_));
  NO2        o1144(.A(ori_ori_n1105_), .B(ori_ori_n162_), .Y(ori_ori_n1173_));
  NOi21      o1145(.An(d), .B(f), .Y(ori_ori_n1174_));
  NA2        o1146(.A(h), .B(ori_ori_n1173_), .Y(ori_ori_n1175_));
  INV        o1147(.A(ori_ori_n1175_), .Y(ori_ori_n1176_));
  NO2        o1148(.A(ori_ori_n1176_), .B(ori_ori_n1172_), .Y(ori_ori_n1177_));
  NA3        o1149(.A(ori_ori_n1177_), .B(ori_ori_n1169_), .C(ori_ori_n1164_), .Y(ori_ori_n1178_));
  NA2        o1150(.A(h), .B(ori_ori_n1114_), .Y(ori_ori_n1179_));
  OAI210     o1151(.A0(ori_ori_n1148_), .A1(ori_ori_n1112_), .B0(ori_ori_n785_), .Y(ori_ori_n1180_));
  NO2        o1152(.A(ori_ori_n917_), .B(ori_ori_n122_), .Y(ori_ori_n1181_));
  NA2        o1153(.A(ori_ori_n1181_), .B(ori_ori_n556_), .Y(ori_ori_n1182_));
  NA3        o1154(.A(ori_ori_n1182_), .B(ori_ori_n1180_), .C(ori_ori_n1179_), .Y(ori_ori_n1183_));
  NA2        o1155(.A(ori_ori_n1128_), .B(ori_ori_n1174_), .Y(ori_ori_n1184_));
  NO2        o1156(.A(ori_ori_n1184_), .B(m), .Y(ori_ori_n1185_));
  NO2        o1157(.A(ori_ori_n142_), .B(ori_ori_n169_), .Y(ori_ori_n1186_));
  OAI210     o1158(.A0(ori_ori_n1186_), .A1(ori_ori_n102_), .B0(ori_ori_n1134_), .Y(ori_ori_n1187_));
  INV        o1159(.A(ori_ori_n1187_), .Y(ori_ori_n1188_));
  NO3        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1185_), .C(ori_ori_n1183_), .Y(ori_ori_n1189_));
  NO2        o1161(.A(ori_ori_n1111_), .B(e), .Y(ori_ori_n1190_));
  NA2        o1162(.A(ori_ori_n1190_), .B(ori_ori_n367_), .Y(ori_ori_n1191_));
  BUFFER     o1163(.A(ori_ori_n122_), .Y(ori_ori_n1192_));
  NO2        o1164(.A(ori_ori_n1192_), .B(ori_ori_n1191_), .Y(ori_ori_n1193_));
  NO2        o1165(.A(ori_ori_n1151_), .B(ori_ori_n323_), .Y(ori_ori_n1194_));
  NO2        o1166(.A(ori_ori_n1194_), .B(ori_ori_n1193_), .Y(ori_ori_n1195_));
  INV        o1167(.A(ori_ori_n1126_), .Y(ori_ori_n1196_));
  INV        o1168(.A(ori_ori_n944_), .Y(ori_ori_n1197_));
  OAI210     o1169(.A0(ori_ori_n1197_), .A1(ori_ori_n60_), .B0(ori_ori_n1196_), .Y(ori_ori_n1198_));
  OR2        o1170(.A(h), .B(ori_ori_n492_), .Y(ori_ori_n1199_));
  NO2        o1171(.A(ori_ori_n1199_), .B(ori_ori_n162_), .Y(ori_ori_n1200_));
  NA2        o1172(.A(ori_ori_n928_), .B(ori_ori_n206_), .Y(ori_ori_n1201_));
  NO2        o1173(.A(ori_ori_n47_), .B(l), .Y(ori_ori_n1202_));
  INV        o1174(.A(ori_ori_n444_), .Y(ori_ori_n1203_));
  NA2        o1175(.A(ori_ori_n1203_), .B(ori_ori_n1202_), .Y(ori_ori_n1204_));
  NA2        o1176(.A(ori_ori_n1204_), .B(ori_ori_n1201_), .Y(ori_ori_n1205_));
  NO3        o1177(.A(ori_ori_n1205_), .B(ori_ori_n1200_), .C(ori_ori_n1198_), .Y(ori_ori_n1206_));
  NA3        o1178(.A(ori_ori_n1206_), .B(ori_ori_n1195_), .C(ori_ori_n1189_), .Y(ori_ori_n1207_));
  NA3        o1179(.A(ori_ori_n850_), .B(ori_ori_n128_), .C(ori_ori_n44_), .Y(ori_ori_n1208_));
  INV        o1180(.A(ori_ori_n1190_), .Y(ori_ori_n1209_));
  NO2        o1181(.A(ori_ori_n1209_), .B(ori_ori_n1171_), .Y(ori_ori_n1210_));
  INV        o1182(.A(ori_ori_n1210_), .Y(ori_ori_n1211_));
  NO2        o1183(.A(ori_ori_n1152_), .B(d), .Y(ori_ori_n1212_));
  INV        o1184(.A(ori_ori_n1212_), .Y(ori_ori_n1213_));
  NA3        o1185(.A(ori_ori_n1213_), .B(ori_ori_n1211_), .C(ori_ori_n1208_), .Y(ori_ori_n1214_));
  OR4        o1186(.A(ori_ori_n1214_), .B(ori_ori_n1207_), .C(ori_ori_n1178_), .D(ori_ori_n1156_), .Y(ori04));
  INV        o1187(.A(ori_ori_n105_), .Y(ori_ori_n1218_));
  INV        o1188(.A(h), .Y(ori_ori_n1219_));
  ZERO       o1189(.Y(ori02));
  ZERO       o1190(.Y(ori03));
  ZERO       o1191(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(g), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  NO2        m0034(.A(mai_mai_n61_), .B(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi21      m0043(.An(e), .B(h), .Y(mai_mai_n72_));
  NAi41      m0044(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n74_));
  INV        m0046(.A(m), .Y(mai_mai_n75_));
  NOi21      m0047(.An(k), .B(l), .Y(mai_mai_n76_));
  AN4        m0048(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n77_));
  NOi31      m0049(.An(h), .B(g), .C(f), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n77_), .Y(mai_mai_n79_));
  NAi32      m0051(.An(m), .Bn(k), .C(j), .Y(mai_mai_n80_));
  NOi32      m0052(.An(h), .Bn(g), .C(f), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n82_));
  INV        m0054(.A(n), .Y(mai_mai_n83_));
  NOi32      m0055(.An(e), .Bn(b), .C(d), .Y(mai_mai_n84_));
  NA2        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  INV        m0057(.A(j), .Y(mai_mai_n86_));
  AN3        m0058(.A(m), .B(k), .C(i), .Y(mai_mai_n87_));
  NA3        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(g), .Y(mai_mai_n88_));
  NAi32      m0060(.An(g), .Bn(f), .C(h), .Y(mai_mai_n89_));
  NAi31      m0061(.An(j), .B(m), .C(l), .Y(mai_mai_n90_));
  NA2        m0062(.A(m), .B(l), .Y(mai_mai_n91_));
  NAi31      m0063(.An(k), .B(j), .C(g), .Y(mai_mai_n92_));
  NO3        m0064(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(f), .Y(mai_mai_n93_));
  AN2        m0065(.A(j), .B(g), .Y(mai_mai_n94_));
  NOi32      m0066(.An(m), .Bn(l), .C(i), .Y(mai_mai_n95_));
  NOi21      m0067(.An(g), .B(i), .Y(mai_mai_n96_));
  NOi32      m0068(.An(m), .Bn(j), .C(k), .Y(mai_mai_n97_));
  AOI220     m0069(.A0(mai_mai_n97_), .A1(mai_mai_n96_), .B0(mai_mai_n95_), .B1(mai_mai_n94_), .Y(mai_mai_n98_));
  NO2        m0070(.A(mai_mai_n98_), .B(f), .Y(mai_mai_n99_));
  NAi41      m0071(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n100_));
  AN2        m0072(.A(e), .B(b), .Y(mai_mai_n101_));
  NOi31      m0073(.An(c), .B(h), .C(f), .Y(mai_mai_n102_));
  NA2        m0074(.A(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  NO3        m0075(.A(mai_mai_n103_), .B(mai_mai_n100_), .C(g), .Y(mai_mai_n104_));
  NOi21      m0076(.An(g), .B(f), .Y(mai_mai_n105_));
  NOi21      m0077(.An(i), .B(h), .Y(mai_mai_n106_));
  NA3        m0078(.A(mai_mai_n106_), .B(mai_mai_n105_), .C(mai_mai_n36_), .Y(mai_mai_n107_));
  INV        m0079(.A(a), .Y(mai_mai_n108_));
  NA2        m0080(.A(mai_mai_n101_), .B(mai_mai_n108_), .Y(mai_mai_n109_));
  INV        m0081(.A(l), .Y(mai_mai_n110_));
  NOi21      m0082(.An(m), .B(n), .Y(mai_mai_n111_));
  AN2        m0083(.A(k), .B(h), .Y(mai_mai_n112_));
  NO2        m0084(.A(mai_mai_n107_), .B(mai_mai_n85_), .Y(mai_mai_n113_));
  INV        m0085(.A(b), .Y(mai_mai_n114_));
  NA2        m0086(.A(l), .B(j), .Y(mai_mai_n115_));
  AN2        m0087(.A(k), .B(i), .Y(mai_mai_n116_));
  NA2        m0088(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NA2        m0089(.A(g), .B(e), .Y(mai_mai_n118_));
  NOi32      m0090(.An(c), .Bn(a), .C(d), .Y(mai_mai_n119_));
  NA2        m0091(.A(mai_mai_n119_), .B(mai_mai_n111_), .Y(mai_mai_n120_));
  NO4        m0092(.A(mai_mai_n120_), .B(mai_mai_n118_), .C(mai_mai_n117_), .D(mai_mai_n114_), .Y(mai_mai_n121_));
  NO3        m0093(.A(mai_mai_n121_), .B(mai_mai_n113_), .C(mai_mai_n104_), .Y(mai_mai_n122_));
  OAI210     m0094(.A0(mai_mai_n98_), .A1(mai_mai_n85_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NOi31      m0095(.An(k), .B(m), .C(j), .Y(mai_mai_n124_));
  NOi31      m0096(.An(k), .B(m), .C(i), .Y(mai_mai_n125_));
  NA3        m0097(.A(mai_mai_n125_), .B(mai_mai_n81_), .C(mai_mai_n77_), .Y(mai_mai_n126_));
  INV        m0098(.A(mai_mai_n126_), .Y(mai_mai_n127_));
  NOi32      m0099(.An(f), .Bn(b), .C(e), .Y(mai_mai_n128_));
  NAi21      m0100(.An(g), .B(h), .Y(mai_mai_n129_));
  NAi21      m0101(.An(m), .B(n), .Y(mai_mai_n130_));
  NAi21      m0102(.An(j), .B(k), .Y(mai_mai_n131_));
  NAi41      m0103(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n132_));
  NAi31      m0104(.An(j), .B(k), .C(h), .Y(mai_mai_n133_));
  NO3        m0105(.A(mai_mai_n133_), .B(mai_mai_n132_), .C(mai_mai_n130_), .Y(mai_mai_n134_));
  INV        m0106(.A(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m0107(.A(k), .B(j), .Y(mai_mai_n136_));
  AN2        m0108(.A(k), .B(j), .Y(mai_mai_n137_));
  NAi21      m0109(.An(c), .B(b), .Y(mai_mai_n138_));
  NA2        m0110(.A(f), .B(d), .Y(mai_mai_n139_));
  NAi31      m0111(.An(f), .B(e), .C(b), .Y(mai_mai_n140_));
  NA2        m0112(.A(d), .B(b), .Y(mai_mai_n141_));
  NAi21      m0113(.An(e), .B(f), .Y(mai_mai_n142_));
  NO2        m0114(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  NA2        m0115(.A(b), .B(a), .Y(mai_mai_n144_));
  NAi21      m0116(.An(e), .B(g), .Y(mai_mai_n145_));
  NAi21      m0117(.An(c), .B(d), .Y(mai_mai_n146_));
  NAi31      m0118(.An(l), .B(k), .C(h), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n130_), .B(mai_mai_n147_), .Y(mai_mai_n148_));
  NAi21      m0120(.An(mai_mai_n127_), .B(mai_mai_n135_), .Y(mai_mai_n149_));
  NAi31      m0121(.An(e), .B(f), .C(b), .Y(mai_mai_n150_));
  NOi21      m0122(.An(g), .B(d), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  NOi21      m0124(.An(h), .B(i), .Y(mai_mai_n153_));
  NOi21      m0125(.An(k), .B(m), .Y(mai_mai_n154_));
  NA3        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .C(n), .Y(mai_mai_n155_));
  NOi21      m0127(.An(mai_mai_n152_), .B(mai_mai_n155_), .Y(mai_mai_n156_));
  NOi21      m0128(.An(h), .B(g), .Y(mai_mai_n157_));
  NO2        m0129(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NAi31      m0131(.An(l), .B(j), .C(h), .Y(mai_mai_n160_));
  NO2        m0132(.A(mai_mai_n160_), .B(mai_mai_n49_), .Y(mai_mai_n161_));
  NA2        m0133(.A(mai_mai_n161_), .B(mai_mai_n67_), .Y(mai_mai_n162_));
  NOi32      m0134(.An(n), .Bn(k), .C(m), .Y(mai_mai_n163_));
  NA2        m0135(.A(l), .B(i), .Y(mai_mai_n164_));
  NA2        m0136(.A(mai_mai_n164_), .B(mai_mai_n163_), .Y(mai_mai_n165_));
  OAI210     m0137(.A0(mai_mai_n165_), .A1(mai_mai_n159_), .B0(mai_mai_n162_), .Y(mai_mai_n166_));
  NAi31      m0138(.An(d), .B(f), .C(c), .Y(mai_mai_n167_));
  NAi31      m0139(.An(e), .B(f), .C(c), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  NA2        m0141(.A(j), .B(h), .Y(mai_mai_n170_));
  OR3        m0142(.A(n), .B(m), .C(k), .Y(mai_mai_n171_));
  NO2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NAi32      m0144(.An(m), .Bn(k), .C(n), .Y(mai_mai_n173_));
  NO2        m0145(.A(mai_mai_n173_), .B(mai_mai_n170_), .Y(mai_mai_n174_));
  AOI220     m0146(.A0(mai_mai_n174_), .A1(mai_mai_n152_), .B0(mai_mai_n172_), .B1(mai_mai_n169_), .Y(mai_mai_n175_));
  NO2        m0147(.A(n), .B(m), .Y(mai_mai_n176_));
  NA2        m0148(.A(mai_mai_n176_), .B(mai_mai_n50_), .Y(mai_mai_n177_));
  NAi21      m0149(.An(f), .B(e), .Y(mai_mai_n178_));
  NA2        m0150(.A(d), .B(c), .Y(mai_mai_n179_));
  NAi21      m0151(.An(d), .B(c), .Y(mai_mai_n180_));
  NAi31      m0152(.An(m), .B(n), .C(b), .Y(mai_mai_n181_));
  NA2        m0153(.A(k), .B(i), .Y(mai_mai_n182_));
  NAi21      m0154(.An(h), .B(f), .Y(mai_mai_n183_));
  NO2        m0155(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  NO2        m0156(.A(mai_mai_n181_), .B(mai_mai_n146_), .Y(mai_mai_n185_));
  NA2        m0157(.A(mai_mai_n185_), .B(mai_mai_n184_), .Y(mai_mai_n186_));
  NOi32      m0158(.An(f), .Bn(c), .C(d), .Y(mai_mai_n187_));
  NOi32      m0159(.An(f), .Bn(c), .C(e), .Y(mai_mai_n188_));
  NO2        m0160(.A(mai_mai_n188_), .B(mai_mai_n187_), .Y(mai_mai_n189_));
  NO3        m0161(.A(n), .B(m), .C(j), .Y(mai_mai_n190_));
  NA2        m0162(.A(mai_mai_n190_), .B(mai_mai_n112_), .Y(mai_mai_n191_));
  AO210      m0163(.A0(mai_mai_n191_), .A1(mai_mai_n177_), .B0(mai_mai_n189_), .Y(mai_mai_n192_));
  NA3        m0164(.A(mai_mai_n192_), .B(mai_mai_n186_), .C(mai_mai_n175_), .Y(mai_mai_n193_));
  OR4        m0165(.A(mai_mai_n193_), .B(mai_mai_n166_), .C(mai_mai_n156_), .D(mai_mai_n149_), .Y(mai_mai_n194_));
  NO4        m0166(.A(mai_mai_n194_), .B(mai_mai_n123_), .C(mai_mai_n82_), .D(mai_mai_n55_), .Y(mai_mai_n195_));
  NA3        m0167(.A(m), .B(mai_mai_n110_), .C(j), .Y(mai_mai_n196_));
  NAi31      m0168(.An(n), .B(h), .C(g), .Y(mai_mai_n197_));
  NO2        m0169(.A(mai_mai_n197_), .B(mai_mai_n196_), .Y(mai_mai_n198_));
  NOi32      m0170(.An(m), .Bn(k), .C(l), .Y(mai_mai_n199_));
  NA3        m0171(.A(mai_mai_n199_), .B(mai_mai_n86_), .C(g), .Y(mai_mai_n200_));
  NO2        m0172(.A(mai_mai_n200_), .B(n), .Y(mai_mai_n201_));
  NOi21      m0173(.An(k), .B(j), .Y(mai_mai_n202_));
  NA4        m0174(.A(mai_mai_n202_), .B(mai_mai_n111_), .C(i), .D(g), .Y(mai_mai_n203_));
  AN2        m0175(.A(i), .B(g), .Y(mai_mai_n204_));
  NA3        m0176(.A(mai_mai_n76_), .B(mai_mai_n204_), .C(mai_mai_n111_), .Y(mai_mai_n205_));
  NA2        m0177(.A(mai_mai_n205_), .B(mai_mai_n203_), .Y(mai_mai_n206_));
  NO3        m0178(.A(mai_mai_n206_), .B(mai_mai_n201_), .C(mai_mai_n198_), .Y(mai_mai_n207_));
  NAi41      m0179(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n208_));
  INV        m0180(.A(mai_mai_n208_), .Y(mai_mai_n209_));
  INV        m0181(.A(f), .Y(mai_mai_n210_));
  INV        m0182(.A(g), .Y(mai_mai_n211_));
  NOi31      m0183(.An(i), .B(j), .C(h), .Y(mai_mai_n212_));
  NOi21      m0184(.An(l), .B(m), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n213_), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  NO2        m0186(.A(mai_mai_n207_), .B(mai_mai_n32_), .Y(mai_mai_n215_));
  NOi21      m0187(.An(n), .B(m), .Y(mai_mai_n216_));
  NOi32      m0188(.An(l), .Bn(i), .C(j), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  OA220      m0190(.A0(mai_mai_n218_), .A1(mai_mai_n103_), .B0(mai_mai_n80_), .B1(mai_mai_n79_), .Y(mai_mai_n219_));
  NAi21      m0191(.An(j), .B(h), .Y(mai_mai_n220_));
  XN2        m0192(.A(i), .B(h), .Y(mai_mai_n221_));
  NA2        m0193(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  NOi31      m0194(.An(k), .B(n), .C(m), .Y(mai_mai_n223_));
  NOi31      m0195(.An(mai_mai_n223_), .B(mai_mai_n179_), .C(mai_mai_n178_), .Y(mai_mai_n224_));
  NA2        m0196(.A(mai_mai_n224_), .B(mai_mai_n222_), .Y(mai_mai_n225_));
  NAi31      m0197(.An(f), .B(e), .C(c), .Y(mai_mai_n226_));
  NO4        m0198(.A(mai_mai_n226_), .B(mai_mai_n171_), .C(mai_mai_n170_), .D(mai_mai_n59_), .Y(mai_mai_n227_));
  NA4        m0199(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n228_));
  NAi32      m0200(.An(m), .Bn(i), .C(k), .Y(mai_mai_n229_));
  NO3        m0201(.A(mai_mai_n229_), .B(mai_mai_n89_), .C(mai_mai_n228_), .Y(mai_mai_n230_));
  INV        m0202(.A(k), .Y(mai_mai_n231_));
  NO2        m0203(.A(mai_mai_n230_), .B(mai_mai_n227_), .Y(mai_mai_n232_));
  NAi21      m0204(.An(n), .B(a), .Y(mai_mai_n233_));
  NO2        m0205(.A(mai_mai_n233_), .B(mai_mai_n141_), .Y(mai_mai_n234_));
  NAi41      m0206(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n235_));
  NO2        m0207(.A(mai_mai_n235_), .B(e), .Y(mai_mai_n236_));
  NO3        m0208(.A(mai_mai_n142_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n237_));
  OAI210     m0209(.A0(mai_mai_n237_), .A1(mai_mai_n236_), .B0(mai_mai_n234_), .Y(mai_mai_n238_));
  AN4        m0210(.A(mai_mai_n238_), .B(mai_mai_n232_), .C(mai_mai_n225_), .D(mai_mai_n219_), .Y(mai_mai_n239_));
  OR2        m0211(.A(h), .B(g), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n240_), .B(mai_mai_n100_), .Y(mai_mai_n241_));
  NA2        m0213(.A(mai_mai_n241_), .B(mai_mai_n128_), .Y(mai_mai_n242_));
  NAi31      m0214(.An(e), .B(d), .C(b), .Y(mai_mai_n243_));
  NA2        m0215(.A(mai_mai_n154_), .B(mai_mai_n106_), .Y(mai_mai_n244_));
  NO2        m0216(.A(n), .B(a), .Y(mai_mai_n245_));
  NAi31      m0217(.An(mai_mai_n235_), .B(mai_mai_n245_), .C(mai_mai_n101_), .Y(mai_mai_n246_));
  NAi21      m0218(.An(h), .B(i), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n176_), .B(k), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n248_), .B(mai_mai_n247_), .Y(mai_mai_n249_));
  NA2        m0221(.A(mai_mai_n249_), .B(mai_mai_n187_), .Y(mai_mai_n250_));
  NA3        m0222(.A(mai_mai_n250_), .B(mai_mai_n246_), .C(mai_mai_n242_), .Y(mai_mai_n251_));
  NOi21      m0223(.An(g), .B(e), .Y(mai_mai_n252_));
  NO2        m0224(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n253_));
  NA2        m0225(.A(mai_mai_n253_), .B(mai_mai_n252_), .Y(mai_mai_n254_));
  NOi32      m0226(.An(l), .Bn(j), .C(i), .Y(mai_mai_n255_));
  AOI210     m0227(.A0(mai_mai_n76_), .A1(mai_mai_n86_), .B0(mai_mai_n255_), .Y(mai_mai_n256_));
  NO2        m0228(.A(mai_mai_n247_), .B(mai_mai_n44_), .Y(mai_mai_n257_));
  NAi21      m0229(.An(f), .B(g), .Y(mai_mai_n258_));
  NO2        m0230(.A(mai_mai_n258_), .B(mai_mai_n65_), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n69_), .B(mai_mai_n115_), .Y(mai_mai_n260_));
  AOI220     m0232(.A0(mai_mai_n260_), .A1(mai_mai_n259_), .B0(mai_mai_n257_), .B1(mai_mai_n67_), .Y(mai_mai_n261_));
  OAI210     m0233(.A0(mai_mai_n256_), .A1(mai_mai_n254_), .B0(mai_mai_n261_), .Y(mai_mai_n262_));
  NO3        m0234(.A(mai_mai_n131_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n263_));
  NOi41      m0235(.An(mai_mai_n239_), .B(mai_mai_n262_), .C(mai_mai_n251_), .D(mai_mai_n215_), .Y(mai_mai_n264_));
  NO4        m0236(.A(mai_mai_n198_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n265_));
  NO2        m0237(.A(mai_mai_n265_), .B(mai_mai_n109_), .Y(mai_mai_n266_));
  NA3        m0238(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n267_));
  NAi21      m0239(.An(h), .B(g), .Y(mai_mai_n268_));
  OR4        m0240(.A(mai_mai_n268_), .B(mai_mai_n267_), .C(mai_mai_n218_), .D(e), .Y(mai_mai_n269_));
  NAi31      m0241(.An(g), .B(k), .C(h), .Y(mai_mai_n270_));
  NO3        m0242(.A(mai_mai_n130_), .B(mai_mai_n270_), .C(l), .Y(mai_mai_n271_));
  NAi31      m0243(.An(e), .B(d), .C(a), .Y(mai_mai_n272_));
  NA2        m0244(.A(mai_mai_n271_), .B(mai_mai_n128_), .Y(mai_mai_n273_));
  NA2        m0245(.A(mai_mai_n273_), .B(mai_mai_n269_), .Y(mai_mai_n274_));
  NA3        m0246(.A(mai_mai_n154_), .B(mai_mai_n153_), .C(mai_mai_n83_), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n275_), .B(mai_mai_n189_), .Y(mai_mai_n276_));
  INV        m0248(.A(mai_mai_n276_), .Y(mai_mai_n277_));
  NA3        m0249(.A(e), .B(c), .C(b), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n60_), .B(mai_mai_n278_), .Y(mai_mai_n279_));
  NAi32      m0251(.An(k), .Bn(i), .C(j), .Y(mai_mai_n280_));
  NAi31      m0252(.An(h), .B(l), .C(i), .Y(mai_mai_n281_));
  NA3        m0253(.A(mai_mai_n281_), .B(mai_mai_n280_), .C(mai_mai_n160_), .Y(mai_mai_n282_));
  NOi21      m0254(.An(mai_mai_n282_), .B(mai_mai_n49_), .Y(mai_mai_n283_));
  OAI210     m0255(.A0(mai_mai_n259_), .A1(mai_mai_n279_), .B0(mai_mai_n283_), .Y(mai_mai_n284_));
  NAi21      m0256(.An(l), .B(k), .Y(mai_mai_n285_));
  NO2        m0257(.A(mai_mai_n285_), .B(mai_mai_n49_), .Y(mai_mai_n286_));
  NOi21      m0258(.An(l), .B(j), .Y(mai_mai_n287_));
  NA2        m0259(.A(mai_mai_n157_), .B(mai_mai_n287_), .Y(mai_mai_n288_));
  NA3        m0260(.A(mai_mai_n116_), .B(mai_mai_n115_), .C(g), .Y(mai_mai_n289_));
  OR3        m0261(.A(mai_mai_n73_), .B(mai_mai_n75_), .C(e), .Y(mai_mai_n290_));
  AOI210     m0262(.A0(mai_mai_n289_), .A1(mai_mai_n288_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  INV        m0263(.A(mai_mai_n291_), .Y(mai_mai_n292_));
  NAi32      m0264(.An(j), .Bn(h), .C(i), .Y(mai_mai_n293_));
  NAi21      m0265(.An(m), .B(l), .Y(mai_mai_n294_));
  NO3        m0266(.A(mai_mai_n294_), .B(mai_mai_n293_), .C(mai_mai_n83_), .Y(mai_mai_n295_));
  NA2        m0267(.A(h), .B(g), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n163_), .B(mai_mai_n45_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  OAI210     m0270(.A0(mai_mai_n298_), .A1(mai_mai_n295_), .B0(mai_mai_n158_), .Y(mai_mai_n299_));
  NA4        m0271(.A(mai_mai_n299_), .B(mai_mai_n292_), .C(mai_mai_n284_), .D(mai_mai_n277_), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n140_), .B(d), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n301_), .B(mai_mai_n53_), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n103_), .B(mai_mai_n100_), .Y(mai_mai_n303_));
  NAi32      m0275(.An(n), .Bn(m), .C(l), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n304_), .B(mai_mai_n293_), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n120_), .B(mai_mai_n114_), .Y(mai_mai_n306_));
  NAi31      m0278(.An(k), .B(l), .C(j), .Y(mai_mai_n307_));
  OAI210     m0279(.A0(mai_mai_n285_), .A1(j), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  NOi21      m0280(.An(mai_mai_n308_), .B(mai_mai_n118_), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n309_), .B(mai_mai_n306_), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n310_), .B(mai_mai_n302_), .Y(mai_mai_n311_));
  NO4        m0283(.A(mai_mai_n311_), .B(mai_mai_n300_), .C(mai_mai_n274_), .D(mai_mai_n266_), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n249_), .B(mai_mai_n188_), .Y(mai_mai_n313_));
  NAi21      m0285(.An(m), .B(k), .Y(mai_mai_n314_));
  NO2        m0286(.A(mai_mai_n221_), .B(mai_mai_n314_), .Y(mai_mai_n315_));
  NAi41      m0287(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n316_));
  NO2        m0288(.A(mai_mai_n316_), .B(mai_mai_n145_), .Y(mai_mai_n317_));
  NA2        m0289(.A(mai_mai_n317_), .B(mai_mai_n315_), .Y(mai_mai_n318_));
  NAi31      m0290(.An(i), .B(l), .C(h), .Y(mai_mai_n319_));
  NO4        m0291(.A(mai_mai_n319_), .B(mai_mai_n145_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n320_));
  NA2        m0292(.A(e), .B(c), .Y(mai_mai_n321_));
  NO3        m0293(.A(mai_mai_n321_), .B(n), .C(d), .Y(mai_mai_n322_));
  NOi21      m0294(.An(f), .B(h), .Y(mai_mai_n323_));
  NA2        m0295(.A(mai_mai_n323_), .B(mai_mai_n116_), .Y(mai_mai_n324_));
  NO2        m0296(.A(mai_mai_n324_), .B(mai_mai_n211_), .Y(mai_mai_n325_));
  NAi31      m0297(.An(d), .B(e), .C(b), .Y(mai_mai_n326_));
  NO2        m0298(.A(mai_mai_n130_), .B(mai_mai_n326_), .Y(mai_mai_n327_));
  NA2        m0299(.A(mai_mai_n327_), .B(mai_mai_n325_), .Y(mai_mai_n328_));
  NAi41      m0300(.An(mai_mai_n320_), .B(mai_mai_n328_), .C(mai_mai_n318_), .D(mai_mai_n313_), .Y(mai_mai_n329_));
  NO4        m0301(.A(mai_mai_n316_), .B(mai_mai_n80_), .C(mai_mai_n72_), .D(mai_mai_n211_), .Y(mai_mai_n330_));
  NA2        m0302(.A(mai_mai_n245_), .B(mai_mai_n101_), .Y(mai_mai_n331_));
  OR2        m0303(.A(mai_mai_n331_), .B(mai_mai_n200_), .Y(mai_mai_n332_));
  NOi31      m0304(.An(l), .B(n), .C(m), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n333_), .B(mai_mai_n212_), .Y(mai_mai_n334_));
  NO2        m0306(.A(mai_mai_n334_), .B(mai_mai_n189_), .Y(mai_mai_n335_));
  NAi32      m0307(.An(mai_mai_n335_), .Bn(mai_mai_n330_), .C(mai_mai_n332_), .Y(mai_mai_n336_));
  NAi32      m0308(.An(m), .Bn(j), .C(k), .Y(mai_mai_n337_));
  NAi41      m0309(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n338_));
  OAI210     m0310(.A0(mai_mai_n208_), .A1(mai_mai_n337_), .B0(mai_mai_n338_), .Y(mai_mai_n339_));
  NOi31      m0311(.An(j), .B(m), .C(k), .Y(mai_mai_n340_));
  NO2        m0312(.A(mai_mai_n124_), .B(mai_mai_n340_), .Y(mai_mai_n341_));
  AN3        m0313(.A(h), .B(g), .C(f), .Y(mai_mai_n342_));
  NAi31      m0314(.An(mai_mai_n341_), .B(mai_mai_n342_), .C(mai_mai_n339_), .Y(mai_mai_n343_));
  NOi32      m0315(.An(m), .Bn(j), .C(l), .Y(mai_mai_n344_));
  NO2        m0316(.A(mai_mai_n344_), .B(mai_mai_n95_), .Y(mai_mai_n345_));
  NO2        m0317(.A(mai_mai_n294_), .B(mai_mai_n293_), .Y(mai_mai_n346_));
  NO2        m0318(.A(mai_mai_n214_), .B(g), .Y(mai_mai_n347_));
  NA2        m0319(.A(mai_mai_n229_), .B(mai_mai_n80_), .Y(mai_mai_n348_));
  NA3        m0320(.A(mai_mai_n348_), .B(mai_mai_n342_), .C(mai_mai_n209_), .Y(mai_mai_n349_));
  NA2        m0321(.A(mai_mai_n349_), .B(mai_mai_n343_), .Y(mai_mai_n350_));
  NA3        m0322(.A(h), .B(g), .C(f), .Y(mai_mai_n351_));
  NA2        m0323(.A(mai_mai_n157_), .B(e), .Y(mai_mai_n352_));
  NO2        m0324(.A(mai_mai_n352_), .B(mai_mai_n41_), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n353_), .B(mai_mai_n306_), .Y(mai_mai_n354_));
  NOi32      m0326(.An(j), .Bn(g), .C(i), .Y(mai_mai_n355_));
  NA3        m0327(.A(mai_mai_n355_), .B(mai_mai_n285_), .C(mai_mai_n111_), .Y(mai_mai_n356_));
  OR2        m0328(.A(mai_mai_n109_), .B(mai_mai_n356_), .Y(mai_mai_n357_));
  NOi32      m0329(.An(e), .Bn(b), .C(a), .Y(mai_mai_n358_));
  AN2        m0330(.A(l), .B(j), .Y(mai_mai_n359_));
  NO2        m0331(.A(mai_mai_n314_), .B(mai_mai_n359_), .Y(mai_mai_n360_));
  NO3        m0332(.A(mai_mai_n316_), .B(mai_mai_n72_), .C(mai_mai_n211_), .Y(mai_mai_n361_));
  NA3        m0333(.A(mai_mai_n205_), .B(mai_mai_n203_), .C(mai_mai_n35_), .Y(mai_mai_n362_));
  AOI220     m0334(.A0(mai_mai_n362_), .A1(mai_mai_n358_), .B0(mai_mai_n361_), .B1(mai_mai_n360_), .Y(mai_mai_n363_));
  NO2        m0335(.A(mai_mai_n326_), .B(n), .Y(mai_mai_n364_));
  NA2        m0336(.A(mai_mai_n204_), .B(k), .Y(mai_mai_n365_));
  NA3        m0337(.A(m), .B(mai_mai_n110_), .C(mai_mai_n210_), .Y(mai_mai_n366_));
  NA4        m0338(.A(mai_mai_n199_), .B(mai_mai_n86_), .C(g), .D(mai_mai_n210_), .Y(mai_mai_n367_));
  OAI210     m0339(.A0(mai_mai_n366_), .A1(mai_mai_n365_), .B0(mai_mai_n367_), .Y(mai_mai_n368_));
  NAi41      m0340(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n369_));
  NA2        m0341(.A(mai_mai_n51_), .B(mai_mai_n111_), .Y(mai_mai_n370_));
  NO2        m0342(.A(mai_mai_n370_), .B(mai_mai_n369_), .Y(mai_mai_n371_));
  AOI220     m0343(.A0(mai_mai_n371_), .A1(b), .B0(mai_mai_n368_), .B1(mai_mai_n364_), .Y(mai_mai_n372_));
  NA4        m0344(.A(mai_mai_n372_), .B(mai_mai_n363_), .C(mai_mai_n357_), .D(mai_mai_n354_), .Y(mai_mai_n373_));
  NO4        m0345(.A(mai_mai_n373_), .B(mai_mai_n350_), .C(mai_mai_n336_), .D(mai_mai_n329_), .Y(mai_mai_n374_));
  NA4        m0346(.A(mai_mai_n374_), .B(mai_mai_n312_), .C(mai_mai_n264_), .D(mai_mai_n195_), .Y(mai10));
  NA3        m0347(.A(m), .B(k), .C(i), .Y(mai_mai_n376_));
  NO3        m0348(.A(mai_mai_n376_), .B(j), .C(mai_mai_n211_), .Y(mai_mai_n377_));
  NOi21      m0349(.An(e), .B(f), .Y(mai_mai_n378_));
  NO4        m0350(.A(mai_mai_n146_), .B(mai_mai_n378_), .C(n), .D(mai_mai_n108_), .Y(mai_mai_n379_));
  NAi31      m0351(.An(b), .B(f), .C(c), .Y(mai_mai_n380_));
  INV        m0352(.A(mai_mai_n380_), .Y(mai_mai_n381_));
  NOi32      m0353(.An(k), .Bn(h), .C(j), .Y(mai_mai_n382_));
  NA2        m0354(.A(mai_mai_n382_), .B(mai_mai_n216_), .Y(mai_mai_n383_));
  NA2        m0355(.A(mai_mai_n155_), .B(mai_mai_n383_), .Y(mai_mai_n384_));
  AOI220     m0356(.A0(mai_mai_n384_), .A1(mai_mai_n381_), .B0(mai_mai_n379_), .B1(mai_mai_n377_), .Y(mai_mai_n385_));
  AN2        m0357(.A(j), .B(h), .Y(mai_mai_n386_));
  NO3        m0358(.A(n), .B(m), .C(k), .Y(mai_mai_n387_));
  NA2        m0359(.A(mai_mai_n387_), .B(mai_mai_n386_), .Y(mai_mai_n388_));
  NO3        m0360(.A(mai_mai_n388_), .B(mai_mai_n146_), .C(mai_mai_n210_), .Y(mai_mai_n389_));
  OR2        m0361(.A(m), .B(k), .Y(mai_mai_n390_));
  NO2        m0362(.A(mai_mai_n170_), .B(mai_mai_n390_), .Y(mai_mai_n391_));
  NA4        m0363(.A(n), .B(f), .C(c), .D(mai_mai_n114_), .Y(mai_mai_n392_));
  NOi21      m0364(.An(mai_mai_n391_), .B(mai_mai_n392_), .Y(mai_mai_n393_));
  NOi32      m0365(.An(d), .Bn(a), .C(c), .Y(mai_mai_n394_));
  NA2        m0366(.A(mai_mai_n394_), .B(mai_mai_n178_), .Y(mai_mai_n395_));
  NAi21      m0367(.An(i), .B(g), .Y(mai_mai_n396_));
  NAi31      m0368(.An(k), .B(m), .C(j), .Y(mai_mai_n397_));
  NO3        m0369(.A(mai_mai_n397_), .B(mai_mai_n396_), .C(n), .Y(mai_mai_n398_));
  NOi21      m0370(.An(mai_mai_n398_), .B(mai_mai_n395_), .Y(mai_mai_n399_));
  NO3        m0371(.A(mai_mai_n399_), .B(mai_mai_n393_), .C(mai_mai_n389_), .Y(mai_mai_n400_));
  NO2        m0372(.A(mai_mai_n392_), .B(mai_mai_n294_), .Y(mai_mai_n401_));
  NOi32      m0373(.An(f), .Bn(d), .C(c), .Y(mai_mai_n402_));
  AOI220     m0374(.A0(mai_mai_n402_), .A1(mai_mai_n305_), .B0(mai_mai_n401_), .B1(mai_mai_n212_), .Y(mai_mai_n403_));
  NA3        m0375(.A(mai_mai_n403_), .B(mai_mai_n400_), .C(mai_mai_n385_), .Y(mai_mai_n404_));
  NO2        m0376(.A(mai_mai_n59_), .B(mai_mai_n114_), .Y(mai_mai_n405_));
  NA2        m0377(.A(mai_mai_n245_), .B(mai_mai_n405_), .Y(mai_mai_n406_));
  INV        m0378(.A(e), .Y(mai_mai_n407_));
  NA2        m0379(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n408_));
  OAI220     m0380(.A0(mai_mai_n408_), .A1(mai_mai_n196_), .B0(mai_mai_n200_), .B1(mai_mai_n407_), .Y(mai_mai_n409_));
  AN2        m0381(.A(g), .B(e), .Y(mai_mai_n410_));
  NA3        m0382(.A(mai_mai_n410_), .B(mai_mai_n199_), .C(i), .Y(mai_mai_n411_));
  OAI210     m0383(.A0(mai_mai_n88_), .A1(mai_mai_n407_), .B0(mai_mai_n411_), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n98_), .B(mai_mai_n407_), .Y(mai_mai_n413_));
  NO3        m0385(.A(mai_mai_n413_), .B(mai_mai_n412_), .C(mai_mai_n409_), .Y(mai_mai_n414_));
  NOi32      m0386(.An(h), .Bn(e), .C(g), .Y(mai_mai_n415_));
  NA3        m0387(.A(mai_mai_n415_), .B(mai_mai_n287_), .C(m), .Y(mai_mai_n416_));
  NOi21      m0388(.An(g), .B(h), .Y(mai_mai_n417_));
  AN3        m0389(.A(m), .B(l), .C(i), .Y(mai_mai_n418_));
  NA3        m0390(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(e), .Y(mai_mai_n419_));
  AN3        m0391(.A(h), .B(g), .C(e), .Y(mai_mai_n420_));
  NA2        m0392(.A(mai_mai_n420_), .B(mai_mai_n95_), .Y(mai_mai_n421_));
  AN3        m0393(.A(mai_mai_n421_), .B(mai_mai_n419_), .C(mai_mai_n416_), .Y(mai_mai_n422_));
  AOI210     m0394(.A0(mai_mai_n422_), .A1(mai_mai_n414_), .B0(mai_mai_n406_), .Y(mai_mai_n423_));
  NA3        m0395(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n424_));
  NO2        m0396(.A(mai_mai_n424_), .B(mai_mai_n406_), .Y(mai_mai_n425_));
  NA3        m0397(.A(mai_mai_n394_), .B(mai_mai_n178_), .C(mai_mai_n83_), .Y(mai_mai_n426_));
  NAi31      m0398(.An(b), .B(c), .C(a), .Y(mai_mai_n427_));
  NO2        m0399(.A(mai_mai_n427_), .B(n), .Y(mai_mai_n428_));
  OAI210     m0400(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n429_));
  NO2        m0401(.A(mai_mai_n429_), .B(mai_mai_n142_), .Y(mai_mai_n430_));
  NA2        m0402(.A(mai_mai_n430_), .B(mai_mai_n428_), .Y(mai_mai_n431_));
  INV        m0403(.A(mai_mai_n431_), .Y(mai_mai_n432_));
  NO4        m0404(.A(mai_mai_n432_), .B(mai_mai_n425_), .C(mai_mai_n423_), .D(mai_mai_n404_), .Y(mai_mai_n433_));
  NA2        m0405(.A(i), .B(g), .Y(mai_mai_n434_));
  NO3        m0406(.A(mai_mai_n272_), .B(mai_mai_n434_), .C(c), .Y(mai_mai_n435_));
  NOi21      m0407(.An(a), .B(n), .Y(mai_mai_n436_));
  NOi21      m0408(.An(d), .B(c), .Y(mai_mai_n437_));
  NA2        m0409(.A(mai_mai_n437_), .B(mai_mai_n436_), .Y(mai_mai_n438_));
  NA3        m0410(.A(i), .B(g), .C(f), .Y(mai_mai_n439_));
  OR2        m0411(.A(mai_mai_n439_), .B(mai_mai_n71_), .Y(mai_mai_n440_));
  NA3        m0412(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(mai_mai_n178_), .Y(mai_mai_n441_));
  AOI210     m0413(.A0(mai_mai_n441_), .A1(mai_mai_n440_), .B0(mai_mai_n438_), .Y(mai_mai_n442_));
  AOI210     m0414(.A0(mai_mai_n435_), .A1(mai_mai_n286_), .B0(mai_mai_n442_), .Y(mai_mai_n443_));
  OR2        m0415(.A(n), .B(m), .Y(mai_mai_n444_));
  NO2        m0416(.A(mai_mai_n444_), .B(mai_mai_n147_), .Y(mai_mai_n445_));
  NO2        m0417(.A(mai_mai_n179_), .B(mai_mai_n142_), .Y(mai_mai_n446_));
  OAI210     m0418(.A0(mai_mai_n445_), .A1(mai_mai_n172_), .B0(mai_mai_n446_), .Y(mai_mai_n447_));
  INV        m0419(.A(mai_mai_n370_), .Y(mai_mai_n448_));
  NA3        m0420(.A(mai_mai_n448_), .B(mai_mai_n358_), .C(d), .Y(mai_mai_n449_));
  NO2        m0421(.A(mai_mai_n427_), .B(mai_mai_n49_), .Y(mai_mai_n450_));
  NAi21      m0422(.An(k), .B(j), .Y(mai_mai_n451_));
  NAi21      m0423(.An(e), .B(d), .Y(mai_mai_n452_));
  INV        m0424(.A(mai_mai_n452_), .Y(mai_mai_n453_));
  NO2        m0425(.A(mai_mai_n248_), .B(mai_mai_n210_), .Y(mai_mai_n454_));
  NA3        m0426(.A(mai_mai_n454_), .B(mai_mai_n453_), .C(mai_mai_n222_), .Y(mai_mai_n455_));
  NA3        m0427(.A(mai_mai_n455_), .B(mai_mai_n449_), .C(mai_mai_n447_), .Y(mai_mai_n456_));
  NO2        m0428(.A(mai_mai_n334_), .B(mai_mai_n210_), .Y(mai_mai_n457_));
  NA2        m0429(.A(mai_mai_n457_), .B(mai_mai_n453_), .Y(mai_mai_n458_));
  NOi31      m0430(.An(n), .B(m), .C(k), .Y(mai_mai_n459_));
  AOI220     m0431(.A0(mai_mai_n459_), .A1(mai_mai_n386_), .B0(mai_mai_n216_), .B1(mai_mai_n50_), .Y(mai_mai_n460_));
  NAi31      m0432(.An(g), .B(f), .C(c), .Y(mai_mai_n461_));
  OR3        m0433(.A(mai_mai_n461_), .B(mai_mai_n460_), .C(e), .Y(mai_mai_n462_));
  NA2        m0434(.A(mai_mai_n462_), .B(mai_mai_n458_), .Y(mai_mai_n463_));
  NOi41      m0435(.An(mai_mai_n443_), .B(mai_mai_n463_), .C(mai_mai_n456_), .D(mai_mai_n262_), .Y(mai_mai_n464_));
  NOi32      m0436(.An(c), .Bn(a), .C(b), .Y(mai_mai_n465_));
  NA2        m0437(.A(mai_mai_n465_), .B(mai_mai_n111_), .Y(mai_mai_n466_));
  INV        m0438(.A(mai_mai_n270_), .Y(mai_mai_n467_));
  AN2        m0439(.A(e), .B(d), .Y(mai_mai_n468_));
  NA2        m0440(.A(mai_mai_n468_), .B(mai_mai_n467_), .Y(mai_mai_n469_));
  NO2        m0441(.A(mai_mai_n129_), .B(mai_mai_n41_), .Y(mai_mai_n470_));
  NO2        m0442(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n471_));
  NOi31      m0443(.An(j), .B(k), .C(i), .Y(mai_mai_n472_));
  NOi21      m0444(.An(mai_mai_n160_), .B(mai_mai_n472_), .Y(mai_mai_n473_));
  NA4        m0445(.A(mai_mai_n319_), .B(mai_mai_n473_), .C(mai_mai_n256_), .D(mai_mai_n117_), .Y(mai_mai_n474_));
  NA2        m0446(.A(mai_mai_n474_), .B(mai_mai_n471_), .Y(mai_mai_n475_));
  AOI210     m0447(.A0(mai_mai_n475_), .A1(mai_mai_n469_), .B0(mai_mai_n466_), .Y(mai_mai_n476_));
  NO2        m0448(.A(mai_mai_n206_), .B(mai_mai_n201_), .Y(mai_mai_n477_));
  NOi21      m0449(.An(a), .B(b), .Y(mai_mai_n478_));
  NA3        m0450(.A(e), .B(d), .C(c), .Y(mai_mai_n479_));
  NAi21      m0451(.An(mai_mai_n479_), .B(mai_mai_n478_), .Y(mai_mai_n480_));
  AOI210     m0452(.A0(mai_mai_n265_), .A1(mai_mai_n477_), .B0(mai_mai_n480_), .Y(mai_mai_n481_));
  NO4        m0453(.A(mai_mai_n183_), .B(mai_mai_n100_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n482_));
  NA2        m0454(.A(mai_mai_n381_), .B(mai_mai_n148_), .Y(mai_mai_n483_));
  OR2        m0455(.A(k), .B(j), .Y(mai_mai_n484_));
  NA2        m0456(.A(l), .B(k), .Y(mai_mai_n485_));
  AOI210     m0457(.A0(mai_mai_n229_), .A1(mai_mai_n337_), .B0(mai_mai_n83_), .Y(mai_mai_n486_));
  INV        m0458(.A(mai_mai_n126_), .Y(mai_mai_n487_));
  NA2        m0459(.A(mai_mai_n394_), .B(mai_mai_n111_), .Y(mai_mai_n488_));
  NO4        m0460(.A(mai_mai_n488_), .B(mai_mai_n92_), .C(mai_mai_n110_), .D(e), .Y(mai_mai_n489_));
  NO3        m0461(.A(mai_mai_n426_), .B(mai_mai_n90_), .C(mai_mai_n129_), .Y(mai_mai_n490_));
  NO4        m0462(.A(mai_mai_n490_), .B(mai_mai_n489_), .C(mai_mai_n487_), .D(mai_mai_n320_), .Y(mai_mai_n491_));
  NA2        m0463(.A(mai_mai_n491_), .B(mai_mai_n483_), .Y(mai_mai_n492_));
  NO4        m0464(.A(mai_mai_n492_), .B(mai_mai_n482_), .C(mai_mai_n481_), .D(mai_mai_n476_), .Y(mai_mai_n493_));
  NA2        m0465(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n494_));
  NOi21      m0466(.An(d), .B(e), .Y(mai_mai_n495_));
  NAi31      m0467(.An(j), .B(l), .C(i), .Y(mai_mai_n496_));
  INV        m0468(.A(mai_mai_n100_), .Y(mai_mai_n497_));
  NO3        m0469(.A(mai_mai_n395_), .B(mai_mai_n345_), .C(mai_mai_n197_), .Y(mai_mai_n498_));
  NO2        m0470(.A(mai_mai_n395_), .B(mai_mai_n370_), .Y(mai_mai_n499_));
  NO3        m0471(.A(mai_mai_n499_), .B(mai_mai_n498_), .C(mai_mai_n303_), .Y(mai_mai_n500_));
  NA3        m0472(.A(mai_mai_n500_), .B(mai_mai_n494_), .C(mai_mai_n239_), .Y(mai_mai_n501_));
  OAI210     m0473(.A0(mai_mai_n125_), .A1(mai_mai_n124_), .B0(n), .Y(mai_mai_n502_));
  NO2        m0474(.A(mai_mai_n502_), .B(mai_mai_n129_), .Y(mai_mai_n503_));
  OA210      m0475(.A0(mai_mai_n241_), .A1(mai_mai_n503_), .B0(mai_mai_n188_), .Y(mai_mai_n504_));
  XO2        m0476(.A(i), .B(h), .Y(mai_mai_n505_));
  NA3        m0477(.A(mai_mai_n505_), .B(mai_mai_n154_), .C(n), .Y(mai_mai_n506_));
  NAi41      m0478(.An(mai_mai_n295_), .B(mai_mai_n506_), .C(mai_mai_n460_), .D(mai_mai_n383_), .Y(mai_mai_n507_));
  NOi32      m0479(.An(mai_mai_n507_), .Bn(mai_mai_n471_), .C(mai_mai_n267_), .Y(mai_mai_n508_));
  NAi31      m0480(.An(c), .B(f), .C(d), .Y(mai_mai_n509_));
  AOI210     m0481(.A0(mai_mai_n275_), .A1(mai_mai_n191_), .B0(mai_mai_n509_), .Y(mai_mai_n510_));
  INV        m0482(.A(mai_mai_n510_), .Y(mai_mai_n511_));
  NA3        m0483(.A(mai_mai_n379_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n512_));
  NA2        m0484(.A(mai_mai_n223_), .B(mai_mai_n106_), .Y(mai_mai_n513_));
  AOI210     m0485(.A0(mai_mai_n513_), .A1(mai_mai_n177_), .B0(mai_mai_n509_), .Y(mai_mai_n514_));
  AOI210     m0486(.A0(mai_mai_n356_), .A1(mai_mai_n35_), .B0(mai_mai_n480_), .Y(mai_mai_n515_));
  NOi31      m0487(.An(mai_mai_n512_), .B(mai_mai_n515_), .C(mai_mai_n514_), .Y(mai_mai_n516_));
  AO220      m0488(.A0(mai_mai_n283_), .A1(mai_mai_n259_), .B0(mai_mai_n161_), .B1(mai_mai_n67_), .Y(mai_mai_n517_));
  NA3        m0489(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n518_));
  NO2        m0490(.A(mai_mai_n518_), .B(mai_mai_n438_), .Y(mai_mai_n519_));
  NO2        m0491(.A(mai_mai_n519_), .B(mai_mai_n291_), .Y(mai_mai_n520_));
  NAi41      m0492(.An(mai_mai_n517_), .B(mai_mai_n520_), .C(mai_mai_n516_), .D(mai_mai_n511_), .Y(mai_mai_n521_));
  NO4        m0493(.A(mai_mai_n521_), .B(mai_mai_n508_), .C(mai_mai_n504_), .D(mai_mai_n501_), .Y(mai_mai_n522_));
  NA4        m0494(.A(mai_mai_n522_), .B(mai_mai_n493_), .C(mai_mai_n464_), .D(mai_mai_n433_), .Y(mai11));
  NO2        m0495(.A(mai_mai_n73_), .B(f), .Y(mai_mai_n524_));
  NA2        m0496(.A(j), .B(g), .Y(mai_mai_n525_));
  NAi31      m0497(.An(i), .B(m), .C(l), .Y(mai_mai_n526_));
  NA3        m0498(.A(m), .B(k), .C(j), .Y(mai_mai_n527_));
  OAI220     m0499(.A0(mai_mai_n527_), .A1(mai_mai_n129_), .B0(mai_mai_n526_), .B1(mai_mai_n525_), .Y(mai_mai_n528_));
  NA2        m0500(.A(mai_mai_n528_), .B(mai_mai_n524_), .Y(mai_mai_n529_));
  NOi32      m0501(.An(e), .Bn(b), .C(f), .Y(mai_mai_n530_));
  NA2        m0502(.A(mai_mai_n255_), .B(mai_mai_n111_), .Y(mai_mai_n531_));
  NA2        m0503(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n532_));
  NO2        m0504(.A(mai_mai_n532_), .B(mai_mai_n297_), .Y(mai_mai_n533_));
  NAi31      m0505(.An(d), .B(e), .C(a), .Y(mai_mai_n534_));
  NO2        m0506(.A(mai_mai_n534_), .B(n), .Y(mai_mai_n535_));
  AOI220     m0507(.A0(mai_mai_n535_), .A1(mai_mai_n99_), .B0(mai_mai_n533_), .B1(mai_mai_n530_), .Y(mai_mai_n536_));
  NAi41      m0508(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n537_));
  AN2        m0509(.A(mai_mai_n537_), .B(mai_mai_n369_), .Y(mai_mai_n538_));
  AOI210     m0510(.A0(mai_mai_n538_), .A1(mai_mai_n395_), .B0(mai_mai_n268_), .Y(mai_mai_n539_));
  NA2        m0511(.A(j), .B(i), .Y(mai_mai_n540_));
  NAi31      m0512(.An(n), .B(m), .C(k), .Y(mai_mai_n541_));
  NO3        m0513(.A(mai_mai_n541_), .B(mai_mai_n540_), .C(mai_mai_n110_), .Y(mai_mai_n542_));
  NO4        m0514(.A(n), .B(d), .C(mai_mai_n114_), .D(a), .Y(mai_mai_n543_));
  OR2        m0515(.A(n), .B(c), .Y(mai_mai_n544_));
  NO2        m0516(.A(mai_mai_n544_), .B(mai_mai_n144_), .Y(mai_mai_n545_));
  NO2        m0517(.A(mai_mai_n545_), .B(mai_mai_n543_), .Y(mai_mai_n546_));
  NOi32      m0518(.An(g), .Bn(f), .C(i), .Y(mai_mai_n547_));
  AOI220     m0519(.A0(mai_mai_n547_), .A1(mai_mai_n97_), .B0(mai_mai_n528_), .B1(f), .Y(mai_mai_n548_));
  NO2        m0520(.A(mai_mai_n270_), .B(mai_mai_n49_), .Y(mai_mai_n549_));
  NO2        m0521(.A(mai_mai_n548_), .B(mai_mai_n546_), .Y(mai_mai_n550_));
  AOI210     m0522(.A0(mai_mai_n542_), .A1(mai_mai_n539_), .B0(mai_mai_n550_), .Y(mai_mai_n551_));
  NA2        m0523(.A(mai_mai_n137_), .B(mai_mai_n34_), .Y(mai_mai_n552_));
  OAI220     m0524(.A0(mai_mai_n552_), .A1(m), .B0(mai_mai_n532_), .B1(mai_mai_n229_), .Y(mai_mai_n553_));
  NOi41      m0525(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n554_));
  NAi32      m0526(.An(e), .Bn(b), .C(c), .Y(mai_mai_n555_));
  OR2        m0527(.A(mai_mai_n555_), .B(mai_mai_n83_), .Y(mai_mai_n556_));
  AN2        m0528(.A(mai_mai_n338_), .B(mai_mai_n316_), .Y(mai_mai_n557_));
  NA2        m0529(.A(mai_mai_n557_), .B(mai_mai_n556_), .Y(mai_mai_n558_));
  OA210      m0530(.A0(mai_mai_n558_), .A1(mai_mai_n554_), .B0(mai_mai_n553_), .Y(mai_mai_n559_));
  OAI220     m0531(.A0(mai_mai_n397_), .A1(mai_mai_n396_), .B0(mai_mai_n526_), .B1(mai_mai_n525_), .Y(mai_mai_n560_));
  NAi31      m0532(.An(d), .B(c), .C(a), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n561_), .B(n), .Y(mai_mai_n562_));
  NA3        m0534(.A(mai_mai_n562_), .B(mai_mai_n560_), .C(e), .Y(mai_mai_n563_));
  NO3        m0535(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n211_), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n226_), .B(mai_mai_n108_), .Y(mai_mai_n565_));
  OAI210     m0537(.A0(mai_mai_n564_), .A1(mai_mai_n398_), .B0(mai_mai_n565_), .Y(mai_mai_n566_));
  NA2        m0538(.A(mai_mai_n566_), .B(mai_mai_n563_), .Y(mai_mai_n567_));
  NO2        m0539(.A(mai_mai_n272_), .B(n), .Y(mai_mai_n568_));
  NO2        m0540(.A(mai_mai_n428_), .B(mai_mai_n568_), .Y(mai_mai_n569_));
  NA2        m0541(.A(mai_mai_n560_), .B(f), .Y(mai_mai_n570_));
  NAi32      m0542(.An(d), .Bn(a), .C(b), .Y(mai_mai_n571_));
  NA2        m0543(.A(h), .B(f), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n572_), .B(mai_mai_n92_), .Y(mai_mai_n573_));
  NO2        m0545(.A(mai_mai_n570_), .B(mai_mai_n569_), .Y(mai_mai_n574_));
  AN3        m0546(.A(j), .B(h), .C(g), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n141_), .B(c), .Y(mai_mai_n576_));
  NA3        m0548(.A(mai_mai_n576_), .B(mai_mai_n575_), .C(mai_mai_n459_), .Y(mai_mai_n577_));
  NA3        m0549(.A(f), .B(d), .C(b), .Y(mai_mai_n578_));
  NO4        m0550(.A(mai_mai_n578_), .B(mai_mai_n173_), .C(mai_mai_n170_), .D(g), .Y(mai_mai_n579_));
  INV        m0551(.A(mai_mai_n577_), .Y(mai_mai_n580_));
  NO4        m0552(.A(mai_mai_n580_), .B(mai_mai_n574_), .C(mai_mai_n567_), .D(mai_mai_n559_), .Y(mai_mai_n581_));
  AN4        m0553(.A(mai_mai_n581_), .B(mai_mai_n551_), .C(mai_mai_n536_), .D(mai_mai_n529_), .Y(mai_mai_n582_));
  INV        m0554(.A(k), .Y(mai_mai_n583_));
  NA3        m0555(.A(l), .B(mai_mai_n583_), .C(i), .Y(mai_mai_n584_));
  INV        m0556(.A(mai_mai_n584_), .Y(mai_mai_n585_));
  NA4        m0557(.A(mai_mai_n394_), .B(mai_mai_n417_), .C(mai_mai_n178_), .D(mai_mai_n111_), .Y(mai_mai_n586_));
  NAi32      m0558(.An(h), .Bn(f), .C(g), .Y(mai_mai_n587_));
  NAi41      m0559(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n588_));
  OAI210     m0560(.A0(mai_mai_n534_), .A1(n), .B0(mai_mai_n588_), .Y(mai_mai_n589_));
  NA2        m0561(.A(mai_mai_n589_), .B(m), .Y(mai_mai_n590_));
  NAi31      m0562(.An(h), .B(g), .C(f), .Y(mai_mai_n591_));
  OR3        m0563(.A(mai_mai_n591_), .B(mai_mai_n272_), .C(mai_mai_n49_), .Y(mai_mai_n592_));
  NA4        m0564(.A(mai_mai_n417_), .B(mai_mai_n119_), .C(mai_mai_n111_), .D(e), .Y(mai_mai_n593_));
  AN2        m0565(.A(mai_mai_n593_), .B(mai_mai_n592_), .Y(mai_mai_n594_));
  OA210      m0566(.A0(mai_mai_n590_), .A1(mai_mai_n587_), .B0(mai_mai_n594_), .Y(mai_mai_n595_));
  NO4        m0567(.A(mai_mai_n591_), .B(mai_mai_n544_), .C(mai_mai_n144_), .D(mai_mai_n75_), .Y(mai_mai_n596_));
  NAi31      m0568(.An(mai_mai_n596_), .B(mai_mai_n595_), .C(mai_mai_n586_), .Y(mai_mai_n597_));
  NAi31      m0569(.An(f), .B(h), .C(g), .Y(mai_mai_n598_));
  NO4        m0570(.A(mai_mai_n307_), .B(mai_mai_n598_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n599_));
  NOi32      m0571(.An(b), .Bn(a), .C(c), .Y(mai_mai_n600_));
  NOi41      m0572(.An(mai_mai_n600_), .B(mai_mai_n351_), .C(mai_mai_n69_), .D(mai_mai_n115_), .Y(mai_mai_n601_));
  OR2        m0573(.A(mai_mai_n601_), .B(mai_mai_n599_), .Y(mai_mai_n602_));
  NOi32      m0574(.An(d), .Bn(a), .C(e), .Y(mai_mai_n603_));
  NA2        m0575(.A(mai_mai_n603_), .B(mai_mai_n111_), .Y(mai_mai_n604_));
  NO2        m0576(.A(n), .B(c), .Y(mai_mai_n605_));
  NA3        m0577(.A(mai_mai_n605_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n606_));
  NAi32      m0578(.An(n), .Bn(f), .C(m), .Y(mai_mai_n607_));
  NA3        m0579(.A(mai_mai_n607_), .B(mai_mai_n606_), .C(mai_mai_n604_), .Y(mai_mai_n608_));
  NOi32      m0580(.An(e), .Bn(a), .C(d), .Y(mai_mai_n609_));
  AOI210     m0581(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n609_), .Y(mai_mai_n610_));
  AOI210     m0582(.A0(mai_mai_n610_), .A1(mai_mai_n210_), .B0(mai_mai_n552_), .Y(mai_mai_n611_));
  AOI210     m0583(.A0(mai_mai_n611_), .A1(mai_mai_n608_), .B0(mai_mai_n602_), .Y(mai_mai_n612_));
  INV        m0584(.A(mai_mai_n612_), .Y(mai_mai_n613_));
  AOI210     m0585(.A0(mai_mai_n597_), .A1(mai_mai_n585_), .B0(mai_mai_n613_), .Y(mai_mai_n614_));
  NO3        m0586(.A(mai_mai_n314_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n615_));
  NA3        m0587(.A(mai_mai_n509_), .B(mai_mai_n168_), .C(mai_mai_n167_), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n461_), .B(mai_mai_n226_), .Y(mai_mai_n617_));
  OR2        m0589(.A(mai_mai_n617_), .B(mai_mai_n616_), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n76_), .B(mai_mai_n111_), .Y(mai_mai_n619_));
  NO2        m0591(.A(mai_mai_n619_), .B(mai_mai_n45_), .Y(mai_mai_n620_));
  AOI220     m0592(.A0(mai_mai_n620_), .A1(mai_mai_n539_), .B0(mai_mai_n618_), .B1(mai_mai_n615_), .Y(mai_mai_n621_));
  NO2        m0593(.A(mai_mai_n621_), .B(mai_mai_n86_), .Y(mai_mai_n622_));
  NA3        m0594(.A(mai_mai_n554_), .B(mai_mai_n340_), .C(mai_mai_n46_), .Y(mai_mai_n623_));
  NOi32      m0595(.An(e), .Bn(c), .C(f), .Y(mai_mai_n624_));
  NOi21      m0596(.An(f), .B(g), .Y(mai_mai_n625_));
  NO2        m0597(.A(mai_mai_n625_), .B(mai_mai_n208_), .Y(mai_mai_n626_));
  AOI220     m0598(.A0(mai_mai_n626_), .A1(mai_mai_n391_), .B0(mai_mai_n624_), .B1(mai_mai_n172_), .Y(mai_mai_n627_));
  NA3        m0599(.A(mai_mai_n627_), .B(mai_mai_n623_), .C(mai_mai_n175_), .Y(mai_mai_n628_));
  AOI210     m0600(.A0(mai_mai_n538_), .A1(mai_mai_n395_), .B0(mai_mai_n296_), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n629_), .B(mai_mai_n260_), .Y(mai_mai_n630_));
  NOi21      m0602(.An(j), .B(l), .Y(mai_mai_n631_));
  NAi21      m0603(.An(k), .B(h), .Y(mai_mai_n632_));
  NO2        m0604(.A(mai_mai_n632_), .B(mai_mai_n258_), .Y(mai_mai_n633_));
  NOi31      m0605(.An(m), .B(n), .C(k), .Y(mai_mai_n634_));
  NA2        m0606(.A(mai_mai_n631_), .B(mai_mai_n634_), .Y(mai_mai_n635_));
  AOI210     m0607(.A0(mai_mai_n395_), .A1(mai_mai_n369_), .B0(mai_mai_n296_), .Y(mai_mai_n636_));
  NAi21      m0608(.An(mai_mai_n635_), .B(mai_mai_n636_), .Y(mai_mai_n637_));
  NO2        m0609(.A(mai_mai_n272_), .B(mai_mai_n49_), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n534_), .B(mai_mai_n49_), .Y(mai_mai_n639_));
  NA2        m0611(.A(mai_mai_n638_), .B(mai_mai_n573_), .Y(mai_mai_n640_));
  NA3        m0612(.A(mai_mai_n640_), .B(mai_mai_n637_), .C(mai_mai_n630_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n106_), .B(mai_mai_n36_), .Y(mai_mai_n642_));
  NO2        m0614(.A(k), .B(mai_mai_n211_), .Y(mai_mai_n643_));
  NO2        m0615(.A(mai_mai_n530_), .B(mai_mai_n358_), .Y(mai_mai_n644_));
  NO2        m0616(.A(mai_mai_n644_), .B(n), .Y(mai_mai_n645_));
  NAi31      m0617(.An(mai_mai_n642_), .B(mai_mai_n645_), .C(mai_mai_n643_), .Y(mai_mai_n646_));
  NO2        m0618(.A(mai_mai_n532_), .B(mai_mai_n173_), .Y(mai_mai_n647_));
  NA3        m0619(.A(mai_mai_n555_), .B(mai_mai_n267_), .C(mai_mai_n140_), .Y(mai_mai_n648_));
  NA2        m0620(.A(mai_mai_n505_), .B(mai_mai_n154_), .Y(mai_mai_n649_));
  NO3        m0621(.A(mai_mai_n392_), .B(mai_mai_n649_), .C(mai_mai_n86_), .Y(mai_mai_n650_));
  AOI210     m0622(.A0(mai_mai_n648_), .A1(mai_mai_n647_), .B0(mai_mai_n650_), .Y(mai_mai_n651_));
  AN3        m0623(.A(f), .B(d), .C(b), .Y(mai_mai_n652_));
  OAI210     m0624(.A0(mai_mai_n652_), .A1(mai_mai_n128_), .B0(n), .Y(mai_mai_n653_));
  NA3        m0625(.A(mai_mai_n505_), .B(mai_mai_n154_), .C(mai_mai_n211_), .Y(mai_mai_n654_));
  AOI210     m0626(.A0(mai_mai_n653_), .A1(mai_mai_n228_), .B0(mai_mai_n654_), .Y(mai_mai_n655_));
  NAi31      m0627(.An(m), .B(n), .C(k), .Y(mai_mai_n656_));
  INV        m0628(.A(mai_mai_n246_), .Y(mai_mai_n657_));
  OAI210     m0629(.A0(mai_mai_n657_), .A1(mai_mai_n655_), .B0(j), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n658_), .B(mai_mai_n651_), .C(mai_mai_n646_), .Y(mai_mai_n659_));
  NO4        m0631(.A(mai_mai_n659_), .B(mai_mai_n641_), .C(mai_mai_n628_), .D(mai_mai_n622_), .Y(mai_mai_n660_));
  NAi31      m0632(.An(g), .B(h), .C(f), .Y(mai_mai_n661_));
  OR3        m0633(.A(mai_mai_n661_), .B(mai_mai_n272_), .C(n), .Y(mai_mai_n662_));
  OA210      m0634(.A0(mai_mai_n534_), .A1(n), .B0(mai_mai_n588_), .Y(mai_mai_n663_));
  NA3        m0635(.A(mai_mai_n415_), .B(mai_mai_n119_), .C(mai_mai_n83_), .Y(mai_mai_n664_));
  OAI210     m0636(.A0(mai_mai_n663_), .A1(mai_mai_n89_), .B0(mai_mai_n664_), .Y(mai_mai_n665_));
  NOi21      m0637(.An(mai_mai_n662_), .B(mai_mai_n665_), .Y(mai_mai_n666_));
  NO2        m0638(.A(mai_mai_n666_), .B(mai_mai_n527_), .Y(mai_mai_n667_));
  NO3        m0639(.A(g), .B(mai_mai_n210_), .C(mai_mai_n56_), .Y(mai_mai_n668_));
  NO2        m0640(.A(mai_mai_n513_), .B(mai_mai_n86_), .Y(mai_mai_n669_));
  OAI210     m0641(.A0(mai_mai_n669_), .A1(mai_mai_n391_), .B0(mai_mai_n668_), .Y(mai_mai_n670_));
  OR2        m0642(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n600_), .B(mai_mai_n342_), .Y(mai_mai_n672_));
  OR2        m0644(.A(mai_mai_n635_), .B(mai_mai_n672_), .Y(mai_mai_n673_));
  NA3        m0645(.A(mai_mai_n524_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n674_));
  AN2        m0646(.A(h), .B(f), .Y(mai_mai_n675_));
  NA2        m0647(.A(mai_mai_n675_), .B(mai_mai_n37_), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n97_), .B(mai_mai_n46_), .Y(mai_mai_n677_));
  OAI220     m0649(.A0(mai_mai_n677_), .A1(mai_mai_n331_), .B0(mai_mai_n676_), .B1(mai_mai_n466_), .Y(mai_mai_n678_));
  AOI210     m0650(.A0(mai_mai_n571_), .A1(mai_mai_n427_), .B0(mai_mai_n49_), .Y(mai_mai_n679_));
  OAI220     m0651(.A0(mai_mai_n591_), .A1(mai_mai_n584_), .B0(mai_mai_n324_), .B1(mai_mai_n525_), .Y(mai_mai_n680_));
  AOI210     m0652(.A0(mai_mai_n680_), .A1(mai_mai_n679_), .B0(mai_mai_n678_), .Y(mai_mai_n681_));
  NA4        m0653(.A(mai_mai_n681_), .B(mai_mai_n674_), .C(mai_mai_n673_), .D(mai_mai_n670_), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n247_), .B(f), .Y(mai_mai_n683_));
  NO2        m0655(.A(mai_mai_n625_), .B(mai_mai_n61_), .Y(mai_mai_n684_));
  NO3        m0656(.A(mai_mai_n684_), .B(mai_mai_n683_), .C(mai_mai_n34_), .Y(mai_mai_n685_));
  NA2        m0657(.A(mai_mai_n327_), .B(mai_mai_n137_), .Y(mai_mai_n686_));
  NA2        m0658(.A(mai_mai_n130_), .B(mai_mai_n49_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n358_), .B(mai_mai_n111_), .Y(mai_mai_n688_));
  OA220      m0660(.A0(mai_mai_n688_), .A1(mai_mai_n552_), .B0(mai_mai_n356_), .B1(mai_mai_n109_), .Y(mai_mai_n689_));
  OAI210     m0661(.A0(mai_mai_n686_), .A1(mai_mai_n685_), .B0(mai_mai_n689_), .Y(mai_mai_n690_));
  NO3        m0662(.A(mai_mai_n402_), .B(mai_mai_n188_), .C(mai_mai_n187_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n691_), .B(mai_mai_n226_), .Y(mai_mai_n692_));
  NA3        m0664(.A(mai_mai_n692_), .B(mai_mai_n249_), .C(j), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n465_), .B(mai_mai_n83_), .Y(mai_mai_n694_));
  NA3        m0666(.A(mai_mai_n693_), .B(mai_mai_n512_), .C(mai_mai_n400_), .Y(mai_mai_n695_));
  NO4        m0667(.A(mai_mai_n695_), .B(mai_mai_n690_), .C(mai_mai_n682_), .D(mai_mai_n667_), .Y(mai_mai_n696_));
  NA4        m0668(.A(mai_mai_n696_), .B(mai_mai_n660_), .C(mai_mai_n614_), .D(mai_mai_n582_), .Y(mai08));
  NO2        m0669(.A(k), .B(h), .Y(mai_mai_n698_));
  AO210      m0670(.A0(mai_mai_n247_), .A1(mai_mai_n451_), .B0(mai_mai_n698_), .Y(mai_mai_n699_));
  NO2        m0671(.A(mai_mai_n699_), .B(mai_mai_n294_), .Y(mai_mai_n700_));
  NA2        m0672(.A(mai_mai_n624_), .B(mai_mai_n83_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n701_), .B(mai_mai_n461_), .Y(mai_mai_n702_));
  AOI210     m0674(.A0(mai_mai_n702_), .A1(mai_mai_n700_), .B0(mai_mai_n490_), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n83_), .B(mai_mai_n108_), .Y(mai_mai_n704_));
  NO2        m0676(.A(mai_mai_n704_), .B(mai_mai_n57_), .Y(mai_mai_n705_));
  NO4        m0677(.A(mai_mai_n376_), .B(mai_mai_n110_), .C(j), .D(mai_mai_n211_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n578_), .B(mai_mai_n228_), .Y(mai_mai_n707_));
  AOI220     m0679(.A0(mai_mai_n707_), .A1(mai_mai_n347_), .B0(mai_mai_n706_), .B1(mai_mai_n705_), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n578_), .A1(mai_mai_n150_), .B0(mai_mai_n83_), .Y(mai_mai_n709_));
  NA4        m0681(.A(mai_mai_n213_), .B(mai_mai_n137_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n710_));
  AN2        m0682(.A(l), .B(k), .Y(mai_mai_n711_));
  NA4        m0683(.A(mai_mai_n711_), .B(mai_mai_n106_), .C(mai_mai_n75_), .D(mai_mai_n211_), .Y(mai_mai_n712_));
  OAI210     m0684(.A0(mai_mai_n710_), .A1(g), .B0(mai_mai_n712_), .Y(mai_mai_n713_));
  NA2        m0685(.A(mai_mai_n713_), .B(mai_mai_n709_), .Y(mai_mai_n714_));
  NA3        m0686(.A(mai_mai_n714_), .B(mai_mai_n708_), .C(mai_mai_n703_), .Y(mai_mai_n715_));
  INV        m0687(.A(mai_mai_n519_), .Y(mai_mai_n716_));
  NO2        m0688(.A(mai_mai_n38_), .B(mai_mai_n210_), .Y(mai_mai_n717_));
  NA2        m0689(.A(mai_mai_n717_), .B(mai_mai_n568_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n716_), .Y(mai_mai_n719_));
  NO2        m0691(.A(mai_mai_n538_), .B(mai_mai_n35_), .Y(mai_mai_n720_));
  INV        m0692(.A(mai_mai_n720_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n699_), .B(mai_mai_n133_), .Y(mai_mai_n722_));
  NA2        m0694(.A(mai_mai_n722_), .B(mai_mai_n401_), .Y(mai_mai_n723_));
  OAI210     m0695(.A0(mai_mai_n721_), .A1(mai_mai_n86_), .B0(mai_mai_n723_), .Y(mai_mai_n724_));
  NA2        m0696(.A(mai_mai_n358_), .B(mai_mai_n43_), .Y(mai_mai_n725_));
  NA3        m0697(.A(mai_mai_n692_), .B(mai_mai_n333_), .C(mai_mai_n382_), .Y(mai_mai_n726_));
  NA2        m0698(.A(mai_mai_n711_), .B(mai_mai_n216_), .Y(mai_mai_n727_));
  NO2        m0699(.A(mai_mai_n727_), .B(mai_mai_n326_), .Y(mai_mai_n728_));
  AOI210     m0700(.A0(mai_mai_n728_), .A1(mai_mai_n683_), .B0(mai_mai_n489_), .Y(mai_mai_n729_));
  NA3        m0701(.A(m), .B(l), .C(k), .Y(mai_mai_n730_));
  AOI210     m0702(.A0(mai_mai_n664_), .A1(mai_mai_n662_), .B0(mai_mai_n730_), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n537_), .B(mai_mai_n268_), .Y(mai_mai_n732_));
  NOi21      m0704(.An(mai_mai_n732_), .B(mai_mai_n531_), .Y(mai_mai_n733_));
  NA4        m0705(.A(mai_mai_n111_), .B(l), .C(k), .D(mai_mai_n86_), .Y(mai_mai_n734_));
  NA3        m0706(.A(mai_mai_n119_), .B(mai_mai_n410_), .C(i), .Y(mai_mai_n735_));
  NO2        m0707(.A(mai_mai_n735_), .B(mai_mai_n734_), .Y(mai_mai_n736_));
  NO3        m0708(.A(mai_mai_n736_), .B(mai_mai_n733_), .C(mai_mai_n731_), .Y(mai_mai_n737_));
  NA4        m0709(.A(mai_mai_n737_), .B(mai_mai_n729_), .C(mai_mai_n726_), .D(mai_mai_n725_), .Y(mai_mai_n738_));
  NO4        m0710(.A(mai_mai_n738_), .B(mai_mai_n724_), .C(mai_mai_n719_), .D(mai_mai_n715_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n626_), .B(mai_mai_n391_), .Y(mai_mai_n740_));
  NOi31      m0712(.An(g), .B(h), .C(f), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n639_), .B(mai_mai_n741_), .Y(mai_mai_n742_));
  AO210      m0714(.A0(mai_mai_n742_), .A1(mai_mai_n592_), .B0(mai_mai_n540_), .Y(mai_mai_n743_));
  NO3        m0715(.A(mai_mai_n395_), .B(mai_mai_n525_), .C(h), .Y(mai_mai_n744_));
  NA2        m0716(.A(mai_mai_n744_), .B(mai_mai_n111_), .Y(mai_mai_n745_));
  NA4        m0717(.A(mai_mai_n745_), .B(mai_mai_n743_), .C(mai_mai_n740_), .D(mai_mai_n246_), .Y(mai_mai_n746_));
  NA2        m0718(.A(mai_mai_n711_), .B(mai_mai_n75_), .Y(mai_mai_n747_));
  NO4        m0719(.A(mai_mai_n691_), .B(mai_mai_n170_), .C(n), .D(i), .Y(mai_mai_n748_));
  NOi21      m0720(.An(h), .B(j), .Y(mai_mai_n749_));
  NA2        m0721(.A(mai_mai_n749_), .B(f), .Y(mai_mai_n750_));
  NO2        m0722(.A(mai_mai_n750_), .B(mai_mai_n243_), .Y(mai_mai_n751_));
  NO2        m0723(.A(mai_mai_n751_), .B(mai_mai_n748_), .Y(mai_mai_n752_));
  OAI220     m0724(.A0(mai_mai_n752_), .A1(mai_mai_n747_), .B0(mai_mai_n594_), .B1(mai_mai_n62_), .Y(mai_mai_n753_));
  AOI210     m0725(.A0(mai_mai_n746_), .A1(l), .B0(mai_mai_n753_), .Y(mai_mai_n754_));
  NO2        m0726(.A(j), .B(i), .Y(mai_mai_n755_));
  NA3        m0727(.A(mai_mai_n755_), .B(mai_mai_n81_), .C(l), .Y(mai_mai_n756_));
  NA2        m0728(.A(mai_mai_n755_), .B(mai_mai_n33_), .Y(mai_mai_n757_));
  NA2        m0729(.A(mai_mai_n420_), .B(mai_mai_n119_), .Y(mai_mai_n758_));
  OR2        m0730(.A(mai_mai_n758_), .B(mai_mai_n757_), .Y(mai_mai_n759_));
  NO3        m0731(.A(mai_mai_n146_), .B(mai_mai_n49_), .C(mai_mai_n108_), .Y(mai_mai_n760_));
  NO3        m0732(.A(mai_mai_n544_), .B(mai_mai_n144_), .C(mai_mai_n75_), .Y(mai_mai_n761_));
  NO3        m0733(.A(mai_mai_n485_), .B(mai_mai_n439_), .C(j), .Y(mai_mai_n762_));
  OAI210     m0734(.A0(mai_mai_n761_), .A1(mai_mai_n760_), .B0(mai_mai_n762_), .Y(mai_mai_n763_));
  OAI210     m0735(.A0(mai_mai_n742_), .A1(mai_mai_n62_), .B0(mai_mai_n763_), .Y(mai_mai_n764_));
  NA2        m0736(.A(k), .B(j), .Y(mai_mai_n765_));
  NO3        m0737(.A(mai_mai_n294_), .B(mai_mai_n765_), .C(mai_mai_n40_), .Y(mai_mai_n766_));
  AOI210     m0738(.A0(mai_mai_n530_), .A1(n), .B0(mai_mai_n554_), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n767_), .B(mai_mai_n557_), .Y(mai_mai_n768_));
  AN3        m0740(.A(mai_mai_n768_), .B(mai_mai_n766_), .C(mai_mai_n96_), .Y(mai_mai_n769_));
  NA2        m0741(.A(mai_mai_n617_), .B(mai_mai_n305_), .Y(mai_mai_n770_));
  INV        m0742(.A(mai_mai_n770_), .Y(mai_mai_n771_));
  NO2        m0743(.A(mai_mai_n294_), .B(mai_mai_n133_), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n772_), .B(mai_mai_n626_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n730_), .B(mai_mai_n89_), .Y(mai_mai_n774_));
  NA2        m0746(.A(mai_mai_n774_), .B(mai_mai_n589_), .Y(mai_mai_n775_));
  NO2        m0747(.A(mai_mai_n591_), .B(mai_mai_n115_), .Y(mai_mai_n776_));
  OAI210     m0748(.A0(mai_mai_n776_), .A1(mai_mai_n762_), .B0(mai_mai_n679_), .Y(mai_mai_n777_));
  NA3        m0749(.A(mai_mai_n777_), .B(mai_mai_n775_), .C(mai_mai_n773_), .Y(mai_mai_n778_));
  OR4        m0750(.A(mai_mai_n778_), .B(mai_mai_n771_), .C(mai_mai_n769_), .D(mai_mai_n764_), .Y(mai_mai_n779_));
  NA3        m0751(.A(mai_mai_n767_), .B(mai_mai_n557_), .C(mai_mai_n556_), .Y(mai_mai_n780_));
  NA4        m0752(.A(mai_mai_n780_), .B(mai_mai_n213_), .C(mai_mai_n451_), .D(mai_mai_n34_), .Y(mai_mai_n781_));
  OAI220     m0753(.A0(mai_mai_n710_), .A1(mai_mai_n701_), .B0(mai_mai_n331_), .B1(mai_mai_n38_), .Y(mai_mai_n782_));
  INV        m0754(.A(mai_mai_n782_), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n547_), .B(mai_mai_n287_), .C(h), .Y(mai_mai_n784_));
  NOi21      m0756(.An(mai_mai_n679_), .B(mai_mai_n784_), .Y(mai_mai_n785_));
  NO2        m0757(.A(mai_mai_n90_), .B(mai_mai_n47_), .Y(mai_mai_n786_));
  OAI220     m0758(.A0(mai_mai_n784_), .A1(mai_mai_n606_), .B0(mai_mai_n756_), .B1(mai_mai_n671_), .Y(mai_mai_n787_));
  AOI210     m0759(.A0(mai_mai_n786_), .A1(mai_mai_n645_), .B0(mai_mai_n787_), .Y(mai_mai_n788_));
  NAi41      m0760(.An(mai_mai_n785_), .B(mai_mai_n788_), .C(mai_mai_n783_), .D(mai_mai_n781_), .Y(mai_mai_n789_));
  OR2        m0761(.A(mai_mai_n774_), .B(mai_mai_n93_), .Y(mai_mai_n790_));
  AOI220     m0762(.A0(mai_mai_n790_), .A1(mai_mai_n234_), .B0(mai_mai_n762_), .B1(mai_mai_n638_), .Y(mai_mai_n791_));
  INV        m0763(.A(mai_mai_n335_), .Y(mai_mai_n792_));
  OAI210     m0764(.A0(mai_mai_n730_), .A1(mai_mai_n661_), .B0(mai_mai_n518_), .Y(mai_mai_n793_));
  AOI220     m0765(.A0(mai_mai_n605_), .A1(mai_mai_n29_), .B0(mai_mai_n465_), .B1(mai_mai_n83_), .Y(mai_mai_n794_));
  INV        m0766(.A(mai_mai_n794_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n784_), .B(mai_mai_n488_), .Y(mai_mai_n796_));
  AOI210     m0768(.A0(mai_mai_n795_), .A1(mai_mai_n793_), .B0(mai_mai_n796_), .Y(mai_mai_n797_));
  NA3        m0769(.A(mai_mai_n797_), .B(mai_mai_n792_), .C(mai_mai_n791_), .Y(mai_mai_n798_));
  NOi41      m0770(.An(mai_mai_n759_), .B(mai_mai_n798_), .C(mai_mai_n789_), .D(mai_mai_n779_), .Y(mai_mai_n799_));
  OR3        m0771(.A(mai_mai_n710_), .B(mai_mai_n228_), .C(g), .Y(mai_mai_n800_));
  NO3        m0772(.A(mai_mai_n341_), .B(mai_mai_n296_), .C(mai_mai_n110_), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n801_), .B(mai_mai_n768_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n803_));
  NO3        m0775(.A(mai_mai_n803_), .B(mai_mai_n757_), .C(mai_mai_n272_), .Y(mai_mai_n804_));
  NO3        m0776(.A(mai_mai_n525_), .B(mai_mai_n91_), .C(h), .Y(mai_mai_n805_));
  AOI210     m0777(.A0(mai_mai_n805_), .A1(mai_mai_n705_), .B0(mai_mai_n804_), .Y(mai_mai_n806_));
  NA4        m0778(.A(mai_mai_n806_), .B(mai_mai_n802_), .C(mai_mai_n800_), .D(mai_mai_n403_), .Y(mai_mai_n807_));
  OR2        m0779(.A(mai_mai_n661_), .B(mai_mai_n90_), .Y(mai_mai_n808_));
  NOi31      m0780(.An(b), .B(d), .C(a), .Y(mai_mai_n809_));
  NO2        m0781(.A(mai_mai_n809_), .B(mai_mai_n603_), .Y(mai_mai_n810_));
  NO2        m0782(.A(mai_mai_n810_), .B(n), .Y(mai_mai_n811_));
  NOi21      m0783(.An(mai_mai_n794_), .B(mai_mai_n811_), .Y(mai_mai_n812_));
  OAI220     m0784(.A0(mai_mai_n812_), .A1(mai_mai_n808_), .B0(mai_mai_n784_), .B1(mai_mai_n604_), .Y(mai_mai_n813_));
  NO2        m0785(.A(mai_mai_n555_), .B(mai_mai_n83_), .Y(mai_mai_n814_));
  NO3        m0786(.A(mai_mai_n625_), .B(mai_mai_n326_), .C(mai_mai_n115_), .Y(mai_mai_n815_));
  NOi21      m0787(.An(mai_mai_n815_), .B(mai_mai_n155_), .Y(mai_mai_n816_));
  AOI210     m0788(.A0(mai_mai_n801_), .A1(mai_mai_n814_), .B0(mai_mai_n816_), .Y(mai_mai_n817_));
  OAI210     m0789(.A0(mai_mai_n710_), .A1(mai_mai_n392_), .B0(mai_mai_n817_), .Y(mai_mai_n818_));
  NO2        m0790(.A(mai_mai_n691_), .B(n), .Y(mai_mai_n819_));
  AOI220     m0791(.A0(mai_mai_n772_), .A1(mai_mai_n668_), .B0(mai_mai_n819_), .B1(mai_mai_n700_), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n321_), .B(mai_mai_n233_), .Y(mai_mai_n821_));
  NA2        m0793(.A(mai_mai_n119_), .B(mai_mai_n83_), .Y(mai_mai_n822_));
  AOI210     m0794(.A0(mai_mai_n424_), .A1(mai_mai_n416_), .B0(mai_mai_n822_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n728_), .B(mai_mai_n34_), .Y(mai_mai_n824_));
  NAi21      m0796(.An(mai_mai_n734_), .B(mai_mai_n435_), .Y(mai_mai_n825_));
  NO2        m0797(.A(mai_mai_n268_), .B(i), .Y(mai_mai_n826_));
  NA2        m0798(.A(mai_mai_n596_), .B(mai_mai_n359_), .Y(mai_mai_n827_));
  AN2        m0799(.A(mai_mai_n827_), .B(mai_mai_n825_), .Y(mai_mai_n828_));
  NAi41      m0800(.An(mai_mai_n823_), .B(mai_mai_n828_), .C(mai_mai_n824_), .D(mai_mai_n820_), .Y(mai_mai_n829_));
  NO4        m0801(.A(mai_mai_n829_), .B(mai_mai_n818_), .C(mai_mai_n813_), .D(mai_mai_n807_), .Y(mai_mai_n830_));
  NA4        m0802(.A(mai_mai_n830_), .B(mai_mai_n799_), .C(mai_mai_n754_), .D(mai_mai_n739_), .Y(mai09));
  INV        m0803(.A(mai_mai_n120_), .Y(mai_mai_n832_));
  NA2        m0804(.A(f), .B(e), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n221_), .B(mai_mai_n110_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n834_), .B(g), .Y(mai_mai_n835_));
  NA4        m0807(.A(mai_mai_n307_), .B(mai_mai_n473_), .C(mai_mai_n256_), .D(mai_mai_n117_), .Y(mai_mai_n836_));
  AOI210     m0808(.A0(mai_mai_n836_), .A1(g), .B0(mai_mai_n470_), .Y(mai_mai_n837_));
  AOI210     m0809(.A0(mai_mai_n837_), .A1(mai_mai_n835_), .B0(mai_mai_n833_), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n445_), .B(e), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n839_), .B(mai_mai_n509_), .Y(mai_mai_n840_));
  AOI210     m0812(.A0(mai_mai_n838_), .A1(mai_mai_n832_), .B0(mai_mai_n840_), .Y(mai_mai_n841_));
  NO2        m0813(.A(mai_mai_n200_), .B(mai_mai_n210_), .Y(mai_mai_n842_));
  NA3        m0814(.A(m), .B(l), .C(i), .Y(mai_mai_n843_));
  OAI220     m0815(.A0(mai_mai_n591_), .A1(mai_mai_n843_), .B0(mai_mai_n351_), .B1(mai_mai_n526_), .Y(mai_mai_n844_));
  NA4        m0816(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(g), .D(f), .Y(mai_mai_n845_));
  NAi31      m0817(.An(mai_mai_n844_), .B(mai_mai_n845_), .C(mai_mai_n440_), .Y(mai_mai_n846_));
  OR2        m0818(.A(mai_mai_n846_), .B(mai_mai_n842_), .Y(mai_mai_n847_));
  NA3        m0819(.A(mai_mai_n808_), .B(mai_mai_n570_), .C(mai_mai_n518_), .Y(mai_mai_n848_));
  OA210      m0820(.A0(mai_mai_n848_), .A1(mai_mai_n847_), .B0(mai_mai_n811_), .Y(mai_mai_n849_));
  INV        m0821(.A(mai_mai_n338_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n851_));
  INV        m0823(.A(mai_mai_n340_), .Y(mai_mai_n852_));
  AOI210     m0824(.A0(mai_mai_n852_), .A1(mai_mai_n851_), .B0(mai_mai_n598_), .Y(mai_mai_n853_));
  INV        m0825(.A(mai_mai_n331_), .Y(mai_mai_n854_));
  NA2        m0826(.A(mai_mai_n342_), .B(mai_mai_n344_), .Y(mai_mai_n855_));
  OAI210     m0827(.A0(mai_mai_n200_), .A1(mai_mai_n210_), .B0(mai_mai_n855_), .Y(mai_mai_n856_));
  AOI220     m0828(.A0(mai_mai_n856_), .A1(mai_mai_n854_), .B0(mai_mai_n853_), .B1(mai_mai_n850_), .Y(mai_mai_n857_));
  NA2        m0829(.A(mai_mai_n164_), .B(mai_mai_n112_), .Y(mai_mai_n858_));
  NA3        m0830(.A(mai_mai_n858_), .B(mai_mai_n699_), .C(mai_mai_n133_), .Y(mai_mai_n859_));
  NA3        m0831(.A(mai_mai_n859_), .B(mai_mai_n185_), .C(mai_mai_n31_), .Y(mai_mai_n860_));
  NA3        m0832(.A(mai_mai_n860_), .B(mai_mai_n857_), .C(mai_mai_n627_), .Y(mai_mai_n861_));
  NO2        m0833(.A(mai_mai_n587_), .B(mai_mai_n496_), .Y(mai_mai_n862_));
  NOi21      m0834(.An(f), .B(d), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n863_), .B(m), .Y(mai_mai_n864_));
  NO2        m0836(.A(mai_mai_n864_), .B(mai_mai_n52_), .Y(mai_mai_n865_));
  NOi32      m0837(.An(g), .Bn(f), .C(d), .Y(mai_mai_n866_));
  NA4        m0838(.A(mai_mai_n866_), .B(mai_mai_n605_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n867_));
  NOi21      m0839(.An(mai_mai_n308_), .B(mai_mai_n867_), .Y(mai_mai_n868_));
  AOI210     m0840(.A0(mai_mai_n865_), .A1(mai_mai_n545_), .B0(mai_mai_n868_), .Y(mai_mai_n869_));
  NA2        m0841(.A(mai_mai_n256_), .B(mai_mai_n117_), .Y(mai_mai_n870_));
  AN2        m0842(.A(f), .B(d), .Y(mai_mai_n871_));
  NA3        m0843(.A(mai_mai_n478_), .B(mai_mai_n871_), .C(mai_mai_n83_), .Y(mai_mai_n872_));
  NO3        m0844(.A(mai_mai_n872_), .B(mai_mai_n75_), .C(mai_mai_n211_), .Y(mai_mai_n873_));
  NO2        m0845(.A(mai_mai_n280_), .B(mai_mai_n56_), .Y(mai_mai_n874_));
  NA2        m0846(.A(mai_mai_n870_), .B(mai_mai_n873_), .Y(mai_mai_n875_));
  NAi31      m0847(.An(mai_mai_n487_), .B(mai_mai_n875_), .C(mai_mai_n869_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n656_), .B(mai_mai_n326_), .Y(mai_mai_n877_));
  AN2        m0849(.A(mai_mai_n877_), .B(mai_mai_n683_), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n878_), .B(mai_mai_n230_), .Y(mai_mai_n879_));
  NA2        m0851(.A(mai_mai_n603_), .B(mai_mai_n83_), .Y(mai_mai_n880_));
  NO2        m0852(.A(mai_mai_n855_), .B(mai_mai_n880_), .Y(mai_mai_n881_));
  NA3        m0853(.A(mai_mai_n154_), .B(mai_mai_n106_), .C(mai_mai_n105_), .Y(mai_mai_n882_));
  OAI220     m0854(.A0(mai_mai_n872_), .A1(mai_mai_n429_), .B0(mai_mai_n338_), .B1(mai_mai_n882_), .Y(mai_mai_n883_));
  NOi41      m0855(.An(mai_mai_n219_), .B(mai_mai_n883_), .C(mai_mai_n881_), .D(mai_mai_n303_), .Y(mai_mai_n884_));
  NA2        m0856(.A(c), .B(mai_mai_n114_), .Y(mai_mai_n885_));
  NO2        m0857(.A(mai_mai_n885_), .B(mai_mai_n407_), .Y(mai_mai_n886_));
  NA3        m0858(.A(mai_mai_n886_), .B(mai_mai_n507_), .C(f), .Y(mai_mai_n887_));
  OR2        m0859(.A(mai_mai_n661_), .B(mai_mai_n541_), .Y(mai_mai_n888_));
  INV        m0860(.A(mai_mai_n888_), .Y(mai_mai_n889_));
  NA2        m0861(.A(mai_mai_n810_), .B(mai_mai_n109_), .Y(mai_mai_n890_));
  NA2        m0862(.A(mai_mai_n890_), .B(mai_mai_n889_), .Y(mai_mai_n891_));
  NA4        m0863(.A(mai_mai_n891_), .B(mai_mai_n887_), .C(mai_mai_n884_), .D(mai_mai_n879_), .Y(mai_mai_n892_));
  NO4        m0864(.A(mai_mai_n892_), .B(mai_mai_n876_), .C(mai_mai_n861_), .D(mai_mai_n849_), .Y(mai_mai_n893_));
  OR2        m0865(.A(mai_mai_n872_), .B(mai_mai_n75_), .Y(mai_mai_n894_));
  NA2        m0866(.A(mai_mai_n110_), .B(j), .Y(mai_mai_n895_));
  NA2        m0867(.A(mai_mai_n834_), .B(g), .Y(mai_mai_n896_));
  AOI210     m0868(.A0(mai_mai_n896_), .A1(mai_mai_n288_), .B0(mai_mai_n894_), .Y(mai_mai_n897_));
  NO2        m0869(.A(mai_mai_n331_), .B(mai_mai_n845_), .Y(mai_mai_n898_));
  NO2        m0870(.A(mai_mai_n226_), .B(mai_mai_n220_), .Y(mai_mai_n899_));
  NA2        m0871(.A(mai_mai_n899_), .B(mai_mai_n223_), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n429_), .B(mai_mai_n833_), .Y(mai_mai_n901_));
  NA2        m0873(.A(mai_mai_n901_), .B(mai_mai_n562_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n902_), .B(mai_mai_n900_), .Y(mai_mai_n903_));
  NA2        m0875(.A(e), .B(d), .Y(mai_mai_n904_));
  OAI220     m0876(.A0(mai_mai_n904_), .A1(c), .B0(mai_mai_n321_), .B1(d), .Y(mai_mai_n905_));
  NA3        m0877(.A(mai_mai_n905_), .B(mai_mai_n454_), .C(mai_mai_n505_), .Y(mai_mai_n906_));
  AOI210     m0878(.A0(mai_mai_n513_), .A1(mai_mai_n177_), .B0(mai_mai_n226_), .Y(mai_mai_n907_));
  INV        m0879(.A(mai_mai_n907_), .Y(mai_mai_n908_));
  NA2        m0880(.A(mai_mai_n280_), .B(mai_mai_n160_), .Y(mai_mai_n909_));
  NA2        m0881(.A(mai_mai_n873_), .B(mai_mai_n909_), .Y(mai_mai_n910_));
  NA3        m0882(.A(mai_mai_n163_), .B(mai_mai_n84_), .C(mai_mai_n34_), .Y(mai_mai_n911_));
  NA4        m0883(.A(mai_mai_n911_), .B(mai_mai_n910_), .C(mai_mai_n908_), .D(mai_mai_n906_), .Y(mai_mai_n912_));
  NO4        m0884(.A(mai_mai_n912_), .B(mai_mai_n903_), .C(mai_mai_n898_), .D(mai_mai_n897_), .Y(mai_mai_n913_));
  NA2        m0885(.A(mai_mai_n850_), .B(mai_mai_n31_), .Y(mai_mai_n914_));
  AO210      m0886(.A0(mai_mai_n914_), .A1(mai_mai_n701_), .B0(mai_mai_n214_), .Y(mai_mai_n915_));
  OAI220     m0887(.A0(mai_mai_n625_), .A1(mai_mai_n61_), .B0(mai_mai_n296_), .B1(j), .Y(mai_mai_n916_));
  AOI220     m0888(.A0(mai_mai_n916_), .A1(mai_mai_n877_), .B0(mai_mai_n615_), .B1(mai_mai_n624_), .Y(mai_mai_n917_));
  OAI210     m0889(.A0(mai_mai_n839_), .A1(mai_mai_n167_), .B0(mai_mai_n917_), .Y(mai_mai_n918_));
  OAI210     m0890(.A0(mai_mai_n834_), .A1(mai_mai_n909_), .B0(mai_mai_n866_), .Y(mai_mai_n919_));
  NO2        m0891(.A(mai_mai_n919_), .B(mai_mai_n606_), .Y(mai_mai_n920_));
  AOI210     m0892(.A0(mai_mai_n116_), .A1(mai_mai_n115_), .B0(mai_mai_n255_), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n921_), .B(mai_mai_n867_), .Y(mai_mai_n922_));
  AO210      m0894(.A0(mai_mai_n854_), .A1(mai_mai_n844_), .B0(mai_mai_n922_), .Y(mai_mai_n923_));
  NOi31      m0895(.An(mai_mai_n545_), .B(mai_mai_n864_), .C(mai_mai_n288_), .Y(mai_mai_n924_));
  NO4        m0896(.A(mai_mai_n924_), .B(mai_mai_n923_), .C(mai_mai_n920_), .D(mai_mai_n918_), .Y(mai_mai_n925_));
  AO220      m0897(.A0(mai_mai_n454_), .A1(mai_mai_n749_), .B0(mai_mai_n172_), .B1(f), .Y(mai_mai_n926_));
  OAI210     m0898(.A0(mai_mai_n926_), .A1(mai_mai_n457_), .B0(mai_mai_n905_), .Y(mai_mai_n927_));
  NO2        m0899(.A(mai_mai_n439_), .B(mai_mai_n71_), .Y(mai_mai_n928_));
  OAI210     m0900(.A0(mai_mai_n848_), .A1(mai_mai_n928_), .B0(mai_mai_n705_), .Y(mai_mai_n929_));
  AN4        m0901(.A(mai_mai_n929_), .B(mai_mai_n927_), .C(mai_mai_n925_), .D(mai_mai_n915_), .Y(mai_mai_n930_));
  NA4        m0902(.A(mai_mai_n930_), .B(mai_mai_n913_), .C(mai_mai_n893_), .D(mai_mai_n841_), .Y(mai12));
  NO2        m0903(.A(mai_mai_n452_), .B(c), .Y(mai_mai_n932_));
  NO4        m0904(.A(mai_mai_n444_), .B(mai_mai_n247_), .C(mai_mai_n583_), .D(mai_mai_n211_), .Y(mai_mai_n933_));
  NA2        m0905(.A(mai_mai_n933_), .B(mai_mai_n932_), .Y(mai_mai_n934_));
  NA2        m0906(.A(mai_mai_n545_), .B(mai_mai_n928_), .Y(mai_mai_n935_));
  NO2        m0907(.A(mai_mai_n452_), .B(mai_mai_n114_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n851_), .B(mai_mai_n351_), .Y(mai_mai_n937_));
  NO2        m0909(.A(mai_mai_n661_), .B(mai_mai_n376_), .Y(mai_mai_n938_));
  AOI220     m0910(.A0(mai_mai_n938_), .A1(mai_mai_n543_), .B0(mai_mai_n937_), .B1(mai_mai_n936_), .Y(mai_mai_n939_));
  NA4        m0911(.A(mai_mai_n939_), .B(mai_mai_n935_), .C(mai_mai_n934_), .D(mai_mai_n443_), .Y(mai_mai_n940_));
  AOI210     m0912(.A0(mai_mai_n229_), .A1(mai_mai_n337_), .B0(mai_mai_n197_), .Y(mai_mai_n941_));
  OR2        m0913(.A(mai_mai_n941_), .B(mai_mai_n933_), .Y(mai_mai_n942_));
  AOI210     m0914(.A0(mai_mai_n334_), .A1(mai_mai_n388_), .B0(mai_mai_n211_), .Y(mai_mai_n943_));
  OAI210     m0915(.A0(mai_mai_n943_), .A1(mai_mai_n942_), .B0(mai_mai_n402_), .Y(mai_mai_n944_));
  NO2        m0916(.A(mai_mai_n642_), .B(mai_mai_n258_), .Y(mai_mai_n945_));
  NO2        m0917(.A(mai_mai_n591_), .B(mai_mai_n843_), .Y(mai_mai_n946_));
  AOI220     m0918(.A0(mai_mai_n946_), .A1(mai_mai_n568_), .B0(mai_mai_n821_), .B1(mai_mai_n945_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n146_), .B(mai_mai_n233_), .Y(mai_mai_n948_));
  NA2        m0920(.A(mai_mai_n947_), .B(mai_mai_n944_), .Y(mai_mai_n949_));
  NA4        m0921(.A(mai_mai_n445_), .B(mai_mai_n437_), .C(mai_mai_n178_), .D(g), .Y(mai_mai_n950_));
  INV        m0922(.A(mai_mai_n950_), .Y(mai_mai_n951_));
  NO3        m0923(.A(mai_mai_n666_), .B(mai_mai_n90_), .C(mai_mai_n45_), .Y(mai_mai_n952_));
  NO4        m0924(.A(mai_mai_n952_), .B(mai_mai_n951_), .C(mai_mai_n949_), .D(mai_mai_n940_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n366_), .B(mai_mai_n365_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n588_), .B(mai_mai_n73_), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n555_), .B(mai_mai_n140_), .Y(mai_mai_n956_));
  NOi21      m0928(.An(mai_mai_n34_), .B(mai_mai_n656_), .Y(mai_mai_n957_));
  AOI220     m0929(.A0(mai_mai_n957_), .A1(mai_mai_n956_), .B0(mai_mai_n955_), .B1(mai_mai_n954_), .Y(mai_mai_n958_));
  OAI210     m0930(.A0(mai_mai_n246_), .A1(mai_mai_n45_), .B0(mai_mai_n958_), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n435_), .B(mai_mai_n260_), .Y(mai_mai_n960_));
  NO3        m0932(.A(mai_mai_n822_), .B(mai_mai_n88_), .C(mai_mai_n407_), .Y(mai_mai_n961_));
  NAi31      m0933(.An(mai_mai_n961_), .B(mai_mai_n960_), .C(mai_mai_n318_), .Y(mai_mai_n962_));
  NO2        m0934(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n502_), .B(mai_mai_n296_), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n964_), .B(mai_mai_n362_), .Y(mai_mai_n965_));
  NO2        m0937(.A(mai_mai_n965_), .B(mai_mai_n140_), .Y(mai_mai_n966_));
  NA2        m0938(.A(mai_mai_n634_), .B(mai_mai_n359_), .Y(mai_mai_n967_));
  OAI210     m0939(.A0(mai_mai_n735_), .A1(mai_mai_n967_), .B0(mai_mai_n363_), .Y(mai_mai_n968_));
  NO4        m0940(.A(mai_mai_n968_), .B(mai_mai_n966_), .C(mai_mai_n962_), .D(mai_mai_n959_), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n346_), .B(g), .Y(mai_mai_n970_));
  NA2        m0942(.A(mai_mai_n157_), .B(i), .Y(mai_mai_n971_));
  NA2        m0943(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n972_));
  OAI220     m0944(.A0(mai_mai_n972_), .A1(mai_mai_n196_), .B0(mai_mai_n971_), .B1(mai_mai_n90_), .Y(mai_mai_n973_));
  AOI210     m0945(.A0(mai_mai_n418_), .A1(mai_mai_n37_), .B0(mai_mai_n973_), .Y(mai_mai_n974_));
  NA2        m0946(.A(mai_mai_n555_), .B(mai_mai_n380_), .Y(mai_mai_n975_));
  AOI210     m0947(.A0(mai_mai_n975_), .A1(n), .B0(mai_mai_n554_), .Y(mai_mai_n976_));
  OAI220     m0948(.A0(mai_mai_n976_), .A1(mai_mai_n970_), .B0(mai_mai_n974_), .B1(mai_mai_n331_), .Y(mai_mai_n977_));
  NO2        m0949(.A(mai_mai_n661_), .B(mai_mai_n496_), .Y(mai_mai_n978_));
  NA3        m0950(.A(mai_mai_n342_), .B(mai_mai_n631_), .C(i), .Y(mai_mai_n979_));
  OAI210     m0951(.A0(mai_mai_n439_), .A1(mai_mai_n307_), .B0(mai_mai_n979_), .Y(mai_mai_n980_));
  OAI220     m0952(.A0(mai_mai_n980_), .A1(mai_mai_n978_), .B0(mai_mai_n679_), .B1(mai_mai_n761_), .Y(mai_mai_n981_));
  OR3        m0953(.A(mai_mai_n307_), .B(mai_mai_n434_), .C(f), .Y(mai_mai_n982_));
  NA3        m0954(.A(mai_mai_n323_), .B(mai_mai_n116_), .C(g), .Y(mai_mai_n983_));
  AOI210     m0955(.A0(mai_mai_n676_), .A1(mai_mai_n983_), .B0(m), .Y(mai_mai_n984_));
  OAI210     m0956(.A0(mai_mai_n984_), .A1(mai_mai_n937_), .B0(mai_mai_n322_), .Y(mai_mai_n985_));
  NA2        m0957(.A(mai_mai_n694_), .B(mai_mai_n880_), .Y(mai_mai_n986_));
  NA2        m0958(.A(mai_mai_n845_), .B(mai_mai_n440_), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n217_), .B(mai_mai_n78_), .Y(mai_mai_n988_));
  NA2        m0960(.A(mai_mai_n988_), .B(mai_mai_n982_), .Y(mai_mai_n989_));
  AOI220     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n253_), .B0(mai_mai_n987_), .B1(mai_mai_n986_), .Y(mai_mai_n990_));
  NA3        m0962(.A(mai_mai_n990_), .B(mai_mai_n985_), .C(mai_mai_n981_), .Y(mai_mai_n991_));
  NO2        m0963(.A(mai_mai_n376_), .B(mai_mai_n89_), .Y(mai_mai_n992_));
  NA2        m0964(.A(mai_mai_n992_), .B(mai_mai_n234_), .Y(mai_mai_n993_));
  NA2        m0965(.A(mai_mai_n665_), .B(mai_mai_n87_), .Y(mai_mai_n994_));
  NO2        m0966(.A(mai_mai_n460_), .B(mai_mai_n211_), .Y(mai_mai_n995_));
  NA2        m0967(.A(mai_mai_n995_), .B(mai_mai_n381_), .Y(mai_mai_n996_));
  NA3        m0968(.A(mai_mai_n996_), .B(mai_mai_n994_), .C(mai_mai_n993_), .Y(mai_mai_n997_));
  OAI210     m0969(.A0(mai_mai_n987_), .A1(mai_mai_n946_), .B0(mai_mai_n543_), .Y(mai_mai_n998_));
  AOI210     m0970(.A0(mai_mai_n419_), .A1(mai_mai_n411_), .B0(mai_mai_n822_), .Y(mai_mai_n999_));
  OAI210     m0971(.A0(mai_mai_n366_), .A1(mai_mai_n365_), .B0(mai_mai_n107_), .Y(mai_mai_n1000_));
  AOI210     m0972(.A0(mai_mai_n1000_), .A1(mai_mai_n535_), .B0(mai_mai_n999_), .Y(mai_mai_n1001_));
  NA2        m0973(.A(mai_mai_n984_), .B(mai_mai_n936_), .Y(mai_mai_n1002_));
  NO3        m0974(.A(mai_mai_n895_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n1003_));
  NA2        m0975(.A(mai_mai_n1003_), .B(mai_mai_n629_), .Y(mai_mai_n1004_));
  NA4        m0976(.A(mai_mai_n1004_), .B(mai_mai_n1002_), .C(mai_mai_n1001_), .D(mai_mai_n998_), .Y(mai_mai_n1005_));
  NO4        m0977(.A(mai_mai_n1005_), .B(mai_mai_n997_), .C(mai_mai_n991_), .D(mai_mai_n977_), .Y(mai_mai_n1006_));
  NAi31      m0978(.An(mai_mai_n138_), .B(mai_mai_n420_), .C(n), .Y(mai_mai_n1007_));
  NO2        m0979(.A(mai_mai_n124_), .B(mai_mai_n340_), .Y(mai_mai_n1008_));
  NO2        m0980(.A(mai_mai_n1008_), .B(mai_mai_n1007_), .Y(mai_mai_n1009_));
  NO3        m0981(.A(mai_mai_n268_), .B(mai_mai_n138_), .C(mai_mai_n407_), .Y(mai_mai_n1010_));
  AOI210     m0982(.A0(mai_mai_n1010_), .A1(mai_mai_n497_), .B0(mai_mai_n1009_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n490_), .B(i), .Y(mai_mai_n1012_));
  NA2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n226_), .B(mai_mai_n168_), .Y(mai_mai_n1014_));
  NO3        m0986(.A(mai_mai_n305_), .B(mai_mai_n445_), .C(mai_mai_n172_), .Y(mai_mai_n1015_));
  NOi31      m0987(.An(mai_mai_n1014_), .B(mai_mai_n1015_), .C(mai_mai_n211_), .Y(mai_mai_n1016_));
  NAi21      m0988(.An(mai_mai_n555_), .B(mai_mai_n995_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n438_), .B(mai_mai_n880_), .Y(mai_mai_n1018_));
  NO3        m0990(.A(mai_mai_n439_), .B(mai_mai_n307_), .C(mai_mai_n75_), .Y(mai_mai_n1019_));
  AOI220     m0991(.A0(mai_mai_n1019_), .A1(mai_mai_n1018_), .B0(mai_mai_n482_), .B1(g), .Y(mai_mai_n1020_));
  NA2        m0992(.A(mai_mai_n1020_), .B(mai_mai_n1017_), .Y(mai_mai_n1021_));
  OAI220     m0993(.A0(mai_mai_n1007_), .A1(mai_mai_n229_), .B0(mai_mai_n979_), .B1(mai_mai_n604_), .Y(mai_mai_n1022_));
  NO2        m0994(.A(mai_mai_n662_), .B(mai_mai_n376_), .Y(mai_mai_n1023_));
  NA2        m0995(.A(mai_mai_n941_), .B(mai_mai_n932_), .Y(mai_mai_n1024_));
  NO3        m0996(.A(mai_mai_n544_), .B(mai_mai_n144_), .C(mai_mai_n210_), .Y(mai_mai_n1025_));
  OAI210     m0997(.A0(mai_mai_n1025_), .A1(mai_mai_n524_), .B0(mai_mai_n377_), .Y(mai_mai_n1026_));
  OAI220     m0998(.A0(mai_mai_n938_), .A1(mai_mai_n946_), .B0(mai_mai_n545_), .B1(mai_mai_n428_), .Y(mai_mai_n1027_));
  NA4        m0999(.A(mai_mai_n1027_), .B(mai_mai_n1026_), .C(mai_mai_n1024_), .D(mai_mai_n623_), .Y(mai_mai_n1028_));
  OAI210     m1000(.A0(mai_mai_n941_), .A1(mai_mai_n933_), .B0(mai_mai_n1014_), .Y(mai_mai_n1029_));
  NA3        m1001(.A(mai_mai_n975_), .B(mai_mai_n486_), .C(mai_mai_n46_), .Y(mai_mai_n1030_));
  AOI210     m1002(.A0(mai_mai_n379_), .A1(mai_mai_n377_), .B0(mai_mai_n330_), .Y(mai_mai_n1031_));
  NA4        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1030_), .C(mai_mai_n1029_), .D(mai_mai_n269_), .Y(mai_mai_n1032_));
  OR4        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1028_), .C(mai_mai_n1023_), .D(mai_mai_n1022_), .Y(mai_mai_n1033_));
  NO4        m1005(.A(mai_mai_n1033_), .B(mai_mai_n1021_), .C(mai_mai_n1016_), .D(mai_mai_n1013_), .Y(mai_mai_n1034_));
  NA4        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1006_), .C(mai_mai_n969_), .D(mai_mai_n953_), .Y(mai13));
  AN2        m1007(.A(c), .B(b), .Y(mai_mai_n1036_));
  NA3        m1008(.A(mai_mai_n245_), .B(mai_mai_n1036_), .C(m), .Y(mai_mai_n1037_));
  NA2        m1009(.A(mai_mai_n495_), .B(f), .Y(mai_mai_n1038_));
  NO4        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1037_), .C(j), .D(mai_mai_n584_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n260_), .B(mai_mai_n1036_), .Y(mai_mai_n1040_));
  NO3        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1038_), .C(mai_mai_n971_), .Y(mai_mai_n1041_));
  NAi32      m1013(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n137_), .B(mai_mai_n45_), .Y(mai_mai_n1043_));
  NO4        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1042_), .C(mai_mai_n591_), .D(mai_mai_n304_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(h), .B(mai_mai_n220_), .Y(mai_mai_n1045_));
  NA2        m1017(.A(mai_mai_n410_), .B(mai_mai_n210_), .Y(mai_mai_n1046_));
  AN2        m1018(.A(d), .B(c), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n1047_), .B(mai_mai_n114_), .Y(mai_mai_n1048_));
  NO4        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1046_), .C(mai_mai_n173_), .D(mai_mai_n164_), .Y(mai_mai_n1049_));
  NA2        m1021(.A(mai_mai_n495_), .B(c), .Y(mai_mai_n1050_));
  NO4        m1022(.A(mai_mai_n1043_), .B(mai_mai_n587_), .C(mai_mai_n1050_), .D(mai_mai_n304_), .Y(mai_mai_n1051_));
  AO210      m1023(.A0(mai_mai_n1049_), .A1(mai_mai_n1045_), .B0(mai_mai_n1051_), .Y(mai_mai_n1052_));
  OR4        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1044_), .C(mai_mai_n1041_), .D(mai_mai_n1039_), .Y(mai_mai_n1053_));
  NAi32      m1025(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1054_));
  NO2        m1026(.A(mai_mai_n1054_), .B(mai_mai_n141_), .Y(mai_mai_n1055_));
  NA2        m1027(.A(mai_mai_n1055_), .B(g), .Y(mai_mai_n1056_));
  OR3        m1028(.A(mai_mai_n220_), .B(mai_mai_n173_), .C(mai_mai_n164_), .Y(mai_mai_n1057_));
  NO2        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1056_), .Y(mai_mai_n1058_));
  NO2        m1030(.A(mai_mai_n1050_), .B(mai_mai_n304_), .Y(mai_mai_n1059_));
  NO2        m1031(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1060_));
  NA2        m1032(.A(mai_mai_n633_), .B(mai_mai_n1060_), .Y(mai_mai_n1061_));
  NOi21      m1033(.An(mai_mai_n1059_), .B(mai_mai_n1061_), .Y(mai_mai_n1062_));
  NO2        m1034(.A(mai_mai_n765_), .B(mai_mai_n110_), .Y(mai_mai_n1063_));
  NOi41      m1035(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1064_));
  NA2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n1063_), .Y(mai_mai_n1065_));
  NO2        m1037(.A(mai_mai_n1065_), .B(mai_mai_n1056_), .Y(mai_mai_n1066_));
  OR3        m1038(.A(e), .B(d), .C(c), .Y(mai_mai_n1067_));
  NA3        m1039(.A(k), .B(j), .C(i), .Y(mai_mai_n1068_));
  NO3        m1040(.A(mai_mai_n1068_), .B(mai_mai_n304_), .C(mai_mai_n89_), .Y(mai_mai_n1069_));
  NOi21      m1041(.An(mai_mai_n1069_), .B(mai_mai_n1067_), .Y(mai_mai_n1070_));
  OR4        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1066_), .C(mai_mai_n1062_), .D(mai_mai_n1058_), .Y(mai_mai_n1071_));
  NA3        m1043(.A(mai_mai_n468_), .B(mai_mai_n333_), .C(mai_mai_n56_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(mai_mai_n1072_), .B(mai_mai_n1061_), .Y(mai_mai_n1073_));
  NO3        m1045(.A(mai_mai_n1072_), .B(mai_mai_n587_), .C(mai_mai_n451_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(f), .B(c), .Y(mai_mai_n1075_));
  NOi21      m1047(.An(mai_mai_n1075_), .B(mai_mai_n444_), .Y(mai_mai_n1076_));
  NA2        m1048(.A(mai_mai_n1076_), .B(mai_mai_n59_), .Y(mai_mai_n1077_));
  OR2        m1049(.A(k), .B(i), .Y(mai_mai_n1078_));
  NO3        m1050(.A(mai_mai_n1078_), .B(mai_mai_n240_), .C(l), .Y(mai_mai_n1079_));
  NOi31      m1051(.An(mai_mai_n1079_), .B(mai_mai_n1077_), .C(j), .Y(mai_mai_n1080_));
  OR3        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1074_), .C(mai_mai_n1073_), .Y(mai_mai_n1081_));
  OR3        m1053(.A(mai_mai_n1081_), .B(mai_mai_n1071_), .C(mai_mai_n1053_), .Y(mai02));
  OR2        m1054(.A(l), .B(k), .Y(mai_mai_n1083_));
  OR3        m1055(.A(h), .B(g), .C(f), .Y(mai_mai_n1084_));
  OR3        m1056(.A(n), .B(m), .C(i), .Y(mai_mai_n1085_));
  NO4        m1057(.A(mai_mai_n1085_), .B(mai_mai_n1084_), .C(mai_mai_n1083_), .D(mai_mai_n1067_), .Y(mai_mai_n1086_));
  NOi31      m1058(.An(e), .B(d), .C(c), .Y(mai_mai_n1087_));
  AOI210     m1059(.A0(mai_mai_n1069_), .A1(mai_mai_n1087_), .B0(mai_mai_n1044_), .Y(mai_mai_n1088_));
  AN3        m1060(.A(g), .B(f), .C(c), .Y(mai_mai_n1089_));
  NA2        m1061(.A(mai_mai_n1089_), .B(mai_mai_n468_), .Y(mai_mai_n1090_));
  OR2        m1062(.A(mai_mai_n1068_), .B(mai_mai_n304_), .Y(mai_mai_n1091_));
  OR2        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1090_), .Y(mai_mai_n1092_));
  NO3        m1064(.A(mai_mai_n1072_), .B(mai_mai_n1043_), .C(mai_mai_n587_), .Y(mai_mai_n1093_));
  NO2        m1065(.A(mai_mai_n1093_), .B(mai_mai_n1058_), .Y(mai_mai_n1094_));
  NA3        m1066(.A(l), .B(k), .C(j), .Y(mai_mai_n1095_));
  NA2        m1067(.A(i), .B(h), .Y(mai_mai_n1096_));
  NO3        m1068(.A(mai_mai_n1096_), .B(mai_mai_n1095_), .C(mai_mai_n130_), .Y(mai_mai_n1097_));
  NO3        m1069(.A(mai_mai_n139_), .B(mai_mai_n278_), .C(mai_mai_n211_), .Y(mai_mai_n1098_));
  AOI210     m1070(.A0(mai_mai_n1098_), .A1(mai_mai_n1097_), .B0(mai_mai_n1062_), .Y(mai_mai_n1099_));
  NA3        m1071(.A(c), .B(b), .C(a), .Y(mai_mai_n1100_));
  NO3        m1072(.A(mai_mai_n1100_), .B(mai_mai_n904_), .C(mai_mai_n210_), .Y(mai_mai_n1101_));
  NO3        m1073(.A(mai_mai_n296_), .B(mai_mai_n49_), .C(mai_mai_n110_), .Y(mai_mai_n1102_));
  AOI210     m1074(.A0(mai_mai_n1102_), .A1(mai_mai_n1101_), .B0(mai_mai_n1073_), .Y(mai_mai_n1103_));
  AN4        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1099_), .C(mai_mai_n1094_), .D(mai_mai_n1092_), .Y(mai_mai_n1104_));
  NO2        m1076(.A(mai_mai_n1048_), .B(mai_mai_n1046_), .Y(mai_mai_n1105_));
  NA2        m1077(.A(mai_mai_n1065_), .B(mai_mai_n1057_), .Y(mai_mai_n1106_));
  AOI210     m1078(.A0(mai_mai_n1106_), .A1(mai_mai_n1105_), .B0(mai_mai_n1039_), .Y(mai_mai_n1107_));
  NAi41      m1079(.An(mai_mai_n1086_), .B(mai_mai_n1107_), .C(mai_mai_n1104_), .D(mai_mai_n1088_), .Y(mai03));
  INV        m1080(.A(mai_mai_n1000_), .Y(mai_mai_n1109_));
  NO2        m1081(.A(mai_mai_n856_), .B(mai_mai_n846_), .Y(mai_mai_n1110_));
  OAI220     m1082(.A0(mai_mai_n1110_), .A1(mai_mai_n694_), .B0(mai_mai_n1109_), .B1(mai_mai_n588_), .Y(mai_mai_n1111_));
  NOi31      m1083(.An(i), .B(k), .C(j), .Y(mai_mai_n1112_));
  NA4        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1087_), .C(mai_mai_n342_), .D(mai_mai_n333_), .Y(mai_mai_n1113_));
  OAI210     m1085(.A0(mai_mai_n822_), .A1(mai_mai_n421_), .B0(mai_mai_n1113_), .Y(mai_mai_n1114_));
  NOi31      m1086(.An(m), .B(n), .C(f), .Y(mai_mai_n1115_));
  NA2        m1087(.A(mai_mai_n1115_), .B(mai_mai_n51_), .Y(mai_mai_n1116_));
  AN2        m1088(.A(e), .B(c), .Y(mai_mai_n1117_));
  NA2        m1089(.A(mai_mai_n1117_), .B(a), .Y(mai_mai_n1118_));
  OAI220     m1090(.A0(mai_mai_n1118_), .A1(mai_mai_n1116_), .B0(mai_mai_n888_), .B1(mai_mai_n427_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n505_), .B(l), .Y(mai_mai_n1120_));
  NOi31      m1092(.An(mai_mai_n866_), .B(mai_mai_n1037_), .C(mai_mai_n1120_), .Y(mai_mai_n1121_));
  NO4        m1093(.A(mai_mai_n1121_), .B(mai_mai_n1119_), .C(mai_mai_n1114_), .D(mai_mai_n999_), .Y(mai_mai_n1122_));
  NO2        m1094(.A(mai_mai_n278_), .B(a), .Y(mai_mai_n1123_));
  INV        m1095(.A(mai_mai_n1044_), .Y(mai_mai_n1124_));
  NO2        m1096(.A(mai_mai_n1096_), .B(mai_mai_n485_), .Y(mai_mai_n1125_));
  NO2        m1097(.A(mai_mai_n86_), .B(g), .Y(mai_mai_n1126_));
  AOI210     m1098(.A0(mai_mai_n1126_), .A1(mai_mai_n1125_), .B0(mai_mai_n1079_), .Y(mai_mai_n1127_));
  OR2        m1099(.A(mai_mai_n1127_), .B(mai_mai_n1077_), .Y(mai_mai_n1128_));
  NA3        m1100(.A(mai_mai_n1128_), .B(mai_mai_n1124_), .C(mai_mai_n1122_), .Y(mai_mai_n1129_));
  NO4        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1111_), .C(mai_mai_n823_), .D(mai_mai_n567_), .Y(mai_mai_n1130_));
  NA2        m1102(.A(c), .B(b), .Y(mai_mai_n1131_));
  NO2        m1103(.A(mai_mai_n704_), .B(mai_mai_n1131_), .Y(mai_mai_n1132_));
  OAI210     m1104(.A0(mai_mai_n864_), .A1(mai_mai_n837_), .B0(mai_mai_n414_), .Y(mai_mai_n1133_));
  OAI210     m1105(.A0(mai_mai_n1133_), .A1(mai_mai_n865_), .B0(mai_mai_n1132_), .Y(mai_mai_n1134_));
  NAi21      m1106(.An(mai_mai_n422_), .B(mai_mai_n1132_), .Y(mai_mai_n1135_));
  NA3        m1107(.A(mai_mai_n428_), .B(mai_mai_n560_), .C(f), .Y(mai_mai_n1136_));
  OAI210     m1108(.A0(mai_mai_n549_), .A1(mai_mai_n39_), .B0(mai_mai_n1123_), .Y(mai_mai_n1137_));
  NA3        m1109(.A(mai_mai_n1137_), .B(mai_mai_n1136_), .C(mai_mai_n1135_), .Y(mai_mai_n1138_));
  NA2        m1110(.A(mai_mai_n256_), .B(mai_mai_n117_), .Y(mai_mai_n1139_));
  OAI210     m1111(.A0(mai_mai_n1139_), .A1(mai_mai_n282_), .B0(g), .Y(mai_mai_n1140_));
  NAi21      m1112(.An(f), .B(d), .Y(mai_mai_n1141_));
  NO2        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1100_), .Y(mai_mai_n1142_));
  INV        m1114(.A(mai_mai_n1142_), .Y(mai_mai_n1143_));
  AOI210     m1115(.A0(mai_mai_n1140_), .A1(mai_mai_n288_), .B0(mai_mai_n1143_), .Y(mai_mai_n1144_));
  AOI210     m1116(.A0(mai_mai_n1144_), .A1(mai_mai_n111_), .B0(mai_mai_n1138_), .Y(mai_mai_n1145_));
  NA2        m1117(.A(mai_mai_n470_), .B(f), .Y(mai_mai_n1146_));
  NO2        m1118(.A(mai_mai_n179_), .B(mai_mai_n233_), .Y(mai_mai_n1147_));
  NA2        m1119(.A(mai_mai_n1147_), .B(m), .Y(mai_mai_n1148_));
  NA3        m1120(.A(mai_mai_n921_), .B(mai_mai_n1120_), .C(mai_mai_n473_), .Y(mai_mai_n1149_));
  OAI210     m1121(.A0(mai_mai_n1149_), .A1(mai_mai_n308_), .B0(mai_mai_n471_), .Y(mai_mai_n1150_));
  AOI210     m1122(.A0(mai_mai_n1150_), .A1(mai_mai_n1146_), .B0(mai_mai_n1148_), .Y(mai_mai_n1151_));
  NA2        m1123(.A(mai_mai_n562_), .B(mai_mai_n409_), .Y(mai_mai_n1152_));
  NA2        m1124(.A(mai_mai_n153_), .B(mai_mai_n33_), .Y(mai_mai_n1153_));
  AOI210     m1125(.A0(mai_mai_n967_), .A1(mai_mai_n1153_), .B0(mai_mai_n211_), .Y(mai_mai_n1154_));
  OAI210     m1126(.A0(mai_mai_n1154_), .A1(mai_mai_n448_), .B0(mai_mai_n1142_), .Y(mai_mai_n1155_));
  NO2        m1127(.A(mai_mai_n370_), .B(mai_mai_n369_), .Y(mai_mai_n1156_));
  AOI210     m1128(.A0(mai_mai_n1147_), .A1(mai_mai_n430_), .B0(mai_mai_n961_), .Y(mai_mai_n1157_));
  NAi41      m1129(.An(mai_mai_n1156_), .B(mai_mai_n1157_), .C(mai_mai_n1155_), .D(mai_mai_n1152_), .Y(mai_mai_n1158_));
  NO2        m1130(.A(mai_mai_n1158_), .B(mai_mai_n1151_), .Y(mai_mai_n1159_));
  NA4        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1145_), .C(mai_mai_n1134_), .D(mai_mai_n1130_), .Y(mai00));
  AOI210     m1132(.A0(mai_mai_n295_), .A1(mai_mai_n211_), .B0(mai_mai_n271_), .Y(mai_mai_n1161_));
  NO2        m1133(.A(mai_mai_n1161_), .B(mai_mai_n578_), .Y(mai_mai_n1162_));
  AOI210     m1134(.A0(mai_mai_n901_), .A1(mai_mai_n948_), .B0(mai_mai_n1114_), .Y(mai_mai_n1163_));
  NO2        m1135(.A(mai_mai_n1093_), .B(mai_mai_n961_), .Y(mai_mai_n1164_));
  NA3        m1136(.A(mai_mai_n1164_), .B(mai_mai_n1163_), .C(mai_mai_n1001_), .Y(mai_mai_n1165_));
  NA2        m1137(.A(mai_mai_n507_), .B(f), .Y(mai_mai_n1166_));
  OAI210     m1138(.A0(mai_mai_n1008_), .A1(mai_mai_n40_), .B0(mai_mai_n649_), .Y(mai_mai_n1167_));
  NA3        m1139(.A(mai_mai_n1167_), .B(mai_mai_n252_), .C(n), .Y(mai_mai_n1168_));
  AOI210     m1140(.A0(mai_mai_n1168_), .A1(mai_mai_n1166_), .B0(mai_mai_n1048_), .Y(mai_mai_n1169_));
  NO4        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1165_), .C(mai_mai_n1162_), .D(mai_mai_n1071_), .Y(mai_mai_n1170_));
  NA2        m1142(.A(mai_mai_n163_), .B(mai_mai_n46_), .Y(mai_mai_n1171_));
  NA3        m1143(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1172_));
  NOi31      m1144(.An(n), .B(m), .C(i), .Y(mai_mai_n1173_));
  NA3        m1145(.A(mai_mai_n1173_), .B(mai_mai_n652_), .C(mai_mai_n51_), .Y(mai_mai_n1174_));
  OAI210     m1146(.A0(mai_mai_n1172_), .A1(mai_mai_n1171_), .B0(mai_mai_n1174_), .Y(mai_mai_n1175_));
  INV        m1147(.A(mai_mai_n577_), .Y(mai_mai_n1176_));
  NO4        m1148(.A(mai_mai_n1176_), .B(mai_mai_n1175_), .C(mai_mai_n1156_), .D(mai_mai_n924_), .Y(mai_mai_n1177_));
  OR2        m1149(.A(mai_mai_n383_), .B(mai_mai_n132_), .Y(mai_mai_n1178_));
  NO2        m1150(.A(h), .B(g), .Y(mai_mai_n1179_));
  INV        m1151(.A(mai_mai_n1178_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n1180_), .B(mai_mai_n262_), .Y(mai_mai_n1181_));
  INV        m1153(.A(mai_mai_n320_), .Y(mai_mai_n1182_));
  INV        m1154(.A(mai_mai_n579_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n1183_), .B(mai_mai_n1182_), .Y(mai_mai_n1184_));
  NO2        m1156(.A(mai_mai_n235_), .B(mai_mai_n178_), .Y(mai_mai_n1185_));
  NA2        m1157(.A(mai_mai_n1185_), .B(mai_mai_n428_), .Y(mai_mai_n1186_));
  NA3        m1158(.A(mai_mai_n176_), .B(mai_mai_n110_), .C(g), .Y(mai_mai_n1187_));
  NA2        m1159(.A(mai_mai_n468_), .B(f), .Y(mai_mai_n1188_));
  NOi31      m1160(.An(mai_mai_n874_), .B(mai_mai_n1188_), .C(mai_mai_n1187_), .Y(mai_mai_n1189_));
  NAi31      m1161(.An(mai_mai_n181_), .B(mai_mai_n862_), .C(mai_mai_n468_), .Y(mai_mai_n1190_));
  NAi31      m1162(.An(mai_mai_n1189_), .B(mai_mai_n1190_), .C(mai_mai_n1186_), .Y(mai_mai_n1191_));
  NO2        m1163(.A(mai_mai_n270_), .B(mai_mai_n75_), .Y(mai_mai_n1192_));
  NO3        m1164(.A(mai_mai_n427_), .B(mai_mai_n833_), .C(n), .Y(mai_mai_n1193_));
  AOI210     m1165(.A0(mai_mai_n1193_), .A1(mai_mai_n1192_), .B0(mai_mai_n1086_), .Y(mai_mai_n1194_));
  NAi31      m1166(.An(mai_mai_n1051_), .B(mai_mai_n1194_), .C(mai_mai_n74_), .Y(mai_mai_n1195_));
  NO4        m1167(.A(mai_mai_n1195_), .B(mai_mai_n1191_), .C(mai_mai_n1184_), .D(mai_mai_n517_), .Y(mai_mai_n1196_));
  AN3        m1168(.A(mai_mai_n1196_), .B(mai_mai_n1181_), .C(mai_mai_n1177_), .Y(mai_mai_n1197_));
  NA2        m1169(.A(mai_mai_n535_), .B(mai_mai_n99_), .Y(mai_mai_n1198_));
  NA3        m1170(.A(mai_mai_n1115_), .B(mai_mai_n609_), .C(mai_mai_n467_), .Y(mai_mai_n1199_));
  NA4        m1171(.A(mai_mai_n1199_), .B(mai_mai_n563_), .C(mai_mai_n1198_), .D(mai_mai_n238_), .Y(mai_mai_n1200_));
  OAI210     m1172(.A0(mai_mai_n466_), .A1(mai_mai_n118_), .B0(mai_mai_n867_), .Y(mai_mai_n1201_));
  AOI220     m1173(.A0(mai_mai_n1201_), .A1(mai_mai_n1149_), .B0(mai_mai_n562_), .B1(mai_mai_n409_), .Y(mai_mai_n1202_));
  OR4        m1174(.A(mai_mai_n1048_), .B(mai_mai_n268_), .C(mai_mai_n218_), .D(e), .Y(mai_mai_n1203_));
  NA2        m1175(.A(n), .B(e), .Y(mai_mai_n1204_));
  NO2        m1176(.A(mai_mai_n1204_), .B(mai_mai_n141_), .Y(mai_mai_n1205_));
  NA2        m1177(.A(mai_mai_n1203_), .B(mai_mai_n1202_), .Y(mai_mai_n1206_));
  AOI210     m1178(.A0(mai_mai_n1205_), .A1(mai_mai_n853_), .B0(mai_mai_n823_), .Y(mai_mai_n1207_));
  AOI220     m1179(.A0(mai_mai_n957_), .A1(mai_mai_n576_), .B0(mai_mai_n652_), .B1(mai_mai_n241_), .Y(mai_mai_n1208_));
  NO2        m1180(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1209_));
  NO3        m1181(.A(mai_mai_n1048_), .B(mai_mai_n1046_), .C(mai_mai_n727_), .Y(mai_mai_n1210_));
  NO2        m1182(.A(mai_mai_n1083_), .B(mai_mai_n130_), .Y(mai_mai_n1211_));
  AN2        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1098_), .Y(mai_mai_n1212_));
  OAI210     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n1210_), .B0(mai_mai_n1209_), .Y(mai_mai_n1213_));
  NA4        m1185(.A(mai_mai_n1213_), .B(mai_mai_n1208_), .C(mai_mai_n1207_), .D(mai_mai_n869_), .Y(mai_mai_n1214_));
  NO4        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1206_), .C(mai_mai_n291_), .D(mai_mai_n1200_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n838_), .B(mai_mai_n760_), .Y(mai_mai_n1216_));
  NA4        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1215_), .C(mai_mai_n1197_), .D(mai_mai_n1170_), .Y(mai01));
  AN2        m1189(.A(mai_mai_n1026_), .B(mai_mai_n1024_), .Y(mai_mai_n1218_));
  NO3        m1190(.A(mai_mai_n804_), .B(mai_mai_n796_), .C(mai_mai_n276_), .Y(mai_mai_n1219_));
  NA2        m1191(.A(mai_mai_n393_), .B(i), .Y(mai_mai_n1220_));
  NA3        m1192(.A(mai_mai_n1220_), .B(mai_mai_n1219_), .C(mai_mai_n1218_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n555_), .B(mai_mai_n267_), .Y(mai_mai_n1222_));
  NA2        m1194(.A(mai_mai_n964_), .B(mai_mai_n1222_), .Y(mai_mai_n1223_));
  NA3        m1195(.A(mai_mai_n1223_), .B(mai_mai_n917_), .C(mai_mai_n332_), .Y(mai_mai_n1224_));
  NA2        m1196(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1225_));
  NA2        m1197(.A(mai_mai_n711_), .B(mai_mai_n94_), .Y(mai_mai_n1226_));
  NO2        m1198(.A(mai_mai_n1226_), .B(mai_mai_n1225_), .Y(mai_mai_n1227_));
  NO2        m1199(.A(mai_mai_n784_), .B(mai_mai_n604_), .Y(mai_mai_n1228_));
  AOI210     m1200(.A0(mai_mai_n1227_), .A1(mai_mai_n638_), .B0(mai_mai_n1228_), .Y(mai_mai_n1229_));
  INV        m1201(.A(mai_mai_n116_), .Y(mai_mai_n1230_));
  OR2        m1202(.A(mai_mai_n1230_), .B(mai_mai_n586_), .Y(mai_mai_n1231_));
  NAi41      m1203(.An(mai_mai_n156_), .B(mai_mai_n1231_), .C(mai_mai_n1229_), .D(mai_mai_n900_), .Y(mai_mai_n1232_));
  NO3        m1204(.A(mai_mai_n785_), .B(mai_mai_n678_), .C(mai_mai_n510_), .Y(mai_mai_n1233_));
  OR2        m1205(.A(mai_mai_n191_), .B(mai_mai_n189_), .Y(mai_mai_n1234_));
  NA3        m1206(.A(mai_mai_n1234_), .B(mai_mai_n1233_), .C(mai_mai_n135_), .Y(mai_mai_n1235_));
  NO4        m1207(.A(mai_mai_n1235_), .B(mai_mai_n1232_), .C(mai_mai_n1224_), .D(mai_mai_n1221_), .Y(mai_mai_n1236_));
  INV        m1208(.A(mai_mai_n203_), .Y(mai_mai_n1237_));
  OAI210     m1209(.A0(mai_mai_n1237_), .A1(mai_mai_n298_), .B0(mai_mai_n530_), .Y(mai_mai_n1238_));
  NA2        m1210(.A(mai_mai_n538_), .B(mai_mai_n395_), .Y(mai_mai_n1239_));
  NOi21      m1211(.An(mai_mai_n564_), .B(mai_mai_n583_), .Y(mai_mai_n1240_));
  NA2        m1212(.A(mai_mai_n1240_), .B(mai_mai_n1239_), .Y(mai_mai_n1241_));
  AOI210     m1213(.A0(mai_mai_n200_), .A1(mai_mai_n88_), .B0(mai_mai_n210_), .Y(mai_mai_n1242_));
  OAI210     m1214(.A0(mai_mai_n811_), .A1(mai_mai_n428_), .B0(mai_mai_n1242_), .Y(mai_mai_n1243_));
  AN3        m1215(.A(m), .B(l), .C(k), .Y(mai_mai_n1244_));
  OAI210     m1216(.A0(mai_mai_n355_), .A1(mai_mai_n34_), .B0(mai_mai_n1244_), .Y(mai_mai_n1245_));
  NA2        m1217(.A(mai_mai_n199_), .B(mai_mai_n34_), .Y(mai_mai_n1246_));
  AO210      m1218(.A0(mai_mai_n1246_), .A1(mai_mai_n1245_), .B0(mai_mai_n331_), .Y(mai_mai_n1247_));
  NA4        m1219(.A(mai_mai_n1247_), .B(mai_mai_n1243_), .C(mai_mai_n1241_), .D(mai_mai_n1238_), .Y(mai_mai_n1248_));
  AOI210     m1220(.A0(mai_mai_n596_), .A1(mai_mai_n116_), .B0(mai_mai_n602_), .Y(mai_mai_n1249_));
  OAI210     m1221(.A0(mai_mai_n1230_), .A1(mai_mai_n595_), .B0(mai_mai_n1249_), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n275_), .B(mai_mai_n191_), .Y(mai_mai_n1251_));
  NA2        m1223(.A(mai_mai_n1251_), .B(mai_mai_n668_), .Y(mai_mai_n1252_));
  NO3        m1224(.A(mai_mai_n822_), .B(mai_mai_n200_), .C(mai_mai_n407_), .Y(mai_mai_n1253_));
  NO2        m1225(.A(mai_mai_n1253_), .B(mai_mai_n961_), .Y(mai_mai_n1254_));
  OAI210     m1226(.A0(mai_mai_n1227_), .A1(mai_mai_n325_), .B0(mai_mai_n679_), .Y(mai_mai_n1255_));
  NA4        m1227(.A(mai_mai_n1255_), .B(mai_mai_n1254_), .C(mai_mai_n1252_), .D(mai_mai_n788_), .Y(mai_mai_n1256_));
  NO3        m1228(.A(mai_mai_n1256_), .B(mai_mai_n1250_), .C(mai_mai_n1248_), .Y(mai_mai_n1257_));
  NA3        m1229(.A(mai_mai_n605_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1258_));
  NO2        m1230(.A(mai_mai_n1258_), .B(mai_mai_n200_), .Y(mai_mai_n1259_));
  AOI210     m1231(.A0(mai_mai_n503_), .A1(mai_mai_n58_), .B0(mai_mai_n1259_), .Y(mai_mai_n1260_));
  OR3        m1232(.A(mai_mai_n1226_), .B(mai_mai_n606_), .C(mai_mai_n1225_), .Y(mai_mai_n1261_));
  INV        m1233(.A(mai_mai_n1175_), .Y(mai_mai_n1262_));
  NA4        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1261_), .C(mai_mai_n1260_), .D(mai_mai_n759_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n971_), .B(mai_mai_n228_), .Y(mai_mai_n1264_));
  NO2        m1236(.A(mai_mai_n972_), .B(mai_mai_n557_), .Y(mai_mai_n1265_));
  OAI210     m1237(.A0(mai_mai_n1265_), .A1(mai_mai_n1264_), .B0(mai_mai_n340_), .Y(mai_mai_n1266_));
  NO3        m1238(.A(mai_mai_n80_), .B(mai_mai_n296_), .C(mai_mai_n45_), .Y(mai_mai_n1267_));
  NA2        m1239(.A(mai_mai_n1267_), .B(mai_mai_n554_), .Y(mai_mai_n1268_));
  NA2        m1240(.A(mai_mai_n1268_), .B(mai_mai_n673_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n367_), .B(mai_mai_n73_), .Y(mai_mai_n1270_));
  INV        m1242(.A(mai_mai_n1270_), .Y(mai_mai_n1271_));
  NA2        m1243(.A(mai_mai_n1267_), .B(mai_mai_n814_), .Y(mai_mai_n1272_));
  NA3        m1244(.A(mai_mai_n1272_), .B(mai_mai_n1271_), .C(mai_mai_n385_), .Y(mai_mai_n1273_));
  NOi41      m1245(.An(mai_mai_n1266_), .B(mai_mai_n1273_), .C(mai_mai_n1269_), .D(mai_mai_n1263_), .Y(mai_mai_n1274_));
  NO2        m1246(.A(mai_mai_n129_), .B(mai_mai_n45_), .Y(mai_mai_n1275_));
  NO2        m1247(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1276_));
  AO220      m1248(.A0(mai_mai_n1276_), .A1(mai_mai_n626_), .B0(mai_mai_n1275_), .B1(mai_mai_n709_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n1277_), .B(mai_mai_n340_), .Y(mai_mai_n1278_));
  NO3        m1250(.A(mai_mai_n1096_), .B(mai_mai_n173_), .C(mai_mai_n86_), .Y(mai_mai_n1279_));
  INV        m1251(.A(mai_mai_n1278_), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n617_), .B(mai_mai_n616_), .Y(mai_mai_n1281_));
  NO4        m1253(.A(mai_mai_n1096_), .B(mai_mai_n1281_), .C(mai_mai_n171_), .D(mai_mai_n86_), .Y(mai_mai_n1282_));
  NO3        m1254(.A(mai_mai_n1282_), .B(mai_mai_n1280_), .C(mai_mai_n641_), .Y(mai_mai_n1283_));
  NA4        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1274_), .C(mai_mai_n1257_), .D(mai_mai_n1236_), .Y(mai06));
  NO2        m1256(.A(mai_mai_n408_), .B(mai_mai_n561_), .Y(mai_mai_n1285_));
  INV        m1257(.A(mai_mai_n734_), .Y(mai_mai_n1286_));
  OAI210     m1258(.A0(mai_mai_n1286_), .A1(mai_mai_n263_), .B0(mai_mai_n1285_), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n220_), .B(mai_mai_n100_), .Y(mai_mai_n1288_));
  OAI210     m1260(.A0(mai_mai_n1288_), .A1(mai_mai_n1279_), .B0(mai_mai_n381_), .Y(mai_mai_n1289_));
  NO3        m1261(.A(mai_mai_n600_), .B(mai_mai_n809_), .C(mai_mai_n603_), .Y(mai_mai_n1290_));
  OR2        m1262(.A(mai_mai_n1290_), .B(mai_mai_n888_), .Y(mai_mai_n1291_));
  NA4        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1289_), .C(mai_mai_n1287_), .D(mai_mai_n1266_), .Y(mai_mai_n1292_));
  NO3        m1264(.A(mai_mai_n1292_), .B(mai_mai_n1269_), .C(mai_mai_n251_), .Y(mai_mai_n1293_));
  NO2        m1265(.A(mai_mai_n296_), .B(mai_mai_n45_), .Y(mai_mai_n1294_));
  AOI210     m1266(.A0(mai_mai_n1294_), .A1(mai_mai_n554_), .B0(mai_mai_n1264_), .Y(mai_mai_n1295_));
  AOI210     m1267(.A0(mai_mai_n1294_), .A1(mai_mai_n558_), .B0(mai_mai_n1277_), .Y(mai_mai_n1296_));
  AOI210     m1268(.A0(mai_mai_n1296_), .A1(mai_mai_n1295_), .B0(mai_mai_n337_), .Y(mai_mai_n1297_));
  OAI210     m1269(.A0(mai_mai_n88_), .A1(mai_mai_n40_), .B0(mai_mai_n677_), .Y(mai_mai_n1298_));
  NA2        m1270(.A(mai_mai_n1298_), .B(mai_mai_n645_), .Y(mai_mai_n1299_));
  NO2        m1271(.A(mai_mai_n513_), .B(mai_mai_n168_), .Y(mai_mai_n1300_));
  NOi21      m1272(.An(mai_mai_n134_), .B(mai_mai_n45_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n610_), .B(mai_mai_n1116_), .Y(mai_mai_n1302_));
  OAI210     m1274(.A0(mai_mai_n461_), .A1(mai_mai_n244_), .B0(mai_mai_n911_), .Y(mai_mai_n1303_));
  NO4        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1302_), .C(mai_mai_n1301_), .D(mai_mai_n1300_), .Y(mai_mai_n1304_));
  OR2        m1276(.A(mai_mai_n601_), .B(mai_mai_n599_), .Y(mai_mai_n1305_));
  NO2        m1277(.A(mai_mai_n366_), .B(mai_mai_n133_), .Y(mai_mai_n1306_));
  INV        m1278(.A(mai_mai_n1305_), .Y(mai_mai_n1307_));
  NA3        m1279(.A(mai_mai_n1307_), .B(mai_mai_n1304_), .C(mai_mai_n1299_), .Y(mai_mai_n1308_));
  NO2        m1280(.A(mai_mai_n750_), .B(mai_mai_n365_), .Y(mai_mai_n1309_));
  NO3        m1281(.A(mai_mai_n679_), .B(mai_mai_n761_), .C(mai_mai_n638_), .Y(mai_mai_n1310_));
  NOi21      m1282(.An(mai_mai_n1309_), .B(mai_mai_n1310_), .Y(mai_mai_n1311_));
  AN2        m1283(.A(mai_mai_n957_), .B(mai_mai_n648_), .Y(mai_mai_n1312_));
  NO4        m1284(.A(mai_mai_n1312_), .B(mai_mai_n1311_), .C(mai_mai_n1308_), .D(mai_mai_n1297_), .Y(mai_mai_n1313_));
  NO2        m1285(.A(mai_mai_n803_), .B(mai_mai_n272_), .Y(mai_mai_n1314_));
  OAI220     m1286(.A0(mai_mai_n734_), .A1(mai_mai_n47_), .B0(mai_mai_n220_), .B1(mai_mai_n619_), .Y(mai_mai_n1315_));
  OAI210     m1287(.A0(mai_mai_n272_), .A1(c), .B0(mai_mai_n644_), .Y(mai_mai_n1316_));
  AOI220     m1288(.A0(mai_mai_n1316_), .A1(mai_mai_n1315_), .B0(mai_mai_n1314_), .B1(mai_mai_n263_), .Y(mai_mai_n1317_));
  OAI220     m1289(.A0(mai_mai_n701_), .A1(mai_mai_n244_), .B0(mai_mai_n509_), .B1(mai_mai_n513_), .Y(mai_mai_n1318_));
  OAI210     m1290(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1319_));
  NO3        m1291(.A(mai_mai_n1319_), .B(mai_mai_n598_), .C(j), .Y(mai_mai_n1320_));
  NOi21      m1292(.An(mai_mai_n1320_), .B(mai_mai_n671_), .Y(mai_mai_n1321_));
  NO3        m1293(.A(mai_mai_n1321_), .B(mai_mai_n1318_), .C(mai_mai_n1119_), .Y(mai_mai_n1322_));
  NA3        m1294(.A(mai_mai_n794_), .B(mai_mai_n438_), .C(mai_mai_n880_), .Y(mai_mai_n1323_));
  NAi31      m1295(.An(mai_mai_n750_), .B(mai_mai_n1323_), .C(mai_mai_n199_), .Y(mai_mai_n1324_));
  NA4        m1296(.A(mai_mai_n1324_), .B(mai_mai_n1322_), .C(mai_mai_n1317_), .D(mai_mai_n1208_), .Y(mai_mai_n1325_));
  NOi31      m1297(.An(mai_mai_n1290_), .B(mai_mai_n465_), .C(mai_mai_n394_), .Y(mai_mai_n1326_));
  OR3        m1298(.A(mai_mai_n1326_), .B(mai_mai_n784_), .C(mai_mai_n541_), .Y(mai_mai_n1327_));
  OR3        m1299(.A(mai_mai_n369_), .B(mai_mai_n220_), .C(mai_mai_n619_), .Y(mai_mai_n1328_));
  AOI210     m1300(.A0(mai_mai_n573_), .A1(mai_mai_n450_), .B0(mai_mai_n371_), .Y(mai_mai_n1329_));
  NA3        m1301(.A(mai_mai_n1329_), .B(mai_mai_n1328_), .C(mai_mai_n1327_), .Y(mai_mai_n1330_));
  AOI220     m1302(.A0(mai_mai_n1309_), .A1(mai_mai_n760_), .B0(mai_mai_n1306_), .B1(mai_mai_n234_), .Y(mai_mai_n1331_));
  AN2        m1303(.A(mai_mai_n933_), .B(mai_mai_n932_), .Y(mai_mai_n1332_));
  NO4        m1304(.A(mai_mai_n1332_), .B(mai_mai_n878_), .C(mai_mai_n499_), .D(mai_mai_n482_), .Y(mai_mai_n1333_));
  NA3        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1331_), .C(mai_mai_n1272_), .Y(mai_mai_n1334_));
  NAi21      m1306(.An(j), .B(i), .Y(mai_mai_n1335_));
  NO4        m1307(.A(mai_mai_n1281_), .B(mai_mai_n1335_), .C(mai_mai_n444_), .D(mai_mai_n231_), .Y(mai_mai_n1336_));
  NO4        m1308(.A(mai_mai_n1336_), .B(mai_mai_n1334_), .C(mai_mai_n1330_), .D(mai_mai_n1325_), .Y(mai_mai_n1337_));
  NA4        m1309(.A(mai_mai_n1337_), .B(mai_mai_n1313_), .C(mai_mai_n1293_), .D(mai_mai_n1283_), .Y(mai07));
  NOi21      m1310(.An(j), .B(k), .Y(mai_mai_n1339_));
  NA4        m1311(.A(mai_mai_n176_), .B(mai_mai_n106_), .C(mai_mai_n1339_), .D(f), .Y(mai_mai_n1340_));
  NAi32      m1312(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1341_));
  NO3        m1313(.A(mai_mai_n1341_), .B(g), .C(f), .Y(mai_mai_n1342_));
  OAI210     m1314(.A0(mai_mai_n319_), .A1(mai_mai_n484_), .B0(mai_mai_n1342_), .Y(mai_mai_n1343_));
  NAi21      m1315(.An(f), .B(c), .Y(mai_mai_n1344_));
  OR2        m1316(.A(e), .B(d), .Y(mai_mai_n1345_));
  OAI220     m1317(.A0(mai_mai_n1345_), .A1(mai_mai_n1344_), .B0(mai_mai_n632_), .B1(mai_mai_n321_), .Y(mai_mai_n1346_));
  NA3        m1318(.A(mai_mai_n1346_), .B(mai_mai_n1060_), .C(mai_mai_n176_), .Y(mai_mai_n1347_));
  NOi31      m1319(.An(n), .B(m), .C(b), .Y(mai_mai_n1348_));
  NO3        m1320(.A(mai_mai_n130_), .B(mai_mai_n451_), .C(h), .Y(mai_mai_n1349_));
  NA3        m1321(.A(mai_mai_n1347_), .B(mai_mai_n1343_), .C(mai_mai_n1340_), .Y(mai_mai_n1350_));
  NOi41      m1322(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1351_));
  NO2        m1323(.A(k), .B(i), .Y(mai_mai_n1352_));
  NA3        m1324(.A(mai_mai_n1352_), .B(mai_mai_n899_), .C(mai_mai_n176_), .Y(mai_mai_n1353_));
  NA2        m1325(.A(mai_mai_n86_), .B(mai_mai_n45_), .Y(mai_mai_n1354_));
  NO2        m1326(.A(mai_mai_n1054_), .B(mai_mai_n444_), .Y(mai_mai_n1355_));
  NA3        m1327(.A(mai_mai_n1355_), .B(mai_mai_n1354_), .C(mai_mai_n211_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n1068_), .B(mai_mai_n304_), .Y(mai_mai_n1357_));
  NA2        m1329(.A(mai_mai_n542_), .B(mai_mai_n81_), .Y(mai_mai_n1358_));
  NA2        m1330(.A(mai_mai_n1209_), .B(mai_mai_n286_), .Y(mai_mai_n1359_));
  NA4        m1331(.A(mai_mai_n1359_), .B(mai_mai_n1358_), .C(mai_mai_n1356_), .D(mai_mai_n1353_), .Y(mai_mai_n1360_));
  NO2        m1332(.A(mai_mai_n1360_), .B(mai_mai_n1350_), .Y(mai_mai_n1361_));
  NO3        m1333(.A(e), .B(d), .C(c), .Y(mai_mai_n1362_));
  NA2        m1334(.A(mai_mai_n1522_), .B(mai_mai_n1362_), .Y(mai_mai_n1363_));
  NO2        m1335(.A(mai_mai_n1363_), .B(mai_mai_n211_), .Y(mai_mai_n1364_));
  OR2        m1336(.A(h), .B(f), .Y(mai_mai_n1365_));
  NO3        m1337(.A(n), .B(m), .C(i), .Y(mai_mai_n1366_));
  OAI210     m1338(.A0(mai_mai_n1117_), .A1(mai_mai_n151_), .B0(mai_mai_n1366_), .Y(mai_mai_n1367_));
  NO2        m1339(.A(mai_mai_n1367_), .B(mai_mai_n1365_), .Y(mai_mai_n1368_));
  NA3        m1340(.A(mai_mai_n698_), .B(mai_mai_n687_), .C(mai_mai_n110_), .Y(mai_mai_n1369_));
  NO2        m1341(.A(mai_mai_n1369_), .B(mai_mai_n45_), .Y(mai_mai_n1370_));
  NO2        m1342(.A(l), .B(k), .Y(mai_mai_n1371_));
  NOi41      m1343(.An(mai_mai_n547_), .B(mai_mai_n1371_), .C(mai_mai_n479_), .D(mai_mai_n444_), .Y(mai_mai_n1372_));
  NO3        m1344(.A(mai_mai_n444_), .B(d), .C(c), .Y(mai_mai_n1373_));
  NO4        m1345(.A(mai_mai_n1372_), .B(mai_mai_n1370_), .C(mai_mai_n1368_), .D(mai_mai_n1364_), .Y(mai_mai_n1374_));
  NO2        m1346(.A(mai_mai_n142_), .B(h), .Y(mai_mai_n1375_));
  NO2        m1347(.A(mai_mai_n1078_), .B(l), .Y(mai_mai_n1376_));
  NO2        m1348(.A(g), .B(c), .Y(mai_mai_n1377_));
  NA3        m1349(.A(mai_mai_n1377_), .B(mai_mai_n139_), .C(mai_mai_n182_), .Y(mai_mai_n1378_));
  NO2        m1350(.A(mai_mai_n1378_), .B(mai_mai_n1376_), .Y(mai_mai_n1379_));
  NA2        m1351(.A(mai_mai_n1379_), .B(mai_mai_n176_), .Y(mai_mai_n1380_));
  NO2        m1352(.A(mai_mai_n452_), .B(a), .Y(mai_mai_n1381_));
  NA3        m1353(.A(mai_mai_n1381_), .B(k), .C(mai_mai_n111_), .Y(mai_mai_n1382_));
  NO2        m1354(.A(i), .B(h), .Y(mai_mai_n1383_));
  AOI210     m1355(.A0(mai_mai_n1141_), .A1(h), .B0(mai_mai_n415_), .Y(mai_mai_n1384_));
  NA2        m1356(.A(mai_mai_n136_), .B(mai_mai_n216_), .Y(mai_mai_n1385_));
  NO2        m1357(.A(mai_mai_n1385_), .B(mai_mai_n1384_), .Y(mai_mai_n1386_));
  NO2        m1358(.A(mai_mai_n757_), .B(mai_mai_n183_), .Y(mai_mai_n1387_));
  NOi31      m1359(.An(m), .B(n), .C(b), .Y(mai_mai_n1388_));
  NOi31      m1360(.An(f), .B(d), .C(c), .Y(mai_mai_n1389_));
  NA2        m1361(.A(mai_mai_n1389_), .B(mai_mai_n1388_), .Y(mai_mai_n1390_));
  INV        m1362(.A(mai_mai_n1390_), .Y(mai_mai_n1391_));
  NO3        m1363(.A(mai_mai_n1391_), .B(mai_mai_n1387_), .C(mai_mai_n1386_), .Y(mai_mai_n1392_));
  NA2        m1364(.A(mai_mai_n1089_), .B(mai_mai_n468_), .Y(mai_mai_n1393_));
  NO4        m1365(.A(mai_mai_n1393_), .B(mai_mai_n1063_), .C(mai_mai_n444_), .D(mai_mai_n45_), .Y(mai_mai_n1394_));
  OAI210     m1366(.A0(mai_mai_n179_), .A1(mai_mai_n525_), .B0(mai_mai_n1064_), .Y(mai_mai_n1395_));
  NO3        m1367(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1396_));
  INV        m1368(.A(mai_mai_n1395_), .Y(mai_mai_n1397_));
  NO2        m1369(.A(mai_mai_n1397_), .B(mai_mai_n1394_), .Y(mai_mai_n1398_));
  AN4        m1370(.A(mai_mai_n1398_), .B(mai_mai_n1392_), .C(mai_mai_n1382_), .D(mai_mai_n1380_), .Y(mai_mai_n1399_));
  NA2        m1371(.A(mai_mai_n1348_), .B(mai_mai_n378_), .Y(mai_mai_n1400_));
  NO2        m1372(.A(mai_mai_n1400_), .B(mai_mai_n1045_), .Y(mai_mai_n1401_));
  NA2        m1373(.A(mai_mai_n1373_), .B(mai_mai_n212_), .Y(mai_mai_n1402_));
  NO2        m1374(.A(mai_mai_n183_), .B(b), .Y(mai_mai_n1403_));
  AOI220     m1375(.A0(mai_mai_n1173_), .A1(mai_mai_n1403_), .B0(mai_mai_n1097_), .B1(mai_mai_n1393_), .Y(mai_mai_n1404_));
  NAi31      m1376(.An(mai_mai_n1401_), .B(mai_mai_n1404_), .C(mai_mai_n1402_), .Y(mai_mai_n1405_));
  NO4        m1377(.A(mai_mai_n130_), .B(g), .C(f), .D(e), .Y(mai_mai_n1406_));
  NA3        m1378(.A(mai_mai_n1352_), .B(mai_mai_n287_), .C(h), .Y(mai_mai_n1407_));
  OR2        m1379(.A(e), .B(a), .Y(mai_mai_n1408_));
  NO2        m1380(.A(mai_mai_n1345_), .B(mai_mai_n1344_), .Y(mai_mai_n1409_));
  AOI210     m1381(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1409_), .Y(mai_mai_n1410_));
  NO2        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1085_), .Y(mai_mai_n1411_));
  NA2        m1383(.A(mai_mai_n1351_), .B(mai_mai_n1371_), .Y(mai_mai_n1412_));
  INV        m1384(.A(mai_mai_n1412_), .Y(mai_mai_n1413_));
  OR3        m1385(.A(mai_mai_n541_), .B(mai_mai_n540_), .C(mai_mai_n110_), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1115_), .B(mai_mai_n407_), .Y(mai_mai_n1415_));
  NO2        m1387(.A(mai_mai_n1415_), .B(mai_mai_n437_), .Y(mai_mai_n1416_));
  AO210      m1388(.A0(mai_mai_n1416_), .A1(mai_mai_n114_), .B0(mai_mai_n1413_), .Y(mai_mai_n1417_));
  NO3        m1389(.A(mai_mai_n1417_), .B(mai_mai_n1411_), .C(mai_mai_n1405_), .Y(mai_mai_n1418_));
  NA4        m1390(.A(mai_mai_n1418_), .B(mai_mai_n1399_), .C(mai_mai_n1374_), .D(mai_mai_n1361_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n390_), .B(j), .Y(mai_mai_n1420_));
  NA3        m1392(.A(mai_mai_n1396_), .B(mai_mai_n1345_), .C(mai_mai_n1115_), .Y(mai_mai_n1421_));
  NAi41      m1393(.An(mai_mai_n1383_), .B(mai_mai_n1076_), .C(mai_mai_n164_), .D(mai_mai_n145_), .Y(mai_mai_n1422_));
  NA2        m1394(.A(mai_mai_n1422_), .B(mai_mai_n1421_), .Y(mai_mai_n1423_));
  NA3        m1395(.A(g), .B(mai_mai_n1420_), .C(mai_mai_n153_), .Y(mai_mai_n1424_));
  INV        m1396(.A(mai_mai_n1424_), .Y(mai_mai_n1425_));
  NO3        m1397(.A(mai_mai_n750_), .B(mai_mai_n171_), .C(mai_mai_n410_), .Y(mai_mai_n1426_));
  NO3        m1398(.A(mai_mai_n1426_), .B(mai_mai_n1425_), .C(mai_mai_n1423_), .Y(mai_mai_n1427_));
  OR2        m1399(.A(n), .B(i), .Y(mai_mai_n1428_));
  OAI210     m1400(.A0(mai_mai_n1428_), .A1(mai_mai_n1075_), .B0(mai_mai_n49_), .Y(mai_mai_n1429_));
  AOI220     m1401(.A0(mai_mai_n1429_), .A1(mai_mai_n1179_), .B0(mai_mai_n826_), .B1(mai_mai_n190_), .Y(mai_mai_n1430_));
  INV        m1402(.A(mai_mai_n1430_), .Y(mai_mai_n1431_));
  NO2        m1403(.A(mai_mai_n130_), .B(l), .Y(mai_mai_n1432_));
  NO2        m1404(.A(mai_mai_n220_), .B(k), .Y(mai_mai_n1433_));
  OAI210     m1405(.A0(mai_mai_n1433_), .A1(mai_mai_n1383_), .B0(mai_mai_n1432_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(mai_mai_n1434_), .B(mai_mai_n31_), .Y(mai_mai_n1435_));
  NO3        m1407(.A(mai_mai_n1414_), .B(mai_mai_n468_), .C(mai_mai_n351_), .Y(mai_mai_n1436_));
  NO3        m1408(.A(mai_mai_n1436_), .B(mai_mai_n1435_), .C(mai_mai_n1431_), .Y(mai_mai_n1437_));
  NO3        m1409(.A(mai_mai_n1100_), .B(mai_mai_n1345_), .C(mai_mai_n49_), .Y(mai_mai_n1438_));
  NO2        m1410(.A(mai_mai_n1085_), .B(h), .Y(mai_mai_n1439_));
  NA3        m1411(.A(mai_mai_n1439_), .B(d), .C(mai_mai_n1046_), .Y(mai_mai_n1440_));
  NO2        m1412(.A(mai_mai_n1440_), .B(c), .Y(mai_mai_n1441_));
  NA2        m1413(.A(mai_mai_n176_), .B(mai_mai_n110_), .Y(mai_mai_n1442_));
  NOi21      m1414(.An(d), .B(f), .Y(mai_mai_n1443_));
  NO2        m1415(.A(mai_mai_n1345_), .B(f), .Y(mai_mai_n1444_));
  INV        m1416(.A(mai_mai_n1441_), .Y(mai_mai_n1445_));
  NA3        m1417(.A(mai_mai_n1445_), .B(mai_mai_n1437_), .C(mai_mai_n1427_), .Y(mai_mai_n1446_));
  NO3        m1418(.A(mai_mai_n1089_), .B(mai_mai_n1075_), .C(mai_mai_n40_), .Y(mai_mai_n1447_));
  NO2        m1419(.A(mai_mai_n468_), .B(mai_mai_n296_), .Y(mai_mai_n1448_));
  OAI210     m1420(.A0(mai_mai_n1448_), .A1(mai_mai_n1447_), .B0(mai_mai_n1357_), .Y(mai_mai_n1449_));
  OAI210     m1421(.A0(mai_mai_n1406_), .A1(mai_mai_n1348_), .B0(mai_mai_n885_), .Y(mai_mai_n1450_));
  NO2        m1422(.A(mai_mai_n1042_), .B(mai_mai_n130_), .Y(mai_mai_n1451_));
  NA2        m1423(.A(mai_mai_n1451_), .B(mai_mai_n625_), .Y(mai_mai_n1452_));
  NA3        m1424(.A(mai_mai_n1452_), .B(mai_mai_n1450_), .C(mai_mai_n1449_), .Y(mai_mai_n1453_));
  NA2        m1425(.A(mai_mai_n1377_), .B(mai_mai_n1443_), .Y(mai_mai_n1454_));
  NO2        m1426(.A(mai_mai_n1454_), .B(m), .Y(mai_mai_n1455_));
  NO2        m1427(.A(mai_mai_n146_), .B(mai_mai_n178_), .Y(mai_mai_n1456_));
  OAI210     m1428(.A0(mai_mai_n1456_), .A1(mai_mai_n108_), .B0(mai_mai_n1388_), .Y(mai_mai_n1457_));
  INV        m1429(.A(mai_mai_n1457_), .Y(mai_mai_n1458_));
  NO3        m1430(.A(mai_mai_n1458_), .B(mai_mai_n1455_), .C(mai_mai_n1453_), .Y(mai_mai_n1459_));
  NO2        m1431(.A(mai_mai_n1344_), .B(e), .Y(mai_mai_n1460_));
  NA2        m1432(.A(mai_mai_n1460_), .B(mai_mai_n405_), .Y(mai_mai_n1461_));
  NA2        m1433(.A(mai_mai_n1126_), .B(mai_mai_n634_), .Y(mai_mai_n1462_));
  OR3        m1434(.A(mai_mai_n1433_), .B(mai_mai_n1209_), .C(mai_mai_n130_), .Y(mai_mai_n1463_));
  OAI220     m1435(.A0(mai_mai_n1463_), .A1(mai_mai_n1461_), .B0(mai_mai_n1462_), .B1(mai_mai_n446_), .Y(mai_mai_n1464_));
  INV        m1436(.A(mai_mai_n1464_), .Y(mai_mai_n1465_));
  NO2        m1437(.A(mai_mai_n178_), .B(c), .Y(mai_mai_n1466_));
  OAI210     m1438(.A0(mai_mai_n1466_), .A1(mai_mai_n1460_), .B0(mai_mai_n176_), .Y(mai_mai_n1467_));
  AOI220     m1439(.A0(mai_mai_n1467_), .A1(mai_mai_n1077_), .B0(mai_mai_n532_), .B1(mai_mai_n365_), .Y(mai_mai_n1468_));
  NA2        m1440(.A(mai_mai_n540_), .B(g), .Y(mai_mai_n1469_));
  AOI210     m1441(.A0(mai_mai_n1469_), .A1(mai_mai_n1373_), .B0(mai_mai_n1438_), .Y(mai_mai_n1470_));
  NO2        m1442(.A(mai_mai_n1408_), .B(f), .Y(mai_mai_n1471_));
  AOI210     m1443(.A0(mai_mai_n1126_), .A1(a), .B0(mai_mai_n1471_), .Y(mai_mai_n1472_));
  OAI220     m1444(.A0(mai_mai_n1472_), .A1(mai_mai_n69_), .B0(mai_mai_n1470_), .B1(mai_mai_n210_), .Y(mai_mai_n1473_));
  AOI210     m1445(.A0(mai_mai_n904_), .A1(mai_mai_n417_), .B0(mai_mai_n102_), .Y(mai_mai_n1474_));
  OR2        m1446(.A(mai_mai_n1474_), .B(mai_mai_n540_), .Y(mai_mai_n1475_));
  NA2        m1447(.A(mai_mai_n1471_), .B(mai_mai_n1354_), .Y(mai_mai_n1476_));
  OAI220     m1448(.A0(mai_mai_n1476_), .A1(mai_mai_n49_), .B0(mai_mai_n1475_), .B1(mai_mai_n171_), .Y(mai_mai_n1477_));
  NA4        m1449(.A(mai_mai_n1098_), .B(mai_mai_n1095_), .C(mai_mai_n216_), .D(mai_mai_n68_), .Y(mai_mai_n1478_));
  NA2        m1450(.A(mai_mai_n1349_), .B(mai_mai_n179_), .Y(mai_mai_n1479_));
  NO2        m1451(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1480_));
  OAI210     m1452(.A0(mai_mai_n1408_), .A1(mai_mai_n863_), .B0(mai_mai_n484_), .Y(mai_mai_n1481_));
  OAI210     m1453(.A0(mai_mai_n1481_), .A1(mai_mai_n1101_), .B0(mai_mai_n1480_), .Y(mai_mai_n1482_));
  NO2        m1454(.A(mai_mai_n247_), .B(g), .Y(mai_mai_n1483_));
  NO2        m1455(.A(m), .B(i), .Y(mai_mai_n1484_));
  BUFFER     m1456(.A(mai_mai_n1484_), .Y(mai_mai_n1485_));
  AOI220     m1457(.A0(mai_mai_n1485_), .A1(mai_mai_n1375_), .B0(mai_mai_n1076_), .B1(mai_mai_n1483_), .Y(mai_mai_n1486_));
  NA4        m1458(.A(mai_mai_n1486_), .B(mai_mai_n1482_), .C(mai_mai_n1479_), .D(mai_mai_n1478_), .Y(mai_mai_n1487_));
  NO4        m1459(.A(mai_mai_n1487_), .B(mai_mai_n1477_), .C(mai_mai_n1473_), .D(mai_mai_n1468_), .Y(mai_mai_n1488_));
  NA3        m1460(.A(mai_mai_n1488_), .B(mai_mai_n1465_), .C(mai_mai_n1459_), .Y(mai_mai_n1489_));
  NA3        m1461(.A(mai_mai_n963_), .B(mai_mai_n136_), .C(mai_mai_n46_), .Y(mai_mai_n1490_));
  AOI210     m1462(.A0(mai_mai_n143_), .A1(c), .B0(mai_mai_n1490_), .Y(mai_mai_n1491_));
  INV        m1463(.A(mai_mai_n180_), .Y(mai_mai_n1492_));
  NA2        m1464(.A(mai_mai_n1492_), .B(mai_mai_n1439_), .Y(mai_mai_n1493_));
  OR2        m1465(.A(mai_mai_n131_), .B(mai_mai_n1400_), .Y(mai_mai_n1494_));
  NA2        m1466(.A(mai_mai_n1494_), .B(mai_mai_n1493_), .Y(mai_mai_n1495_));
  NO2        m1467(.A(mai_mai_n1495_), .B(mai_mai_n1491_), .Y(mai_mai_n1496_));
  AOI210     m1468(.A0(mai_mai_n151_), .A1(mai_mai_n56_), .B0(mai_mai_n1460_), .Y(mai_mai_n1497_));
  NO2        m1469(.A(mai_mai_n1497_), .B(mai_mai_n1442_), .Y(mai_mai_n1498_));
  NOi21      m1470(.An(mai_mai_n1349_), .B(e), .Y(mai_mai_n1499_));
  NO2        m1471(.A(mai_mai_n1499_), .B(mai_mai_n1498_), .Y(mai_mai_n1500_));
  AN2        m1472(.A(mai_mai_n1098_), .B(mai_mai_n1083_), .Y(mai_mai_n1501_));
  AOI220     m1473(.A0(mai_mai_n1484_), .A1(mai_mai_n643_), .B0(mai_mai_n1060_), .B1(mai_mai_n154_), .Y(mai_mai_n1502_));
  NOi31      m1474(.An(mai_mai_n30_), .B(mai_mai_n1502_), .C(n), .Y(mai_mai_n1503_));
  AOI210     m1475(.A0(mai_mai_n1501_), .A1(mai_mai_n1173_), .B0(mai_mai_n1503_), .Y(mai_mai_n1504_));
  NA2        m1476(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1505_));
  NO2        m1477(.A(mai_mai_n1352_), .B(mai_mai_n116_), .Y(mai_mai_n1506_));
  OAI220     m1478(.A0(mai_mai_n1506_), .A1(mai_mai_n1400_), .B0(mai_mai_n1415_), .B1(mai_mai_n1505_), .Y(mai_mai_n1507_));
  INV        m1479(.A(mai_mai_n1507_), .Y(mai_mai_n1508_));
  NA4        m1480(.A(mai_mai_n1508_), .B(mai_mai_n1504_), .C(mai_mai_n1500_), .D(mai_mai_n1496_), .Y(mai_mai_n1509_));
  OR4        m1481(.A(mai_mai_n1509_), .B(mai_mai_n1489_), .C(mai_mai_n1446_), .D(mai_mai_n1419_), .Y(mai04));
  NOi31      m1482(.An(mai_mai_n1406_), .B(mai_mai_n1407_), .C(mai_mai_n1048_), .Y(mai_mai_n1511_));
  NA2        m1483(.A(mai_mai_n1444_), .B(mai_mai_n826_), .Y(mai_mai_n1512_));
  NO3        m1484(.A(mai_mai_n1512_), .B(mai_mai_n1037_), .C(mai_mai_n485_), .Y(mai_mai_n1513_));
  OR3        m1485(.A(mai_mai_n1513_), .B(mai_mai_n1511_), .C(mai_mai_n1066_), .Y(mai_mai_n1514_));
  NO2        m1486(.A(mai_mai_n1354_), .B(mai_mai_n89_), .Y(mai_mai_n1515_));
  AOI210     m1487(.A0(mai_mai_n1515_), .A1(mai_mai_n1059_), .B0(mai_mai_n1189_), .Y(mai_mai_n1516_));
  NA2        m1488(.A(mai_mai_n1516_), .B(mai_mai_n1213_), .Y(mai_mai_n1517_));
  NO4        m1489(.A(mai_mai_n1517_), .B(mai_mai_n1514_), .C(mai_mai_n1074_), .D(mai_mai_n1053_), .Y(mai_mai_n1518_));
  NA4        m1490(.A(mai_mai_n1518_), .B(mai_mai_n1128_), .C(mai_mai_n1113_), .D(mai_mai_n1104_), .Y(mai05));
  INV        m1491(.A(m), .Y(mai_mai_n1522_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(g), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(g), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(g), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO4        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .D(men_men_n92_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO3        u0081(.A(men_men_n109_), .B(men_men_n106_), .C(g), .Y(men_men_n110_));
  NOi21      u0082(.An(g), .B(f), .Y(men_men_n111_));
  NOi21      u0083(.An(i), .B(h), .Y(men_men_n112_));
  NA3        u0084(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n36_), .Y(men_men_n113_));
  INV        u0085(.A(a), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n107_), .B(men_men_n114_), .Y(men_men_n115_));
  INV        u0087(.A(l), .Y(men_men_n116_));
  NOi21      u0088(.An(m), .B(n), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(h), .Y(men_men_n118_));
  NO2        u0090(.A(men_men_n113_), .B(men_men_n88_), .Y(men_men_n119_));
  INV        u0091(.A(b), .Y(men_men_n120_));
  NA2        u0092(.A(l), .B(j), .Y(men_men_n121_));
  AN2        u0093(.A(k), .B(i), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NA2        u0095(.A(g), .B(e), .Y(men_men_n124_));
  NOi32      u0096(.An(c), .Bn(a), .C(d), .Y(men_men_n125_));
  NA2        u0097(.A(men_men_n125_), .B(men_men_n117_), .Y(men_men_n126_));
  NO4        u0098(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .D(men_men_n120_), .Y(men_men_n127_));
  NO3        u0099(.A(men_men_n127_), .B(men_men_n119_), .C(men_men_n110_), .Y(men_men_n128_));
  OAI210     u0100(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n128_), .Y(men_men_n129_));
  NOi31      u0101(.An(k), .B(m), .C(j), .Y(men_men_n130_));
  NA3        u0102(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n131_));
  NOi31      u0103(.An(k), .B(m), .C(i), .Y(men_men_n132_));
  NA3        u0104(.A(men_men_n132_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n134_));
  NOi32      u0106(.An(f), .Bn(b), .C(e), .Y(men_men_n135_));
  NAi21      u0107(.An(g), .B(h), .Y(men_men_n136_));
  NAi21      u0108(.An(m), .B(n), .Y(men_men_n137_));
  NAi21      u0109(.An(j), .B(k), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NAi41      u0111(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n140_));
  NAi31      u0112(.An(j), .B(k), .C(h), .Y(men_men_n141_));
  NO3        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n137_), .Y(men_men_n142_));
  AOI210     u0114(.A0(men_men_n139_), .A1(men_men_n135_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u0115(.A(k), .B(j), .Y(men_men_n144_));
  NO2        u0116(.A(men_men_n144_), .B(men_men_n137_), .Y(men_men_n145_));
  AN2        u0117(.A(k), .B(j), .Y(men_men_n146_));
  NAi21      u0118(.An(c), .B(b), .Y(men_men_n147_));
  NA2        u0119(.A(f), .B(d), .Y(men_men_n148_));
  NO4        u0120(.A(men_men_n148_), .B(men_men_n147_), .C(men_men_n146_), .D(men_men_n136_), .Y(men_men_n149_));
  NA2        u0121(.A(h), .B(c), .Y(men_men_n150_));
  NAi31      u0122(.An(f), .B(e), .C(b), .Y(men_men_n151_));
  NA2        u0123(.A(men_men_n149_), .B(men_men_n145_), .Y(men_men_n152_));
  NA2        u0124(.A(d), .B(b), .Y(men_men_n153_));
  NAi21      u0125(.An(e), .B(f), .Y(men_men_n154_));
  NO2        u0126(.A(men_men_n154_), .B(men_men_n153_), .Y(men_men_n155_));
  NA2        u0127(.A(b), .B(a), .Y(men_men_n156_));
  NAi21      u0128(.An(e), .B(g), .Y(men_men_n157_));
  NAi21      u0129(.An(c), .B(d), .Y(men_men_n158_));
  NAi31      u0130(.An(l), .B(k), .C(h), .Y(men_men_n159_));
  NO2        u0131(.A(men_men_n137_), .B(men_men_n159_), .Y(men_men_n160_));
  NA2        u0132(.A(men_men_n160_), .B(men_men_n155_), .Y(men_men_n161_));
  NAi41      u0133(.An(men_men_n134_), .B(men_men_n161_), .C(men_men_n152_), .D(men_men_n143_), .Y(men_men_n162_));
  NAi31      u0134(.An(e), .B(f), .C(b), .Y(men_men_n163_));
  NOi21      u0135(.An(g), .B(d), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NOi21      u0137(.An(h), .B(i), .Y(men_men_n166_));
  NOi21      u0138(.An(k), .B(m), .Y(men_men_n167_));
  NA3        u0139(.A(men_men_n167_), .B(men_men_n166_), .C(n), .Y(men_men_n168_));
  NOi21      u0140(.An(h), .B(g), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NAi31      u0143(.An(l), .B(j), .C(h), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n49_), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n67_), .Y(men_men_n174_));
  NOi32      u0146(.An(n), .Bn(k), .C(m), .Y(men_men_n175_));
  NA2        u0147(.A(l), .B(i), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OAI210     u0149(.A0(men_men_n177_), .A1(men_men_n171_), .B0(men_men_n174_), .Y(men_men_n178_));
  NAi31      u0150(.An(d), .B(f), .C(c), .Y(men_men_n179_));
  NAi31      u0151(.An(e), .B(f), .C(c), .Y(men_men_n180_));
  NA2        u0152(.A(men_men_n180_), .B(men_men_n179_), .Y(men_men_n181_));
  NA2        u0153(.A(j), .B(h), .Y(men_men_n182_));
  OR3        u0154(.A(n), .B(m), .C(k), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  NAi32      u0156(.An(m), .Bn(k), .C(n), .Y(men_men_n185_));
  NO2        u0157(.A(men_men_n185_), .B(men_men_n182_), .Y(men_men_n186_));
  AOI220     u0158(.A0(men_men_n186_), .A1(men_men_n165_), .B0(men_men_n184_), .B1(men_men_n181_), .Y(men_men_n187_));
  NO2        u0159(.A(n), .B(m), .Y(men_men_n188_));
  NA2        u0160(.A(men_men_n188_), .B(men_men_n50_), .Y(men_men_n189_));
  NAi21      u0161(.An(f), .B(e), .Y(men_men_n190_));
  NA2        u0162(.A(d), .B(c), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi21      u0164(.An(men_men_n192_), .B(men_men_n189_), .Y(men_men_n193_));
  NAi21      u0165(.An(d), .B(c), .Y(men_men_n194_));
  NAi31      u0166(.An(m), .B(n), .C(b), .Y(men_men_n195_));
  NA2        u0167(.A(k), .B(i), .Y(men_men_n196_));
  NAi21      u0168(.An(h), .B(f), .Y(men_men_n197_));
  NO2        u0169(.A(men_men_n195_), .B(men_men_n158_), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(d), .Y(men_men_n199_));
  NOi32      u0171(.An(f), .Bn(c), .C(e), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n200_), .B(men_men_n199_), .Y(men_men_n201_));
  NO3        u0173(.A(n), .B(m), .C(j), .Y(men_men_n202_));
  NA2        u0174(.A(men_men_n202_), .B(men_men_n118_), .Y(men_men_n203_));
  AO210      u0175(.A0(men_men_n203_), .A1(men_men_n189_), .B0(men_men_n201_), .Y(men_men_n204_));
  NAi31      u0176(.An(men_men_n193_), .B(men_men_n204_), .C(men_men_n187_), .Y(men_men_n205_));
  OR3        u0177(.A(men_men_n205_), .B(men_men_n178_), .C(men_men_n162_), .Y(men_men_n206_));
  NO4        u0178(.A(men_men_n206_), .B(men_men_n129_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n207_));
  NA3        u0179(.A(m), .B(men_men_n116_), .C(j), .Y(men_men_n208_));
  NAi31      u0180(.An(n), .B(h), .C(g), .Y(men_men_n209_));
  NO2        u0181(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  NOi32      u0182(.An(m), .Bn(k), .C(l), .Y(men_men_n211_));
  NA3        u0183(.A(men_men_n211_), .B(men_men_n89_), .C(g), .Y(men_men_n212_));
  NO2        u0184(.A(men_men_n212_), .B(n), .Y(men_men_n213_));
  NOi21      u0185(.An(k), .B(j), .Y(men_men_n214_));
  NA4        u0186(.A(men_men_n214_), .B(men_men_n117_), .C(i), .D(g), .Y(men_men_n215_));
  AN2        u0187(.A(i), .B(g), .Y(men_men_n216_));
  NA3        u0188(.A(men_men_n76_), .B(men_men_n216_), .C(men_men_n117_), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n215_), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n213_), .C(men_men_n210_), .Y(men_men_n219_));
  NAi41      u0191(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n220_));
  INV        u0192(.A(men_men_n220_), .Y(men_men_n221_));
  INV        u0193(.A(f), .Y(men_men_n222_));
  INV        u0194(.A(g), .Y(men_men_n223_));
  NOi31      u0195(.An(i), .B(j), .C(h), .Y(men_men_n224_));
  NOi21      u0196(.An(l), .B(m), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NO3        u0198(.A(men_men_n226_), .B(men_men_n223_), .C(men_men_n222_), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n221_), .Y(men_men_n228_));
  OAI210     u0200(.A0(men_men_n219_), .A1(men_men_n32_), .B0(men_men_n228_), .Y(men_men_n229_));
  NOi21      u0201(.An(n), .B(m), .Y(men_men_n230_));
  NOi32      u0202(.An(l), .Bn(i), .C(j), .Y(men_men_n231_));
  NA2        u0203(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  OA220      u0204(.A0(men_men_n232_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n233_));
  NAi21      u0205(.An(j), .B(h), .Y(men_men_n234_));
  XN2        u0206(.A(i), .B(h), .Y(men_men_n235_));
  NA2        u0207(.A(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  NOi31      u0208(.An(k), .B(n), .C(m), .Y(men_men_n237_));
  NOi31      u0209(.An(men_men_n237_), .B(men_men_n191_), .C(men_men_n190_), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n238_), .B(men_men_n236_), .Y(men_men_n239_));
  NAi31      u0211(.An(f), .B(e), .C(c), .Y(men_men_n240_));
  NO4        u0212(.A(men_men_n240_), .B(men_men_n183_), .C(men_men_n182_), .D(men_men_n59_), .Y(men_men_n241_));
  NA4        u0213(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n242_));
  NAi32      u0214(.An(m), .Bn(i), .C(k), .Y(men_men_n243_));
  NO3        u0215(.A(men_men_n243_), .B(men_men_n93_), .C(men_men_n242_), .Y(men_men_n244_));
  INV        u0216(.A(k), .Y(men_men_n245_));
  NO2        u0217(.A(men_men_n244_), .B(men_men_n241_), .Y(men_men_n246_));
  NAi21      u0218(.An(n), .B(a), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n247_), .B(men_men_n153_), .Y(men_men_n248_));
  NAi41      u0220(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(e), .Y(men_men_n250_));
  NO3        u0222(.A(men_men_n154_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n251_));
  OAI210     u0223(.A0(men_men_n251_), .A1(men_men_n250_), .B0(men_men_n248_), .Y(men_men_n252_));
  AN4        u0224(.A(men_men_n252_), .B(men_men_n246_), .C(men_men_n239_), .D(men_men_n233_), .Y(men_men_n253_));
  OR2        u0225(.A(h), .B(g), .Y(men_men_n254_));
  NAi41      u0226(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n255_));
  NO2        u0227(.A(men_men_n255_), .B(men_men_n222_), .Y(men_men_n256_));
  NA2        u0228(.A(men_men_n167_), .B(men_men_n112_), .Y(men_men_n257_));
  NAi21      u0229(.An(men_men_n257_), .B(men_men_n256_), .Y(men_men_n258_));
  NO2        u0230(.A(n), .B(a), .Y(men_men_n259_));
  NAi31      u0231(.An(men_men_n249_), .B(men_men_n259_), .C(men_men_n107_), .Y(men_men_n260_));
  AN2        u0232(.A(men_men_n260_), .B(men_men_n258_), .Y(men_men_n261_));
  NAi21      u0233(.An(h), .B(i), .Y(men_men_n262_));
  NA2        u0234(.A(men_men_n188_), .B(k), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n263_), .B(men_men_n262_), .Y(men_men_n264_));
  NA2        u0236(.A(men_men_n264_), .B(men_men_n199_), .Y(men_men_n265_));
  NA2        u0237(.A(men_men_n265_), .B(men_men_n261_), .Y(men_men_n266_));
  NOi21      u0238(.An(g), .B(e), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n268_));
  NA2        u0240(.A(men_men_n268_), .B(men_men_n267_), .Y(men_men_n269_));
  NOi32      u0241(.An(l), .Bn(j), .C(i), .Y(men_men_n270_));
  AOI210     u0242(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n270_), .Y(men_men_n271_));
  NO2        u0243(.A(men_men_n262_), .B(men_men_n44_), .Y(men_men_n272_));
  NAi21      u0244(.An(f), .B(g), .Y(men_men_n273_));
  NO2        u0245(.A(men_men_n273_), .B(men_men_n65_), .Y(men_men_n274_));
  NO2        u0246(.A(men_men_n69_), .B(men_men_n121_), .Y(men_men_n275_));
  AOI220     u0247(.A0(men_men_n275_), .A1(men_men_n274_), .B0(men_men_n272_), .B1(men_men_n67_), .Y(men_men_n276_));
  OAI210     u0248(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n276_), .Y(men_men_n277_));
  NO3        u0249(.A(men_men_n138_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n278_));
  NOi41      u0250(.An(men_men_n253_), .B(men_men_n277_), .C(men_men_n266_), .D(men_men_n229_), .Y(men_men_n279_));
  NO4        u0251(.A(men_men_n210_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n280_));
  NO2        u0252(.A(men_men_n280_), .B(men_men_n115_), .Y(men_men_n281_));
  NA3        u0253(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n282_));
  NAi21      u0254(.An(h), .B(g), .Y(men_men_n283_));
  OR4        u0255(.A(men_men_n283_), .B(men_men_n282_), .C(men_men_n232_), .D(e), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n257_), .B(men_men_n273_), .Y(men_men_n285_));
  NA2        u0257(.A(men_men_n285_), .B(men_men_n78_), .Y(men_men_n286_));
  NAi31      u0258(.An(g), .B(k), .C(h), .Y(men_men_n287_));
  NO3        u0259(.A(men_men_n137_), .B(men_men_n287_), .C(l), .Y(men_men_n288_));
  NAi31      u0260(.An(e), .B(d), .C(a), .Y(men_men_n289_));
  NA2        u0261(.A(men_men_n288_), .B(men_men_n135_), .Y(men_men_n290_));
  NA3        u0262(.A(men_men_n290_), .B(men_men_n286_), .C(men_men_n284_), .Y(men_men_n291_));
  NA4        u0263(.A(men_men_n167_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n121_), .Y(men_men_n292_));
  NA3        u0264(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n86_), .Y(men_men_n293_));
  NO2        u0265(.A(men_men_n293_), .B(men_men_n201_), .Y(men_men_n294_));
  NOi21      u0266(.An(men_men_n292_), .B(men_men_n294_), .Y(men_men_n295_));
  NA3        u0267(.A(e), .B(c), .C(b), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n60_), .B(men_men_n296_), .Y(men_men_n297_));
  NAi32      u0269(.An(k), .Bn(i), .C(j), .Y(men_men_n298_));
  NAi31      u0270(.An(h), .B(l), .C(i), .Y(men_men_n299_));
  NA3        u0271(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n172_), .Y(men_men_n300_));
  NOi21      u0272(.An(men_men_n300_), .B(men_men_n49_), .Y(men_men_n301_));
  OAI210     u0273(.A0(men_men_n274_), .A1(men_men_n297_), .B0(men_men_n301_), .Y(men_men_n302_));
  NAi21      u0274(.An(l), .B(k), .Y(men_men_n303_));
  NO2        u0275(.A(men_men_n303_), .B(men_men_n49_), .Y(men_men_n304_));
  NOi21      u0276(.An(l), .B(j), .Y(men_men_n305_));
  NA2        u0277(.A(men_men_n169_), .B(men_men_n305_), .Y(men_men_n306_));
  NA3        u0278(.A(men_men_n122_), .B(men_men_n121_), .C(g), .Y(men_men_n307_));
  OR3        u0279(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n308_));
  AOI210     u0280(.A0(men_men_n307_), .A1(men_men_n306_), .B0(men_men_n308_), .Y(men_men_n309_));
  INV        u0281(.A(men_men_n309_), .Y(men_men_n310_));
  NAi32      u0282(.An(j), .Bn(h), .C(i), .Y(men_men_n311_));
  NAi21      u0283(.An(m), .B(l), .Y(men_men_n312_));
  NO3        u0284(.A(men_men_n312_), .B(men_men_n311_), .C(men_men_n86_), .Y(men_men_n313_));
  NA2        u0285(.A(h), .B(g), .Y(men_men_n314_));
  NA2        u0286(.A(men_men_n175_), .B(men_men_n45_), .Y(men_men_n315_));
  NO2        u0287(.A(men_men_n315_), .B(men_men_n314_), .Y(men_men_n316_));
  OAI210     u0288(.A0(men_men_n316_), .A1(men_men_n313_), .B0(men_men_n170_), .Y(men_men_n317_));
  NA4        u0289(.A(men_men_n317_), .B(men_men_n310_), .C(men_men_n302_), .D(men_men_n295_), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n151_), .B(d), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n320_));
  NAi32      u0292(.An(n), .Bn(m), .C(l), .Y(men_men_n321_));
  NO2        u0293(.A(men_men_n321_), .B(men_men_n311_), .Y(men_men_n322_));
  NA2        u0294(.A(men_men_n322_), .B(men_men_n192_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n126_), .B(men_men_n120_), .Y(men_men_n324_));
  NAi31      u0296(.An(k), .B(l), .C(j), .Y(men_men_n325_));
  OAI210     u0297(.A0(men_men_n303_), .A1(j), .B0(men_men_n325_), .Y(men_men_n326_));
  NOi21      u0298(.An(men_men_n326_), .B(men_men_n124_), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n327_), .B(men_men_n324_), .Y(men_men_n328_));
  NA2        u0300(.A(men_men_n328_), .B(men_men_n323_), .Y(men_men_n329_));
  NO4        u0301(.A(men_men_n329_), .B(men_men_n318_), .C(men_men_n291_), .D(men_men_n281_), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n264_), .B(men_men_n200_), .Y(men_men_n331_));
  NAi21      u0303(.An(m), .B(k), .Y(men_men_n332_));
  NO2        u0304(.A(men_men_n235_), .B(men_men_n332_), .Y(men_men_n333_));
  NAi31      u0305(.An(i), .B(l), .C(h), .Y(men_men_n334_));
  NO4        u0306(.A(men_men_n334_), .B(men_men_n157_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n335_));
  NA2        u0307(.A(e), .B(c), .Y(men_men_n336_));
  NO3        u0308(.A(men_men_n336_), .B(n), .C(d), .Y(men_men_n337_));
  NOi21      u0309(.An(f), .B(h), .Y(men_men_n338_));
  NAi31      u0310(.An(d), .B(e), .C(b), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n137_), .B(men_men_n339_), .Y(men_men_n340_));
  NAi21      u0312(.An(men_men_n335_), .B(men_men_n331_), .Y(men_men_n341_));
  NA2        u0313(.A(men_men_n259_), .B(men_men_n107_), .Y(men_men_n342_));
  OR2        u0314(.A(men_men_n342_), .B(men_men_n212_), .Y(men_men_n343_));
  NOi31      u0315(.An(l), .B(n), .C(m), .Y(men_men_n344_));
  NA2        u0316(.A(men_men_n344_), .B(men_men_n224_), .Y(men_men_n345_));
  NO2        u0317(.A(men_men_n345_), .B(men_men_n201_), .Y(men_men_n346_));
  NAi21      u0318(.An(men_men_n346_), .B(men_men_n343_), .Y(men_men_n347_));
  NAi32      u0319(.An(m), .Bn(j), .C(k), .Y(men_men_n348_));
  NAi41      u0320(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n349_));
  NOi31      u0321(.An(j), .B(m), .C(k), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n130_), .B(men_men_n350_), .Y(men_men_n351_));
  AN3        u0323(.A(h), .B(g), .C(f), .Y(men_men_n352_));
  NOi32      u0324(.An(m), .Bn(j), .C(l), .Y(men_men_n353_));
  NO2        u0325(.A(men_men_n353_), .B(men_men_n100_), .Y(men_men_n354_));
  NAi32      u0326(.An(men_men_n354_), .Bn(men_men_n209_), .C(men_men_n319_), .Y(men_men_n355_));
  NO2        u0327(.A(men_men_n312_), .B(men_men_n311_), .Y(men_men_n356_));
  NO2        u0328(.A(men_men_n226_), .B(g), .Y(men_men_n357_));
  NO2        u0329(.A(men_men_n163_), .B(men_men_n86_), .Y(men_men_n358_));
  AOI220     u0330(.A0(men_men_n358_), .A1(men_men_n357_), .B0(men_men_n256_), .B1(men_men_n356_), .Y(men_men_n359_));
  NA2        u0331(.A(men_men_n243_), .B(men_men_n81_), .Y(men_men_n360_));
  NA3        u0332(.A(men_men_n360_), .B(men_men_n352_), .C(men_men_n221_), .Y(men_men_n361_));
  NA3        u0333(.A(men_men_n361_), .B(men_men_n359_), .C(men_men_n355_), .Y(men_men_n362_));
  NA3        u0334(.A(h), .B(g), .C(f), .Y(men_men_n363_));
  NO2        u0335(.A(men_men_n363_), .B(men_men_n77_), .Y(men_men_n364_));
  NA2        u0336(.A(men_men_n349_), .B(men_men_n220_), .Y(men_men_n365_));
  NA2        u0337(.A(men_men_n169_), .B(e), .Y(men_men_n366_));
  NO2        u0338(.A(men_men_n366_), .B(men_men_n41_), .Y(men_men_n367_));
  AOI220     u0339(.A0(men_men_n367_), .A1(men_men_n324_), .B0(men_men_n365_), .B1(men_men_n364_), .Y(men_men_n368_));
  NOi32      u0340(.An(j), .Bn(g), .C(i), .Y(men_men_n369_));
  NA3        u0341(.A(men_men_n369_), .B(men_men_n303_), .C(men_men_n117_), .Y(men_men_n370_));
  AO210      u0342(.A0(men_men_n115_), .A1(men_men_n32_), .B0(men_men_n370_), .Y(men_men_n371_));
  NOi32      u0343(.An(e), .Bn(b), .C(a), .Y(men_men_n372_));
  AN2        u0344(.A(l), .B(j), .Y(men_men_n373_));
  NA3        u0345(.A(men_men_n217_), .B(men_men_n215_), .C(men_men_n35_), .Y(men_men_n374_));
  NA2        u0346(.A(men_men_n374_), .B(men_men_n372_), .Y(men_men_n375_));
  NO2        u0347(.A(men_men_n339_), .B(n), .Y(men_men_n376_));
  NA2        u0348(.A(men_men_n216_), .B(k), .Y(men_men_n377_));
  NA3        u0349(.A(m), .B(men_men_n116_), .C(men_men_n222_), .Y(men_men_n378_));
  NA4        u0350(.A(men_men_n211_), .B(men_men_n89_), .C(g), .D(men_men_n222_), .Y(men_men_n379_));
  OAI210     u0351(.A0(men_men_n378_), .A1(men_men_n377_), .B0(men_men_n379_), .Y(men_men_n380_));
  NAi41      u0352(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n51_), .B(men_men_n117_), .Y(men_men_n382_));
  NO2        u0354(.A(men_men_n382_), .B(men_men_n381_), .Y(men_men_n383_));
  AOI220     u0355(.A0(men_men_n383_), .A1(b), .B0(men_men_n380_), .B1(men_men_n376_), .Y(men_men_n384_));
  NA4        u0356(.A(men_men_n384_), .B(men_men_n375_), .C(men_men_n371_), .D(men_men_n368_), .Y(men_men_n385_));
  NO4        u0357(.A(men_men_n385_), .B(men_men_n362_), .C(men_men_n347_), .D(men_men_n341_), .Y(men_men_n386_));
  NA4        u0358(.A(men_men_n386_), .B(men_men_n330_), .C(men_men_n279_), .D(men_men_n207_), .Y(men10));
  NA3        u0359(.A(m), .B(k), .C(i), .Y(men_men_n388_));
  NO3        u0360(.A(men_men_n388_), .B(j), .C(men_men_n223_), .Y(men_men_n389_));
  NOi21      u0361(.An(e), .B(f), .Y(men_men_n390_));
  NO4        u0362(.A(men_men_n158_), .B(men_men_n390_), .C(n), .D(men_men_n114_), .Y(men_men_n391_));
  NAi31      u0363(.An(b), .B(f), .C(c), .Y(men_men_n392_));
  INV        u0364(.A(men_men_n392_), .Y(men_men_n393_));
  NOi32      u0365(.An(k), .Bn(h), .C(j), .Y(men_men_n394_));
  NA2        u0366(.A(men_men_n394_), .B(men_men_n230_), .Y(men_men_n395_));
  NA2        u0367(.A(men_men_n168_), .B(men_men_n395_), .Y(men_men_n396_));
  AOI220     u0368(.A0(men_men_n396_), .A1(men_men_n393_), .B0(men_men_n391_), .B1(men_men_n389_), .Y(men_men_n397_));
  AN2        u0369(.A(j), .B(h), .Y(men_men_n398_));
  NO3        u0370(.A(n), .B(m), .C(k), .Y(men_men_n399_));
  NA2        u0371(.A(men_men_n399_), .B(men_men_n398_), .Y(men_men_n400_));
  NO3        u0372(.A(men_men_n400_), .B(men_men_n158_), .C(men_men_n222_), .Y(men_men_n401_));
  OR2        u0373(.A(m), .B(k), .Y(men_men_n402_));
  NO2        u0374(.A(men_men_n182_), .B(men_men_n402_), .Y(men_men_n403_));
  NA4        u0375(.A(n), .B(f), .C(c), .D(men_men_n120_), .Y(men_men_n404_));
  NOi21      u0376(.An(men_men_n403_), .B(men_men_n404_), .Y(men_men_n405_));
  NOi32      u0377(.An(d), .Bn(a), .C(c), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n406_), .B(men_men_n190_), .Y(men_men_n407_));
  NAi21      u0379(.An(i), .B(g), .Y(men_men_n408_));
  NAi31      u0380(.An(k), .B(m), .C(j), .Y(men_men_n409_));
  NO3        u0381(.A(men_men_n409_), .B(men_men_n408_), .C(n), .Y(men_men_n410_));
  NOi21      u0382(.An(men_men_n410_), .B(men_men_n407_), .Y(men_men_n411_));
  NO3        u0383(.A(men_men_n411_), .B(men_men_n405_), .C(men_men_n401_), .Y(men_men_n412_));
  NO2        u0384(.A(men_men_n404_), .B(men_men_n312_), .Y(men_men_n413_));
  NOi32      u0385(.An(f), .Bn(d), .C(c), .Y(men_men_n414_));
  AOI220     u0386(.A0(men_men_n414_), .A1(men_men_n322_), .B0(men_men_n413_), .B1(men_men_n224_), .Y(men_men_n415_));
  NA3        u0387(.A(men_men_n415_), .B(men_men_n412_), .C(men_men_n397_), .Y(men_men_n416_));
  NO2        u0388(.A(men_men_n59_), .B(men_men_n120_), .Y(men_men_n417_));
  NA2        u0389(.A(men_men_n259_), .B(men_men_n417_), .Y(men_men_n418_));
  INV        u0390(.A(e), .Y(men_men_n419_));
  NA2        u0391(.A(men_men_n46_), .B(e), .Y(men_men_n420_));
  OAI220     u0392(.A0(men_men_n420_), .A1(men_men_n208_), .B0(men_men_n212_), .B1(men_men_n419_), .Y(men_men_n421_));
  AN2        u0393(.A(g), .B(e), .Y(men_men_n422_));
  NA3        u0394(.A(men_men_n422_), .B(men_men_n211_), .C(i), .Y(men_men_n423_));
  INV        u0395(.A(men_men_n423_), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n103_), .B(men_men_n419_), .Y(men_men_n425_));
  NO3        u0397(.A(men_men_n425_), .B(men_men_n424_), .C(men_men_n421_), .Y(men_men_n426_));
  NOi32      u0398(.An(h), .Bn(e), .C(g), .Y(men_men_n427_));
  NA3        u0399(.A(men_men_n427_), .B(men_men_n305_), .C(m), .Y(men_men_n428_));
  NOi21      u0400(.An(g), .B(h), .Y(men_men_n429_));
  AN3        u0401(.A(m), .B(l), .C(i), .Y(men_men_n430_));
  NA3        u0402(.A(men_men_n430_), .B(men_men_n429_), .C(e), .Y(men_men_n431_));
  AN3        u0403(.A(h), .B(g), .C(e), .Y(men_men_n432_));
  NA2        u0404(.A(men_men_n432_), .B(men_men_n100_), .Y(men_men_n433_));
  NO2        u0405(.A(men_men_n426_), .B(men_men_n418_), .Y(men_men_n434_));
  NA3        u0406(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n435_));
  NO2        u0407(.A(men_men_n435_), .B(men_men_n418_), .Y(men_men_n436_));
  NA3        u0408(.A(men_men_n406_), .B(men_men_n190_), .C(men_men_n86_), .Y(men_men_n437_));
  NAi31      u0409(.An(b), .B(c), .C(a), .Y(men_men_n438_));
  NO2        u0410(.A(men_men_n438_), .B(n), .Y(men_men_n439_));
  OAI210     u0411(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n440_), .B(men_men_n154_), .Y(men_men_n441_));
  NA2        u0413(.A(men_men_n441_), .B(men_men_n439_), .Y(men_men_n442_));
  INV        u0414(.A(men_men_n442_), .Y(men_men_n443_));
  NO4        u0415(.A(men_men_n443_), .B(men_men_n436_), .C(men_men_n434_), .D(men_men_n416_), .Y(men_men_n444_));
  NA2        u0416(.A(i), .B(g), .Y(men_men_n445_));
  NO3        u0417(.A(men_men_n289_), .B(men_men_n445_), .C(c), .Y(men_men_n446_));
  NOi21      u0418(.An(a), .B(n), .Y(men_men_n447_));
  NOi21      u0419(.An(d), .B(c), .Y(men_men_n448_));
  NA2        u0420(.A(men_men_n448_), .B(men_men_n447_), .Y(men_men_n449_));
  NA3        u0421(.A(i), .B(g), .C(f), .Y(men_men_n450_));
  OR2        u0422(.A(men_men_n450_), .B(men_men_n71_), .Y(men_men_n451_));
  NA3        u0423(.A(men_men_n430_), .B(men_men_n429_), .C(men_men_n190_), .Y(men_men_n452_));
  AOI210     u0424(.A0(men_men_n452_), .A1(men_men_n451_), .B0(men_men_n449_), .Y(men_men_n453_));
  AOI210     u0425(.A0(men_men_n446_), .A1(men_men_n304_), .B0(men_men_n453_), .Y(men_men_n454_));
  OR2        u0426(.A(n), .B(m), .Y(men_men_n455_));
  NO2        u0427(.A(men_men_n455_), .B(men_men_n159_), .Y(men_men_n456_));
  NO2        u0428(.A(men_men_n191_), .B(men_men_n154_), .Y(men_men_n457_));
  OAI210     u0429(.A0(men_men_n456_), .A1(men_men_n184_), .B0(men_men_n457_), .Y(men_men_n458_));
  INV        u0430(.A(men_men_n382_), .Y(men_men_n459_));
  NA3        u0431(.A(men_men_n459_), .B(men_men_n372_), .C(d), .Y(men_men_n460_));
  NO2        u0432(.A(men_men_n438_), .B(men_men_n49_), .Y(men_men_n461_));
  NO3        u0433(.A(men_men_n66_), .B(men_men_n116_), .C(e), .Y(men_men_n462_));
  NAi21      u0434(.An(k), .B(j), .Y(men_men_n463_));
  NA3        u0435(.A(i), .B(men_men_n462_), .C(men_men_n461_), .Y(men_men_n464_));
  NAi21      u0436(.An(e), .B(d), .Y(men_men_n465_));
  INV        u0437(.A(men_men_n465_), .Y(men_men_n466_));
  NO2        u0438(.A(men_men_n263_), .B(men_men_n222_), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n467_), .B(men_men_n466_), .C(men_men_n236_), .Y(men_men_n468_));
  NA4        u0440(.A(men_men_n468_), .B(men_men_n464_), .C(men_men_n460_), .D(men_men_n458_), .Y(men_men_n469_));
  NO2        u0441(.A(men_men_n345_), .B(men_men_n222_), .Y(men_men_n470_));
  NA2        u0442(.A(men_men_n470_), .B(men_men_n466_), .Y(men_men_n471_));
  NOi31      u0443(.An(n), .B(m), .C(k), .Y(men_men_n472_));
  AOI220     u0444(.A0(men_men_n472_), .A1(men_men_n398_), .B0(men_men_n230_), .B1(men_men_n50_), .Y(men_men_n473_));
  NAi31      u0445(.An(g), .B(f), .C(c), .Y(men_men_n474_));
  NA2        u0446(.A(men_men_n471_), .B(men_men_n323_), .Y(men_men_n475_));
  NOi41      u0447(.An(men_men_n454_), .B(men_men_n475_), .C(men_men_n469_), .D(men_men_n277_), .Y(men_men_n476_));
  NOi32      u0448(.An(c), .Bn(a), .C(b), .Y(men_men_n477_));
  NA2        u0449(.A(men_men_n477_), .B(men_men_n117_), .Y(men_men_n478_));
  AN2        u0450(.A(e), .B(d), .Y(men_men_n479_));
  INV        u0451(.A(men_men_n154_), .Y(men_men_n480_));
  NO2        u0452(.A(men_men_n136_), .B(men_men_n41_), .Y(men_men_n481_));
  NO2        u0453(.A(men_men_n66_), .B(e), .Y(men_men_n482_));
  NOi31      u0454(.An(j), .B(k), .C(i), .Y(men_men_n483_));
  NOi21      u0455(.An(men_men_n172_), .B(men_men_n483_), .Y(men_men_n484_));
  NA4        u0456(.A(men_men_n334_), .B(men_men_n484_), .C(men_men_n271_), .D(men_men_n123_), .Y(men_men_n485_));
  AOI220     u0457(.A0(men_men_n485_), .A1(men_men_n482_), .B0(men_men_n481_), .B1(men_men_n480_), .Y(men_men_n486_));
  NO2        u0458(.A(men_men_n486_), .B(men_men_n478_), .Y(men_men_n487_));
  NO2        u0459(.A(men_men_n218_), .B(men_men_n213_), .Y(men_men_n488_));
  NOi21      u0460(.An(a), .B(b), .Y(men_men_n489_));
  NA3        u0461(.A(e), .B(d), .C(c), .Y(men_men_n490_));
  NAi21      u0462(.An(men_men_n490_), .B(men_men_n489_), .Y(men_men_n491_));
  NO2        u0463(.A(men_men_n437_), .B(men_men_n212_), .Y(men_men_n492_));
  NOi21      u0464(.An(men_men_n491_), .B(men_men_n492_), .Y(men_men_n493_));
  AOI210     u0465(.A0(men_men_n280_), .A1(men_men_n488_), .B0(men_men_n493_), .Y(men_men_n494_));
  NO4        u0466(.A(men_men_n197_), .B(men_men_n106_), .C(men_men_n56_), .D(b), .Y(men_men_n495_));
  NA2        u0467(.A(men_men_n393_), .B(men_men_n160_), .Y(men_men_n496_));
  OR2        u0468(.A(k), .B(j), .Y(men_men_n497_));
  NA2        u0469(.A(l), .B(k), .Y(men_men_n498_));
  NA3        u0470(.A(men_men_n498_), .B(men_men_n497_), .C(men_men_n230_), .Y(men_men_n499_));
  AOI210     u0471(.A0(men_men_n243_), .A1(men_men_n348_), .B0(men_men_n86_), .Y(men_men_n500_));
  NOi21      u0472(.An(men_men_n499_), .B(men_men_n500_), .Y(men_men_n501_));
  OR3        u0473(.A(men_men_n501_), .B(men_men_n150_), .C(men_men_n140_), .Y(men_men_n502_));
  NA3        u0474(.A(men_men_n292_), .B(men_men_n133_), .C(men_men_n131_), .Y(men_men_n503_));
  NA2        u0475(.A(men_men_n406_), .B(men_men_n117_), .Y(men_men_n504_));
  NO4        u0476(.A(men_men_n504_), .B(men_men_n97_), .C(men_men_n116_), .D(e), .Y(men_men_n505_));
  NO3        u0477(.A(men_men_n437_), .B(men_men_n94_), .C(men_men_n136_), .Y(men_men_n506_));
  NO4        u0478(.A(men_men_n506_), .B(men_men_n505_), .C(men_men_n503_), .D(men_men_n335_), .Y(men_men_n507_));
  NA3        u0479(.A(men_men_n507_), .B(men_men_n502_), .C(men_men_n496_), .Y(men_men_n508_));
  NO4        u0480(.A(men_men_n508_), .B(men_men_n495_), .C(men_men_n494_), .D(men_men_n487_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n510_));
  NOi21      u0482(.An(d), .B(e), .Y(men_men_n511_));
  NO2        u0483(.A(men_men_n197_), .B(men_men_n56_), .Y(men_men_n512_));
  NAi31      u0484(.An(j), .B(l), .C(i), .Y(men_men_n513_));
  OAI210     u0485(.A0(men_men_n513_), .A1(men_men_n137_), .B0(men_men_n106_), .Y(men_men_n514_));
  NA3        u0486(.A(men_men_n514_), .B(men_men_n512_), .C(men_men_n511_), .Y(men_men_n515_));
  NO3        u0487(.A(men_men_n407_), .B(men_men_n354_), .C(men_men_n209_), .Y(men_men_n516_));
  NO2        u0488(.A(men_men_n407_), .B(men_men_n382_), .Y(men_men_n517_));
  NO4        u0489(.A(men_men_n517_), .B(men_men_n516_), .C(men_men_n193_), .D(men_men_n320_), .Y(men_men_n518_));
  NA4        u0490(.A(men_men_n518_), .B(men_men_n515_), .C(men_men_n510_), .D(men_men_n253_), .Y(men_men_n519_));
  OAI210     u0491(.A0(men_men_n132_), .A1(men_men_n130_), .B0(n), .Y(men_men_n520_));
  NO2        u0492(.A(men_men_n520_), .B(men_men_n136_), .Y(men_men_n521_));
  OA210      u0493(.A0(men_men_n313_), .A1(men_men_n521_), .B0(men_men_n200_), .Y(men_men_n522_));
  XO2        u0494(.A(i), .B(h), .Y(men_men_n523_));
  NA3        u0495(.A(men_men_n523_), .B(men_men_n167_), .C(n), .Y(men_men_n524_));
  NAi41      u0496(.An(men_men_n313_), .B(men_men_n524_), .C(men_men_n473_), .D(men_men_n395_), .Y(men_men_n525_));
  NAi31      u0497(.An(c), .B(f), .C(d), .Y(men_men_n526_));
  AOI210     u0498(.A0(men_men_n293_), .A1(men_men_n203_), .B0(men_men_n526_), .Y(men_men_n527_));
  NOi21      u0499(.An(men_men_n84_), .B(men_men_n527_), .Y(men_men_n528_));
  NA3        u0500(.A(men_men_n391_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n529_));
  NA2        u0501(.A(men_men_n237_), .B(men_men_n112_), .Y(men_men_n530_));
  AOI210     u0502(.A0(men_men_n530_), .A1(men_men_n189_), .B0(men_men_n526_), .Y(men_men_n531_));
  AOI210     u0503(.A0(men_men_n370_), .A1(men_men_n35_), .B0(men_men_n491_), .Y(men_men_n532_));
  NOi31      u0504(.An(men_men_n529_), .B(men_men_n532_), .C(men_men_n531_), .Y(men_men_n533_));
  AO220      u0505(.A0(men_men_n301_), .A1(men_men_n274_), .B0(men_men_n173_), .B1(men_men_n67_), .Y(men_men_n534_));
  NA3        u0506(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n535_), .B(men_men_n449_), .Y(men_men_n536_));
  NO2        u0508(.A(men_men_n536_), .B(men_men_n309_), .Y(men_men_n537_));
  NAi41      u0509(.An(men_men_n534_), .B(men_men_n537_), .C(men_men_n533_), .D(men_men_n528_), .Y(men_men_n538_));
  NO3        u0510(.A(men_men_n538_), .B(men_men_n522_), .C(men_men_n519_), .Y(men_men_n539_));
  NA4        u0511(.A(men_men_n539_), .B(men_men_n509_), .C(men_men_n476_), .D(men_men_n444_), .Y(men11));
  NO2        u0512(.A(men_men_n73_), .B(f), .Y(men_men_n541_));
  NA2        u0513(.A(j), .B(g), .Y(men_men_n542_));
  NAi31      u0514(.An(i), .B(m), .C(l), .Y(men_men_n543_));
  NA3        u0515(.A(m), .B(k), .C(j), .Y(men_men_n544_));
  OAI220     u0516(.A0(men_men_n544_), .A1(men_men_n136_), .B0(men_men_n543_), .B1(men_men_n542_), .Y(men_men_n545_));
  NA2        u0517(.A(men_men_n545_), .B(men_men_n541_), .Y(men_men_n546_));
  NOi32      u0518(.An(e), .Bn(b), .C(f), .Y(men_men_n547_));
  NA2        u0519(.A(men_men_n270_), .B(men_men_n117_), .Y(men_men_n548_));
  NA2        u0520(.A(men_men_n46_), .B(j), .Y(men_men_n549_));
  NO2        u0521(.A(men_men_n549_), .B(men_men_n315_), .Y(men_men_n550_));
  NAi31      u0522(.An(d), .B(e), .C(a), .Y(men_men_n551_));
  NO2        u0523(.A(men_men_n551_), .B(n), .Y(men_men_n552_));
  AOI220     u0524(.A0(men_men_n552_), .A1(men_men_n104_), .B0(men_men_n550_), .B1(men_men_n547_), .Y(men_men_n553_));
  NAi41      u0525(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n554_));
  AN2        u0526(.A(men_men_n554_), .B(men_men_n381_), .Y(men_men_n555_));
  AOI210     u0527(.A0(men_men_n555_), .A1(men_men_n407_), .B0(men_men_n283_), .Y(men_men_n556_));
  NA2        u0528(.A(j), .B(i), .Y(men_men_n557_));
  NAi31      u0529(.An(n), .B(m), .C(k), .Y(men_men_n558_));
  NO3        u0530(.A(men_men_n558_), .B(men_men_n557_), .C(men_men_n116_), .Y(men_men_n559_));
  NO4        u0531(.A(n), .B(d), .C(men_men_n120_), .D(a), .Y(men_men_n560_));
  OR2        u0532(.A(n), .B(c), .Y(men_men_n561_));
  NO2        u0533(.A(men_men_n561_), .B(men_men_n156_), .Y(men_men_n562_));
  NO2        u0534(.A(men_men_n562_), .B(men_men_n560_), .Y(men_men_n563_));
  NOi32      u0535(.An(g), .Bn(f), .C(i), .Y(men_men_n564_));
  AOI220     u0536(.A0(men_men_n564_), .A1(men_men_n102_), .B0(men_men_n545_), .B1(f), .Y(men_men_n565_));
  NO2        u0537(.A(men_men_n287_), .B(men_men_n49_), .Y(men_men_n566_));
  NO2        u0538(.A(men_men_n565_), .B(men_men_n563_), .Y(men_men_n567_));
  AOI210     u0539(.A0(men_men_n559_), .A1(men_men_n556_), .B0(men_men_n567_), .Y(men_men_n568_));
  NA2        u0540(.A(men_men_n146_), .B(men_men_n34_), .Y(men_men_n569_));
  OAI220     u0541(.A0(men_men_n569_), .A1(m), .B0(men_men_n549_), .B1(men_men_n243_), .Y(men_men_n570_));
  NOi41      u0542(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n571_));
  NAi32      u0543(.An(e), .Bn(b), .C(c), .Y(men_men_n572_));
  OR2        u0544(.A(men_men_n572_), .B(men_men_n86_), .Y(men_men_n573_));
  NA2        u0545(.A(men_men_n349_), .B(men_men_n573_), .Y(men_men_n574_));
  OA210      u0546(.A0(men_men_n574_), .A1(men_men_n571_), .B0(men_men_n570_), .Y(men_men_n575_));
  OAI220     u0547(.A0(men_men_n409_), .A1(men_men_n408_), .B0(men_men_n543_), .B1(men_men_n542_), .Y(men_men_n576_));
  NAi31      u0548(.An(d), .B(c), .C(a), .Y(men_men_n577_));
  NO2        u0549(.A(men_men_n577_), .B(n), .Y(men_men_n578_));
  NA3        u0550(.A(men_men_n578_), .B(men_men_n576_), .C(e), .Y(men_men_n579_));
  NO3        u0551(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n223_), .Y(men_men_n580_));
  NO2        u0552(.A(men_men_n240_), .B(men_men_n114_), .Y(men_men_n581_));
  OAI210     u0553(.A0(men_men_n580_), .A1(men_men_n410_), .B0(men_men_n581_), .Y(men_men_n582_));
  NA2        u0554(.A(men_men_n582_), .B(men_men_n579_), .Y(men_men_n583_));
  NO2        u0555(.A(men_men_n289_), .B(n), .Y(men_men_n584_));
  NO2        u0556(.A(men_men_n439_), .B(men_men_n584_), .Y(men_men_n585_));
  NA2        u0557(.A(men_men_n576_), .B(f), .Y(men_men_n586_));
  NAi32      u0558(.An(d), .Bn(a), .C(b), .Y(men_men_n587_));
  NO2        u0559(.A(men_men_n587_), .B(men_men_n49_), .Y(men_men_n588_));
  NA2        u0560(.A(h), .B(f), .Y(men_men_n589_));
  NO2        u0561(.A(men_men_n589_), .B(men_men_n97_), .Y(men_men_n590_));
  NO3        u0562(.A(men_men_n185_), .B(men_men_n182_), .C(g), .Y(men_men_n591_));
  AOI220     u0563(.A0(men_men_n591_), .A1(men_men_n58_), .B0(men_men_n590_), .B1(men_men_n588_), .Y(men_men_n592_));
  OAI210     u0564(.A0(men_men_n586_), .A1(men_men_n585_), .B0(men_men_n592_), .Y(men_men_n593_));
  AN3        u0565(.A(j), .B(h), .C(g), .Y(men_men_n594_));
  NA3        u0566(.A(f), .B(d), .C(b), .Y(men_men_n595_));
  NO4        u0567(.A(men_men_n595_), .B(men_men_n185_), .C(men_men_n182_), .D(g), .Y(men_men_n596_));
  NO4        u0568(.A(men_men_n596_), .B(men_men_n593_), .C(men_men_n583_), .D(men_men_n575_), .Y(men_men_n597_));
  AN4        u0569(.A(men_men_n597_), .B(men_men_n568_), .C(men_men_n553_), .D(men_men_n546_), .Y(men_men_n598_));
  INV        u0570(.A(k), .Y(men_men_n599_));
  NA3        u0571(.A(l), .B(men_men_n599_), .C(i), .Y(men_men_n600_));
  INV        u0572(.A(men_men_n600_), .Y(men_men_n601_));
  NA4        u0573(.A(men_men_n406_), .B(men_men_n429_), .C(men_men_n190_), .D(men_men_n117_), .Y(men_men_n602_));
  NAi32      u0574(.An(h), .Bn(f), .C(g), .Y(men_men_n603_));
  NAi41      u0575(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n604_));
  OAI210     u0576(.A0(men_men_n551_), .A1(n), .B0(men_men_n604_), .Y(men_men_n605_));
  NA2        u0577(.A(men_men_n605_), .B(m), .Y(men_men_n606_));
  NAi31      u0578(.An(h), .B(g), .C(f), .Y(men_men_n607_));
  OR3        u0579(.A(men_men_n607_), .B(men_men_n289_), .C(men_men_n49_), .Y(men_men_n608_));
  NA4        u0580(.A(men_men_n429_), .B(men_men_n125_), .C(men_men_n117_), .D(e), .Y(men_men_n609_));
  AN2        u0581(.A(men_men_n609_), .B(men_men_n608_), .Y(men_men_n610_));
  OA210      u0582(.A0(men_men_n606_), .A1(men_men_n603_), .B0(men_men_n610_), .Y(men_men_n611_));
  NO3        u0583(.A(men_men_n603_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n612_));
  NO4        u0584(.A(men_men_n607_), .B(men_men_n561_), .C(men_men_n156_), .D(men_men_n75_), .Y(men_men_n613_));
  OR2        u0585(.A(men_men_n613_), .B(men_men_n612_), .Y(men_men_n614_));
  NAi31      u0586(.An(men_men_n614_), .B(men_men_n611_), .C(men_men_n602_), .Y(men_men_n615_));
  NAi31      u0587(.An(f), .B(h), .C(g), .Y(men_men_n616_));
  NO4        u0588(.A(men_men_n325_), .B(men_men_n616_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n617_));
  NOi32      u0589(.An(b), .Bn(a), .C(c), .Y(men_men_n618_));
  NOi41      u0590(.An(men_men_n618_), .B(men_men_n363_), .C(men_men_n69_), .D(men_men_n121_), .Y(men_men_n619_));
  OR2        u0591(.A(men_men_n619_), .B(men_men_n617_), .Y(men_men_n620_));
  NOi32      u0592(.An(d), .Bn(a), .C(e), .Y(men_men_n621_));
  NA2        u0593(.A(men_men_n621_), .B(men_men_n117_), .Y(men_men_n622_));
  NO2        u0594(.A(n), .B(c), .Y(men_men_n623_));
  NA3        u0595(.A(men_men_n623_), .B(men_men_n29_), .C(m), .Y(men_men_n624_));
  NAi32      u0596(.An(n), .Bn(f), .C(m), .Y(men_men_n625_));
  NA3        u0597(.A(men_men_n625_), .B(men_men_n624_), .C(men_men_n622_), .Y(men_men_n626_));
  NOi32      u0598(.An(e), .Bn(a), .C(d), .Y(men_men_n627_));
  AOI210     u0599(.A0(men_men_n29_), .A1(d), .B0(men_men_n627_), .Y(men_men_n628_));
  AOI210     u0600(.A0(men_men_n628_), .A1(men_men_n222_), .B0(men_men_n569_), .Y(men_men_n629_));
  AOI210     u0601(.A0(men_men_n629_), .A1(men_men_n626_), .B0(men_men_n620_), .Y(men_men_n630_));
  OAI210     u0602(.A0(men_men_n258_), .A1(men_men_n89_), .B0(men_men_n630_), .Y(men_men_n631_));
  AOI210     u0603(.A0(men_men_n615_), .A1(men_men_n601_), .B0(men_men_n631_), .Y(men_men_n632_));
  NO3        u0604(.A(men_men_n332_), .B(men_men_n61_), .C(n), .Y(men_men_n633_));
  NA3        u0605(.A(men_men_n526_), .B(men_men_n180_), .C(men_men_n179_), .Y(men_men_n634_));
  NA2        u0606(.A(men_men_n474_), .B(men_men_n240_), .Y(men_men_n635_));
  OR2        u0607(.A(men_men_n635_), .B(men_men_n634_), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n76_), .B(men_men_n117_), .Y(men_men_n637_));
  NO2        u0609(.A(men_men_n637_), .B(men_men_n45_), .Y(men_men_n638_));
  AOI220     u0610(.A0(men_men_n638_), .A1(men_men_n556_), .B0(men_men_n636_), .B1(men_men_n633_), .Y(men_men_n639_));
  NO2        u0611(.A(men_men_n639_), .B(men_men_n89_), .Y(men_men_n640_));
  NA3        u0612(.A(men_men_n571_), .B(men_men_n350_), .C(men_men_n46_), .Y(men_men_n641_));
  NOi32      u0613(.An(e), .Bn(c), .C(f), .Y(men_men_n642_));
  NOi21      u0614(.An(f), .B(g), .Y(men_men_n643_));
  NO2        u0615(.A(men_men_n643_), .B(men_men_n220_), .Y(men_men_n644_));
  AOI220     u0616(.A0(men_men_n644_), .A1(men_men_n403_), .B0(men_men_n642_), .B1(men_men_n184_), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n645_), .B(men_men_n641_), .C(men_men_n187_), .Y(men_men_n646_));
  AOI210     u0618(.A0(men_men_n555_), .A1(men_men_n407_), .B0(men_men_n314_), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n647_), .B(men_men_n275_), .Y(men_men_n648_));
  NOi21      u0620(.An(j), .B(l), .Y(men_men_n649_));
  NAi21      u0621(.An(k), .B(h), .Y(men_men_n650_));
  NO2        u0622(.A(men_men_n650_), .B(men_men_n273_), .Y(men_men_n651_));
  NA2        u0623(.A(men_men_n651_), .B(men_men_n649_), .Y(men_men_n652_));
  OR2        u0624(.A(men_men_n652_), .B(men_men_n606_), .Y(men_men_n653_));
  NOi31      u0625(.An(m), .B(n), .C(k), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n649_), .B(men_men_n654_), .Y(men_men_n655_));
  AOI210     u0627(.A0(men_men_n407_), .A1(men_men_n381_), .B0(men_men_n314_), .Y(men_men_n656_));
  NAi21      u0628(.An(men_men_n655_), .B(men_men_n656_), .Y(men_men_n657_));
  NO2        u0629(.A(men_men_n289_), .B(men_men_n49_), .Y(men_men_n658_));
  NO2        u0630(.A(men_men_n325_), .B(men_men_n616_), .Y(men_men_n659_));
  NO2        u0631(.A(men_men_n551_), .B(men_men_n49_), .Y(men_men_n660_));
  AOI220     u0632(.A0(men_men_n660_), .A1(men_men_n659_), .B0(men_men_n658_), .B1(men_men_n590_), .Y(men_men_n661_));
  NA4        u0633(.A(men_men_n661_), .B(men_men_n657_), .C(men_men_n653_), .D(men_men_n648_), .Y(men_men_n662_));
  NA2        u0634(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n663_));
  NO2        u0635(.A(k), .B(men_men_n223_), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n547_), .B(men_men_n372_), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n549_), .B(men_men_n185_), .Y(men_men_n666_));
  NA3        u0638(.A(men_men_n572_), .B(men_men_n282_), .C(men_men_n151_), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n523_), .B(men_men_n167_), .Y(men_men_n668_));
  NO3        u0640(.A(men_men_n404_), .B(men_men_n668_), .C(men_men_n89_), .Y(men_men_n669_));
  AOI210     u0641(.A0(men_men_n667_), .A1(men_men_n666_), .B0(men_men_n669_), .Y(men_men_n670_));
  AN3        u0642(.A(f), .B(d), .C(b), .Y(men_men_n671_));
  NA3        u0643(.A(men_men_n523_), .B(men_men_n167_), .C(men_men_n223_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n242_), .B(men_men_n672_), .Y(men_men_n673_));
  NAi31      u0645(.An(m), .B(n), .C(k), .Y(men_men_n674_));
  OR2        u0646(.A(men_men_n140_), .B(men_men_n61_), .Y(men_men_n675_));
  OAI210     u0647(.A0(men_men_n675_), .A1(men_men_n674_), .B0(men_men_n260_), .Y(men_men_n676_));
  OAI210     u0648(.A0(men_men_n676_), .A1(men_men_n673_), .B0(j), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n677_), .B(men_men_n670_), .Y(men_men_n678_));
  NO4        u0650(.A(men_men_n678_), .B(men_men_n662_), .C(men_men_n646_), .D(men_men_n640_), .Y(men_men_n679_));
  NA2        u0651(.A(men_men_n391_), .B(men_men_n169_), .Y(men_men_n680_));
  NAi31      u0652(.An(g), .B(h), .C(f), .Y(men_men_n681_));
  OR3        u0653(.A(men_men_n681_), .B(men_men_n289_), .C(n), .Y(men_men_n682_));
  OA210      u0654(.A0(men_men_n551_), .A1(n), .B0(men_men_n604_), .Y(men_men_n683_));
  NA3        u0655(.A(men_men_n427_), .B(men_men_n125_), .C(men_men_n86_), .Y(men_men_n684_));
  OAI210     u0656(.A0(men_men_n683_), .A1(men_men_n93_), .B0(men_men_n684_), .Y(men_men_n685_));
  NOi21      u0657(.An(men_men_n682_), .B(men_men_n685_), .Y(men_men_n686_));
  AOI210     u0658(.A0(men_men_n686_), .A1(men_men_n680_), .B0(men_men_n544_), .Y(men_men_n687_));
  NO3        u0659(.A(g), .B(men_men_n222_), .C(men_men_n56_), .Y(men_men_n688_));
  NAi21      u0660(.An(h), .B(j), .Y(men_men_n689_));
  NO2        u0661(.A(men_men_n530_), .B(men_men_n89_), .Y(men_men_n690_));
  OAI210     u0662(.A0(men_men_n690_), .A1(men_men_n403_), .B0(men_men_n688_), .Y(men_men_n691_));
  OR2        u0663(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n692_));
  NA2        u0664(.A(men_men_n618_), .B(men_men_n352_), .Y(men_men_n693_));
  OA220      u0665(.A0(men_men_n655_), .A1(men_men_n693_), .B0(men_men_n652_), .B1(men_men_n692_), .Y(men_men_n694_));
  NA3        u0666(.A(men_men_n541_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n695_));
  AN2        u0667(.A(h), .B(f), .Y(men_men_n696_));
  NA2        u0668(.A(men_men_n696_), .B(men_men_n37_), .Y(men_men_n697_));
  AOI210     u0669(.A0(men_men_n587_), .A1(men_men_n438_), .B0(men_men_n49_), .Y(men_men_n698_));
  NA3        u0670(.A(men_men_n695_), .B(men_men_n694_), .C(men_men_n691_), .Y(men_men_n699_));
  NO2        u0671(.A(men_men_n262_), .B(f), .Y(men_men_n700_));
  NO2        u0672(.A(men_men_n643_), .B(men_men_n61_), .Y(men_men_n701_));
  NO2        u0673(.A(men_men_n701_), .B(men_men_n700_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n340_), .B(men_men_n146_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n137_), .B(men_men_n49_), .Y(men_men_n704_));
  AOI220     u0676(.A0(men_men_n704_), .A1(men_men_n547_), .B0(men_men_n372_), .B1(men_men_n117_), .Y(men_men_n705_));
  OA220      u0677(.A0(men_men_n705_), .A1(men_men_n569_), .B0(men_men_n370_), .B1(men_men_n115_), .Y(men_men_n706_));
  OAI210     u0678(.A0(men_men_n703_), .A1(men_men_n702_), .B0(men_men_n706_), .Y(men_men_n707_));
  NO3        u0679(.A(men_men_n414_), .B(men_men_n200_), .C(men_men_n199_), .Y(men_men_n708_));
  NA2        u0680(.A(men_men_n708_), .B(men_men_n240_), .Y(men_men_n709_));
  NA3        u0681(.A(men_men_n709_), .B(men_men_n264_), .C(j), .Y(men_men_n710_));
  NO3        u0682(.A(men_men_n474_), .B(men_men_n182_), .C(i), .Y(men_men_n711_));
  NA2        u0683(.A(men_men_n477_), .B(men_men_n86_), .Y(men_men_n712_));
  NO4        u0684(.A(men_men_n544_), .B(men_men_n712_), .C(men_men_n136_), .D(men_men_n222_), .Y(men_men_n713_));
  INV        u0685(.A(men_men_n713_), .Y(men_men_n714_));
  NA4        u0686(.A(men_men_n714_), .B(men_men_n710_), .C(men_men_n529_), .D(men_men_n412_), .Y(men_men_n715_));
  NO4        u0687(.A(men_men_n715_), .B(men_men_n707_), .C(men_men_n699_), .D(men_men_n687_), .Y(men_men_n716_));
  NA4        u0688(.A(men_men_n716_), .B(men_men_n679_), .C(men_men_n632_), .D(men_men_n598_), .Y(men08));
  NO2        u0689(.A(k), .B(h), .Y(men_men_n718_));
  AO210      u0690(.A0(men_men_n262_), .A1(men_men_n463_), .B0(men_men_n718_), .Y(men_men_n719_));
  NO2        u0691(.A(men_men_n719_), .B(men_men_n312_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n642_), .B(men_men_n86_), .Y(men_men_n721_));
  NA2        u0693(.A(men_men_n721_), .B(men_men_n474_), .Y(men_men_n722_));
  AOI210     u0694(.A0(men_men_n722_), .A1(men_men_n720_), .B0(men_men_n506_), .Y(men_men_n723_));
  NA2        u0695(.A(men_men_n86_), .B(men_men_n114_), .Y(men_men_n724_));
  NO2        u0696(.A(men_men_n724_), .B(men_men_n57_), .Y(men_men_n725_));
  NA2        u0697(.A(men_men_n595_), .B(men_men_n242_), .Y(men_men_n726_));
  NA2        u0698(.A(men_men_n726_), .B(men_men_n357_), .Y(men_men_n727_));
  AOI210     u0699(.A0(men_men_n595_), .A1(men_men_n163_), .B0(men_men_n86_), .Y(men_men_n728_));
  NA4        u0700(.A(men_men_n225_), .B(men_men_n146_), .C(men_men_n45_), .D(h), .Y(men_men_n729_));
  AN2        u0701(.A(l), .B(k), .Y(men_men_n730_));
  NA4        u0702(.A(men_men_n730_), .B(men_men_n112_), .C(men_men_n75_), .D(men_men_n223_), .Y(men_men_n731_));
  NA3        u0703(.A(men_men_n727_), .B(men_men_n723_), .C(men_men_n359_), .Y(men_men_n732_));
  AN2        u0704(.A(men_men_n552_), .B(men_men_n98_), .Y(men_men_n733_));
  NO4        u0705(.A(men_men_n182_), .B(men_men_n402_), .C(men_men_n116_), .D(g), .Y(men_men_n734_));
  AOI210     u0706(.A0(men_men_n734_), .A1(men_men_n726_), .B0(men_men_n536_), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n38_), .B(men_men_n222_), .Y(men_men_n736_));
  AOI220     u0708(.A0(men_men_n644_), .A1(men_men_n356_), .B0(men_men_n736_), .B1(men_men_n584_), .Y(men_men_n737_));
  NAi31      u0709(.An(men_men_n733_), .B(men_men_n737_), .C(men_men_n735_), .Y(men_men_n738_));
  NO2        u0710(.A(men_men_n555_), .B(men_men_n35_), .Y(men_men_n739_));
  OAI210     u0711(.A0(men_men_n572_), .A1(men_men_n47_), .B0(men_men_n675_), .Y(men_men_n740_));
  NO2        u0712(.A(men_men_n498_), .B(men_men_n137_), .Y(men_men_n741_));
  AOI210     u0713(.A0(men_men_n741_), .A1(men_men_n740_), .B0(men_men_n739_), .Y(men_men_n742_));
  NO3        u0714(.A(men_men_n332_), .B(men_men_n136_), .C(men_men_n41_), .Y(men_men_n743_));
  NAi21      u0715(.An(men_men_n743_), .B(men_men_n731_), .Y(men_men_n744_));
  NA2        u0716(.A(men_men_n719_), .B(men_men_n141_), .Y(men_men_n745_));
  AOI220     u0717(.A0(men_men_n745_), .A1(men_men_n413_), .B0(men_men_n744_), .B1(men_men_n78_), .Y(men_men_n746_));
  OAI210     u0718(.A0(men_men_n742_), .A1(men_men_n89_), .B0(men_men_n746_), .Y(men_men_n747_));
  NA3        u0719(.A(men_men_n709_), .B(men_men_n344_), .C(men_men_n394_), .Y(men_men_n748_));
  NA2        u0720(.A(men_men_n730_), .B(men_men_n230_), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n749_), .B(men_men_n339_), .Y(men_men_n750_));
  AOI210     u0722(.A0(men_men_n750_), .A1(men_men_n700_), .B0(men_men_n505_), .Y(men_men_n751_));
  NA3        u0723(.A(m), .B(l), .C(k), .Y(men_men_n752_));
  AOI210     u0724(.A0(men_men_n684_), .A1(men_men_n682_), .B0(men_men_n752_), .Y(men_men_n753_));
  NO2        u0725(.A(men_men_n554_), .B(men_men_n283_), .Y(men_men_n754_));
  NOi21      u0726(.An(men_men_n754_), .B(men_men_n548_), .Y(men_men_n755_));
  NA4        u0727(.A(men_men_n117_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n756_));
  NA3        u0728(.A(men_men_n125_), .B(men_men_n422_), .C(i), .Y(men_men_n757_));
  NO2        u0729(.A(men_men_n757_), .B(men_men_n756_), .Y(men_men_n758_));
  NO3        u0730(.A(men_men_n758_), .B(men_men_n755_), .C(men_men_n753_), .Y(men_men_n759_));
  NA3        u0731(.A(men_men_n759_), .B(men_men_n751_), .C(men_men_n748_), .Y(men_men_n760_));
  NO4        u0732(.A(men_men_n760_), .B(men_men_n747_), .C(men_men_n738_), .D(men_men_n732_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n644_), .B(men_men_n403_), .Y(men_men_n762_));
  NOi31      u0734(.An(g), .B(h), .C(f), .Y(men_men_n763_));
  NA2        u0735(.A(men_men_n660_), .B(men_men_n763_), .Y(men_men_n764_));
  AO210      u0736(.A0(men_men_n764_), .A1(men_men_n608_), .B0(men_men_n557_), .Y(men_men_n765_));
  NO3        u0737(.A(men_men_n407_), .B(men_men_n542_), .C(h), .Y(men_men_n766_));
  AOI210     u0738(.A0(men_men_n766_), .A1(men_men_n117_), .B0(men_men_n517_), .Y(men_men_n767_));
  NA4        u0739(.A(men_men_n767_), .B(men_men_n765_), .C(men_men_n762_), .D(men_men_n261_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n730_), .B(men_men_n75_), .Y(men_men_n769_));
  NO4        u0741(.A(men_men_n708_), .B(men_men_n182_), .C(n), .D(i), .Y(men_men_n770_));
  NOi21      u0742(.An(h), .B(j), .Y(men_men_n771_));
  NA2        u0743(.A(men_men_n771_), .B(f), .Y(men_men_n772_));
  NO2        u0744(.A(men_men_n772_), .B(men_men_n255_), .Y(men_men_n773_));
  NO3        u0745(.A(men_men_n773_), .B(men_men_n770_), .C(men_men_n711_), .Y(men_men_n774_));
  OAI220     u0746(.A0(men_men_n774_), .A1(men_men_n769_), .B0(men_men_n610_), .B1(men_men_n62_), .Y(men_men_n775_));
  AOI210     u0747(.A0(men_men_n768_), .A1(l), .B0(men_men_n775_), .Y(men_men_n776_));
  NO2        u0748(.A(j), .B(i), .Y(men_men_n777_));
  NA3        u0749(.A(men_men_n777_), .B(men_men_n82_), .C(l), .Y(men_men_n778_));
  NA2        u0750(.A(men_men_n777_), .B(men_men_n33_), .Y(men_men_n779_));
  NA2        u0751(.A(men_men_n432_), .B(men_men_n125_), .Y(men_men_n780_));
  OA220      u0752(.A0(men_men_n780_), .A1(men_men_n779_), .B0(men_men_n778_), .B1(men_men_n606_), .Y(men_men_n781_));
  NO3        u0753(.A(men_men_n158_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n782_));
  NO3        u0754(.A(men_men_n561_), .B(men_men_n156_), .C(men_men_n75_), .Y(men_men_n783_));
  NO3        u0755(.A(men_men_n498_), .B(men_men_n450_), .C(j), .Y(men_men_n784_));
  OAI210     u0756(.A0(men_men_n783_), .A1(men_men_n782_), .B0(men_men_n784_), .Y(men_men_n785_));
  OAI210     u0757(.A0(men_men_n764_), .A1(men_men_n62_), .B0(men_men_n785_), .Y(men_men_n786_));
  NA2        u0758(.A(k), .B(j), .Y(men_men_n787_));
  AOI210     u0759(.A0(men_men_n547_), .A1(n), .B0(men_men_n571_), .Y(men_men_n788_));
  NA2        u0760(.A(men_men_n788_), .B(men_men_n349_), .Y(men_men_n789_));
  NO3        u0761(.A(men_men_n182_), .B(men_men_n402_), .C(men_men_n116_), .Y(men_men_n790_));
  AOI220     u0762(.A0(men_men_n790_), .A1(men_men_n256_), .B0(men_men_n635_), .B1(men_men_n322_), .Y(men_men_n791_));
  NAi31      u0763(.An(men_men_n628_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n792_), .B(men_men_n791_), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n312_), .B(men_men_n141_), .Y(men_men_n794_));
  AOI220     u0766(.A0(men_men_n794_), .A1(men_men_n644_), .B0(men_men_n743_), .B1(men_men_n728_), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n784_), .B(men_men_n698_), .Y(men_men_n796_));
  NA2        u0768(.A(men_men_n796_), .B(men_men_n795_), .Y(men_men_n797_));
  OR3        u0769(.A(men_men_n797_), .B(men_men_n793_), .C(men_men_n786_), .Y(men_men_n798_));
  NA3        u0770(.A(men_men_n788_), .B(men_men_n349_), .C(men_men_n573_), .Y(men_men_n799_));
  NA4        u0771(.A(men_men_n799_), .B(men_men_n225_), .C(men_men_n463_), .D(men_men_n34_), .Y(men_men_n800_));
  NO4        u0772(.A(men_men_n498_), .B(men_men_n445_), .C(j), .D(f), .Y(men_men_n801_));
  NO2        u0773(.A(men_men_n729_), .B(men_men_n721_), .Y(men_men_n802_));
  AOI210     u0774(.A0(men_men_n801_), .A1(men_men_n268_), .B0(men_men_n802_), .Y(men_men_n803_));
  NA3        u0775(.A(men_men_n564_), .B(men_men_n305_), .C(h), .Y(men_men_n804_));
  NOi21      u0776(.An(men_men_n698_), .B(men_men_n804_), .Y(men_men_n805_));
  OAI220     u0777(.A0(men_men_n804_), .A1(men_men_n624_), .B0(men_men_n778_), .B1(men_men_n692_), .Y(men_men_n806_));
  INV        u0778(.A(men_men_n806_), .Y(men_men_n807_));
  NAi41      u0779(.An(men_men_n805_), .B(men_men_n807_), .C(men_men_n803_), .D(men_men_n800_), .Y(men_men_n808_));
  AOI220     u0780(.A0(men_men_n98_), .A1(men_men_n248_), .B0(men_men_n784_), .B1(men_men_n658_), .Y(men_men_n809_));
  NO2        u0781(.A(men_men_n683_), .B(men_men_n75_), .Y(men_men_n810_));
  AOI210     u0782(.A0(men_men_n801_), .A1(men_men_n810_), .B0(men_men_n346_), .Y(men_men_n811_));
  OAI210     u0783(.A0(men_men_n752_), .A1(men_men_n681_), .B0(men_men_n535_), .Y(men_men_n812_));
  NA3        u0784(.A(men_men_n259_), .B(men_men_n59_), .C(b), .Y(men_men_n813_));
  AOI220     u0785(.A0(men_men_n623_), .A1(men_men_n29_), .B0(men_men_n477_), .B1(men_men_n86_), .Y(men_men_n814_));
  NA2        u0786(.A(men_men_n814_), .B(men_men_n813_), .Y(men_men_n815_));
  NO2        u0787(.A(men_men_n804_), .B(men_men_n504_), .Y(men_men_n816_));
  AOI210     u0788(.A0(men_men_n815_), .A1(men_men_n812_), .B0(men_men_n816_), .Y(men_men_n817_));
  NA3        u0789(.A(men_men_n817_), .B(men_men_n811_), .C(men_men_n809_), .Y(men_men_n818_));
  NOi41      u0790(.An(men_men_n781_), .B(men_men_n818_), .C(men_men_n808_), .D(men_men_n798_), .Y(men_men_n819_));
  OR2        u0791(.A(men_men_n729_), .B(men_men_n242_), .Y(men_men_n820_));
  NO3        u0792(.A(men_men_n351_), .B(men_men_n314_), .C(men_men_n116_), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n821_), .B(men_men_n789_), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n823_));
  NO3        u0795(.A(men_men_n823_), .B(men_men_n779_), .C(men_men_n289_), .Y(men_men_n824_));
  NO3        u0796(.A(men_men_n542_), .B(men_men_n96_), .C(h), .Y(men_men_n825_));
  AOI210     u0797(.A0(men_men_n825_), .A1(men_men_n725_), .B0(men_men_n824_), .Y(men_men_n826_));
  NA4        u0798(.A(men_men_n826_), .B(men_men_n822_), .C(men_men_n820_), .D(men_men_n415_), .Y(men_men_n827_));
  OR2        u0799(.A(men_men_n681_), .B(men_men_n94_), .Y(men_men_n828_));
  NOi31      u0800(.An(b), .B(d), .C(a), .Y(men_men_n829_));
  NO2        u0801(.A(men_men_n829_), .B(men_men_n621_), .Y(men_men_n830_));
  NO2        u0802(.A(men_men_n830_), .B(n), .Y(men_men_n831_));
  NOi21      u0803(.An(men_men_n814_), .B(men_men_n831_), .Y(men_men_n832_));
  OAI220     u0804(.A0(men_men_n832_), .A1(men_men_n828_), .B0(men_men_n804_), .B1(men_men_n622_), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n572_), .B(men_men_n86_), .Y(men_men_n834_));
  NO3        u0806(.A(men_men_n643_), .B(men_men_n339_), .C(men_men_n121_), .Y(men_men_n835_));
  NOi21      u0807(.An(men_men_n835_), .B(men_men_n168_), .Y(men_men_n836_));
  AOI210     u0808(.A0(men_men_n821_), .A1(men_men_n834_), .B0(men_men_n836_), .Y(men_men_n837_));
  OAI210     u0809(.A0(men_men_n729_), .A1(men_men_n404_), .B0(men_men_n837_), .Y(men_men_n838_));
  NO2        u0810(.A(men_men_n708_), .B(n), .Y(men_men_n839_));
  AOI220     u0811(.A0(men_men_n794_), .A1(men_men_n688_), .B0(men_men_n839_), .B1(men_men_n720_), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n336_), .B(men_men_n247_), .Y(men_men_n841_));
  OAI210     u0813(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n841_), .Y(men_men_n842_));
  NA2        u0814(.A(men_men_n125_), .B(men_men_n86_), .Y(men_men_n843_));
  AOI210     u0815(.A0(men_men_n435_), .A1(men_men_n428_), .B0(men_men_n843_), .Y(men_men_n844_));
  NAi21      u0816(.An(men_men_n844_), .B(men_men_n842_), .Y(men_men_n845_));
  NA2        u0817(.A(men_men_n750_), .B(men_men_n34_), .Y(men_men_n846_));
  NAi21      u0818(.An(men_men_n756_), .B(men_men_n446_), .Y(men_men_n847_));
  NO2        u0819(.A(men_men_n283_), .B(i), .Y(men_men_n848_));
  NA2        u0820(.A(men_men_n734_), .B(men_men_n358_), .Y(men_men_n849_));
  OAI210     u0821(.A0(men_men_n613_), .A1(men_men_n612_), .B0(men_men_n373_), .Y(men_men_n850_));
  AN3        u0822(.A(men_men_n850_), .B(men_men_n849_), .C(men_men_n847_), .Y(men_men_n851_));
  NAi41      u0823(.An(men_men_n845_), .B(men_men_n851_), .C(men_men_n846_), .D(men_men_n840_), .Y(men_men_n852_));
  NO4        u0824(.A(men_men_n852_), .B(men_men_n838_), .C(men_men_n833_), .D(men_men_n827_), .Y(men_men_n853_));
  NA4        u0825(.A(men_men_n853_), .B(men_men_n819_), .C(men_men_n776_), .D(men_men_n761_), .Y(men09));
  INV        u0826(.A(men_men_n126_), .Y(men_men_n855_));
  NA2        u0827(.A(f), .B(e), .Y(men_men_n856_));
  NO2        u0828(.A(men_men_n235_), .B(men_men_n116_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n857_), .B(g), .Y(men_men_n858_));
  NA4        u0830(.A(men_men_n325_), .B(men_men_n484_), .C(men_men_n271_), .D(men_men_n123_), .Y(men_men_n859_));
  AOI210     u0831(.A0(men_men_n859_), .A1(g), .B0(men_men_n481_), .Y(men_men_n860_));
  AOI210     u0832(.A0(men_men_n860_), .A1(men_men_n858_), .B0(men_men_n856_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n456_), .B(e), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n861_), .B(men_men_n855_), .Y(men_men_n863_));
  NO2        u0835(.A(men_men_n212_), .B(men_men_n222_), .Y(men_men_n864_));
  NA3        u0836(.A(m), .B(l), .C(i), .Y(men_men_n865_));
  OAI220     u0837(.A0(men_men_n607_), .A1(men_men_n865_), .B0(men_men_n363_), .B1(men_men_n543_), .Y(men_men_n866_));
  NA4        u0838(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n867_));
  NAi31      u0839(.An(men_men_n866_), .B(men_men_n867_), .C(men_men_n451_), .Y(men_men_n868_));
  OR2        u0840(.A(men_men_n868_), .B(men_men_n864_), .Y(men_men_n869_));
  NA3        u0841(.A(men_men_n828_), .B(men_men_n586_), .C(men_men_n535_), .Y(men_men_n870_));
  OA210      u0842(.A0(men_men_n870_), .A1(men_men_n869_), .B0(men_men_n831_), .Y(men_men_n871_));
  INV        u0843(.A(men_men_n349_), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n873_));
  NOi31      u0845(.An(k), .B(m), .C(l), .Y(men_men_n874_));
  NO2        u0846(.A(men_men_n350_), .B(men_men_n874_), .Y(men_men_n875_));
  AOI210     u0847(.A0(men_men_n875_), .A1(men_men_n873_), .B0(men_men_n616_), .Y(men_men_n876_));
  NA2        u0848(.A(men_men_n813_), .B(men_men_n342_), .Y(men_men_n877_));
  NA2        u0849(.A(men_men_n352_), .B(men_men_n353_), .Y(men_men_n878_));
  OAI210     u0850(.A0(men_men_n212_), .A1(men_men_n222_), .B0(men_men_n878_), .Y(men_men_n879_));
  AOI220     u0851(.A0(men_men_n879_), .A1(men_men_n877_), .B0(men_men_n876_), .B1(men_men_n872_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n176_), .B(men_men_n118_), .Y(men_men_n881_));
  NA3        u0853(.A(men_men_n881_), .B(men_men_n719_), .C(men_men_n141_), .Y(men_men_n882_));
  NA3        u0854(.A(men_men_n882_), .B(men_men_n198_), .C(men_men_n31_), .Y(men_men_n883_));
  NA4        u0855(.A(men_men_n883_), .B(men_men_n880_), .C(men_men_n645_), .D(men_men_n84_), .Y(men_men_n884_));
  NO2        u0856(.A(men_men_n603_), .B(men_men_n513_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n885_), .B(men_men_n198_), .Y(men_men_n886_));
  NOi21      u0858(.An(f), .B(d), .Y(men_men_n887_));
  NA2        u0859(.A(men_men_n887_), .B(m), .Y(men_men_n888_));
  NO2        u0860(.A(men_men_n888_), .B(men_men_n52_), .Y(men_men_n889_));
  NOi32      u0861(.An(g), .Bn(f), .C(d), .Y(men_men_n890_));
  NA4        u0862(.A(men_men_n890_), .B(men_men_n623_), .C(men_men_n29_), .D(m), .Y(men_men_n891_));
  NOi21      u0863(.An(men_men_n326_), .B(men_men_n891_), .Y(men_men_n892_));
  AOI210     u0864(.A0(men_men_n889_), .A1(men_men_n562_), .B0(men_men_n892_), .Y(men_men_n893_));
  NA3        u0865(.A(men_men_n325_), .B(men_men_n271_), .C(men_men_n123_), .Y(men_men_n894_));
  AN2        u0866(.A(f), .B(d), .Y(men_men_n895_));
  NA3        u0867(.A(men_men_n489_), .B(men_men_n895_), .C(men_men_n86_), .Y(men_men_n896_));
  NO3        u0868(.A(men_men_n896_), .B(men_men_n75_), .C(men_men_n223_), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n298_), .B(men_men_n56_), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n894_), .B(men_men_n897_), .Y(men_men_n899_));
  NAi41      u0871(.An(men_men_n503_), .B(men_men_n899_), .C(men_men_n893_), .D(men_men_n886_), .Y(men_men_n900_));
  NO4        u0872(.A(men_men_n643_), .B(men_men_n137_), .C(men_men_n339_), .D(men_men_n159_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n674_), .B(men_men_n339_), .Y(men_men_n902_));
  AN2        u0874(.A(men_men_n902_), .B(men_men_n700_), .Y(men_men_n903_));
  NO3        u0875(.A(men_men_n903_), .B(men_men_n901_), .C(men_men_n244_), .Y(men_men_n904_));
  NA2        u0876(.A(men_men_n621_), .B(men_men_n86_), .Y(men_men_n905_));
  NO2        u0877(.A(men_men_n878_), .B(men_men_n905_), .Y(men_men_n906_));
  NO2        u0878(.A(men_men_n896_), .B(men_men_n440_), .Y(men_men_n907_));
  NOi41      u0879(.An(men_men_n233_), .B(men_men_n907_), .C(men_men_n906_), .D(men_men_n320_), .Y(men_men_n908_));
  NA2        u0880(.A(c), .B(men_men_n120_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n909_), .B(men_men_n419_), .Y(men_men_n910_));
  NA3        u0882(.A(men_men_n910_), .B(men_men_n525_), .C(f), .Y(men_men_n911_));
  OR2        u0883(.A(men_men_n681_), .B(men_men_n558_), .Y(men_men_n912_));
  INV        u0884(.A(men_men_n912_), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n830_), .B(men_men_n115_), .Y(men_men_n914_));
  NA2        u0886(.A(men_men_n914_), .B(men_men_n913_), .Y(men_men_n915_));
  NA4        u0887(.A(men_men_n915_), .B(men_men_n911_), .C(men_men_n908_), .D(men_men_n904_), .Y(men_men_n916_));
  NO4        u0888(.A(men_men_n916_), .B(men_men_n900_), .C(men_men_n884_), .D(men_men_n871_), .Y(men_men_n917_));
  OR2        u0889(.A(men_men_n896_), .B(men_men_n75_), .Y(men_men_n918_));
  NA2        u0890(.A(men_men_n116_), .B(j), .Y(men_men_n919_));
  NA2        u0891(.A(men_men_n857_), .B(g), .Y(men_men_n920_));
  AOI210     u0892(.A0(men_men_n920_), .A1(men_men_n306_), .B0(men_men_n918_), .Y(men_men_n921_));
  NO2        u0893(.A(men_men_n342_), .B(men_men_n867_), .Y(men_men_n922_));
  NO2        u0894(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n923_));
  NO2        u0895(.A(men_men_n240_), .B(men_men_n234_), .Y(men_men_n924_));
  AOI220     u0896(.A0(men_men_n924_), .A1(men_men_n237_), .B0(men_men_n319_), .B1(men_men_n923_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n440_), .B(men_men_n856_), .Y(men_men_n926_));
  NA2        u0898(.A(men_men_n926_), .B(men_men_n578_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n927_), .B(men_men_n925_), .Y(men_men_n928_));
  NA2        u0900(.A(e), .B(d), .Y(men_men_n929_));
  OAI220     u0901(.A0(men_men_n929_), .A1(c), .B0(men_men_n336_), .B1(d), .Y(men_men_n930_));
  NA3        u0902(.A(men_men_n930_), .B(men_men_n467_), .C(men_men_n523_), .Y(men_men_n931_));
  AOI210     u0903(.A0(men_men_n530_), .A1(men_men_n189_), .B0(men_men_n240_), .Y(men_men_n932_));
  AOI210     u0904(.A0(men_men_n644_), .A1(men_men_n356_), .B0(men_men_n932_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n298_), .B(men_men_n172_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n897_), .B(men_men_n934_), .Y(men_men_n935_));
  NA3        u0907(.A(men_men_n935_), .B(men_men_n933_), .C(men_men_n931_), .Y(men_men_n936_));
  NO4        u0908(.A(men_men_n936_), .B(men_men_n928_), .C(men_men_n922_), .D(men_men_n921_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n872_), .B(men_men_n31_), .Y(men_men_n938_));
  AO210      u0910(.A0(men_men_n938_), .A1(men_men_n721_), .B0(men_men_n226_), .Y(men_men_n939_));
  OAI220     u0911(.A0(men_men_n643_), .A1(men_men_n61_), .B0(men_men_n314_), .B1(j), .Y(men_men_n940_));
  AOI220     u0912(.A0(men_men_n940_), .A1(men_men_n902_), .B0(men_men_n633_), .B1(men_men_n642_), .Y(men_men_n941_));
  OAI210     u0913(.A0(men_men_n862_), .A1(men_men_n179_), .B0(men_men_n941_), .Y(men_men_n942_));
  OAI210     u0914(.A0(men_men_n857_), .A1(men_men_n934_), .B0(men_men_n890_), .Y(men_men_n943_));
  NO2        u0915(.A(men_men_n943_), .B(men_men_n624_), .Y(men_men_n944_));
  AOI210     u0916(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n270_), .Y(men_men_n945_));
  NO2        u0917(.A(men_men_n945_), .B(men_men_n891_), .Y(men_men_n946_));
  BUFFER     u0918(.A(men_men_n946_), .Y(men_men_n947_));
  NOi31      u0919(.An(men_men_n562_), .B(men_men_n888_), .C(men_men_n306_), .Y(men_men_n948_));
  NO4        u0920(.A(men_men_n948_), .B(men_men_n947_), .C(men_men_n944_), .D(men_men_n942_), .Y(men_men_n949_));
  AO220      u0921(.A0(men_men_n467_), .A1(men_men_n771_), .B0(men_men_n184_), .B1(f), .Y(men_men_n950_));
  OAI210     u0922(.A0(men_men_n950_), .A1(men_men_n470_), .B0(men_men_n930_), .Y(men_men_n951_));
  NO2        u0923(.A(men_men_n450_), .B(men_men_n71_), .Y(men_men_n952_));
  OAI210     u0924(.A0(men_men_n870_), .A1(men_men_n952_), .B0(men_men_n725_), .Y(men_men_n953_));
  AN4        u0925(.A(men_men_n953_), .B(men_men_n951_), .C(men_men_n949_), .D(men_men_n939_), .Y(men_men_n954_));
  NA4        u0926(.A(men_men_n954_), .B(men_men_n937_), .C(men_men_n917_), .D(men_men_n863_), .Y(men12));
  NO2        u0927(.A(men_men_n465_), .B(c), .Y(men_men_n956_));
  NO4        u0928(.A(men_men_n455_), .B(men_men_n262_), .C(men_men_n599_), .D(men_men_n223_), .Y(men_men_n957_));
  NA2        u0929(.A(men_men_n957_), .B(men_men_n956_), .Y(men_men_n958_));
  NA2        u0930(.A(men_men_n562_), .B(men_men_n952_), .Y(men_men_n959_));
  NO2        u0931(.A(men_men_n465_), .B(men_men_n120_), .Y(men_men_n960_));
  NO2        u0932(.A(men_men_n873_), .B(men_men_n363_), .Y(men_men_n961_));
  NO2        u0933(.A(men_men_n681_), .B(men_men_n388_), .Y(men_men_n962_));
  AOI220     u0934(.A0(men_men_n962_), .A1(men_men_n560_), .B0(men_men_n961_), .B1(men_men_n960_), .Y(men_men_n963_));
  NA4        u0935(.A(men_men_n963_), .B(men_men_n959_), .C(men_men_n958_), .D(men_men_n454_), .Y(men_men_n964_));
  AOI210     u0936(.A0(men_men_n243_), .A1(men_men_n348_), .B0(men_men_n209_), .Y(men_men_n965_));
  OR2        u0937(.A(men_men_n965_), .B(men_men_n957_), .Y(men_men_n966_));
  AOI210     u0938(.A0(men_men_n345_), .A1(men_men_n400_), .B0(men_men_n223_), .Y(men_men_n967_));
  OAI210     u0939(.A0(men_men_n967_), .A1(men_men_n966_), .B0(men_men_n414_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n663_), .B(men_men_n273_), .Y(men_men_n969_));
  NO2        u0941(.A(men_men_n607_), .B(men_men_n865_), .Y(men_men_n970_));
  AOI220     u0942(.A0(men_men_n970_), .A1(men_men_n584_), .B0(men_men_n841_), .B1(men_men_n969_), .Y(men_men_n971_));
  NO2        u0943(.A(men_men_n158_), .B(men_men_n247_), .Y(men_men_n972_));
  NA3        u0944(.A(men_men_n972_), .B(men_men_n250_), .C(i), .Y(men_men_n973_));
  NA3        u0945(.A(men_men_n973_), .B(men_men_n971_), .C(men_men_n968_), .Y(men_men_n974_));
  OR2        u0946(.A(men_men_n337_), .B(men_men_n960_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n975_), .B(men_men_n364_), .Y(men_men_n976_));
  NO3        u0948(.A(men_men_n137_), .B(men_men_n159_), .C(men_men_n223_), .Y(men_men_n977_));
  NA2        u0949(.A(men_men_n977_), .B(men_men_n547_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n978_), .B(men_men_n976_), .Y(men_men_n979_));
  NO3        u0951(.A(men_men_n686_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n980_));
  NO4        u0952(.A(men_men_n980_), .B(men_men_n979_), .C(men_men_n974_), .D(men_men_n964_), .Y(men_men_n981_));
  NO2        u0953(.A(men_men_n378_), .B(men_men_n377_), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n604_), .B(men_men_n73_), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n572_), .B(men_men_n151_), .Y(men_men_n984_));
  NOi21      u0956(.An(men_men_n34_), .B(men_men_n674_), .Y(men_men_n985_));
  AOI220     u0957(.A0(men_men_n985_), .A1(men_men_n984_), .B0(men_men_n983_), .B1(men_men_n982_), .Y(men_men_n986_));
  OAI210     u0958(.A0(men_men_n260_), .A1(men_men_n45_), .B0(men_men_n986_), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n446_), .B(men_men_n275_), .Y(men_men_n988_));
  NO3        u0960(.A(men_men_n843_), .B(men_men_n91_), .C(men_men_n419_), .Y(men_men_n989_));
  NAi21      u0961(.An(men_men_n989_), .B(men_men_n988_), .Y(men_men_n990_));
  NO2        u0962(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n991_));
  NO2        u0963(.A(men_men_n520_), .B(men_men_n314_), .Y(men_men_n992_));
  INV        u0964(.A(men_men_n992_), .Y(men_men_n993_));
  NO2        u0965(.A(men_men_n993_), .B(men_men_n151_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n654_), .B(men_men_n373_), .Y(men_men_n995_));
  OAI210     u0967(.A0(men_men_n757_), .A1(men_men_n995_), .B0(men_men_n375_), .Y(men_men_n996_));
  NO4        u0968(.A(men_men_n996_), .B(men_men_n994_), .C(men_men_n990_), .D(men_men_n987_), .Y(men_men_n997_));
  NA2        u0969(.A(men_men_n356_), .B(g), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n169_), .B(i), .Y(men_men_n999_));
  NO2        u0971(.A(men_men_n151_), .B(men_men_n86_), .Y(men_men_n1000_));
  OR2        u0972(.A(men_men_n1000_), .B(men_men_n571_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n572_), .B(men_men_n392_), .Y(men_men_n1002_));
  AOI210     u0974(.A0(men_men_n1002_), .A1(n), .B0(men_men_n1001_), .Y(men_men_n1003_));
  NO2        u0975(.A(men_men_n1003_), .B(men_men_n998_), .Y(men_men_n1004_));
  NO2        u0976(.A(men_men_n681_), .B(men_men_n513_), .Y(men_men_n1005_));
  NA3        u0977(.A(men_men_n352_), .B(men_men_n649_), .C(i), .Y(men_men_n1006_));
  OAI210     u0978(.A0(men_men_n450_), .A1(men_men_n325_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  OAI220     u0979(.A0(men_men_n1007_), .A1(men_men_n1005_), .B0(men_men_n698_), .B1(men_men_n783_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n627_), .B(men_men_n117_), .Y(men_men_n1009_));
  OR3        u0981(.A(men_men_n325_), .B(men_men_n445_), .C(f), .Y(men_men_n1010_));
  NA3        u0982(.A(men_men_n649_), .B(men_men_n82_), .C(i), .Y(men_men_n1011_));
  OA220      u0983(.A0(men_men_n1011_), .A1(men_men_n1009_), .B0(men_men_n1010_), .B1(men_men_n606_), .Y(men_men_n1012_));
  NA3        u0984(.A(men_men_n338_), .B(men_men_n122_), .C(g), .Y(men_men_n1013_));
  AOI210     u0985(.A0(men_men_n697_), .A1(men_men_n1013_), .B0(m), .Y(men_men_n1014_));
  OAI210     u0986(.A0(men_men_n1014_), .A1(men_men_n961_), .B0(men_men_n337_), .Y(men_men_n1015_));
  NA2        u0987(.A(men_men_n712_), .B(men_men_n905_), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n867_), .B(men_men_n451_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n231_), .B(men_men_n79_), .Y(men_men_n1018_));
  NA3        u0990(.A(men_men_n1018_), .B(men_men_n1011_), .C(men_men_n1010_), .Y(men_men_n1019_));
  AOI220     u0991(.A0(men_men_n1019_), .A1(men_men_n268_), .B0(men_men_n1017_), .B1(men_men_n1016_), .Y(men_men_n1020_));
  NA4        u0992(.A(men_men_n1020_), .B(men_men_n1015_), .C(men_men_n1012_), .D(men_men_n1008_), .Y(men_men_n1021_));
  NA2        u0993(.A(men_men_n969_), .B(men_men_n248_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n685_), .B(men_men_n90_), .Y(men_men_n1023_));
  NO2        u0995(.A(men_men_n473_), .B(men_men_n223_), .Y(men_men_n1024_));
  AOI220     u0996(.A0(men_men_n1024_), .A1(men_men_n393_), .B0(men_men_n975_), .B1(men_men_n227_), .Y(men_men_n1025_));
  AOI220     u0997(.A0(men_men_n962_), .A1(men_men_n972_), .B0(men_men_n605_), .B1(men_men_n92_), .Y(men_men_n1026_));
  NA4        u0998(.A(men_men_n1026_), .B(men_men_n1025_), .C(men_men_n1023_), .D(men_men_n1022_), .Y(men_men_n1027_));
  NA2        u0999(.A(men_men_n1017_), .B(men_men_n560_), .Y(men_men_n1028_));
  AOI210     u1000(.A0(men_men_n431_), .A1(men_men_n423_), .B0(men_men_n843_), .Y(men_men_n1029_));
  OAI210     u1001(.A0(men_men_n378_), .A1(men_men_n377_), .B0(men_men_n113_), .Y(men_men_n1030_));
  AOI210     u1002(.A0(men_men_n1030_), .A1(men_men_n552_), .B0(men_men_n1029_), .Y(men_men_n1031_));
  NA2        u1003(.A(men_men_n1014_), .B(men_men_n960_), .Y(men_men_n1032_));
  NO3        u1004(.A(men_men_n919_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1033_));
  AOI220     u1005(.A0(men_men_n1033_), .A1(men_men_n647_), .B0(men_men_n666_), .B1(men_men_n547_), .Y(men_men_n1034_));
  NA4        u1006(.A(men_men_n1034_), .B(men_men_n1032_), .C(men_men_n1031_), .D(men_men_n1028_), .Y(men_men_n1035_));
  NO4        u1007(.A(men_men_n1035_), .B(men_men_n1027_), .C(men_men_n1021_), .D(men_men_n1004_), .Y(men_men_n1036_));
  NAi31      u1008(.An(men_men_n147_), .B(men_men_n432_), .C(n), .Y(men_men_n1037_));
  NO3        u1009(.A(men_men_n130_), .B(men_men_n350_), .C(men_men_n874_), .Y(men_men_n1038_));
  NO2        u1010(.A(men_men_n1038_), .B(men_men_n1037_), .Y(men_men_n1039_));
  NO3        u1011(.A(men_men_n283_), .B(men_men_n147_), .C(men_men_n419_), .Y(men_men_n1040_));
  AOI210     u1012(.A0(men_men_n1040_), .A1(men_men_n514_), .B0(men_men_n1039_), .Y(men_men_n1041_));
  NA2        u1013(.A(men_men_n506_), .B(i), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n1042_), .B(men_men_n1041_), .Y(men_men_n1043_));
  NA2        u1015(.A(men_men_n240_), .B(men_men_n180_), .Y(men_men_n1044_));
  NO3        u1016(.A(men_men_n322_), .B(men_men_n456_), .C(men_men_n184_), .Y(men_men_n1045_));
  NOi31      u1017(.An(men_men_n1044_), .B(men_men_n1045_), .C(men_men_n223_), .Y(men_men_n1046_));
  NAi21      u1018(.An(men_men_n572_), .B(men_men_n1024_), .Y(men_men_n1047_));
  NA2        u1019(.A(men_men_n449_), .B(men_men_n905_), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n450_), .B(men_men_n325_), .C(men_men_n75_), .Y(men_men_n1049_));
  AOI220     u1021(.A0(men_men_n1049_), .A1(men_men_n1048_), .B0(men_men_n495_), .B1(g), .Y(men_men_n1050_));
  NA2        u1022(.A(men_men_n1050_), .B(men_men_n1047_), .Y(men_men_n1051_));
  OAI220     u1023(.A0(men_men_n1037_), .A1(men_men_n243_), .B0(men_men_n1006_), .B1(men_men_n622_), .Y(men_men_n1052_));
  NO2        u1024(.A(men_men_n682_), .B(men_men_n388_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n965_), .B(men_men_n956_), .Y(men_men_n1054_));
  NO3        u1026(.A(men_men_n561_), .B(men_men_n156_), .C(men_men_n222_), .Y(men_men_n1055_));
  OAI210     u1027(.A0(men_men_n1055_), .A1(men_men_n541_), .B0(men_men_n389_), .Y(men_men_n1056_));
  OAI220     u1028(.A0(men_men_n962_), .A1(men_men_n970_), .B0(men_men_n562_), .B1(men_men_n439_), .Y(men_men_n1057_));
  NA4        u1029(.A(men_men_n1057_), .B(men_men_n1056_), .C(men_men_n1054_), .D(men_men_n641_), .Y(men_men_n1058_));
  OAI210     u1030(.A0(men_men_n965_), .A1(men_men_n957_), .B0(men_men_n1044_), .Y(men_men_n1059_));
  NA3        u1031(.A(men_men_n1002_), .B(men_men_n500_), .C(men_men_n46_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n391_), .B(men_men_n389_), .Y(men_men_n1061_));
  NA4        u1033(.A(men_men_n1061_), .B(men_men_n1060_), .C(men_men_n1059_), .D(men_men_n284_), .Y(men_men_n1062_));
  OR4        u1034(.A(men_men_n1062_), .B(men_men_n1058_), .C(men_men_n1053_), .D(men_men_n1052_), .Y(men_men_n1063_));
  NO4        u1035(.A(men_men_n1063_), .B(men_men_n1051_), .C(men_men_n1046_), .D(men_men_n1043_), .Y(men_men_n1064_));
  NA4        u1036(.A(men_men_n1064_), .B(men_men_n1036_), .C(men_men_n997_), .D(men_men_n981_), .Y(men13));
  NA2        u1037(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1066_));
  AN2        u1038(.A(c), .B(b), .Y(men_men_n1067_));
  NA3        u1039(.A(men_men_n259_), .B(men_men_n1067_), .C(m), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n511_), .B(f), .Y(men_men_n1069_));
  NO4        u1041(.A(men_men_n1069_), .B(men_men_n1068_), .C(men_men_n1066_), .D(men_men_n600_), .Y(men_men_n1070_));
  NA2        u1042(.A(men_men_n275_), .B(men_men_n1067_), .Y(men_men_n1071_));
  NO4        u1043(.A(men_men_n1071_), .B(men_men_n1069_), .C(men_men_n999_), .D(a), .Y(men_men_n1072_));
  NAi32      u1044(.An(d), .Bn(c), .C(e), .Y(men_men_n1073_));
  NA2        u1045(.A(men_men_n146_), .B(men_men_n45_), .Y(men_men_n1074_));
  NO4        u1046(.A(men_men_n1074_), .B(men_men_n1073_), .C(men_men_n607_), .D(men_men_n321_), .Y(men_men_n1075_));
  NA2        u1047(.A(men_men_n689_), .B(men_men_n234_), .Y(men_men_n1076_));
  NA2        u1048(.A(men_men_n422_), .B(men_men_n222_), .Y(men_men_n1077_));
  AN2        u1049(.A(d), .B(c), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n1078_), .B(men_men_n120_), .Y(men_men_n1079_));
  NO4        u1051(.A(men_men_n1079_), .B(men_men_n1077_), .C(men_men_n185_), .D(men_men_n176_), .Y(men_men_n1080_));
  NA2        u1052(.A(men_men_n511_), .B(c), .Y(men_men_n1081_));
  NO4        u1053(.A(men_men_n1074_), .B(men_men_n603_), .C(men_men_n1081_), .D(men_men_n321_), .Y(men_men_n1082_));
  AO210      u1054(.A0(men_men_n1080_), .A1(men_men_n1076_), .B0(men_men_n1082_), .Y(men_men_n1083_));
  OR4        u1055(.A(men_men_n1083_), .B(men_men_n1075_), .C(men_men_n1072_), .D(men_men_n1070_), .Y(men_men_n1084_));
  NAi32      u1056(.An(f), .Bn(e), .C(c), .Y(men_men_n1085_));
  NO2        u1057(.A(men_men_n1085_), .B(men_men_n153_), .Y(men_men_n1086_));
  NA2        u1058(.A(men_men_n1086_), .B(g), .Y(men_men_n1087_));
  OR3        u1059(.A(men_men_n234_), .B(men_men_n185_), .C(men_men_n176_), .Y(men_men_n1088_));
  NO2        u1060(.A(men_men_n1088_), .B(men_men_n1087_), .Y(men_men_n1089_));
  NO2        u1061(.A(men_men_n1081_), .B(men_men_n321_), .Y(men_men_n1090_));
  NO2        u1062(.A(j), .B(men_men_n45_), .Y(men_men_n1091_));
  NA2        u1063(.A(men_men_n651_), .B(men_men_n1091_), .Y(men_men_n1092_));
  NOi21      u1064(.An(men_men_n1090_), .B(men_men_n1092_), .Y(men_men_n1093_));
  NO2        u1065(.A(men_men_n787_), .B(men_men_n116_), .Y(men_men_n1094_));
  NOi41      u1066(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1095_));
  NA2        u1067(.A(men_men_n1095_), .B(men_men_n1094_), .Y(men_men_n1096_));
  NO2        u1068(.A(men_men_n1096_), .B(men_men_n1087_), .Y(men_men_n1097_));
  OR3        u1069(.A(e), .B(d), .C(c), .Y(men_men_n1098_));
  NA3        u1070(.A(k), .B(j), .C(i), .Y(men_men_n1099_));
  NO3        u1071(.A(men_men_n1099_), .B(men_men_n321_), .C(men_men_n93_), .Y(men_men_n1100_));
  NOi21      u1072(.An(men_men_n1100_), .B(men_men_n1098_), .Y(men_men_n1101_));
  OR4        u1073(.A(men_men_n1101_), .B(men_men_n1097_), .C(men_men_n1093_), .D(men_men_n1089_), .Y(men_men_n1102_));
  NA3        u1074(.A(men_men_n479_), .B(men_men_n344_), .C(men_men_n56_), .Y(men_men_n1103_));
  NO2        u1075(.A(men_men_n1103_), .B(men_men_n1092_), .Y(men_men_n1104_));
  NO4        u1076(.A(men_men_n1103_), .B(men_men_n603_), .C(men_men_n463_), .D(men_men_n45_), .Y(men_men_n1105_));
  NO2        u1077(.A(f), .B(c), .Y(men_men_n1106_));
  NOi21      u1078(.An(men_men_n1106_), .B(men_men_n455_), .Y(men_men_n1107_));
  NA2        u1079(.A(men_men_n1107_), .B(men_men_n59_), .Y(men_men_n1108_));
  OR2        u1080(.A(k), .B(i), .Y(men_men_n1109_));
  NO3        u1081(.A(men_men_n1109_), .B(men_men_n254_), .C(l), .Y(men_men_n1110_));
  NOi31      u1082(.An(men_men_n1110_), .B(men_men_n1108_), .C(j), .Y(men_men_n1111_));
  OR3        u1083(.A(men_men_n1111_), .B(men_men_n1105_), .C(men_men_n1104_), .Y(men_men_n1112_));
  OR3        u1084(.A(men_men_n1112_), .B(men_men_n1102_), .C(men_men_n1084_), .Y(men02));
  OR2        u1085(.A(l), .B(k), .Y(men_men_n1114_));
  OR3        u1086(.A(h), .B(g), .C(f), .Y(men_men_n1115_));
  OR3        u1087(.A(n), .B(m), .C(i), .Y(men_men_n1116_));
  NO4        u1088(.A(men_men_n1116_), .B(men_men_n1115_), .C(men_men_n1114_), .D(men_men_n1098_), .Y(men_men_n1117_));
  NOi31      u1089(.An(e), .B(d), .C(c), .Y(men_men_n1118_));
  AOI210     u1090(.A0(men_men_n1100_), .A1(men_men_n1118_), .B0(men_men_n1075_), .Y(men_men_n1119_));
  AN3        u1091(.A(g), .B(f), .C(c), .Y(men_men_n1120_));
  NA3        u1092(.A(men_men_n1120_), .B(men_men_n479_), .C(h), .Y(men_men_n1121_));
  OR2        u1093(.A(men_men_n1099_), .B(men_men_n321_), .Y(men_men_n1122_));
  OR2        u1094(.A(men_men_n1122_), .B(men_men_n1121_), .Y(men_men_n1123_));
  NO3        u1095(.A(men_men_n1103_), .B(men_men_n1074_), .C(men_men_n603_), .Y(men_men_n1124_));
  NO2        u1096(.A(men_men_n1124_), .B(men_men_n1089_), .Y(men_men_n1125_));
  NA3        u1097(.A(l), .B(k), .C(j), .Y(men_men_n1126_));
  NA2        u1098(.A(i), .B(h), .Y(men_men_n1127_));
  NO3        u1099(.A(men_men_n1127_), .B(men_men_n1126_), .C(men_men_n137_), .Y(men_men_n1128_));
  NO3        u1100(.A(men_men_n148_), .B(men_men_n296_), .C(men_men_n223_), .Y(men_men_n1129_));
  AOI210     u1101(.A0(men_men_n1129_), .A1(men_men_n1128_), .B0(men_men_n1093_), .Y(men_men_n1130_));
  NA3        u1102(.A(c), .B(b), .C(a), .Y(men_men_n1131_));
  NO3        u1103(.A(men_men_n1131_), .B(men_men_n929_), .C(men_men_n222_), .Y(men_men_n1132_));
  NO4        u1104(.A(men_men_n1099_), .B(men_men_n314_), .C(men_men_n49_), .D(men_men_n116_), .Y(men_men_n1133_));
  AOI210     u1105(.A0(men_men_n1133_), .A1(men_men_n1132_), .B0(men_men_n1104_), .Y(men_men_n1134_));
  AN4        u1106(.A(men_men_n1134_), .B(men_men_n1130_), .C(men_men_n1125_), .D(men_men_n1123_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n1079_), .B(men_men_n1077_), .Y(men_men_n1136_));
  NA2        u1108(.A(men_men_n1096_), .B(men_men_n1088_), .Y(men_men_n1137_));
  AOI210     u1109(.A0(men_men_n1137_), .A1(men_men_n1136_), .B0(men_men_n1070_), .Y(men_men_n1138_));
  NAi41      u1110(.An(men_men_n1117_), .B(men_men_n1138_), .C(men_men_n1135_), .D(men_men_n1119_), .Y(men03));
  NO2        u1111(.A(men_men_n543_), .B(men_men_n616_), .Y(men_men_n1140_));
  NA4        u1112(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n222_), .Y(men_men_n1141_));
  NA4        u1113(.A(men_men_n594_), .B(m), .C(men_men_n116_), .D(men_men_n222_), .Y(men_men_n1142_));
  NA3        u1114(.A(men_men_n1142_), .B(men_men_n379_), .C(men_men_n1141_), .Y(men_men_n1143_));
  NO3        u1115(.A(men_men_n1143_), .B(men_men_n1140_), .C(men_men_n1030_), .Y(men_men_n1144_));
  NOi41      u1116(.An(men_men_n828_), .B(men_men_n879_), .C(men_men_n868_), .D(men_men_n736_), .Y(men_men_n1145_));
  OAI220     u1117(.A0(men_men_n1145_), .A1(men_men_n712_), .B0(men_men_n1144_), .B1(men_men_n604_), .Y(men_men_n1146_));
  NA4        u1118(.A(i), .B(men_men_n1118_), .C(men_men_n352_), .D(men_men_n344_), .Y(men_men_n1147_));
  OAI210     u1119(.A0(men_men_n843_), .A1(men_men_n433_), .B0(men_men_n1147_), .Y(men_men_n1148_));
  NOi31      u1120(.An(m), .B(n), .C(f), .Y(men_men_n1149_));
  NA2        u1121(.A(men_men_n1149_), .B(men_men_n51_), .Y(men_men_n1150_));
  AN2        u1122(.A(e), .B(c), .Y(men_men_n1151_));
  NO2        u1123(.A(men_men_n912_), .B(men_men_n438_), .Y(men_men_n1152_));
  NA2        u1124(.A(men_men_n523_), .B(l), .Y(men_men_n1153_));
  NOi31      u1125(.An(men_men_n890_), .B(men_men_n1068_), .C(men_men_n1153_), .Y(men_men_n1154_));
  NO4        u1126(.A(men_men_n1154_), .B(men_men_n1152_), .C(men_men_n1148_), .D(men_men_n1029_), .Y(men_men_n1155_));
  NO2        u1127(.A(men_men_n296_), .B(a), .Y(men_men_n1156_));
  INV        u1128(.A(men_men_n1075_), .Y(men_men_n1157_));
  NO2        u1129(.A(men_men_n1127_), .B(men_men_n498_), .Y(men_men_n1158_));
  NO2        u1130(.A(men_men_n89_), .B(g), .Y(men_men_n1159_));
  AOI210     u1131(.A0(men_men_n1159_), .A1(men_men_n1158_), .B0(men_men_n1110_), .Y(men_men_n1160_));
  OR2        u1132(.A(men_men_n1160_), .B(men_men_n1108_), .Y(men_men_n1161_));
  NA3        u1133(.A(men_men_n1161_), .B(men_men_n1157_), .C(men_men_n1155_), .Y(men_men_n1162_));
  NO4        u1134(.A(men_men_n1162_), .B(men_men_n1146_), .C(men_men_n845_), .D(men_men_n583_), .Y(men_men_n1163_));
  NA2        u1135(.A(c), .B(b), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n724_), .B(men_men_n1164_), .Y(men_men_n1165_));
  OAI210     u1137(.A0(men_men_n888_), .A1(men_men_n860_), .B0(men_men_n426_), .Y(men_men_n1166_));
  OAI210     u1138(.A0(men_men_n1166_), .A1(men_men_n889_), .B0(men_men_n1165_), .Y(men_men_n1167_));
  NA3        u1139(.A(men_men_n439_), .B(men_men_n576_), .C(f), .Y(men_men_n1168_));
  OAI210     u1140(.A0(men_men_n566_), .A1(men_men_n39_), .B0(men_men_n1156_), .Y(men_men_n1169_));
  NA2        u1141(.A(men_men_n1169_), .B(men_men_n1168_), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n271_), .B(men_men_n123_), .Y(men_men_n1171_));
  OAI210     u1143(.A0(men_men_n1171_), .A1(men_men_n300_), .B0(g), .Y(men_men_n1172_));
  NAi21      u1144(.An(f), .B(d), .Y(men_men_n1173_));
  NO2        u1145(.A(men_men_n1173_), .B(men_men_n1131_), .Y(men_men_n1174_));
  INV        u1146(.A(men_men_n1174_), .Y(men_men_n1175_));
  AOI210     u1147(.A0(men_men_n1172_), .A1(men_men_n306_), .B0(men_men_n1175_), .Y(men_men_n1176_));
  AOI210     u1148(.A0(men_men_n1176_), .A1(men_men_n117_), .B0(men_men_n1170_), .Y(men_men_n1177_));
  NA2        u1149(.A(men_men_n481_), .B(men_men_n480_), .Y(men_men_n1178_));
  NO2        u1150(.A(men_men_n191_), .B(men_men_n247_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n1179_), .B(m), .Y(men_men_n1180_));
  NA3        u1152(.A(men_men_n945_), .B(men_men_n1153_), .C(men_men_n484_), .Y(men_men_n1181_));
  OAI210     u1153(.A0(men_men_n1181_), .A1(men_men_n326_), .B0(men_men_n482_), .Y(men_men_n1182_));
  AOI210     u1154(.A0(men_men_n1182_), .A1(men_men_n1178_), .B0(men_men_n1180_), .Y(men_men_n1183_));
  NA2        u1155(.A(men_men_n578_), .B(men_men_n421_), .Y(men_men_n1184_));
  NA2        u1156(.A(men_men_n166_), .B(men_men_n33_), .Y(men_men_n1185_));
  AOI210     u1157(.A0(men_men_n995_), .A1(men_men_n1185_), .B0(men_men_n223_), .Y(men_men_n1186_));
  OAI210     u1158(.A0(men_men_n1186_), .A1(men_men_n459_), .B0(men_men_n1174_), .Y(men_men_n1187_));
  NO2        u1159(.A(men_men_n382_), .B(men_men_n381_), .Y(men_men_n1188_));
  AOI210     u1160(.A0(men_men_n1179_), .A1(men_men_n441_), .B0(men_men_n989_), .Y(men_men_n1189_));
  NAi41      u1161(.An(men_men_n1188_), .B(men_men_n1189_), .C(men_men_n1187_), .D(men_men_n1184_), .Y(men_men_n1190_));
  NO2        u1162(.A(men_men_n1190_), .B(men_men_n1183_), .Y(men_men_n1191_));
  NA4        u1163(.A(men_men_n1191_), .B(men_men_n1177_), .C(men_men_n1167_), .D(men_men_n1163_), .Y(men00));
  AOI210     u1164(.A0(men_men_n313_), .A1(men_men_n223_), .B0(men_men_n288_), .Y(men_men_n1193_));
  NO2        u1165(.A(men_men_n1193_), .B(men_men_n595_), .Y(men_men_n1194_));
  AOI210     u1166(.A0(men_men_n926_), .A1(men_men_n972_), .B0(men_men_n1148_), .Y(men_men_n1195_));
  NO3        u1167(.A(men_men_n1124_), .B(men_men_n989_), .C(men_men_n733_), .Y(men_men_n1196_));
  NA3        u1168(.A(men_men_n1196_), .B(men_men_n1195_), .C(men_men_n1031_), .Y(men_men_n1197_));
  NA2        u1169(.A(men_men_n525_), .B(f), .Y(men_men_n1198_));
  OAI210     u1170(.A0(men_men_n1038_), .A1(men_men_n40_), .B0(men_men_n668_), .Y(men_men_n1199_));
  NA3        u1171(.A(men_men_n1199_), .B(men_men_n267_), .C(n), .Y(men_men_n1200_));
  AOI210     u1172(.A0(men_men_n1200_), .A1(men_men_n1198_), .B0(men_men_n1079_), .Y(men_men_n1201_));
  NO4        u1173(.A(men_men_n1201_), .B(men_men_n1197_), .C(men_men_n1194_), .D(men_men_n1102_), .Y(men_men_n1202_));
  NA3        u1174(.A(men_men_n175_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1203_));
  NA3        u1175(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1204_));
  NOi31      u1176(.An(n), .B(m), .C(i), .Y(men_men_n1205_));
  NA3        u1177(.A(men_men_n1205_), .B(men_men_n671_), .C(men_men_n51_), .Y(men_men_n1206_));
  OAI210     u1178(.A0(men_men_n1204_), .A1(men_men_n1203_), .B0(men_men_n1206_), .Y(men_men_n1207_));
  NO3        u1179(.A(men_men_n1207_), .B(men_men_n1188_), .C(men_men_n948_), .Y(men_men_n1208_));
  NO4        u1180(.A(men_men_n501_), .B(men_men_n366_), .C(men_men_n1164_), .D(men_men_n59_), .Y(men_men_n1209_));
  NA3        u1181(.A(men_men_n394_), .B(men_men_n230_), .C(g), .Y(men_men_n1210_));
  OR2        u1182(.A(men_men_n395_), .B(men_men_n140_), .Y(men_men_n1211_));
  NO2        u1183(.A(h), .B(g), .Y(men_men_n1212_));
  NA4        u1184(.A(men_men_n514_), .B(men_men_n479_), .C(men_men_n1212_), .D(men_men_n1067_), .Y(men_men_n1213_));
  OAI220     u1185(.A0(men_men_n543_), .A1(men_men_n616_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1214_));
  NA2        u1186(.A(men_men_n1214_), .B(men_men_n552_), .Y(men_men_n1215_));
  AOI220     u1187(.A0(men_men_n333_), .A1(men_men_n256_), .B0(men_men_n186_), .B1(men_men_n155_), .Y(men_men_n1216_));
  NA4        u1188(.A(men_men_n1216_), .B(men_men_n1215_), .C(men_men_n1213_), .D(men_men_n1211_), .Y(men_men_n1217_));
  NO3        u1189(.A(men_men_n1217_), .B(men_men_n1209_), .C(men_men_n277_), .Y(men_men_n1218_));
  INV        u1190(.A(men_men_n335_), .Y(men_men_n1219_));
  AOI210     u1191(.A0(men_men_n256_), .A1(men_men_n356_), .B0(men_men_n596_), .Y(men_men_n1220_));
  NA3        u1192(.A(men_men_n1220_), .B(men_men_n1219_), .C(men_men_n161_), .Y(men_men_n1221_));
  NA3        u1193(.A(men_men_n188_), .B(men_men_n116_), .C(g), .Y(men_men_n1222_));
  NA3        u1194(.A(men_men_n479_), .B(men_men_n40_), .C(f), .Y(men_men_n1223_));
  NOi31      u1195(.An(men_men_n898_), .B(men_men_n1223_), .C(men_men_n1222_), .Y(men_men_n1224_));
  NAi31      u1196(.An(men_men_n195_), .B(men_men_n885_), .C(men_men_n479_), .Y(men_men_n1225_));
  NAi21      u1197(.An(men_men_n1224_), .B(men_men_n1225_), .Y(men_men_n1226_));
  NO2        u1198(.A(men_men_n287_), .B(men_men_n75_), .Y(men_men_n1227_));
  NO3        u1199(.A(men_men_n438_), .B(men_men_n856_), .C(n), .Y(men_men_n1228_));
  AOI210     u1200(.A0(men_men_n1228_), .A1(men_men_n1227_), .B0(men_men_n1117_), .Y(men_men_n1229_));
  NAi31      u1201(.An(men_men_n1082_), .B(men_men_n1229_), .C(men_men_n74_), .Y(men_men_n1230_));
  NO4        u1202(.A(men_men_n1230_), .B(men_men_n1226_), .C(men_men_n1221_), .D(men_men_n534_), .Y(men_men_n1231_));
  AN3        u1203(.A(men_men_n1231_), .B(men_men_n1218_), .C(men_men_n1208_), .Y(men_men_n1232_));
  NA2        u1204(.A(men_men_n552_), .B(men_men_n104_), .Y(men_men_n1233_));
  NA3        u1205(.A(men_men_n579_), .B(men_men_n1233_), .C(men_men_n252_), .Y(men_men_n1234_));
  NA2        u1206(.A(men_men_n1143_), .B(men_men_n552_), .Y(men_men_n1235_));
  NA4        u1207(.A(men_men_n671_), .B(men_men_n214_), .C(men_men_n230_), .D(men_men_n169_), .Y(men_men_n1236_));
  NA3        u1208(.A(men_men_n1236_), .B(men_men_n1235_), .C(men_men_n310_), .Y(men_men_n1237_));
  OAI210     u1209(.A0(men_men_n478_), .A1(men_men_n124_), .B0(men_men_n891_), .Y(men_men_n1238_));
  AOI220     u1210(.A0(men_men_n1238_), .A1(men_men_n1181_), .B0(men_men_n578_), .B1(men_men_n421_), .Y(men_men_n1239_));
  OR4        u1211(.A(men_men_n1079_), .B(men_men_n283_), .C(men_men_n232_), .D(e), .Y(men_men_n1240_));
  NO2        u1212(.A(men_men_n226_), .B(men_men_n223_), .Y(men_men_n1241_));
  NA2        u1213(.A(n), .B(e), .Y(men_men_n1242_));
  NO2        u1214(.A(men_men_n1242_), .B(men_men_n153_), .Y(men_men_n1243_));
  AOI220     u1215(.A0(men_men_n1243_), .A1(men_men_n285_), .B0(men_men_n872_), .B1(men_men_n1241_), .Y(men_men_n1244_));
  OAI210     u1216(.A0(men_men_n367_), .A1(men_men_n327_), .B0(men_men_n461_), .Y(men_men_n1245_));
  NA4        u1217(.A(men_men_n1245_), .B(men_men_n1244_), .C(men_men_n1240_), .D(men_men_n1239_), .Y(men_men_n1246_));
  AOI210     u1218(.A0(men_men_n1243_), .A1(men_men_n876_), .B0(men_men_n844_), .Y(men_men_n1247_));
  NO2        u1219(.A(men_men_n68_), .B(h), .Y(men_men_n1248_));
  NO3        u1220(.A(men_men_n1079_), .B(men_men_n1077_), .C(men_men_n749_), .Y(men_men_n1249_));
  INV        u1221(.A(men_men_n137_), .Y(men_men_n1250_));
  AN2        u1222(.A(men_men_n1250_), .B(men_men_n1129_), .Y(men_men_n1251_));
  OAI210     u1223(.A0(men_men_n1251_), .A1(men_men_n1249_), .B0(men_men_n1248_), .Y(men_men_n1252_));
  NA3        u1224(.A(men_men_n1252_), .B(men_men_n1247_), .C(men_men_n893_), .Y(men_men_n1253_));
  NO4        u1225(.A(men_men_n1253_), .B(men_men_n1246_), .C(men_men_n1237_), .D(men_men_n1234_), .Y(men_men_n1254_));
  NA2        u1226(.A(men_men_n861_), .B(men_men_n782_), .Y(men_men_n1255_));
  NA4        u1227(.A(men_men_n1255_), .B(men_men_n1254_), .C(men_men_n1232_), .D(men_men_n1202_), .Y(men01));
  AN2        u1228(.A(men_men_n1056_), .B(men_men_n1054_), .Y(men_men_n1257_));
  NO4        u1229(.A(men_men_n824_), .B(men_men_n816_), .C(men_men_n492_), .D(men_men_n294_), .Y(men_men_n1258_));
  NA2        u1230(.A(men_men_n405_), .B(i), .Y(men_men_n1259_));
  NA3        u1231(.A(men_men_n1259_), .B(men_men_n1258_), .C(men_men_n1257_), .Y(men_men_n1260_));
  NA2        u1232(.A(men_men_n605_), .B(men_men_n92_), .Y(men_men_n1261_));
  INV        u1233(.A(men_men_n572_), .Y(men_men_n1262_));
  NA2        u1234(.A(men_men_n992_), .B(men_men_n1262_), .Y(men_men_n1263_));
  NA4        u1235(.A(men_men_n1263_), .B(men_men_n1261_), .C(men_men_n941_), .D(men_men_n343_), .Y(men_men_n1264_));
  NA2        u1236(.A(men_men_n45_), .B(f), .Y(men_men_n1265_));
  NA2        u1237(.A(men_men_n730_), .B(men_men_n99_), .Y(men_men_n1266_));
  NO2        u1238(.A(men_men_n1266_), .B(men_men_n1265_), .Y(men_men_n1267_));
  OAI210     u1239(.A0(men_men_n804_), .A1(men_men_n622_), .B0(men_men_n1236_), .Y(men_men_n1268_));
  AOI210     u1240(.A0(men_men_n1267_), .A1(men_men_n658_), .B0(men_men_n1268_), .Y(men_men_n1269_));
  INV        u1241(.A(men_men_n122_), .Y(men_men_n1270_));
  OA220      u1242(.A0(men_men_n1270_), .A1(men_men_n602_), .B0(men_men_n683_), .B1(men_men_n379_), .Y(men_men_n1271_));
  NA3        u1243(.A(men_men_n1271_), .B(men_men_n1269_), .C(men_men_n925_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n805_), .B(men_men_n527_), .Y(men_men_n1273_));
  NA4        u1245(.A(men_men_n730_), .B(men_men_n99_), .C(men_men_n45_), .D(men_men_n222_), .Y(men_men_n1274_));
  OA220      u1246(.A0(men_men_n1274_), .A1(men_men_n692_), .B0(men_men_n203_), .B1(men_men_n201_), .Y(men_men_n1275_));
  NA3        u1247(.A(men_men_n1275_), .B(men_men_n1273_), .C(men_men_n143_), .Y(men_men_n1276_));
  NO4        u1248(.A(men_men_n1276_), .B(men_men_n1272_), .C(men_men_n1264_), .D(men_men_n1260_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n1210_), .B(men_men_n215_), .Y(men_men_n1278_));
  OAI210     u1250(.A0(men_men_n1278_), .A1(men_men_n316_), .B0(men_men_n547_), .Y(men_men_n1279_));
  NA2        u1251(.A(men_men_n555_), .B(men_men_n407_), .Y(men_men_n1280_));
  NOi21      u1252(.An(men_men_n580_), .B(men_men_n599_), .Y(men_men_n1281_));
  NA2        u1253(.A(men_men_n1281_), .B(men_men_n1280_), .Y(men_men_n1282_));
  AOI210     u1254(.A0(men_men_n212_), .A1(men_men_n91_), .B0(men_men_n222_), .Y(men_men_n1283_));
  OAI210     u1255(.A0(men_men_n831_), .A1(men_men_n439_), .B0(men_men_n1283_), .Y(men_men_n1284_));
  AN3        u1256(.A(m), .B(l), .C(k), .Y(men_men_n1285_));
  OAI210     u1257(.A0(men_men_n369_), .A1(men_men_n34_), .B0(men_men_n1285_), .Y(men_men_n1286_));
  NA2        u1258(.A(men_men_n211_), .B(men_men_n34_), .Y(men_men_n1287_));
  AO210      u1259(.A0(men_men_n1287_), .A1(men_men_n1286_), .B0(men_men_n342_), .Y(men_men_n1288_));
  NA4        u1260(.A(men_men_n1288_), .B(men_men_n1284_), .C(men_men_n1282_), .D(men_men_n1279_), .Y(men_men_n1289_));
  AOI210     u1261(.A0(men_men_n614_), .A1(men_men_n122_), .B0(men_men_n620_), .Y(men_men_n1290_));
  OAI210     u1262(.A0(men_men_n1270_), .A1(men_men_n611_), .B0(men_men_n1290_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n293_), .B(men_men_n203_), .Y(men_men_n1292_));
  NA2        u1264(.A(men_men_n1292_), .B(men_men_n688_), .Y(men_men_n1293_));
  NO3        u1265(.A(men_men_n843_), .B(men_men_n212_), .C(men_men_n419_), .Y(men_men_n1294_));
  NO2        u1266(.A(men_men_n1294_), .B(men_men_n989_), .Y(men_men_n1295_));
  NA3        u1267(.A(men_men_n1295_), .B(men_men_n1293_), .C(men_men_n807_), .Y(men_men_n1296_));
  NO3        u1268(.A(men_men_n1296_), .B(men_men_n1291_), .C(men_men_n1289_), .Y(men_men_n1297_));
  NA3        u1269(.A(men_men_n623_), .B(men_men_n29_), .C(f), .Y(men_men_n1298_));
  NO2        u1270(.A(men_men_n1298_), .B(men_men_n212_), .Y(men_men_n1299_));
  AOI210     u1271(.A0(men_men_n521_), .A1(men_men_n58_), .B0(men_men_n1299_), .Y(men_men_n1300_));
  OR3        u1272(.A(men_men_n1266_), .B(men_men_n624_), .C(men_men_n1265_), .Y(men_men_n1301_));
  NO2        u1273(.A(men_men_n1274_), .B(men_men_n1009_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n215_), .B(men_men_n115_), .Y(men_men_n1303_));
  NO3        u1275(.A(men_men_n1303_), .B(men_men_n1302_), .C(men_men_n1207_), .Y(men_men_n1304_));
  NA4        u1276(.A(men_men_n1304_), .B(men_men_n1301_), .C(men_men_n1300_), .D(men_men_n781_), .Y(men_men_n1305_));
  NO2        u1277(.A(men_men_n999_), .B(men_men_n242_), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n590_), .B(men_men_n588_), .Y(men_men_n1307_));
  NO3        u1279(.A(men_men_n81_), .B(men_men_n314_), .C(men_men_n45_), .Y(men_men_n1308_));
  NA2        u1280(.A(men_men_n1308_), .B(men_men_n571_), .Y(men_men_n1309_));
  NA3        u1281(.A(men_men_n1309_), .B(men_men_n1307_), .C(men_men_n694_), .Y(men_men_n1310_));
  NO2        u1282(.A(men_men_n379_), .B(men_men_n73_), .Y(men_men_n1311_));
  INV        u1283(.A(men_men_n1311_), .Y(men_men_n1312_));
  NA2        u1284(.A(men_men_n1312_), .B(men_men_n397_), .Y(men_men_n1313_));
  NO3        u1285(.A(men_men_n1313_), .B(men_men_n1310_), .C(men_men_n1305_), .Y(men_men_n1314_));
  NO2        u1286(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1315_));
  NO2        u1287(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1316_));
  AO220      u1288(.A0(men_men_n1316_), .A1(men_men_n644_), .B0(men_men_n1315_), .B1(men_men_n728_), .Y(men_men_n1317_));
  NA2        u1289(.A(men_men_n1317_), .B(men_men_n350_), .Y(men_men_n1318_));
  INV        u1290(.A(men_men_n140_), .Y(men_men_n1319_));
  NO3        u1291(.A(men_men_n1127_), .B(men_men_n185_), .C(men_men_n89_), .Y(men_men_n1320_));
  AOI220     u1292(.A0(men_men_n1320_), .A1(men_men_n1319_), .B0(men_men_n1308_), .B1(men_men_n1000_), .Y(men_men_n1321_));
  NA2        u1293(.A(men_men_n1321_), .B(men_men_n1318_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n635_), .B(men_men_n634_), .Y(men_men_n1323_));
  NO4        u1295(.A(men_men_n1127_), .B(men_men_n1323_), .C(men_men_n183_), .D(men_men_n89_), .Y(men_men_n1324_));
  NO3        u1296(.A(men_men_n1324_), .B(men_men_n1322_), .C(men_men_n662_), .Y(men_men_n1325_));
  NA4        u1297(.A(men_men_n1325_), .B(men_men_n1314_), .C(men_men_n1297_), .D(men_men_n1277_), .Y(men06));
  NO2        u1298(.A(men_men_n420_), .B(men_men_n577_), .Y(men_men_n1327_));
  INV        u1299(.A(men_men_n756_), .Y(men_men_n1328_));
  OAI210     u1300(.A0(men_men_n1328_), .A1(men_men_n278_), .B0(men_men_n1327_), .Y(men_men_n1329_));
  NO2        u1301(.A(men_men_n234_), .B(men_men_n106_), .Y(men_men_n1330_));
  OAI210     u1302(.A0(men_men_n1330_), .A1(men_men_n1320_), .B0(men_men_n393_), .Y(men_men_n1331_));
  NO3        u1303(.A(men_men_n618_), .B(men_men_n829_), .C(men_men_n621_), .Y(men_men_n1332_));
  OR2        u1304(.A(men_men_n1332_), .B(men_men_n912_), .Y(men_men_n1333_));
  NA3        u1305(.A(men_men_n1333_), .B(men_men_n1331_), .C(men_men_n1329_), .Y(men_men_n1334_));
  NO3        u1306(.A(men_men_n1334_), .B(men_men_n1310_), .C(men_men_n266_), .Y(men_men_n1335_));
  NO2        u1307(.A(men_men_n314_), .B(men_men_n45_), .Y(men_men_n1336_));
  AOI210     u1308(.A0(men_men_n1336_), .A1(men_men_n1001_), .B0(men_men_n1306_), .Y(men_men_n1337_));
  AOI210     u1309(.A0(men_men_n1336_), .A1(men_men_n574_), .B0(men_men_n1317_), .Y(men_men_n1338_));
  AOI210     u1310(.A0(men_men_n1338_), .A1(men_men_n1337_), .B0(men_men_n348_), .Y(men_men_n1339_));
  NO2        u1311(.A(men_men_n530_), .B(men_men_n180_), .Y(men_men_n1340_));
  NOi21      u1312(.An(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n628_), .B(men_men_n1150_), .Y(men_men_n1342_));
  NO2        u1314(.A(men_men_n474_), .B(men_men_n257_), .Y(men_men_n1343_));
  NO4        u1315(.A(men_men_n1343_), .B(men_men_n1342_), .C(men_men_n1341_), .D(men_men_n1340_), .Y(men_men_n1344_));
  OR2        u1316(.A(men_men_n619_), .B(men_men_n617_), .Y(men_men_n1345_));
  NO2        u1317(.A(men_men_n378_), .B(men_men_n141_), .Y(men_men_n1346_));
  AOI210     u1318(.A0(men_men_n1346_), .A1(men_men_n605_), .B0(men_men_n1345_), .Y(men_men_n1347_));
  NA2        u1319(.A(men_men_n1347_), .B(men_men_n1344_), .Y(men_men_n1348_));
  NO2        u1320(.A(men_men_n772_), .B(men_men_n377_), .Y(men_men_n1349_));
  NO3        u1321(.A(men_men_n698_), .B(men_men_n783_), .C(men_men_n658_), .Y(men_men_n1350_));
  NOi21      u1322(.An(men_men_n1349_), .B(men_men_n1350_), .Y(men_men_n1351_));
  AN2        u1323(.A(men_men_n985_), .B(men_men_n667_), .Y(men_men_n1352_));
  NO4        u1324(.A(men_men_n1352_), .B(men_men_n1351_), .C(men_men_n1348_), .D(men_men_n1339_), .Y(men_men_n1353_));
  NO2        u1325(.A(men_men_n823_), .B(men_men_n289_), .Y(men_men_n1354_));
  OAI220     u1326(.A0(men_men_n756_), .A1(men_men_n47_), .B0(men_men_n234_), .B1(men_men_n637_), .Y(men_men_n1355_));
  OAI210     u1327(.A0(men_men_n289_), .A1(c), .B0(men_men_n665_), .Y(men_men_n1356_));
  AOI220     u1328(.A0(men_men_n1356_), .A1(men_men_n1355_), .B0(men_men_n1354_), .B1(men_men_n278_), .Y(men_men_n1357_));
  NO3        u1329(.A(men_men_n254_), .B(men_men_n106_), .C(men_men_n296_), .Y(men_men_n1358_));
  OAI220     u1330(.A0(men_men_n721_), .A1(men_men_n257_), .B0(men_men_n526_), .B1(men_men_n530_), .Y(men_men_n1359_));
  OAI210     u1331(.A0(l), .A1(i), .B0(k), .Y(men_men_n1360_));
  NO3        u1332(.A(men_men_n1360_), .B(men_men_n616_), .C(j), .Y(men_men_n1361_));
  NOi21      u1333(.An(men_men_n1361_), .B(men_men_n692_), .Y(men_men_n1362_));
  NO4        u1334(.A(men_men_n1362_), .B(men_men_n1359_), .C(men_men_n1358_), .D(men_men_n1152_), .Y(men_men_n1363_));
  NA4        u1335(.A(men_men_n814_), .B(men_men_n813_), .C(men_men_n449_), .D(men_men_n905_), .Y(men_men_n1364_));
  NAi31      u1336(.An(men_men_n772_), .B(men_men_n1364_), .C(men_men_n211_), .Y(men_men_n1365_));
  NA3        u1337(.A(men_men_n1365_), .B(men_men_n1363_), .C(men_men_n1357_), .Y(men_men_n1366_));
  NOi31      u1338(.An(men_men_n1332_), .B(men_men_n477_), .C(men_men_n406_), .Y(men_men_n1367_));
  OR3        u1339(.A(men_men_n1367_), .B(men_men_n804_), .C(men_men_n558_), .Y(men_men_n1368_));
  OR3        u1340(.A(men_men_n381_), .B(men_men_n234_), .C(men_men_n637_), .Y(men_men_n1369_));
  INV        u1341(.A(men_men_n383_), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n1361_), .B(men_men_n810_), .Y(men_men_n1371_));
  NA4        u1343(.A(men_men_n1371_), .B(men_men_n1370_), .C(men_men_n1369_), .D(men_men_n1368_), .Y(men_men_n1372_));
  AOI220     u1344(.A0(men_men_n1349_), .A1(men_men_n782_), .B0(men_men_n1346_), .B1(men_men_n248_), .Y(men_men_n1373_));
  AN2        u1345(.A(men_men_n957_), .B(men_men_n956_), .Y(men_men_n1374_));
  NO4        u1346(.A(men_men_n1374_), .B(men_men_n903_), .C(men_men_n517_), .D(men_men_n495_), .Y(men_men_n1375_));
  NA2        u1347(.A(men_men_n1375_), .B(men_men_n1373_), .Y(men_men_n1376_));
  NAi21      u1348(.An(j), .B(i), .Y(men_men_n1377_));
  NO4        u1349(.A(men_men_n1323_), .B(men_men_n1377_), .C(men_men_n455_), .D(men_men_n245_), .Y(men_men_n1378_));
  NO4        u1350(.A(men_men_n1378_), .B(men_men_n1376_), .C(men_men_n1372_), .D(men_men_n1366_), .Y(men_men_n1379_));
  NA4        u1351(.A(men_men_n1379_), .B(men_men_n1353_), .C(men_men_n1335_), .D(men_men_n1325_), .Y(men07));
  NOi21      u1352(.An(j), .B(k), .Y(men_men_n1381_));
  NAi32      u1353(.An(m), .Bn(b), .C(n), .Y(men_men_n1382_));
  NO3        u1354(.A(men_men_n1382_), .B(g), .C(f), .Y(men_men_n1383_));
  OAI210     u1355(.A0(men_men_n334_), .A1(men_men_n497_), .B0(men_men_n1383_), .Y(men_men_n1384_));
  NAi21      u1356(.An(f), .B(c), .Y(men_men_n1385_));
  OR2        u1357(.A(e), .B(d), .Y(men_men_n1386_));
  NOi31      u1358(.An(n), .B(m), .C(b), .Y(men_men_n1387_));
  NO3        u1359(.A(men_men_n137_), .B(men_men_n463_), .C(h), .Y(men_men_n1388_));
  INV        u1360(.A(men_men_n1384_), .Y(men_men_n1389_));
  NOi41      u1361(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1390_));
  NA3        u1362(.A(men_men_n1390_), .B(men_men_n895_), .C(men_men_n422_), .Y(men_men_n1391_));
  NO2        u1363(.A(men_men_n1391_), .B(men_men_n56_), .Y(men_men_n1392_));
  NA2        u1364(.A(men_men_n1129_), .B(men_men_n230_), .Y(men_men_n1393_));
  NO2        u1365(.A(men_men_n1393_), .B(men_men_n61_), .Y(men_men_n1394_));
  NO2        u1366(.A(k), .B(i), .Y(men_men_n1395_));
  NA3        u1367(.A(men_men_n1395_), .B(men_men_n924_), .C(men_men_n188_), .Y(men_men_n1396_));
  NA2        u1368(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1397_));
  NO2        u1369(.A(men_men_n1085_), .B(men_men_n455_), .Y(men_men_n1398_));
  NA3        u1370(.A(men_men_n1398_), .B(men_men_n1397_), .C(men_men_n223_), .Y(men_men_n1399_));
  NO2        u1371(.A(men_men_n1099_), .B(men_men_n321_), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n1248_), .B(men_men_n304_), .Y(men_men_n1401_));
  NA3        u1373(.A(men_men_n1401_), .B(men_men_n1399_), .C(men_men_n1396_), .Y(men_men_n1402_));
  NO4        u1374(.A(men_men_n1402_), .B(men_men_n1394_), .C(men_men_n1392_), .D(men_men_n1389_), .Y(men_men_n1403_));
  NO3        u1375(.A(e), .B(d), .C(c), .Y(men_men_n1404_));
  OAI210     u1376(.A0(men_men_n137_), .A1(men_men_n223_), .B0(men_men_n625_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1405_), .B(men_men_n1404_), .Y(men_men_n1406_));
  INV        u1378(.A(men_men_n1406_), .Y(men_men_n1407_));
  OR2        u1379(.A(h), .B(f), .Y(men_men_n1408_));
  NO3        u1380(.A(n), .B(m), .C(i), .Y(men_men_n1409_));
  OAI210     u1381(.A0(men_men_n1151_), .A1(men_men_n164_), .B0(men_men_n1409_), .Y(men_men_n1410_));
  NO2        u1382(.A(i), .B(g), .Y(men_men_n1411_));
  OR3        u1383(.A(men_men_n1411_), .B(men_men_n1382_), .C(men_men_n72_), .Y(men_men_n1412_));
  OAI220     u1384(.A0(men_men_n1412_), .A1(men_men_n497_), .B0(men_men_n1410_), .B1(men_men_n1408_), .Y(men_men_n1413_));
  NA3        u1385(.A(men_men_n718_), .B(men_men_n704_), .C(men_men_n116_), .Y(men_men_n1414_));
  NA3        u1386(.A(men_men_n1387_), .B(men_men_n1094_), .C(men_men_n696_), .Y(men_men_n1415_));
  AOI210     u1387(.A0(men_men_n1415_), .A1(men_men_n1414_), .B0(men_men_n45_), .Y(men_men_n1416_));
  NA2        u1388(.A(men_men_n1409_), .B(men_men_n664_), .Y(men_men_n1417_));
  NO2        u1389(.A(l), .B(k), .Y(men_men_n1418_));
  NO3        u1390(.A(men_men_n455_), .B(d), .C(c), .Y(men_men_n1419_));
  NO3        u1391(.A(men_men_n1416_), .B(men_men_n1413_), .C(men_men_n1407_), .Y(men_men_n1420_));
  NO2        u1392(.A(men_men_n154_), .B(h), .Y(men_men_n1421_));
  NO2        u1393(.A(men_men_n1109_), .B(l), .Y(men_men_n1422_));
  NO2        u1394(.A(g), .B(c), .Y(men_men_n1423_));
  NA3        u1395(.A(men_men_n1423_), .B(men_men_n148_), .C(men_men_n196_), .Y(men_men_n1424_));
  NO2        u1396(.A(men_men_n1424_), .B(men_men_n1422_), .Y(men_men_n1425_));
  NA2        u1397(.A(men_men_n1425_), .B(men_men_n188_), .Y(men_men_n1426_));
  NO2        u1398(.A(men_men_n465_), .B(a), .Y(men_men_n1427_));
  NA3        u1399(.A(men_men_n1427_), .B(men_men_n1595_), .C(men_men_n117_), .Y(men_men_n1428_));
  NO2        u1400(.A(i), .B(h), .Y(men_men_n1429_));
  NA2        u1401(.A(men_men_n1429_), .B(men_men_n230_), .Y(men_men_n1430_));
  AOI210     u1402(.A0(men_men_n1173_), .A1(h), .B0(men_men_n427_), .Y(men_men_n1431_));
  NA2        u1403(.A(men_men_n144_), .B(men_men_n230_), .Y(men_men_n1432_));
  AOI210     u1404(.A0(men_men_n267_), .A1(men_men_n120_), .B0(men_men_n547_), .Y(men_men_n1433_));
  OAI220     u1405(.A0(men_men_n1433_), .A1(men_men_n1430_), .B0(men_men_n1432_), .B1(men_men_n1431_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n779_), .B(men_men_n197_), .Y(men_men_n1435_));
  NOi31      u1407(.An(m), .B(n), .C(b), .Y(men_men_n1436_));
  NOi31      u1408(.An(f), .B(d), .C(c), .Y(men_men_n1437_));
  NA2        u1409(.A(men_men_n1437_), .B(men_men_n1436_), .Y(men_men_n1438_));
  INV        u1410(.A(men_men_n1438_), .Y(men_men_n1439_));
  NO3        u1411(.A(men_men_n1439_), .B(men_men_n1435_), .C(men_men_n1434_), .Y(men_men_n1440_));
  NA2        u1412(.A(men_men_n1120_), .B(men_men_n479_), .Y(men_men_n1441_));
  NO4        u1413(.A(men_men_n1441_), .B(men_men_n1094_), .C(men_men_n455_), .D(men_men_n45_), .Y(men_men_n1442_));
  OAI210     u1414(.A0(men_men_n191_), .A1(men_men_n542_), .B0(men_men_n1095_), .Y(men_men_n1443_));
  NO3        u1415(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1444_));
  INV        u1416(.A(men_men_n1443_), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n1445_), .B(men_men_n1442_), .Y(men_men_n1446_));
  AN4        u1418(.A(men_men_n1446_), .B(men_men_n1440_), .C(men_men_n1428_), .D(men_men_n1426_), .Y(men_men_n1447_));
  NA2        u1419(.A(men_men_n1387_), .B(men_men_n390_), .Y(men_men_n1448_));
  NO2        u1420(.A(men_men_n1448_), .B(men_men_n1076_), .Y(men_men_n1449_));
  NA2        u1421(.A(men_men_n1419_), .B(men_men_n224_), .Y(men_men_n1450_));
  NO2        u1422(.A(men_men_n197_), .B(b), .Y(men_men_n1451_));
  AOI220     u1423(.A0(men_men_n1205_), .A1(men_men_n1451_), .B0(men_men_n1128_), .B1(men_men_n1441_), .Y(men_men_n1452_));
  NO2        u1424(.A(i), .B(men_men_n222_), .Y(men_men_n1453_));
  NA4        u1425(.A(men_men_n1179_), .B(men_men_n1453_), .C(men_men_n107_), .D(m), .Y(men_men_n1454_));
  NAi41      u1426(.An(men_men_n1449_), .B(men_men_n1454_), .C(men_men_n1452_), .D(men_men_n1450_), .Y(men_men_n1455_));
  NO4        u1427(.A(men_men_n137_), .B(g), .C(f), .D(e), .Y(men_men_n1456_));
  NA3        u1428(.A(men_men_n1395_), .B(men_men_n305_), .C(h), .Y(men_men_n1457_));
  NA2        u1429(.A(men_men_n202_), .B(men_men_n101_), .Y(men_men_n1458_));
  OR2        u1430(.A(e), .B(a), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n30_), .B(h), .Y(men_men_n1460_));
  NO2        u1432(.A(men_men_n1460_), .B(men_men_n1116_), .Y(men_men_n1461_));
  NOi41      u1433(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1462_));
  NA2        u1434(.A(men_men_n1462_), .B(men_men_n117_), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n1390_), .B(men_men_n1418_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n1464_), .B(men_men_n1463_), .Y(men_men_n1465_));
  OR3        u1437(.A(men_men_n558_), .B(men_men_n557_), .C(men_men_n116_), .Y(men_men_n1466_));
  NA2        u1438(.A(men_men_n1149_), .B(men_men_n419_), .Y(men_men_n1467_));
  OAI220     u1439(.A0(men_men_n1467_), .A1(men_men_n448_), .B0(men_men_n1466_), .B1(men_men_n314_), .Y(men_men_n1468_));
  AO210      u1440(.A0(men_men_n1468_), .A1(men_men_n120_), .B0(men_men_n1465_), .Y(men_men_n1469_));
  NO3        u1441(.A(men_men_n1469_), .B(men_men_n1461_), .C(men_men_n1455_), .Y(men_men_n1470_));
  NA4        u1442(.A(men_men_n1470_), .B(men_men_n1447_), .C(men_men_n1420_), .D(men_men_n1403_), .Y(men_men_n1471_));
  NO2        u1443(.A(men_men_n1164_), .B(men_men_n114_), .Y(men_men_n1472_));
  NA2        u1444(.A(men_men_n390_), .B(men_men_n56_), .Y(men_men_n1473_));
  AOI210     u1445(.A0(men_men_n1473_), .A1(men_men_n1085_), .B0(men_men_n1417_), .Y(men_men_n1474_));
  NA2        u1446(.A(men_men_n224_), .B(men_men_n188_), .Y(men_men_n1475_));
  AOI210     u1447(.A0(men_men_n1475_), .A1(men_men_n1222_), .B0(men_men_n1473_), .Y(men_men_n1476_));
  NO2        u1448(.A(men_men_n1121_), .B(men_men_n1116_), .Y(men_men_n1477_));
  NO3        u1449(.A(men_men_n1477_), .B(men_men_n1476_), .C(men_men_n1474_), .Y(men_men_n1478_));
  NO2        u1450(.A(men_men_n402_), .B(j), .Y(men_men_n1479_));
  NA3        u1451(.A(men_men_n1444_), .B(men_men_n1386_), .C(men_men_n1149_), .Y(men_men_n1480_));
  NAi41      u1452(.An(men_men_n1429_), .B(men_men_n1107_), .C(men_men_n176_), .D(men_men_n157_), .Y(men_men_n1481_));
  NA2        u1453(.A(men_men_n1481_), .B(men_men_n1480_), .Y(men_men_n1482_));
  NA3        u1454(.A(g), .B(men_men_n1479_), .C(men_men_n166_), .Y(men_men_n1483_));
  INV        u1455(.A(men_men_n1483_), .Y(men_men_n1484_));
  NO3        u1456(.A(men_men_n772_), .B(men_men_n183_), .C(men_men_n422_), .Y(men_men_n1485_));
  NO3        u1457(.A(men_men_n1485_), .B(men_men_n1484_), .C(men_men_n1482_), .Y(men_men_n1486_));
  NO3        u1458(.A(men_men_n1116_), .B(men_men_n599_), .C(g), .Y(men_men_n1487_));
  NOi21      u1459(.An(men_men_n1475_), .B(men_men_n1487_), .Y(men_men_n1488_));
  AOI210     u1460(.A0(men_men_n1488_), .A1(men_men_n1458_), .B0(men_men_n1085_), .Y(men_men_n1489_));
  OR2        u1461(.A(n), .B(i), .Y(men_men_n1490_));
  OAI210     u1462(.A0(men_men_n1490_), .A1(men_men_n1106_), .B0(men_men_n49_), .Y(men_men_n1491_));
  AOI220     u1463(.A0(men_men_n1491_), .A1(men_men_n1212_), .B0(men_men_n848_), .B1(men_men_n202_), .Y(men_men_n1492_));
  INV        u1464(.A(men_men_n1492_), .Y(men_men_n1493_));
  OAI220     u1465(.A0(men_men_n689_), .A1(g), .B0(men_men_n234_), .B1(c), .Y(men_men_n1494_));
  AOI210     u1466(.A0(men_men_n1451_), .A1(men_men_n41_), .B0(men_men_n1494_), .Y(men_men_n1495_));
  NO2        u1467(.A(men_men_n234_), .B(k), .Y(men_men_n1496_));
  NO2        u1468(.A(men_men_n1495_), .B(men_men_n185_), .Y(men_men_n1497_));
  NO3        u1469(.A(men_men_n1497_), .B(men_men_n1493_), .C(men_men_n1489_), .Y(men_men_n1498_));
  INV        u1470(.A(men_men_n49_), .Y(men_men_n1499_));
  NO3        u1471(.A(men_men_n1131_), .B(men_men_n1386_), .C(men_men_n49_), .Y(men_men_n1500_));
  NA2        u1472(.A(men_men_n1132_), .B(men_men_n1499_), .Y(men_men_n1501_));
  NO2        u1473(.A(men_men_n1116_), .B(h), .Y(men_men_n1502_));
  NA3        u1474(.A(men_men_n1502_), .B(d), .C(men_men_n1077_), .Y(men_men_n1503_));
  OAI220     u1475(.A0(men_men_n1503_), .A1(c), .B0(men_men_n1501_), .B1(j), .Y(men_men_n1504_));
  NA3        u1476(.A(men_men_n1472_), .B(men_men_n479_), .C(f), .Y(men_men_n1505_));
  NA2        u1477(.A(men_men_n188_), .B(men_men_n116_), .Y(men_men_n1506_));
  NO2        u1478(.A(men_men_n1381_), .B(men_men_n42_), .Y(men_men_n1507_));
  AOI210     u1479(.A0(men_men_n117_), .A1(men_men_n40_), .B0(men_men_n1507_), .Y(men_men_n1508_));
  NO2        u1480(.A(men_men_n1508_), .B(men_men_n1505_), .Y(men_men_n1509_));
  AOI210     u1481(.A0(men_men_n542_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1510_));
  NA2        u1482(.A(men_men_n1510_), .B(men_men_n1427_), .Y(men_men_n1511_));
  NO2        u1483(.A(men_men_n1377_), .B(men_men_n183_), .Y(men_men_n1512_));
  NOi21      u1484(.An(d), .B(f), .Y(men_men_n1513_));
  NO3        u1485(.A(men_men_n1437_), .B(men_men_n1513_), .C(men_men_n40_), .Y(men_men_n1514_));
  NA2        u1486(.A(men_men_n1514_), .B(men_men_n1512_), .Y(men_men_n1515_));
  NO2        u1487(.A(men_men_n1386_), .B(f), .Y(men_men_n1516_));
  NA2        u1488(.A(men_men_n1427_), .B(men_men_n1507_), .Y(men_men_n1517_));
  NO2        u1489(.A(men_men_n314_), .B(c), .Y(men_men_n1518_));
  NA2        u1490(.A(men_men_n1518_), .B(men_men_n559_), .Y(men_men_n1519_));
  NA4        u1491(.A(men_men_n1519_), .B(men_men_n1517_), .C(men_men_n1515_), .D(men_men_n1511_), .Y(men_men_n1520_));
  NO3        u1492(.A(men_men_n1520_), .B(men_men_n1509_), .C(men_men_n1504_), .Y(men_men_n1521_));
  NA4        u1493(.A(men_men_n1521_), .B(men_men_n1498_), .C(men_men_n1486_), .D(men_men_n1478_), .Y(men_men_n1522_));
  NO3        u1494(.A(men_men_n1120_), .B(men_men_n1106_), .C(men_men_n40_), .Y(men_men_n1523_));
  OAI220     u1495(.A0(men_men_n479_), .A1(men_men_n314_), .B0(men_men_n136_), .B1(men_men_n59_), .Y(men_men_n1524_));
  OAI210     u1496(.A0(men_men_n1524_), .A1(men_men_n1523_), .B0(men_men_n1400_), .Y(men_men_n1525_));
  OAI210     u1497(.A0(men_men_n1456_), .A1(men_men_n1387_), .B0(men_men_n909_), .Y(men_men_n1526_));
  OAI220     u1498(.A0(men_men_n1073_), .A1(men_men_n137_), .B0(men_men_n689_), .B1(men_men_n183_), .Y(men_men_n1527_));
  NA2        u1499(.A(men_men_n1527_), .B(men_men_n643_), .Y(men_men_n1528_));
  NA3        u1500(.A(men_men_n1528_), .B(men_men_n1526_), .C(men_men_n1525_), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1423_), .B(men_men_n1513_), .Y(men_men_n1530_));
  NO2        u1502(.A(men_men_n1530_), .B(m), .Y(men_men_n1531_));
  NA3        u1503(.A(men_men_n1129_), .B(men_men_n112_), .C(men_men_n230_), .Y(men_men_n1532_));
  OAI220     u1504(.A0(men_men_n158_), .A1(men_men_n190_), .B0(men_men_n463_), .B1(g), .Y(men_men_n1533_));
  OAI210     u1505(.A0(men_men_n1533_), .A1(men_men_n114_), .B0(men_men_n1436_), .Y(men_men_n1534_));
  NA2        u1506(.A(men_men_n1534_), .B(men_men_n1532_), .Y(men_men_n1535_));
  NO3        u1507(.A(men_men_n1535_), .B(men_men_n1531_), .C(men_men_n1529_), .Y(men_men_n1536_));
  NO2        u1508(.A(men_men_n1385_), .B(e), .Y(men_men_n1537_));
  NA2        u1509(.A(men_men_n1537_), .B(men_men_n417_), .Y(men_men_n1538_));
  NA2        u1510(.A(men_men_n1159_), .B(men_men_n654_), .Y(men_men_n1539_));
  OR3        u1511(.A(men_men_n1496_), .B(men_men_n1248_), .C(men_men_n137_), .Y(men_men_n1540_));
  OAI220     u1512(.A0(men_men_n1540_), .A1(men_men_n1538_), .B0(men_men_n1539_), .B1(men_men_n457_), .Y(men_men_n1541_));
  NO3        u1513(.A(men_men_n1466_), .B(men_men_n363_), .C(a), .Y(men_men_n1542_));
  NO2        u1514(.A(men_men_n1542_), .B(men_men_n1541_), .Y(men_men_n1543_));
  NO2        u1515(.A(men_men_n190_), .B(c), .Y(men_men_n1544_));
  OAI210     u1516(.A0(men_men_n1544_), .A1(men_men_n1537_), .B0(men_men_n188_), .Y(men_men_n1545_));
  AOI220     u1517(.A0(men_men_n1545_), .A1(men_men_n1108_), .B0(men_men_n549_), .B1(men_men_n377_), .Y(men_men_n1546_));
  NA2        u1518(.A(men_men_n557_), .B(g), .Y(men_men_n1547_));
  AOI210     u1519(.A0(men_men_n1547_), .A1(men_men_n1419_), .B0(men_men_n1500_), .Y(men_men_n1548_));
  NO2        u1520(.A(men_men_n1548_), .B(men_men_n222_), .Y(men_men_n1549_));
  AOI210     u1521(.A0(men_men_n929_), .A1(men_men_n429_), .B0(men_men_n108_), .Y(men_men_n1550_));
  OR2        u1522(.A(men_men_n1550_), .B(men_men_n557_), .Y(men_men_n1551_));
  NO2        u1523(.A(men_men_n1551_), .B(men_men_n183_), .Y(men_men_n1552_));
  NA2        u1524(.A(men_men_n1388_), .B(men_men_n191_), .Y(men_men_n1553_));
  NO2        u1525(.A(men_men_n49_), .B(l), .Y(men_men_n1554_));
  OAI210     u1526(.A0(men_men_n1459_), .A1(men_men_n887_), .B0(men_men_n497_), .Y(men_men_n1555_));
  OAI210     u1527(.A0(men_men_n1555_), .A1(men_men_n1132_), .B0(men_men_n1554_), .Y(men_men_n1556_));
  NO2        u1528(.A(m), .B(i), .Y(men_men_n1557_));
  BUFFER     u1529(.A(men_men_n1557_), .Y(men_men_n1558_));
  NA2        u1530(.A(men_men_n1558_), .B(men_men_n1421_), .Y(men_men_n1559_));
  NA3        u1531(.A(men_men_n1559_), .B(men_men_n1556_), .C(men_men_n1553_), .Y(men_men_n1560_));
  NO4        u1532(.A(men_men_n1560_), .B(men_men_n1552_), .C(men_men_n1549_), .D(men_men_n1546_), .Y(men_men_n1561_));
  NA3        u1533(.A(men_men_n1561_), .B(men_men_n1543_), .C(men_men_n1536_), .Y(men_men_n1562_));
  NA3        u1534(.A(men_men_n991_), .B(men_men_n144_), .C(men_men_n46_), .Y(men_men_n1563_));
  NO2        u1535(.A(men_men_n155_), .B(men_men_n1563_), .Y(men_men_n1564_));
  INV        u1536(.A(men_men_n194_), .Y(men_men_n1565_));
  NA2        u1537(.A(men_men_n1565_), .B(men_men_n1502_), .Y(men_men_n1566_));
  AO210      u1538(.A0(men_men_n138_), .A1(l), .B0(men_men_n1448_), .Y(men_men_n1567_));
  NO2        u1539(.A(men_men_n72_), .B(c), .Y(men_men_n1568_));
  NO4        u1540(.A(men_men_n1408_), .B(men_men_n195_), .C(men_men_n463_), .D(men_men_n45_), .Y(men_men_n1569_));
  AOI210     u1541(.A0(men_men_n1512_), .A1(men_men_n1568_), .B0(men_men_n1569_), .Y(men_men_n1570_));
  NA3        u1542(.A(men_men_n1570_), .B(men_men_n1567_), .C(men_men_n1566_), .Y(men_men_n1571_));
  NO2        u1543(.A(men_men_n1571_), .B(men_men_n1564_), .Y(men_men_n1572_));
  NO4        u1544(.A(men_men_n234_), .B(men_men_n195_), .C(men_men_n267_), .D(k), .Y(men_men_n1573_));
  AOI210     u1545(.A0(men_men_n164_), .A1(men_men_n56_), .B0(men_men_n1537_), .Y(men_men_n1574_));
  NO2        u1546(.A(men_men_n1574_), .B(men_men_n1506_), .Y(men_men_n1575_));
  NO2        u1547(.A(men_men_n1563_), .B(men_men_n114_), .Y(men_men_n1576_));
  NO3        u1548(.A(men_men_n1576_), .B(men_men_n1575_), .C(men_men_n1573_), .Y(men_men_n1577_));
  NO2        u1549(.A(men_men_n1505_), .B(men_men_n69_), .Y(men_men_n1578_));
  NA2        u1550(.A(men_men_n59_), .B(a), .Y(men_men_n1579_));
  NO2        u1551(.A(men_men_n1467_), .B(men_men_n1579_), .Y(men_men_n1580_));
  NO2        u1552(.A(men_men_n1580_), .B(men_men_n1578_), .Y(men_men_n1581_));
  NA3        u1553(.A(men_men_n1581_), .B(men_men_n1577_), .C(men_men_n1572_), .Y(men_men_n1582_));
  OR4        u1554(.A(men_men_n1582_), .B(men_men_n1562_), .C(men_men_n1522_), .D(men_men_n1471_), .Y(men04));
  NOi31      u1555(.An(men_men_n1456_), .B(men_men_n1457_), .C(men_men_n1079_), .Y(men_men_n1584_));
  NA2        u1556(.A(men_men_n1516_), .B(men_men_n848_), .Y(men_men_n1585_));
  NO4        u1557(.A(men_men_n1585_), .B(men_men_n1068_), .C(men_men_n498_), .D(j), .Y(men_men_n1586_));
  OR3        u1558(.A(men_men_n1586_), .B(men_men_n1584_), .C(men_men_n1097_), .Y(men_men_n1587_));
  NO3        u1559(.A(men_men_n1397_), .B(men_men_n93_), .C(k), .Y(men_men_n1588_));
  AOI210     u1560(.A0(men_men_n1588_), .A1(men_men_n1090_), .B0(men_men_n1224_), .Y(men_men_n1589_));
  NA2        u1561(.A(men_men_n1589_), .B(men_men_n1252_), .Y(men_men_n1590_));
  NO4        u1562(.A(men_men_n1590_), .B(men_men_n1587_), .C(men_men_n1105_), .D(men_men_n1084_), .Y(men_men_n1591_));
  NA4        u1563(.A(men_men_n1591_), .B(men_men_n1161_), .C(men_men_n1147_), .D(men_men_n1135_), .Y(men05));
  INV        u1564(.A(i), .Y(men_men_n1595_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule