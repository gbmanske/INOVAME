// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n133_, new_new_n134_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n987_,
    new_new_n988_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(mai1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA3        g031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  OAI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi31      g042(.An(new_new_n64_), .B(new_new_n62_), .C(new_new_n58_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(new_new_n78_), .B(new_new_n55_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n80_), .B(new_new_n60_), .Y(new_new_n82_));
  INV        g060(.A(i_6_), .Y(new_new_n83_));
  OR4        g061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n84_), .Y(new_new_n85_));
  NO2        g063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n85_), .B(new_new_n86_), .Y(new_new_n87_));
  OAI210     g065(.A0(new_new_n82_), .A1(new_new_n79_), .B0(new_new_n87_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n60_), .Y(new_new_n91_));
  NA2        g069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  INV        g070(.A(new_new_n91_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n88_), .B0(new_new_n77_), .Y(new_new_n94_));
  AN3        g072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n95_));
  NAi21      g073(.An(i_6_), .B(i_11_), .Y(new_new_n96_));
  NO2        g074(.A(i_5_), .B(i_8_), .Y(new_new_n97_));
  NOi21      g075(.An(new_new_n97_), .B(new_new_n96_), .Y(new_new_n98_));
  AOI220     g076(.A0(new_new_n98_), .A1(new_new_n59_), .B0(new_new_n95_), .B1(new_new_n32_), .Y(new_new_n99_));
  INV        g077(.A(i_7_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n47_), .B(new_new_n100_), .Y(new_new_n101_));
  NO2        g079(.A(i_0_), .B(i_5_), .Y(new_new_n102_));
  NO2        g080(.A(new_new_n102_), .B(new_new_n83_), .Y(new_new_n103_));
  NA2        g081(.A(i_12_), .B(i_3_), .Y(new_new_n104_));
  INV        g082(.A(new_new_n104_), .Y(new_new_n105_));
  NA3        g083(.A(new_new_n105_), .B(new_new_n103_), .C(new_new_n101_), .Y(new_new_n106_));
  NAi21      g084(.An(i_7_), .B(i_11_), .Y(new_new_n107_));
  NO3        g085(.A(new_new_n107_), .B(new_new_n89_), .C(new_new_n51_), .Y(new_new_n108_));
  AN2        g086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g088(.A(new_new_n77_), .B(new_new_n55_), .Y(new_new_n111_));
  NO2        g089(.A(i_8_), .B(new_new_n100_), .Y(new_new_n112_));
  NA2        g090(.A(i_12_), .B(i_7_), .Y(new_new_n113_));
  NA2        g091(.A(i_11_), .B(i_12_), .Y(new_new_n114_));
  NAi41      g092(.An(new_new_n108_), .B(new_new_n114_), .C(new_new_n106_), .D(new_new_n99_), .Y(new_new_n115_));
  NOi21      g093(.An(i_1_), .B(i_5_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(i_11_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n100_), .B(new_new_n37_), .Y(new_new_n118_));
  NA2        g096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n118_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n47_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n122_));
  NAi21      g100(.An(i_3_), .B(i_8_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n59_), .Y(new_new_n124_));
  NOi31      g102(.An(new_new_n124_), .B(new_new_n122_), .C(new_new_n121_), .Y(new_new_n125_));
  NO2        g103(.A(i_1_), .B(new_new_n83_), .Y(new_new_n126_));
  NO2        g104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  OAI220     g106(.A0(new_new_n128_), .A1(new_new_n107_), .B0(new_new_n125_), .B1(new_new_n117_), .Y(new_new_n129_));
  NO3        g107(.A(new_new_n129_), .B(new_new_n115_), .C(new_new_n94_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n76_), .Y(mai2));
  NO2        g109(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n132_));
  NA2        g110(.A(i_6_), .B(new_new_n25_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n132_), .Y(new_new_n134_));
  NA4        g112(.A(new_new_n134_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(mai0));
  AN2        g113(.A(i_8_), .B(i_7_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_6_), .Y(new_new_n137_));
  NO2        g115(.A(i_12_), .B(i_13_), .Y(new_new_n138_));
  NAi21      g116(.An(i_5_), .B(i_11_), .Y(new_new_n139_));
  NOi21      g117(.An(new_new_n138_), .B(new_new_n139_), .Y(new_new_n140_));
  NO2        g118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NA2        g119(.A(i_2_), .B(i_3_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n142_), .B(i_4_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n140_), .Y(new_new_n144_));
  AN2        g122(.A(new_new_n138_), .B(new_new_n80_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(new_new_n27_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n70_), .B(new_new_n47_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n40_), .Y(new_new_n156_));
  NO2        g134(.A(i_3_), .B(i_5_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  OAI210     g137(.A0(new_new_n159_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n160_), .B(new_new_n150_), .Y(new_new_n161_));
  AOI210     g139(.A0(new_new_n161_), .A1(new_new_n144_), .B0(new_new_n137_), .Y(new_new_n162_));
  NA3        g140(.A(new_new_n70_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n163_));
  NA2        g141(.A(i_3_), .B(new_new_n48_), .Y(new_new_n164_));
  NOi21      g142(.An(i_4_), .B(i_9_), .Y(new_new_n165_));
  NOi21      g143(.An(i_11_), .B(i_13_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  NO2        g145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA3        g148(.A(new_new_n170_), .B(new_new_n168_), .C(new_new_n80_), .Y(new_new_n171_));
  AOI210     g149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n163_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n70_), .B(new_new_n60_), .Y(new_new_n173_));
  INV        g151(.A(new_new_n173_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n36_), .B(i_5_), .Y(new_new_n175_));
  NAi31      g153(.An(new_new_n175_), .B(new_new_n145_), .C(i_11_), .Y(new_new_n176_));
  NA2        g154(.A(i_3_), .B(i_5_), .Y(new_new_n177_));
  OR2        g155(.A(new_new_n177_), .B(new_new_n167_), .Y(new_new_n178_));
  AOI210     g156(.A0(new_new_n178_), .A1(new_new_n176_), .B0(new_new_n174_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n70_), .B(i_5_), .Y(new_new_n180_));
  NO2        g158(.A(i_13_), .B(i_10_), .Y(new_new_n181_));
  NA3        g159(.A(new_new_n181_), .B(new_new_n180_), .C(new_new_n45_), .Y(new_new_n182_));
  NO2        g160(.A(i_2_), .B(i_1_), .Y(new_new_n183_));
  NA2        g161(.A(new_new_n183_), .B(i_3_), .Y(new_new_n184_));
  NAi21      g162(.An(i_4_), .B(i_12_), .Y(new_new_n185_));
  NO3        g163(.A(new_new_n184_), .B(new_new_n182_), .C(new_new_n25_), .Y(new_new_n186_));
  NO3        g164(.A(new_new_n186_), .B(new_new_n179_), .C(new_new_n172_), .Y(new_new_n187_));
  INV        g165(.A(i_8_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n188_), .B(i_7_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n189_), .B(i_6_), .Y(new_new_n190_));
  NO3        g168(.A(i_3_), .B(new_new_n83_), .C(new_new_n48_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(new_new_n112_), .Y(new_new_n192_));
  NO3        g170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n194_));
  NO3        g172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n195_));
  OAI210     g173(.A0(new_new_n95_), .A1(i_12_), .B0(new_new_n195_), .Y(new_new_n196_));
  AOI210     g174(.A0(new_new_n196_), .A1(new_new_n194_), .B0(new_new_n192_), .Y(new_new_n197_));
  NO2        g175(.A(i_3_), .B(i_8_), .Y(new_new_n198_));
  NO3        g176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n102_), .B(new_new_n55_), .Y(new_new_n200_));
  NO2        g178(.A(i_13_), .B(i_9_), .Y(new_new_n201_));
  NA3        g179(.A(new_new_n201_), .B(i_6_), .C(new_new_n188_), .Y(new_new_n202_));
  NAi21      g180(.An(i_12_), .B(i_3_), .Y(new_new_n203_));
  OR2        g181(.A(new_new_n203_), .B(new_new_n202_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n45_), .B(i_5_), .Y(new_new_n205_));
  NO3        g183(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n206_));
  NA2        g184(.A(new_new_n206_), .B(new_new_n205_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n207_), .B(new_new_n204_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n208_), .B(new_new_n197_), .Y(new_new_n209_));
  OAI220     g187(.A0(new_new_n209_), .A1(i_4_), .B0(new_new_n190_), .B1(new_new_n187_), .Y(new_new_n210_));
  NAi21      g188(.An(i_12_), .B(i_7_), .Y(new_new_n211_));
  NA3        g189(.A(i_13_), .B(new_new_n188_), .C(i_10_), .Y(new_new_n212_));
  NA2        g190(.A(i_0_), .B(i_5_), .Y(new_new_n213_));
  NAi31      g191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n36_), .B(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n47_), .B(new_new_n60_), .Y(new_new_n217_));
  INV        g195(.A(i_13_), .Y(new_new_n218_));
  NO2        g196(.A(i_12_), .B(new_new_n218_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n37_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n177_), .B(i_4_), .Y(new_new_n221_));
  NA2        g199(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n222_));
  OR2        g200(.A(i_8_), .B(i_7_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n223_), .B(new_new_n83_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n51_), .B(i_1_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  INV        g204(.A(i_12_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n45_), .B(new_new_n227_), .Y(new_new_n228_));
  NO3        g206(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n229_));
  NA2        g207(.A(i_2_), .B(i_1_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n226_), .B(new_new_n222_), .Y(new_new_n231_));
  NO3        g209(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n232_));
  NAi21      g210(.An(i_4_), .B(i_3_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n233_), .B(new_new_n72_), .Y(new_new_n234_));
  NO2        g212(.A(i_0_), .B(i_6_), .Y(new_new_n235_));
  NOi41      g213(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n230_), .B(new_new_n177_), .Y(new_new_n238_));
  NAi21      g216(.An(new_new_n237_), .B(new_new_n238_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n239_), .Y(new_new_n240_));
  AOI210     g218(.A0(new_new_n240_), .A1(new_new_n40_), .B0(new_new_n231_), .Y(new_new_n241_));
  NO2        g219(.A(i_11_), .B(new_new_n218_), .Y(new_new_n242_));
  NOi21      g220(.An(i_1_), .B(i_6_), .Y(new_new_n243_));
  NAi21      g221(.An(i_3_), .B(i_7_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n227_), .B(i_9_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n70_), .B(i_5_), .Y(new_new_n247_));
  NA3        g225(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n223_), .B(new_new_n37_), .Y(new_new_n249_));
  NA2        g227(.A(i_12_), .B(i_6_), .Y(new_new_n250_));
  OR2        g228(.A(i_13_), .B(i_9_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n233_), .B(i_2_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n242_), .B(i_9_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n148_), .B(new_new_n60_), .Y(new_new_n254_));
  NO3        g232(.A(i_11_), .B(new_new_n218_), .C(new_new_n25_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n244_), .B(i_8_), .Y(new_new_n256_));
  NA3        g234(.A(i_5_), .B(new_new_n256_), .C(new_new_n255_), .Y(new_new_n257_));
  NO3        g235(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n258_));
  NA3        g236(.A(new_new_n258_), .B(new_new_n249_), .C(new_new_n219_), .Y(new_new_n259_));
  AOI210     g237(.A0(new_new_n259_), .A1(new_new_n257_), .B0(new_new_n254_), .Y(new_new_n260_));
  INV        g238(.A(new_new_n260_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n261_), .B(new_new_n241_), .Y(new_new_n262_));
  NO3        g240(.A(i_12_), .B(new_new_n218_), .C(new_new_n37_), .Y(new_new_n263_));
  INV        g241(.A(new_new_n263_), .Y(new_new_n264_));
  NA2        g242(.A(i_8_), .B(new_new_n100_), .Y(new_new_n265_));
  NOi21      g243(.An(new_new_n157_), .B(new_new_n83_), .Y(new_new_n266_));
  NO3        g244(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n267_));
  AOI220     g245(.A0(new_new_n267_), .A1(new_new_n191_), .B0(new_new_n266_), .B1(new_new_n225_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n268_), .B(new_new_n265_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n230_), .B(i_0_), .Y(new_new_n270_));
  NA2        g248(.A(i_0_), .B(i_1_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n271_), .B(i_2_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n56_), .B(i_6_), .Y(new_new_n273_));
  NA3        g251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n157_), .Y(new_new_n274_));
  OAI210     g252(.A0(new_new_n159_), .A1(new_new_n137_), .B0(new_new_n274_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n275_), .B(new_new_n269_), .Y(new_new_n276_));
  NO2        g254(.A(i_3_), .B(i_10_), .Y(new_new_n277_));
  NA3        g255(.A(new_new_n277_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n278_));
  NO2        g256(.A(i_2_), .B(new_new_n100_), .Y(new_new_n279_));
  NA2        g257(.A(i_1_), .B(new_new_n36_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(i_8_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n281_), .B(new_new_n279_), .Y(new_new_n282_));
  AN2        g260(.A(i_3_), .B(i_10_), .Y(new_new_n283_));
  NA4        g261(.A(new_new_n283_), .B(new_new_n193_), .C(new_new_n170_), .D(new_new_n168_), .Y(new_new_n284_));
  NO2        g262(.A(i_5_), .B(new_new_n37_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n286_));
  OR2        g264(.A(new_new_n282_), .B(new_new_n278_), .Y(new_new_n287_));
  OAI220     g265(.A0(new_new_n287_), .A1(i_6_), .B0(new_new_n276_), .B1(new_new_n264_), .Y(new_new_n288_));
  NO4        g266(.A(new_new_n288_), .B(new_new_n262_), .C(new_new_n210_), .D(new_new_n162_), .Y(new_new_n289_));
  NO3        g267(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n290_));
  INV        g268(.A(new_new_n56_), .Y(new_new_n291_));
  NA2        g269(.A(new_new_n270_), .B(new_new_n291_), .Y(new_new_n292_));
  NO3        g270(.A(i_6_), .B(new_new_n188_), .C(i_7_), .Y(new_new_n293_));
  INV        g271(.A(new_new_n293_), .Y(new_new_n294_));
  AOI210     g272(.A0(new_new_n294_), .A1(new_new_n292_), .B0(new_new_n164_), .Y(new_new_n295_));
  NO2        g273(.A(i_2_), .B(i_3_), .Y(new_new_n296_));
  OR2        g274(.A(i_0_), .B(i_5_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n213_), .B(new_new_n297_), .Y(new_new_n298_));
  NA4        g276(.A(new_new_n298_), .B(new_new_n224_), .C(new_new_n296_), .D(i_1_), .Y(new_new_n299_));
  NA3        g277(.A(new_new_n270_), .B(new_new_n266_), .C(new_new_n112_), .Y(new_new_n300_));
  NAi21      g278(.An(i_8_), .B(i_7_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(i_6_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n151_), .B(new_new_n47_), .Y(new_new_n303_));
  NA3        g281(.A(new_new_n303_), .B(new_new_n302_), .C(new_new_n157_), .Y(new_new_n304_));
  NA3        g282(.A(new_new_n304_), .B(new_new_n300_), .C(new_new_n299_), .Y(new_new_n305_));
  OAI210     g283(.A0(new_new_n305_), .A1(new_new_n295_), .B0(i_4_), .Y(new_new_n306_));
  NO2        g284(.A(i_12_), .B(i_10_), .Y(new_new_n307_));
  NOi21      g285(.An(i_5_), .B(i_0_), .Y(new_new_n308_));
  NA4        g286(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n309_));
  NO2        g287(.A(i_6_), .B(i_8_), .Y(new_new_n310_));
  NOi21      g288(.An(i_0_), .B(i_2_), .Y(new_new_n311_));
  AN2        g289(.A(new_new_n311_), .B(new_new_n310_), .Y(new_new_n312_));
  NO2        g290(.A(i_1_), .B(i_7_), .Y(new_new_n313_));
  AO220      g291(.A0(new_new_n313_), .A1(new_new_n312_), .B0(new_new_n302_), .B1(new_new_n225_), .Y(new_new_n314_));
  NA3        g292(.A(new_new_n314_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n315_), .B(new_new_n306_), .Y(new_new_n316_));
  NO3        g294(.A(new_new_n223_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n317_));
  NO3        g295(.A(new_new_n301_), .B(i_2_), .C(i_1_), .Y(new_new_n318_));
  OAI210     g296(.A0(new_new_n318_), .A1(new_new_n317_), .B0(i_6_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n319_), .B(new_new_n298_), .Y(new_new_n320_));
  NOi21      g298(.An(new_new_n147_), .B(new_new_n103_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n321_), .B(new_new_n119_), .Y(new_new_n322_));
  OAI210     g300(.A0(new_new_n322_), .A1(new_new_n320_), .B0(i_3_), .Y(new_new_n323_));
  INV        g301(.A(new_new_n81_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n271_), .B(new_new_n78_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n325_), .B(new_new_n127_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n92_), .B(new_new_n188_), .Y(new_new_n327_));
  NA2        g305(.A(new_new_n327_), .B(new_new_n60_), .Y(new_new_n328_));
  AOI210     g306(.A0(new_new_n328_), .A1(new_new_n326_), .B0(new_new_n324_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n188_), .B(i_9_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n330_), .B(new_new_n200_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n331_), .B(new_new_n47_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n332_), .B(new_new_n329_), .Y(new_new_n333_));
  AOI210     g311(.A0(new_new_n333_), .A1(new_new_n323_), .B0(new_new_n156_), .Y(new_new_n334_));
  AOI210     g312(.A0(new_new_n316_), .A1(new_new_n290_), .B0(new_new_n334_), .Y(new_new_n335_));
  NOi32      g313(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n336_));
  INV        g314(.A(new_new_n336_), .Y(new_new_n337_));
  NAi21      g315(.An(i_1_), .B(i_5_), .Y(new_new_n338_));
  NAi41      g316(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n339_));
  OAI220     g317(.A0(new_new_n339_), .A1(new_new_n338_), .B0(new_new_n214_), .B1(new_new_n153_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n153_), .B(new_new_n151_), .Y(new_new_n341_));
  NOi32      g319(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n342_));
  NAi21      g320(.An(i_6_), .B(i_1_), .Y(new_new_n343_));
  NA3        g321(.A(new_new_n343_), .B(new_new_n342_), .C(new_new_n47_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n344_), .B(i_0_), .Y(new_new_n345_));
  OR3        g323(.A(new_new_n345_), .B(new_new_n341_), .C(new_new_n340_), .Y(new_new_n346_));
  NO2        g324(.A(i_1_), .B(new_new_n100_), .Y(new_new_n347_));
  NAi21      g325(.An(i_3_), .B(i_4_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(i_9_), .Y(new_new_n349_));
  AN2        g327(.A(i_6_), .B(i_7_), .Y(new_new_n350_));
  NA2        g328(.A(i_2_), .B(i_7_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n348_), .B(i_10_), .Y(new_new_n352_));
  AOI210     g330(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n353_));
  OAI210     g331(.A0(new_new_n353_), .A1(new_new_n183_), .B0(new_new_n352_), .Y(new_new_n354_));
  AOI220     g332(.A0(new_new_n352_), .A1(new_new_n313_), .B0(new_new_n229_), .B1(new_new_n183_), .Y(new_new_n355_));
  AOI210     g333(.A0(new_new_n355_), .A1(new_new_n354_), .B0(i_5_), .Y(new_new_n356_));
  NO3        g334(.A(new_new_n356_), .B(new_new_n346_), .C(new_new_n987_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(new_new_n337_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n359_));
  AN2        g337(.A(i_12_), .B(i_5_), .Y(new_new_n360_));
  NO2        g338(.A(i_11_), .B(i_6_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n233_), .B(i_5_), .Y(new_new_n362_));
  NO2        g340(.A(i_5_), .B(i_10_), .Y(new_new_n363_));
  AOI220     g341(.A0(new_new_n363_), .A1(new_new_n252_), .B0(new_new_n362_), .B1(new_new_n193_), .Y(new_new_n364_));
  NA2        g342(.A(new_new_n138_), .B(new_new_n46_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n365_), .B(new_new_n364_), .Y(new_new_n366_));
  NA2        g344(.A(new_new_n366_), .B(new_new_n359_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n368_));
  NO3        g346(.A(new_new_n83_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n369_));
  NO2        g347(.A(i_3_), .B(new_new_n100_), .Y(new_new_n370_));
  NO2        g348(.A(i_11_), .B(i_12_), .Y(new_new_n371_));
  NA3        g349(.A(new_new_n112_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n372_));
  NO2        g350(.A(new_new_n372_), .B(new_new_n214_), .Y(new_new_n373_));
  NAi21      g351(.An(i_13_), .B(i_0_), .Y(new_new_n374_));
  INV        g352(.A(new_new_n374_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n373_), .B(new_new_n375_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n376_), .B(new_new_n367_), .Y(new_new_n377_));
  NO3        g355(.A(i_1_), .B(i_12_), .C(new_new_n83_), .Y(new_new_n378_));
  NO2        g356(.A(i_0_), .B(i_11_), .Y(new_new_n379_));
  AN2        g357(.A(i_1_), .B(i_6_), .Y(new_new_n380_));
  NOi21      g358(.An(i_2_), .B(i_12_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n381_), .B(new_new_n380_), .Y(new_new_n382_));
  INV        g360(.A(new_new_n382_), .Y(new_new_n383_));
  NA2        g361(.A(new_new_n136_), .B(i_9_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n384_), .B(i_4_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n383_), .B(new_new_n385_), .Y(new_new_n386_));
  NAi21      g364(.An(i_9_), .B(i_4_), .Y(new_new_n387_));
  OR2        g365(.A(i_13_), .B(i_10_), .Y(new_new_n388_));
  NO3        g366(.A(new_new_n388_), .B(new_new_n114_), .C(new_new_n387_), .Y(new_new_n389_));
  OR2        g367(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n100_), .B(new_new_n25_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n263_), .B(new_new_n391_), .Y(new_new_n392_));
  NA2        g370(.A(i_5_), .B(new_new_n206_), .Y(new_new_n393_));
  OAI220     g371(.A0(new_new_n393_), .A1(new_new_n390_), .B0(new_new_n392_), .B1(new_new_n321_), .Y(new_new_n394_));
  INV        g372(.A(new_new_n394_), .Y(new_new_n395_));
  AOI210     g373(.A0(new_new_n395_), .A1(new_new_n386_), .B0(new_new_n26_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n300_), .B(new_new_n299_), .Y(new_new_n397_));
  AOI220     g375(.A0(new_new_n273_), .A1(new_new_n267_), .B0(new_new_n270_), .B1(new_new_n291_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n164_), .Y(new_new_n399_));
  AOI220     g377(.A0(i_3_), .A1(new_new_n272_), .B0(new_new_n258_), .B1(new_new_n206_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(new_new_n265_), .Y(new_new_n401_));
  NO3        g379(.A(new_new_n401_), .B(new_new_n399_), .C(new_new_n397_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n191_), .B(new_new_n95_), .Y(new_new_n403_));
  NA3        g381(.A(new_new_n303_), .B(new_new_n157_), .C(new_new_n83_), .Y(new_new_n404_));
  AOI210     g382(.A0(new_new_n404_), .A1(new_new_n403_), .B0(new_new_n301_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n188_), .B(i_10_), .Y(new_new_n406_));
  NA3        g384(.A(new_new_n247_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n273_), .B(new_new_n225_), .Y(new_new_n408_));
  OAI220     g386(.A0(new_new_n408_), .A1(new_new_n177_), .B0(new_new_n407_), .B1(new_new_n406_), .Y(new_new_n409_));
  NA3        g387(.A(new_new_n313_), .B(new_new_n312_), .C(i_5_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n293_), .B(new_new_n298_), .Y(new_new_n411_));
  OAI210     g389(.A0(new_new_n411_), .A1(new_new_n184_), .B0(new_new_n410_), .Y(new_new_n412_));
  NO3        g390(.A(new_new_n412_), .B(new_new_n409_), .C(new_new_n405_), .Y(new_new_n413_));
  AOI210     g391(.A0(new_new_n413_), .A1(new_new_n402_), .B0(new_new_n253_), .Y(new_new_n414_));
  NO4        g392(.A(new_new_n414_), .B(new_new_n396_), .C(new_new_n377_), .D(new_new_n358_), .Y(new_new_n415_));
  NO2        g393(.A(new_new_n70_), .B(i_13_), .Y(new_new_n416_));
  NO2        g394(.A(i_10_), .B(i_9_), .Y(new_new_n417_));
  NAi21      g395(.An(i_12_), .B(i_8_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n418_), .B(i_3_), .Y(new_new_n419_));
  INV        g397(.A(i_0_), .Y(new_new_n420_));
  NO3        g398(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n250_), .B(new_new_n96_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n422_), .B(new_new_n421_), .Y(new_new_n423_));
  NA2        g401(.A(i_8_), .B(i_9_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n263_), .B(new_new_n200_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(new_new_n424_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n242_), .B(new_new_n285_), .Y(new_new_n427_));
  NO3        g405(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n428_));
  INV        g406(.A(new_new_n428_), .Y(new_new_n429_));
  NA3        g407(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n430_));
  NO2        g408(.A(new_new_n429_), .B(new_new_n427_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n431_), .B(new_new_n426_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n272_), .B(new_new_n107_), .Y(new_new_n433_));
  OR2        g411(.A(new_new_n433_), .B(new_new_n202_), .Y(new_new_n434_));
  OA210      g412(.A0(new_new_n331_), .A1(new_new_n100_), .B0(new_new_n274_), .Y(new_new_n435_));
  OA220      g413(.A0(new_new_n435_), .A1(new_new_n156_), .B0(new_new_n434_), .B1(new_new_n222_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n95_), .B(i_13_), .Y(new_new_n437_));
  NO2        g415(.A(i_2_), .B(i_13_), .Y(new_new_n438_));
  NO3        g416(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n439_));
  NO2        g417(.A(i_6_), .B(i_7_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n439_), .Y(new_new_n441_));
  NO2        g419(.A(i_11_), .B(i_1_), .Y(new_new_n442_));
  OR2        g420(.A(i_11_), .B(i_8_), .Y(new_new_n443_));
  NOi21      g421(.An(i_2_), .B(i_7_), .Y(new_new_n444_));
  NAi31      g422(.An(new_new_n443_), .B(new_new_n444_), .C(i_0_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n388_), .B(i_6_), .Y(new_new_n446_));
  NA3        g424(.A(new_new_n446_), .B(i_1_), .C(new_new_n72_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n447_), .B(new_new_n445_), .Y(new_new_n448_));
  NO2        g426(.A(i_3_), .B(new_new_n188_), .Y(new_new_n449_));
  NO2        g427(.A(i_6_), .B(i_10_), .Y(new_new_n450_));
  NA4        g428(.A(new_new_n450_), .B(new_new_n290_), .C(new_new_n449_), .D(new_new_n227_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n451_), .B(new_new_n149_), .Y(new_new_n452_));
  NA3        g430(.A(new_new_n236_), .B(new_new_n166_), .C(new_new_n127_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n151_), .B(i_3_), .Y(new_new_n455_));
  NAi31      g433(.An(new_new_n454_), .B(new_new_n455_), .C(new_new_n219_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n368_), .B(new_new_n173_), .C(new_new_n143_), .Y(new_new_n457_));
  NA3        g435(.A(new_new_n457_), .B(new_new_n456_), .C(new_new_n453_), .Y(new_new_n458_));
  NO3        g436(.A(new_new_n458_), .B(new_new_n452_), .C(new_new_n448_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n421_), .B(new_new_n360_), .Y(new_new_n460_));
  NAi21      g438(.An(new_new_n212_), .B(new_new_n371_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n26_), .B(i_5_), .Y(new_new_n462_));
  NO2        g440(.A(i_0_), .B(new_new_n83_), .Y(new_new_n463_));
  NA3        g441(.A(new_new_n463_), .B(new_new_n462_), .C(new_new_n136_), .Y(new_new_n464_));
  OR3        g442(.A(new_new_n280_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n465_));
  NO2        g443(.A(new_new_n465_), .B(new_new_n464_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n27_), .B(i_10_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n290_), .B(new_new_n229_), .Y(new_new_n468_));
  OAI220     g446(.A0(new_new_n468_), .A1(new_new_n407_), .B0(new_new_n467_), .B1(new_new_n437_), .Y(new_new_n469_));
  NA4        g447(.A(new_new_n283_), .B(new_new_n217_), .C(new_new_n70_), .D(new_new_n227_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n441_), .Y(new_new_n471_));
  NO3        g449(.A(new_new_n471_), .B(new_new_n469_), .C(new_new_n466_), .Y(new_new_n472_));
  NA4        g450(.A(new_new_n472_), .B(new_new_n459_), .C(new_new_n436_), .D(new_new_n432_), .Y(new_new_n473_));
  NA3        g451(.A(new_new_n283_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n474_));
  OAI210     g452(.A0(new_new_n278_), .A1(new_new_n175_), .B0(new_new_n474_), .Y(new_new_n475_));
  AN2        g453(.A(new_new_n267_), .B(new_new_n224_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n476_), .B(new_new_n475_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n290_), .B(new_new_n158_), .Y(new_new_n478_));
  OAI210     g456(.A0(new_new_n478_), .A1(new_new_n222_), .B0(new_new_n284_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(new_new_n302_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n360_), .B(new_new_n218_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n336_), .B(new_new_n70_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n350_), .B(new_new_n342_), .Y(new_new_n483_));
  OR2        g461(.A(new_new_n481_), .B(new_new_n483_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n36_), .B(i_8_), .Y(new_new_n485_));
  NAi41      g463(.An(new_new_n482_), .B(new_new_n450_), .C(new_new_n485_), .D(new_new_n47_), .Y(new_new_n486_));
  AOI210     g464(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n389_), .Y(new_new_n487_));
  NA3        g465(.A(new_new_n487_), .B(new_new_n486_), .C(new_new_n484_), .Y(new_new_n488_));
  INV        g466(.A(new_new_n488_), .Y(new_new_n489_));
  AOI210     g467(.A0(new_new_n189_), .A1(i_9_), .B0(new_new_n249_), .Y(new_new_n490_));
  NO2        g468(.A(new_new_n490_), .B(new_new_n194_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n177_), .B(new_new_n83_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n492_), .B(new_new_n491_), .Y(new_new_n493_));
  NA4        g471(.A(new_new_n493_), .B(new_new_n489_), .C(new_new_n480_), .D(new_new_n477_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n362_), .B(new_new_n272_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n163_), .B(new_new_n495_), .Y(new_new_n496_));
  NO2        g474(.A(i_12_), .B(new_new_n188_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n497_), .B(new_new_n218_), .Y(new_new_n498_));
  NO3        g476(.A(i_6_), .B(new_new_n498_), .C(new_new_n433_), .Y(new_new_n499_));
  NOi31      g477(.An(new_new_n293_), .B(new_new_n388_), .C(new_new_n38_), .Y(new_new_n500_));
  OAI210     g478(.A0(new_new_n500_), .A1(new_new_n499_), .B0(new_new_n496_), .Y(new_new_n501_));
  NO2        g479(.A(i_8_), .B(i_7_), .Y(new_new_n502_));
  INV        g480(.A(i_5_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n503_), .B(new_new_n217_), .Y(new_new_n504_));
  AOI220     g482(.A0(new_new_n303_), .A1(new_new_n40_), .B0(new_new_n225_), .B1(new_new_n201_), .Y(new_new_n505_));
  OAI220     g483(.A0(new_new_n505_), .A1(new_new_n177_), .B0(new_new_n504_), .B1(new_new_n233_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n45_), .B(i_10_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(i_6_), .Y(new_new_n508_));
  NA3        g486(.A(new_new_n508_), .B(new_new_n506_), .C(new_new_n502_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n437_), .B(new_new_n128_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n510_), .B(new_new_n249_), .Y(new_new_n511_));
  NOi31      g489(.An(new_new_n270_), .B(new_new_n278_), .C(new_new_n175_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n512_), .B(new_new_n428_), .Y(new_new_n513_));
  NA4        g491(.A(new_new_n513_), .B(new_new_n511_), .C(new_new_n509_), .D(new_new_n501_), .Y(new_new_n514_));
  NA3        g492(.A(new_new_n213_), .B(new_new_n68_), .C(new_new_n45_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n263_), .B(new_new_n81_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n515_), .A1(new_new_n326_), .B0(new_new_n516_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n273_), .B(new_new_n267_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(new_new_n167_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n417_), .B(new_new_n215_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n520_), .B(new_new_n521_), .Y(new_new_n522_));
  AOI210     g500(.A0(new_new_n343_), .A1(new_new_n47_), .B0(new_new_n347_), .Y(new_new_n523_));
  NA2        g501(.A(i_0_), .B(new_new_n48_), .Y(new_new_n524_));
  NA3        g502(.A(new_new_n497_), .B(new_new_n255_), .C(new_new_n524_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n523_), .B(new_new_n525_), .Y(new_new_n526_));
  NO4        g504(.A(new_new_n526_), .B(new_new_n522_), .C(new_new_n519_), .D(new_new_n517_), .Y(new_new_n527_));
  NO4        g505(.A(new_new_n243_), .B(new_new_n43_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n528_));
  NO3        g506(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n223_), .B(new_new_n36_), .Y(new_new_n530_));
  AN2        g508(.A(new_new_n530_), .B(new_new_n529_), .Y(new_new_n531_));
  OA210      g509(.A0(new_new_n531_), .A1(new_new_n528_), .B0(new_new_n336_), .Y(new_new_n532_));
  NO2        g510(.A(new_new_n388_), .B(i_1_), .Y(new_new_n533_));
  NOi31      g511(.An(new_new_n533_), .B(new_new_n422_), .C(new_new_n70_), .Y(new_new_n534_));
  AN4        g512(.A(new_new_n534_), .B(new_new_n385_), .C(new_new_n462_), .D(i_2_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n398_), .B(new_new_n171_), .Y(new_new_n536_));
  NO3        g514(.A(new_new_n536_), .B(new_new_n535_), .C(new_new_n532_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n113_), .B(new_new_n23_), .Y(new_new_n538_));
  NA2        g516(.A(new_new_n293_), .B(new_new_n158_), .Y(new_new_n539_));
  AOI220     g517(.A0(new_new_n539_), .A1(new_new_n408_), .B0(new_new_n178_), .B1(new_new_n176_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n193_), .B(new_new_n37_), .Y(new_new_n541_));
  NOi31      g519(.An(new_new_n140_), .B(new_new_n541_), .C(new_new_n309_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n542_), .B(new_new_n540_), .Y(new_new_n543_));
  INV        g521(.A(new_new_n296_), .Y(new_new_n544_));
  NO2        g522(.A(i_12_), .B(new_new_n83_), .Y(new_new_n545_));
  NA3        g523(.A(new_new_n545_), .B(new_new_n255_), .C(new_new_n524_), .Y(new_new_n546_));
  NA3        g524(.A(new_new_n361_), .B(new_new_n263_), .C(new_new_n213_), .Y(new_new_n547_));
  AOI210     g525(.A0(new_new_n547_), .A1(new_new_n546_), .B0(new_new_n544_), .Y(new_new_n548_));
  NA2        g526(.A(new_new_n168_), .B(i_0_), .Y(new_new_n549_));
  NO3        g527(.A(new_new_n549_), .B(new_new_n319_), .C(new_new_n278_), .Y(new_new_n550_));
  OR2        g528(.A(i_2_), .B(i_5_), .Y(new_new_n551_));
  OR2        g529(.A(new_new_n551_), .B(new_new_n380_), .Y(new_new_n552_));
  AOI210     g530(.A0(new_new_n351_), .A1(new_new_n235_), .B0(new_new_n193_), .Y(new_new_n553_));
  AOI210     g531(.A0(new_new_n553_), .A1(new_new_n552_), .B0(new_new_n461_), .Y(new_new_n554_));
  NO3        g532(.A(new_new_n554_), .B(new_new_n550_), .C(new_new_n548_), .Y(new_new_n555_));
  NA4        g533(.A(new_new_n555_), .B(new_new_n543_), .C(new_new_n537_), .D(new_new_n527_), .Y(new_new_n556_));
  NO4        g534(.A(new_new_n556_), .B(new_new_n514_), .C(new_new_n494_), .D(new_new_n473_), .Y(new_new_n557_));
  NA4        g535(.A(new_new_n557_), .B(new_new_n415_), .C(new_new_n335_), .D(new_new_n289_), .Y(mai7));
  NO2        g536(.A(new_new_n92_), .B(new_new_n52_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n107_), .B(new_new_n89_), .Y(new_new_n560_));
  NA2        g538(.A(i_3_), .B(new_new_n560_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n450_), .B(new_new_n81_), .Y(new_new_n562_));
  NA2        g540(.A(i_11_), .B(new_new_n188_), .Y(new_new_n563_));
  NA2        g541(.A(new_new_n138_), .B(new_new_n563_), .Y(new_new_n564_));
  OAI210     g542(.A0(new_new_n564_), .A1(new_new_n562_), .B0(new_new_n561_), .Y(new_new_n565_));
  NA3        g543(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n227_), .B(i_4_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n567_), .B(i_8_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n104_), .B(new_new_n566_), .Y(new_new_n569_));
  NA2        g547(.A(i_2_), .B(new_new_n83_), .Y(new_new_n570_));
  OAI210     g548(.A0(new_new_n86_), .A1(new_new_n198_), .B0(new_new_n199_), .Y(new_new_n571_));
  NO2        g549(.A(i_7_), .B(new_new_n37_), .Y(new_new_n572_));
  NA2        g550(.A(i_4_), .B(i_8_), .Y(new_new_n573_));
  NO3        g551(.A(new_new_n569_), .B(new_new_n565_), .C(new_new_n559_), .Y(new_new_n574_));
  AOI210     g552(.A0(new_new_n123_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n575_));
  AOI210     g553(.A0(new_new_n575_), .A1(new_new_n227_), .B0(new_new_n155_), .Y(new_new_n576_));
  OR2        g554(.A(i_6_), .B(i_10_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n577_), .B(new_new_n23_), .Y(new_new_n578_));
  OR3        g556(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n579_));
  NO3        g557(.A(new_new_n579_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n580_));
  INV        g558(.A(new_new_n195_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n580_), .B(new_new_n578_), .Y(new_new_n582_));
  OA220      g560(.A0(new_new_n582_), .A1(new_new_n544_), .B0(new_new_n576_), .B1(new_new_n251_), .Y(new_new_n583_));
  AOI210     g561(.A0(new_new_n583_), .A1(new_new_n574_), .B0(new_new_n60_), .Y(new_new_n584_));
  NOi21      g562(.An(i_11_), .B(i_7_), .Y(new_new_n585_));
  AO210      g563(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n586_), .B(new_new_n585_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n587_), .B(new_new_n201_), .Y(new_new_n588_));
  NA3        g566(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n588_), .B(new_new_n60_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n85_), .B(new_new_n60_), .Y(new_new_n591_));
  AO210      g569(.A0(new_new_n591_), .A1(new_new_n355_), .B0(new_new_n41_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n219_), .B(new_new_n60_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n60_), .B(i_9_), .Y(new_new_n594_));
  NO2        g572(.A(i_1_), .B(i_12_), .Y(new_new_n595_));
  NA3        g573(.A(new_new_n595_), .B(new_new_n109_), .C(new_new_n24_), .Y(new_new_n596_));
  BUFFER     g574(.A(new_new_n596_), .Y(new_new_n597_));
  NA3        g575(.A(new_new_n597_), .B(new_new_n593_), .C(new_new_n592_), .Y(new_new_n598_));
  OAI210     g576(.A0(new_new_n598_), .A1(new_new_n590_), .B0(i_6_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n589_), .B(new_new_n107_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n600_), .B(new_new_n545_), .Y(new_new_n601_));
  NO2        g579(.A(i_6_), .B(i_11_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n601_), .B(new_new_n423_), .Y(new_new_n603_));
  NO4        g581(.A(new_new_n211_), .B(new_new_n123_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n604_), .B(new_new_n594_), .Y(new_new_n605_));
  INV        g583(.A(new_new_n605_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n502_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n607_));
  INV        g585(.A(i_2_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n132_), .B(i_9_), .Y(new_new_n609_));
  NA3        g587(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n47_), .B(i_1_), .Y(new_new_n611_));
  NA3        g589(.A(new_new_n611_), .B(new_new_n250_), .C(new_new_n45_), .Y(new_new_n612_));
  OAI220     g590(.A0(new_new_n612_), .A1(new_new_n610_), .B0(new_new_n609_), .B1(new_new_n608_), .Y(new_new_n613_));
  NA3        g591(.A(new_new_n594_), .B(new_new_n296_), .C(i_6_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n614_), .B(new_new_n23_), .Y(new_new_n615_));
  AOI210     g593(.A0(new_new_n442_), .A1(new_new_n391_), .B0(new_new_n232_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n616_), .B(new_new_n570_), .Y(new_new_n617_));
  NAi21      g595(.An(new_new_n607_), .B(new_new_n91_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n611_), .B(new_new_n250_), .Y(new_new_n619_));
  NO2        g597(.A(i_11_), .B(new_new_n37_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n24_), .Y(new_new_n621_));
  OAI210     g599(.A0(new_new_n621_), .A1(new_new_n619_), .B0(new_new_n618_), .Y(new_new_n622_));
  OR4        g600(.A(new_new_n622_), .B(new_new_n617_), .C(new_new_n615_), .D(new_new_n613_), .Y(new_new_n623_));
  NO3        g601(.A(new_new_n623_), .B(new_new_n606_), .C(new_new_n603_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n227_), .B(new_new_n100_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n585_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n626_), .B(i_1_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n627_), .B(new_new_n579_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n387_), .B(new_new_n83_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n628_), .B(new_new_n47_), .Y(new_new_n630_));
  NA2        g608(.A(i_3_), .B(new_new_n188_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n113_), .Y(new_new_n632_));
  AN2        g610(.A(new_new_n632_), .B(new_new_n508_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n223_), .B(new_new_n45_), .Y(new_new_n634_));
  NO3        g612(.A(new_new_n634_), .B(new_new_n286_), .C(new_new_n228_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n114_), .B(new_new_n37_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n636_), .B(i_6_), .Y(new_new_n637_));
  NO2        g615(.A(new_new_n83_), .B(i_9_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n60_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n639_), .B(new_new_n595_), .Y(new_new_n640_));
  NO4        g618(.A(new_new_n640_), .B(new_new_n637_), .C(new_new_n635_), .D(i_4_), .Y(new_new_n641_));
  NA2        g619(.A(i_1_), .B(i_3_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n424_), .B(new_new_n92_), .Y(new_new_n643_));
  INV        g621(.A(new_new_n643_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n642_), .Y(new_new_n645_));
  NO3        g623(.A(new_new_n645_), .B(new_new_n641_), .C(new_new_n633_), .Y(new_new_n646_));
  NA4        g624(.A(new_new_n646_), .B(new_new_n630_), .C(new_new_n624_), .D(new_new_n599_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n350_), .B(new_new_n349_), .Y(new_new_n648_));
  INV        g626(.A(new_new_n648_), .Y(new_new_n649_));
  NA2        g627(.A(new_new_n649_), .B(i_1_), .Y(new_new_n650_));
  AOI210     g628(.A0(new_new_n250_), .A1(new_new_n96_), .B0(i_1_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n348_), .B(i_2_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n652_), .B(new_new_n651_), .Y(new_new_n653_));
  OAI210     g631(.A0(new_new_n614_), .A1(new_new_n418_), .B0(new_new_n653_), .Y(new_new_n654_));
  INV        g632(.A(new_new_n654_), .Y(new_new_n655_));
  AOI210     g633(.A0(new_new_n655_), .A1(new_new_n650_), .B0(i_13_), .Y(new_new_n656_));
  OR2        g634(.A(i_11_), .B(i_7_), .Y(new_new_n657_));
  NA3        g635(.A(new_new_n657_), .B(new_new_n105_), .C(new_new_n132_), .Y(new_new_n658_));
  AOI220     g636(.A0(new_new_n438_), .A1(new_new_n155_), .B0(i_2_), .B1(new_new_n132_), .Y(new_new_n659_));
  OAI210     g637(.A0(new_new_n659_), .A1(new_new_n45_), .B0(new_new_n658_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n52_), .B(i_12_), .Y(new_new_n661_));
  INV        g639(.A(new_new_n661_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n444_), .B(new_new_n24_), .Y(new_new_n663_));
  AOI220     g641(.A0(new_new_n663_), .A1(new_new_n629_), .B0(new_new_n236_), .B1(new_new_n126_), .Y(new_new_n664_));
  OAI220     g642(.A0(new_new_n664_), .A1(new_new_n41_), .B0(new_new_n662_), .B1(new_new_n92_), .Y(new_new_n665_));
  AOI210     g643(.A0(new_new_n660_), .A1(new_new_n310_), .B0(new_new_n665_), .Y(new_new_n666_));
  INV        g644(.A(new_new_n113_), .Y(new_new_n667_));
  AOI220     g645(.A0(new_new_n667_), .A1(new_new_n69_), .B0(new_new_n361_), .B1(new_new_n611_), .Y(new_new_n668_));
  NO2        g646(.A(new_new_n668_), .B(new_new_n233_), .Y(new_new_n669_));
  AOI210     g647(.A0(new_new_n418_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n670_));
  NOi31      g648(.An(new_new_n670_), .B(new_new_n562_), .C(new_new_n45_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n122_), .B(i_13_), .Y(new_new_n672_));
  NO2        g650(.A(new_new_n610_), .B(new_new_n113_), .Y(new_new_n673_));
  INV        g651(.A(new_new_n673_), .Y(new_new_n674_));
  OAI220     g652(.A0(new_new_n674_), .A1(new_new_n68_), .B0(new_new_n672_), .B1(new_new_n651_), .Y(new_new_n675_));
  NO3        g653(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n100_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n26_), .B(new_new_n188_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n677_), .B(i_7_), .Y(new_new_n678_));
  NO3        g656(.A(new_new_n444_), .B(new_new_n227_), .C(new_new_n83_), .Y(new_new_n679_));
  AOI210     g657(.A0(new_new_n679_), .A1(new_new_n678_), .B0(new_new_n676_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n91_), .B(new_new_n101_), .Y(new_new_n681_));
  OAI220     g659(.A0(new_new_n681_), .A1(new_new_n568_), .B0(new_new_n680_), .B1(new_new_n581_), .Y(new_new_n682_));
  NO4        g660(.A(new_new_n682_), .B(new_new_n675_), .C(new_new_n671_), .D(new_new_n669_), .Y(new_new_n683_));
  OR2        g661(.A(i_11_), .B(i_6_), .Y(new_new_n684_));
  NA3        g662(.A(new_new_n567_), .B(new_new_n677_), .C(i_7_), .Y(new_new_n685_));
  AOI210     g663(.A0(new_new_n685_), .A1(new_new_n674_), .B0(new_new_n684_), .Y(new_new_n686_));
  NA3        g664(.A(new_new_n381_), .B(new_new_n572_), .C(new_new_n96_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n602_), .B(i_13_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n101_), .B(new_new_n677_), .Y(new_new_n689_));
  NAi21      g667(.An(i_11_), .B(i_12_), .Y(new_new_n690_));
  NOi41      g668(.An(new_new_n110_), .B(new_new_n690_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n691_));
  NO3        g669(.A(new_new_n444_), .B(new_new_n545_), .C(new_new_n573_), .Y(new_new_n692_));
  AOI220     g670(.A0(new_new_n692_), .A1(new_new_n290_), .B0(new_new_n691_), .B1(new_new_n689_), .Y(new_new_n693_));
  NA3        g671(.A(new_new_n693_), .B(new_new_n688_), .C(new_new_n687_), .Y(new_new_n694_));
  OAI210     g672(.A0(new_new_n694_), .A1(new_new_n686_), .B0(new_new_n60_), .Y(new_new_n695_));
  NO2        g673(.A(i_2_), .B(i_12_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n347_), .B(new_new_n696_), .Y(new_new_n697_));
  NO3        g675(.A(i_9_), .B(i_3_), .C(new_new_n567_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n698_), .B(new_new_n347_), .Y(new_new_n699_));
  NO2        g677(.A(new_new_n123_), .B(i_2_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n700_), .B(new_new_n595_), .Y(new_new_n701_));
  NA3        g679(.A(new_new_n701_), .B(new_new_n699_), .C(new_new_n697_), .Y(new_new_n702_));
  NA3        g680(.A(new_new_n702_), .B(new_new_n46_), .C(new_new_n218_), .Y(new_new_n703_));
  NA4        g681(.A(new_new_n703_), .B(new_new_n695_), .C(new_new_n683_), .D(new_new_n666_), .Y(new_new_n704_));
  OR4        g682(.A(new_new_n704_), .B(new_new_n656_), .C(new_new_n647_), .D(new_new_n584_), .Y(mai5));
  NA2        g683(.A(new_new_n626_), .B(new_new_n252_), .Y(new_new_n706_));
  AN2        g684(.A(new_new_n24_), .B(i_10_), .Y(new_new_n707_));
  NA3        g685(.A(new_new_n707_), .B(new_new_n696_), .C(new_new_n107_), .Y(new_new_n708_));
  NO2        g686(.A(new_new_n568_), .B(i_11_), .Y(new_new_n709_));
  NA2        g687(.A(new_new_n86_), .B(new_new_n709_), .Y(new_new_n710_));
  NA3        g688(.A(new_new_n710_), .B(new_new_n708_), .C(new_new_n706_), .Y(new_new_n711_));
  NO3        g689(.A(i_11_), .B(new_new_n227_), .C(i_13_), .Y(new_new_n712_));
  NO2        g690(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n713_));
  NA2        g691(.A(i_12_), .B(i_8_), .Y(new_new_n714_));
  OAI210     g692(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n714_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n417_), .Y(new_new_n716_));
  AOI220     g694(.A0(new_new_n296_), .A1(new_new_n538_), .B0(new_new_n715_), .B1(new_new_n713_), .Y(new_new_n717_));
  INV        g695(.A(new_new_n717_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n718_), .B(new_new_n711_), .Y(new_new_n719_));
  INV        g697(.A(new_new_n166_), .Y(new_new_n720_));
  INV        g698(.A(new_new_n236_), .Y(new_new_n721_));
  OAI210     g699(.A0(new_new_n652_), .A1(new_new_n419_), .B0(new_new_n110_), .Y(new_new_n722_));
  AOI210     g700(.A0(new_new_n722_), .A1(new_new_n721_), .B0(new_new_n720_), .Y(new_new_n723_));
  NO2        g701(.A(new_new_n424_), .B(new_new_n26_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n724_), .B(new_new_n391_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(i_2_), .Y(new_new_n726_));
  INV        g704(.A(new_new_n726_), .Y(new_new_n727_));
  AOI210     g705(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n388_), .Y(new_new_n728_));
  AOI210     g706(.A0(new_new_n728_), .A1(new_new_n727_), .B0(new_new_n723_), .Y(new_new_n729_));
  NO2        g707(.A(new_new_n185_), .B(new_new_n120_), .Y(new_new_n730_));
  OAI210     g708(.A0(new_new_n730_), .A1(new_new_n713_), .B0(i_2_), .Y(new_new_n731_));
  INV        g709(.A(new_new_n167_), .Y(new_new_n732_));
  NO3        g710(.A(new_new_n586_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n733_));
  AOI210     g711(.A0(new_new_n732_), .A1(new_new_n86_), .B0(new_new_n733_), .Y(new_new_n734_));
  AOI210     g712(.A0(new_new_n734_), .A1(new_new_n731_), .B0(new_new_n188_), .Y(new_new_n735_));
  OA210      g713(.A0(new_new_n587_), .A1(new_new_n121_), .B0(i_13_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n195_), .B(new_new_n198_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n145_), .B(new_new_n563_), .Y(new_new_n738_));
  AOI210     g716(.A0(new_new_n738_), .A1(new_new_n737_), .B0(new_new_n351_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n203_), .A1(new_new_n142_), .B0(new_new_n485_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n740_), .B(new_new_n391_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n101_), .B(new_new_n45_), .Y(new_new_n742_));
  INV        g720(.A(new_new_n279_), .Y(new_new_n743_));
  NA4        g721(.A(new_new_n743_), .B(new_new_n283_), .C(new_new_n119_), .D(new_new_n43_), .Y(new_new_n744_));
  OAI210     g722(.A0(new_new_n744_), .A1(new_new_n742_), .B0(new_new_n741_), .Y(new_new_n745_));
  NO4        g723(.A(new_new_n745_), .B(new_new_n739_), .C(new_new_n736_), .D(new_new_n735_), .Y(new_new_n746_));
  NA2        g724(.A(new_new_n538_), .B(new_new_n28_), .Y(new_new_n747_));
  NA2        g725(.A(new_new_n712_), .B(new_new_n256_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n748_), .B(new_new_n747_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n59_), .B(i_12_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n750_), .B(new_new_n121_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n751_), .B(new_new_n563_), .Y(new_new_n752_));
  AOI220     g730(.A0(new_new_n752_), .A1(new_new_n36_), .B0(new_new_n749_), .B1(new_new_n47_), .Y(new_new_n753_));
  NA4        g731(.A(new_new_n753_), .B(new_new_n746_), .C(new_new_n729_), .D(new_new_n719_), .Y(mai6));
  NO3        g732(.A(new_new_n246_), .B(new_new_n285_), .C(i_1_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n180_), .B(new_new_n133_), .Y(new_new_n756_));
  OAI210     g734(.A0(new_new_n756_), .A1(new_new_n755_), .B0(new_new_n700_), .Y(new_new_n757_));
  NA4        g735(.A(new_new_n363_), .B(new_new_n449_), .C(new_new_n68_), .D(new_new_n100_), .Y(new_new_n758_));
  INV        g736(.A(new_new_n758_), .Y(new_new_n759_));
  NO2        g737(.A(new_new_n214_), .B(new_new_n454_), .Y(new_new_n760_));
  NO2        g738(.A(i_11_), .B(i_9_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n759_), .B(new_new_n308_), .Y(new_new_n762_));
  AO210      g740(.A0(new_new_n762_), .A1(new_new_n757_), .B0(i_12_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n352_), .B(new_new_n313_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n545_), .B(new_new_n60_), .Y(new_new_n765_));
  BUFFER     g743(.A(new_new_n591_), .Y(new_new_n766_));
  NA3        g744(.A(new_new_n766_), .B(new_new_n765_), .C(new_new_n764_), .Y(new_new_n767_));
  INV        g745(.A(new_new_n192_), .Y(new_new_n768_));
  AOI220     g746(.A0(new_new_n768_), .A1(new_new_n761_), .B0(new_new_n767_), .B1(new_new_n70_), .Y(new_new_n769_));
  INV        g747(.A(new_new_n307_), .Y(new_new_n770_));
  NA2        g748(.A(new_new_n72_), .B(new_new_n126_), .Y(new_new_n771_));
  INV        g749(.A(new_new_n119_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n772_), .B(new_new_n47_), .Y(new_new_n773_));
  AOI210     g751(.A0(new_new_n773_), .A1(new_new_n771_), .B0(new_new_n770_), .Y(new_new_n774_));
  NO2        g752(.A(new_new_n243_), .B(i_9_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n775_), .B(new_new_n750_), .Y(new_new_n776_));
  AOI210     g754(.A0(new_new_n776_), .A1(new_new_n483_), .B0(new_new_n180_), .Y(new_new_n777_));
  NAi32      g755(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n778_));
  NO2        g756(.A(new_new_n684_), .B(new_new_n778_), .Y(new_new_n779_));
  OR3        g757(.A(new_new_n779_), .B(new_new_n777_), .C(new_new_n774_), .Y(new_new_n780_));
  NO2        g758(.A(new_new_n657_), .B(i_2_), .Y(new_new_n781_));
  NA2        g759(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n782_));
  NO2        g760(.A(new_new_n782_), .B(new_new_n380_), .Y(new_new_n783_));
  NA2        g761(.A(new_new_n783_), .B(new_new_n781_), .Y(new_new_n784_));
  OR2        g762(.A(new_new_n587_), .B(new_new_n419_), .Y(new_new_n785_));
  NA3        g763(.A(new_new_n785_), .B(new_new_n141_), .C(new_new_n66_), .Y(new_new_n786_));
  OR2        g764(.A(new_new_n716_), .B(new_new_n36_), .Y(new_new_n787_));
  NA3        g765(.A(new_new_n787_), .B(new_new_n786_), .C(new_new_n784_), .Y(new_new_n788_));
  OAI210     g766(.A0(i_6_), .A1(i_11_), .B0(new_new_n84_), .Y(new_new_n789_));
  AOI220     g767(.A0(new_new_n789_), .A1(new_new_n529_), .B0(new_new_n760_), .B1(new_new_n678_), .Y(new_new_n790_));
  NA2        g768(.A(new_new_n369_), .B(new_new_n67_), .Y(new_new_n791_));
  NA3        g769(.A(new_new_n791_), .B(new_new_n790_), .C(new_new_n571_), .Y(new_new_n792_));
  BUFFER     g770(.A(new_new_n85_), .Y(new_new_n793_));
  NA3        g771(.A(new_new_n793_), .B(new_new_n450_), .C(new_new_n213_), .Y(new_new_n794_));
  AOI210     g772(.A0(new_new_n419_), .A1(new_new_n417_), .B0(new_new_n528_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n577_), .B(new_new_n101_), .Y(new_new_n796_));
  OAI210     g774(.A0(new_new_n796_), .A1(new_new_n111_), .B0(new_new_n379_), .Y(new_new_n797_));
  INV        g775(.A(new_new_n552_), .Y(new_new_n798_));
  NA3        g776(.A(new_new_n798_), .B(new_new_n307_), .C(i_7_), .Y(new_new_n799_));
  NA4        g777(.A(new_new_n799_), .B(new_new_n797_), .C(new_new_n795_), .D(new_new_n794_), .Y(new_new_n800_));
  NO4        g778(.A(new_new_n800_), .B(new_new_n792_), .C(new_new_n788_), .D(new_new_n780_), .Y(new_new_n801_));
  NA4        g779(.A(new_new_n801_), .B(new_new_n769_), .C(new_new_n763_), .D(new_new_n357_), .Y(mai3));
  NA2        g780(.A(i_6_), .B(i_7_), .Y(new_new_n803_));
  NO2        g781(.A(new_new_n803_), .B(i_0_), .Y(new_new_n804_));
  NO2        g782(.A(i_11_), .B(new_new_n227_), .Y(new_new_n805_));
  OAI210     g783(.A0(new_new_n804_), .A1(new_new_n270_), .B0(new_new_n805_), .Y(new_new_n806_));
  NO2        g784(.A(new_new_n806_), .B(new_new_n188_), .Y(new_new_n807_));
  NO3        g785(.A(new_new_n420_), .B(new_new_n89_), .C(new_new_n45_), .Y(new_new_n808_));
  OA210      g786(.A0(new_new_n808_), .A1(new_new_n807_), .B0(new_new_n168_), .Y(new_new_n809_));
  NA2        g787(.A(new_new_n381_), .B(new_new_n46_), .Y(new_new_n810_));
  AN2        g788(.A(new_new_n422_), .B(new_new_n53_), .Y(new_new_n811_));
  INV        g789(.A(new_new_n811_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n812_), .B(new_new_n48_), .Y(new_new_n813_));
  NO4        g791(.A(new_new_n353_), .B(new_new_n360_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n670_), .B(new_new_n638_), .Y(new_new_n815_));
  NA2        g793(.A(new_new_n311_), .B(i_5_), .Y(new_new_n816_));
  OAI220     g794(.A0(new_new_n816_), .A1(new_new_n815_), .B0(new_new_n988_), .B1(new_new_n60_), .Y(new_new_n817_));
  NOi21      g795(.An(i_5_), .B(i_9_), .Y(new_new_n818_));
  NA2        g796(.A(new_new_n818_), .B(new_new_n416_), .Y(new_new_n819_));
  BUFFER     g797(.A(new_new_n250_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n820_), .B(new_new_n442_), .Y(new_new_n821_));
  NO3        g799(.A(new_new_n384_), .B(new_new_n250_), .C(new_new_n70_), .Y(new_new_n822_));
  NO2        g800(.A(new_new_n169_), .B(new_new_n142_), .Y(new_new_n823_));
  AOI210     g801(.A0(new_new_n823_), .A1(new_new_n235_), .B0(new_new_n822_), .Y(new_new_n824_));
  OAI220     g802(.A0(new_new_n824_), .A1(new_new_n175_), .B0(new_new_n821_), .B1(new_new_n819_), .Y(new_new_n825_));
  NO4        g803(.A(new_new_n825_), .B(new_new_n817_), .C(new_new_n813_), .D(new_new_n809_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n180_), .B(new_new_n24_), .Y(new_new_n827_));
  NO2        g805(.A(new_new_n636_), .B(new_new_n560_), .Y(new_new_n828_));
  NO2        g806(.A(new_new_n828_), .B(new_new_n827_), .Y(new_new_n829_));
  INV        g807(.A(new_new_n829_), .Y(new_new_n830_));
  NO2        g808(.A(new_new_n363_), .B(new_new_n271_), .Y(new_new_n831_));
  NA2        g809(.A(new_new_n831_), .B(new_new_n673_), .Y(new_new_n832_));
  NO4        g810(.A(new_new_n551_), .B(new_new_n211_), .C(new_new_n388_), .D(new_new_n380_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n833_), .B(i_11_), .Y(new_new_n834_));
  AN2        g812(.A(new_new_n95_), .B(new_new_n234_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n712_), .B(new_new_n308_), .Y(new_new_n836_));
  AOI210     g814(.A0(new_new_n450_), .A1(new_new_n86_), .B0(new_new_n55_), .Y(new_new_n837_));
  OAI220     g815(.A0(new_new_n837_), .A1(new_new_n836_), .B0(new_new_n621_), .B1(new_new_n504_), .Y(new_new_n838_));
  NO2        g816(.A(new_new_n245_), .B(new_new_n147_), .Y(new_new_n839_));
  INV        g817(.A(new_new_n507_), .Y(new_new_n840_));
  NO4        g818(.A(new_new_n113_), .B(new_new_n55_), .C(new_new_n631_), .D(i_5_), .Y(new_new_n841_));
  AO220      g819(.A0(new_new_n841_), .A1(new_new_n840_), .B0(new_new_n839_), .B1(i_6_), .Y(new_new_n842_));
  AOI220     g820(.A0(new_new_n311_), .A1(new_new_n97_), .B0(new_new_n180_), .B1(new_new_n81_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n533_), .B(i_4_), .Y(new_new_n844_));
  INV        g822(.A(new_new_n183_), .Y(new_new_n845_));
  OAI220     g823(.A0(new_new_n845_), .A1(new_new_n836_), .B0(new_new_n844_), .B1(new_new_n843_), .Y(new_new_n846_));
  NO4        g824(.A(new_new_n846_), .B(new_new_n842_), .C(new_new_n838_), .D(new_new_n835_), .Y(new_new_n847_));
  NA4        g825(.A(new_new_n847_), .B(new_new_n834_), .C(new_new_n832_), .D(new_new_n830_), .Y(new_new_n848_));
  NA2        g826(.A(i_11_), .B(i_9_), .Y(new_new_n849_));
  NO2        g827(.A(new_new_n48_), .B(i_7_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n368_), .B(new_new_n173_), .Y(new_new_n851_));
  NA2        g829(.A(new_new_n851_), .B(new_new_n154_), .Y(new_new_n852_));
  NO2        g830(.A(new_new_n849_), .B(new_new_n70_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n169_), .B(i_0_), .Y(new_new_n854_));
  INV        g832(.A(new_new_n854_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n440_), .B(new_new_n221_), .Y(new_new_n856_));
  AOI210     g834(.A0(new_new_n350_), .A1(new_new_n42_), .B0(new_new_n378_), .Y(new_new_n857_));
  OAI220     g835(.A0(new_new_n857_), .A1(new_new_n819_), .B0(new_new_n856_), .B1(new_new_n855_), .Y(new_new_n858_));
  NO2        g836(.A(new_new_n858_), .B(new_new_n852_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n620_), .B(new_new_n116_), .Y(new_new_n860_));
  NO2        g838(.A(i_6_), .B(new_new_n860_), .Y(new_new_n861_));
  AOI210     g839(.A0(new_new_n418_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n862_));
  NA2        g840(.A(new_new_n166_), .B(new_new_n102_), .Y(new_new_n863_));
  NOi32      g841(.An(new_new_n862_), .Bn(new_new_n183_), .C(new_new_n863_), .Y(new_new_n864_));
  NA2        g842(.A(new_new_n572_), .B(new_new_n308_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n865_), .B(new_new_n810_), .Y(new_new_n866_));
  NO3        g844(.A(new_new_n866_), .B(new_new_n864_), .C(new_new_n861_), .Y(new_new_n867_));
  NOi21      g845(.An(i_7_), .B(i_5_), .Y(new_new_n868_));
  OR2        g846(.A(new_new_n863_), .B(new_new_n483_), .Y(new_new_n869_));
  NO3        g847(.A(new_new_n374_), .B(new_new_n339_), .C(new_new_n338_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n248_), .B(new_new_n297_), .Y(new_new_n871_));
  INV        g849(.A(new_new_n690_), .Y(new_new_n872_));
  AOI210     g850(.A0(new_new_n872_), .A1(new_new_n871_), .B0(new_new_n870_), .Y(new_new_n873_));
  NA4        g851(.A(new_new_n873_), .B(new_new_n869_), .C(new_new_n867_), .D(new_new_n859_), .Y(new_new_n874_));
  AN2        g852(.A(new_new_n310_), .B(new_new_n308_), .Y(new_new_n875_));
  AN2        g853(.A(new_new_n875_), .B(new_new_n823_), .Y(new_new_n876_));
  INV        g854(.A(new_new_n876_), .Y(new_new_n877_));
  OA210      g855(.A0(new_new_n440_), .A1(new_new_n217_), .B0(new_new_n439_), .Y(new_new_n878_));
  NA2        g856(.A(new_new_n853_), .B(new_new_n283_), .Y(new_new_n879_));
  OAI210     g857(.A0(i_2_), .A1(new_new_n182_), .B0(new_new_n879_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n880_), .B(new_new_n440_), .Y(new_new_n881_));
  NAi21      g859(.An(i_9_), .B(i_5_), .Y(new_new_n882_));
  NO2        g860(.A(new_new_n882_), .B(new_new_n374_), .Y(new_new_n883_));
  NO2        g861(.A(new_new_n566_), .B(new_new_n104_), .Y(new_new_n884_));
  AOI220     g862(.A0(new_new_n884_), .A1(i_0_), .B0(new_new_n883_), .B1(new_new_n587_), .Y(new_new_n885_));
  NO2        g863(.A(new_new_n885_), .B(new_new_n83_), .Y(new_new_n886_));
  NO2        g864(.A(new_new_n886_), .B(new_new_n488_), .Y(new_new_n887_));
  NA3        g865(.A(new_new_n887_), .B(new_new_n881_), .C(new_new_n877_), .Y(new_new_n888_));
  NO3        g866(.A(new_new_n888_), .B(new_new_n874_), .C(new_new_n848_), .Y(new_new_n889_));
  NO2        g867(.A(i_0_), .B(new_new_n690_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n70_), .B(new_new_n45_), .Y(new_new_n891_));
  INV        g869(.A(new_new_n891_), .Y(new_new_n892_));
  NO3        g870(.A(new_new_n104_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n893_));
  AO220      g871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n890_), .B1(new_new_n168_), .Y(new_new_n894_));
  AOI210     g872(.A0(new_new_n765_), .A1(new_new_n648_), .B0(new_new_n863_), .Y(new_new_n895_));
  AOI210     g873(.A0(new_new_n894_), .A1(new_new_n327_), .B0(new_new_n895_), .Y(new_new_n896_));
  NA2        g874(.A(new_new_n700_), .B(new_new_n140_), .Y(new_new_n897_));
  INV        g875(.A(new_new_n897_), .Y(new_new_n898_));
  NA3        g876(.A(new_new_n898_), .B(new_new_n638_), .C(new_new_n70_), .Y(new_new_n899_));
  NA3        g877(.A(new_new_n804_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n900_));
  NA2        g878(.A(new_new_n805_), .B(i_9_), .Y(new_new_n901_));
  AOI210     g879(.A0(new_new_n900_), .A1(new_new_n464_), .B0(new_new_n901_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n235_), .B(new_new_n220_), .Y(new_new_n903_));
  NO2        g881(.A(new_new_n903_), .B(new_new_n147_), .Y(new_new_n904_));
  NO2        g882(.A(new_new_n904_), .B(new_new_n902_), .Y(new_new_n905_));
  NA3        g883(.A(new_new_n905_), .B(new_new_n899_), .C(new_new_n896_), .Y(new_new_n906_));
  NA2        g884(.A(new_new_n875_), .B(new_new_n351_), .Y(new_new_n907_));
  AOI210     g885(.A0(new_new_n278_), .A1(new_new_n156_), .B0(new_new_n907_), .Y(new_new_n908_));
  NA3        g886(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n909_));
  NA2        g887(.A(new_new_n850_), .B(new_new_n455_), .Y(new_new_n910_));
  AOI210     g888(.A0(new_new_n909_), .A1(new_new_n156_), .B0(new_new_n910_), .Y(new_new_n911_));
  NO2        g889(.A(new_new_n911_), .B(new_new_n908_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n534_), .B(new_new_n72_), .Y(new_new_n913_));
  NO3        g891(.A(new_new_n205_), .B(new_new_n360_), .C(i_0_), .Y(new_new_n914_));
  OAI210     g892(.A0(new_new_n914_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n915_));
  INV        g893(.A(new_new_n213_), .Y(new_new_n916_));
  OAI220     g894(.A0(new_new_n498_), .A1(new_new_n133_), .B0(i_12_), .B1(new_new_n581_), .Y(new_new_n917_));
  NA3        g895(.A(new_new_n917_), .B(new_new_n370_), .C(new_new_n916_), .Y(new_new_n918_));
  NA4        g896(.A(new_new_n918_), .B(new_new_n915_), .C(new_new_n913_), .D(new_new_n912_), .Y(new_new_n919_));
  INV        g897(.A(new_new_n108_), .Y(new_new_n920_));
  AOI220     g898(.A0(new_new_n868_), .A1(new_new_n455_), .B0(new_new_n804_), .B1(new_new_n157_), .Y(new_new_n921_));
  NA2        g899(.A(new_new_n330_), .B(new_new_n170_), .Y(new_new_n922_));
  OA220      g900(.A0(new_new_n922_), .A1(new_new_n921_), .B0(new_new_n920_), .B1(i_5_), .Y(new_new_n923_));
  AOI210     g901(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n924_));
  NA2        g902(.A(new_new_n924_), .B(new_new_n878_), .Y(new_new_n925_));
  NA3        g903(.A(new_new_n578_), .B(new_new_n180_), .C(new_new_n81_), .Y(new_new_n926_));
  INV        g904(.A(new_new_n926_), .Y(new_new_n927_));
  NO3        g905(.A(new_new_n810_), .B(new_new_n52_), .C(new_new_n48_), .Y(new_new_n928_));
  NA2        g906(.A(new_new_n460_), .B(new_new_n453_), .Y(new_new_n929_));
  NO3        g907(.A(new_new_n929_), .B(new_new_n928_), .C(new_new_n927_), .Y(new_new_n930_));
  NA3        g908(.A(new_new_n363_), .B(new_new_n166_), .C(new_new_n165_), .Y(new_new_n931_));
  NA3        g909(.A(new_new_n850_), .B(new_new_n270_), .C(new_new_n220_), .Y(new_new_n932_));
  NA2        g910(.A(new_new_n932_), .B(new_new_n931_), .Y(new_new_n933_));
  NOi31      g911(.An(new_new_n362_), .B(new_new_n891_), .C(new_new_n230_), .Y(new_new_n934_));
  NO3        g912(.A(new_new_n849_), .B(new_new_n213_), .C(new_new_n185_), .Y(new_new_n935_));
  NO3        g913(.A(new_new_n935_), .B(new_new_n934_), .C(new_new_n933_), .Y(new_new_n936_));
  NA4        g914(.A(new_new_n936_), .B(new_new_n930_), .C(new_new_n925_), .D(new_new_n923_), .Y(new_new_n937_));
  INV        g915(.A(new_new_n580_), .Y(new_new_n938_));
  NO3        g916(.A(new_new_n938_), .B(new_new_n524_), .C(new_new_n324_), .Y(new_new_n939_));
  INV        g917(.A(new_new_n939_), .Y(new_new_n940_));
  NA2        g918(.A(new_new_n759_), .B(new_new_n170_), .Y(new_new_n941_));
  NA3        g919(.A(new_new_n97_), .B(i_10_), .C(i_11_), .Y(new_new_n942_));
  NO2        g920(.A(new_new_n942_), .B(new_new_n149_), .Y(new_new_n943_));
  NA2        g921(.A(new_new_n868_), .B(new_new_n438_), .Y(new_new_n944_));
  NO2        g922(.A(new_new_n944_), .B(new_new_n639_), .Y(new_new_n945_));
  AOI210     g923(.A0(new_new_n945_), .A1(new_new_n854_), .B0(new_new_n943_), .Y(new_new_n946_));
  NA3        g924(.A(new_new_n946_), .B(new_new_n941_), .C(new_new_n940_), .Y(new_new_n947_));
  NO4        g925(.A(new_new_n947_), .B(new_new_n937_), .C(new_new_n919_), .D(new_new_n906_), .Y(new_new_n948_));
  NA2        g926(.A(new_new_n781_), .B(new_new_n37_), .Y(new_new_n949_));
  NA3        g927(.A(new_new_n862_), .B(new_new_n347_), .C(i_5_), .Y(new_new_n950_));
  NA3        g928(.A(new_new_n950_), .B(new_new_n949_), .C(new_new_n576_), .Y(new_new_n951_));
  NA2        g929(.A(new_new_n951_), .B(new_new_n201_), .Y(new_new_n952_));
  AN2        g930(.A(new_new_n657_), .B(new_new_n348_), .Y(new_new_n953_));
  NA2        g931(.A(new_new_n181_), .B(new_new_n183_), .Y(new_new_n954_));
  AO210      g932(.A0(new_new_n953_), .A1(new_new_n33_), .B0(new_new_n954_), .Y(new_new_n955_));
  OAI210     g933(.A0(new_new_n580_), .A1(new_new_n578_), .B0(new_new_n296_), .Y(new_new_n956_));
  NAi31      g934(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n957_));
  NO2        g935(.A(new_new_n67_), .B(new_new_n957_), .Y(new_new_n958_));
  INV        g936(.A(new_new_n958_), .Y(new_new_n959_));
  NA3        g937(.A(new_new_n959_), .B(new_new_n956_), .C(new_new_n955_), .Y(new_new_n960_));
  NO2        g938(.A(new_new_n430_), .B(new_new_n250_), .Y(new_new_n961_));
  NO4        g939(.A(new_new_n223_), .B(new_new_n139_), .C(new_new_n642_), .D(new_new_n37_), .Y(new_new_n962_));
  NO3        g940(.A(new_new_n962_), .B(new_new_n961_), .C(new_new_n833_), .Y(new_new_n963_));
  OAI210     g941(.A0(new_new_n942_), .A1(new_new_n142_), .B0(new_new_n963_), .Y(new_new_n964_));
  AOI210     g942(.A0(new_new_n960_), .A1(new_new_n48_), .B0(new_new_n964_), .Y(new_new_n965_));
  AOI210     g943(.A0(new_new_n965_), .A1(new_new_n952_), .B0(new_new_n70_), .Y(new_new_n966_));
  NO2        g944(.A(new_new_n531_), .B(new_new_n356_), .Y(new_new_n967_));
  NO2        g945(.A(new_new_n967_), .B(new_new_n720_), .Y(new_new_n968_));
  NA2        g946(.A(new_new_n248_), .B(new_new_n54_), .Y(new_new_n969_));
  AOI220     g947(.A0(new_new_n969_), .A1(new_new_n73_), .B0(new_new_n325_), .B1(new_new_n246_), .Y(new_new_n970_));
  NO2        g948(.A(new_new_n970_), .B(new_new_n227_), .Y(new_new_n971_));
  INV        g949(.A(new_new_n971_), .Y(new_new_n972_));
  NA2        g950(.A(new_new_n573_), .B(new_new_n211_), .Y(new_new_n973_));
  OAI210     g951(.A0(new_new_n973_), .A1(new_new_n862_), .B0(new_new_n201_), .Y(new_new_n974_));
  NA2        g952(.A(new_new_n158_), .B(i_5_), .Y(new_new_n975_));
  NO2        g953(.A(new_new_n974_), .B(new_new_n975_), .Y(new_new_n976_));
  NO4        g954(.A(new_new_n882_), .B(new_new_n443_), .C(new_new_n244_), .D(new_new_n243_), .Y(new_new_n977_));
  NO2        g955(.A(new_new_n977_), .B(new_new_n528_), .Y(new_new_n978_));
  INV        g956(.A(new_new_n340_), .Y(new_new_n979_));
  AOI210     g957(.A0(new_new_n979_), .A1(new_new_n978_), .B0(new_new_n41_), .Y(new_new_n980_));
  NO2        g958(.A(new_new_n980_), .B(new_new_n976_), .Y(new_new_n981_));
  OAI210     g959(.A0(new_new_n972_), .A1(i_4_), .B0(new_new_n981_), .Y(new_new_n982_));
  NO3        g960(.A(new_new_n982_), .B(new_new_n968_), .C(new_new_n966_), .Y(new_new_n983_));
  NA4        g961(.A(new_new_n983_), .B(new_new_n948_), .C(new_new_n889_), .D(new_new_n826_), .Y(mai4));
  INV        g962(.A(new_new_n237_), .Y(new_new_n987_));
  INV        g963(.A(new_new_n814_), .Y(new_new_n988_));
endmodule


