//Benchmark atmr_intb_466_0.25

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n268_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n302_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n327_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  INV        o035(.A(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n59_));
  NO2        o037(.A(ori_ori_n29_), .B(ori_ori_n58_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n61_));
  OAI210     o039(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n61_), .Y(ori_ori_n62_));
  AOI220     o040(.A0(ori_ori_n62_), .A1(ori_ori_n55_), .B0(ori_ori_n60_), .B1(ori_ori_n31_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(x05), .Y(ori_ori_n64_));
  NA2        o042(.A(x09), .B(x05), .Y(ori_ori_n65_));
  NA2        o043(.A(x10), .B(x06), .Y(ori_ori_n66_));
  NA3        o044(.A(ori_ori_n66_), .B(ori_ori_n65_), .C(ori_ori_n28_), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n67_), .B(x03), .Y(ori_ori_n68_));
  NOi31      o046(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n69_));
  NO2        o047(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n70_), .B(ori_ori_n36_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n70_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n72_));
  AOI210     o050(.A0(ori_ori_n71_), .A1(ori_ori_n48_), .B0(ori_ori_n72_), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n74_));
  NO2        o052(.A(x08), .B(x01), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n35_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n73_), .Y(ori_ori_n77_));
  AN2        o055(.A(ori_ori_n77_), .B(ori_ori_n68_), .Y(ori_ori_n78_));
  INV        o056(.A(ori_ori_n76_), .Y(ori_ori_n79_));
  NA2        o057(.A(x11), .B(x00), .Y(ori_ori_n80_));
  NO2        o058(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n81_));
  NOi21      o059(.An(ori_ori_n80_), .B(ori_ori_n81_), .Y(ori_ori_n82_));
  INV        o060(.A(ori_ori_n82_), .Y(ori_ori_n83_));
  NOi21      o061(.An(x01), .B(x10), .Y(ori_ori_n84_));
  NO2        o062(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n85_));
  NO3        o063(.A(ori_ori_n85_), .B(ori_ori_n84_), .C(x06), .Y(ori_ori_n86_));
  NA2        o064(.A(ori_ori_n86_), .B(ori_ori_n27_), .Y(ori_ori_n87_));
  OAI210     o065(.A0(ori_ori_n83_), .A1(x07), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  NO3        o066(.A(ori_ori_n88_), .B(ori_ori_n78_), .C(ori_ori_n64_), .Y(ori01));
  INV        o067(.A(x12), .Y(ori_ori_n90_));
  INV        o068(.A(x13), .Y(ori_ori_n91_));
  NO2        o069(.A(x10), .B(x01), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(ori_ori_n92_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n95_));
  NOi21      o073(.An(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n96_));
  NA2        o074(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n97_));
  NO2        o075(.A(ori_ori_n97_), .B(x05), .Y(ori_ori_n98_));
  INV        o076(.A(ori_ori_n96_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n66_), .Y(ori_ori_n100_));
  NA2        o078(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n101_));
  NA2        o079(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n102_), .B(ori_ori_n101_), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n105_));
  NA3        o083(.A(ori_ori_n105_), .B(ori_ori_n104_), .C(x13), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n107_));
  NOi21      o085(.An(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n108_));
  NO3        o086(.A(ori_ori_n108_), .B(x06), .C(x03), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n109_), .B(ori_ori_n100_), .Y(ori_ori_n110_));
  NA2        o088(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n111_));
  OAI210     o089(.A0(ori_ori_n75_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n115_));
  AOI210     o093(.A0(ori_ori_n115_), .A1(ori_ori_n49_), .B0(ori_ori_n114_), .Y(ori_ori_n116_));
  AN2        o094(.A(ori_ori_n116_), .B(ori_ori_n113_), .Y(ori_ori_n117_));
  NO2        o095(.A(x09), .B(x05), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(ori_ori_n47_), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n94_), .B(ori_ori_n49_), .Y(ori_ori_n120_));
  NA2        o098(.A(x09), .B(x00), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n95_), .B(ori_ori_n121_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n120_), .B(ori_ori_n117_), .Y(ori_ori_n123_));
  NO2        o101(.A(x03), .B(x02), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n76_), .B(ori_ori_n91_), .Y(ori_ori_n125_));
  OAI210     o103(.A0(ori_ori_n125_), .A1(ori_ori_n96_), .B0(ori_ori_n124_), .Y(ori_ori_n126_));
  OA210      o104(.A0(ori_ori_n123_), .A1(x11), .B0(ori_ori_n126_), .Y(ori_ori_n127_));
  OAI210     o105(.A0(ori_ori_n110_), .A1(ori_ori_n23_), .B0(ori_ori_n127_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n94_), .B(ori_ori_n40_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n129_), .B(ori_ori_n41_), .Y(ori_ori_n130_));
  NO2        o108(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n131_));
  AOI210     o109(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n130_), .B(ori_ori_n132_), .Y(ori_ori_n133_));
  NA2        o111(.A(x10), .B(x05), .Y(ori_ori_n134_));
  NO2        o112(.A(x09), .B(x01), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n95_), .B(x08), .Y(ori_ori_n136_));
  NOi21      o114(.An(x09), .B(x00), .Y(ori_ori_n137_));
  NO3        o115(.A(ori_ori_n74_), .B(ori_ori_n137_), .C(ori_ori_n47_), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n138_), .B(ori_ori_n102_), .Y(ori_ori_n139_));
  NA2        o117(.A(x06), .B(x05), .Y(ori_ori_n140_));
  OAI210     o118(.A0(ori_ori_n140_), .A1(ori_ori_n35_), .B0(ori_ori_n90_), .Y(ori_ori_n141_));
  AOI210     o119(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n141_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n142_), .B(ori_ori_n139_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n91_), .B(x12), .Y(ori_ori_n144_));
  AOI210     o122(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n144_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n146_), .B(x02), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n145_), .B(ori_ori_n143_), .Y(ori_ori_n148_));
  NA2        o126(.A(ori_ori_n148_), .B(ori_ori_n133_), .Y(ori_ori_n149_));
  AOI210     o127(.A0(ori_ori_n128_), .A1(ori_ori_n90_), .B0(ori_ori_n149_), .Y(ori_ori_n150_));
  INV        o128(.A(ori_ori_n67_), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n151_), .B(ori_ori_n113_), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n153_), .B(ori_ori_n112_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n152_), .B(x12), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n84_), .B(x06), .Y(ori_ori_n156_));
  AOI210     o134(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n157_));
  NO3        o135(.A(ori_ori_n157_), .B(ori_ori_n156_), .C(ori_ori_n41_), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n115_), .Y(ori_ori_n159_));
  OAI210     o137(.A0(ori_ori_n159_), .A1(ori_ori_n158_), .B0(x02), .Y(ori_ori_n160_));
  AOI210     o138(.A0(ori_ori_n160_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n161_));
  OAI210     o139(.A0(ori_ori_n155_), .A1(ori_ori_n53_), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  INV        o140(.A(ori_ori_n115_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n164_));
  NO2        o142(.A(ori_ori_n70_), .B(ori_ori_n36_), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n91_), .B(x03), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n167_));
  NOi21      o145(.An(x13), .B(x04), .Y(ori_ori_n168_));
  NO3        o146(.A(ori_ori_n168_), .B(ori_ori_n69_), .C(ori_ori_n137_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n169_), .B(x05), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n170_), .B(ori_ori_n167_), .Y(ori_ori_n171_));
  OAI210     o149(.A0(ori_ori_n297_), .A1(ori_ori_n163_), .B0(ori_ori_n171_), .Y(ori_ori_n172_));
  INV        o150(.A(ori_ori_n81_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n173_), .B(x12), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n175_));
  NO2        o153(.A(x06), .B(x00), .Y(ori_ori_n176_));
  INV        o154(.A(ori_ori_n66_), .Y(ori_ori_n177_));
  NO2        o155(.A(ori_ori_n177_), .B(x05), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n179_), .B(x03), .Y(ori_ori_n180_));
  OR2        o158(.A(ori_ori_n180_), .B(ori_ori_n178_), .Y(ori_ori_n181_));
  NA2        o159(.A(x13), .B(ori_ori_n90_), .Y(ori_ori_n182_));
  NA3        o160(.A(ori_ori_n182_), .B(ori_ori_n141_), .C(ori_ori_n82_), .Y(ori_ori_n183_));
  OAI210     o161(.A0(ori_ori_n181_), .A1(ori_ori_n175_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  AOI210     o162(.A0(ori_ori_n174_), .A1(ori_ori_n172_), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n185_), .A1(ori_ori_n162_), .B0(x07), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n65_), .B(ori_ori_n29_), .Y(ori_ori_n187_));
  NOi31      o165(.An(ori_ori_n111_), .B(ori_ori_n168_), .C(ori_ori_n137_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n188_), .B(ori_ori_n187_), .Y(ori_ori_n189_));
  NO2        o167(.A(x12), .B(x02), .Y(ori_ori_n190_));
  INV        o168(.A(ori_ori_n190_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n191_), .B(ori_ori_n173_), .Y(ori_ori_n192_));
  OA210      o170(.A0(ori_ori_n69_), .A1(ori_ori_n189_), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n194_), .B(x01), .Y(ori_ori_n195_));
  INV        o173(.A(ori_ori_n195_), .Y(ori_ori_n196_));
  AOI210     o174(.A0(ori_ori_n196_), .A1(ori_ori_n106_), .B0(ori_ori_n29_), .Y(ori_ori_n197_));
  NO3        o175(.A(ori_ori_n80_), .B(x12), .C(x03), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n197_), .B(ori_ori_n198_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n200_));
  NO3        o178(.A(ori_ori_n200_), .B(ori_ori_n157_), .C(ori_ori_n29_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n175_), .B(ori_ori_n28_), .Y(ori_ori_n202_));
  OAI210     o180(.A0(ori_ori_n201_), .A1(ori_ori_n163_), .B0(ori_ori_n202_), .Y(ori_ori_n203_));
  NA2        o181(.A(ori_ori_n203_), .B(ori_ori_n199_), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n204_), .B(ori_ori_n193_), .C(ori_ori_n186_), .Y(ori_ori_n205_));
  OAI210     o183(.A0(ori_ori_n150_), .A1(ori_ori_n57_), .B0(ori_ori_n205_), .Y(ori02));
  AOI210     o184(.A0(ori_ori_n111_), .A1(ori_ori_n76_), .B0(ori_ori_n104_), .Y(ori_ori_n207_));
  NOi21      o185(.An(ori_ori_n169_), .B(ori_ori_n135_), .Y(ori_ori_n208_));
  NO2        o186(.A(ori_ori_n208_), .B(ori_ori_n32_), .Y(ori_ori_n209_));
  OAI210     o187(.A0(ori_ori_n209_), .A1(ori_ori_n207_), .B0(ori_ori_n134_), .Y(ori_ori_n210_));
  INV        o188(.A(ori_ori_n134_), .Y(ori_ori_n211_));
  AOI220     o189(.A0(ori_ori_n157_), .A1(ori_ori_n211_), .B0(ori_ori_n125_), .B1(ori_ori_n124_), .Y(ori_ori_n212_));
  AOI210     o190(.A0(ori_ori_n212_), .A1(ori_ori_n210_), .B0(ori_ori_n48_), .Y(ori_ori_n213_));
  NO2        o191(.A(x05), .B(x02), .Y(ori_ori_n214_));
  OAI210     o192(.A0(ori_ori_n154_), .A1(ori_ori_n137_), .B0(ori_ori_n214_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n215_), .B(ori_ori_n115_), .Y(ori_ori_n216_));
  NAi21      o194(.An(ori_ori_n170_), .B(ori_ori_n297_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n179_), .B(ori_ori_n47_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  AN2        o197(.A(ori_ori_n166_), .B(ori_ori_n165_), .Y(ori_ori_n220_));
  BUFFER     o198(.A(ori_ori_n119_), .Y(ori_ori_n221_));
  AOI210     o199(.A0(ori_ori_n221_), .A1(ori_ori_n112_), .B0(x06), .Y(ori_ori_n222_));
  OAI210     o200(.A0(ori_ori_n222_), .A1(ori_ori_n220_), .B0(ori_ori_n85_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n223_), .B(ori_ori_n219_), .Y(ori_ori_n224_));
  NO3        o202(.A(ori_ori_n224_), .B(ori_ori_n216_), .C(ori_ori_n213_), .Y(ori_ori_n225_));
  INV        o203(.A(x13), .Y(ori_ori_n226_));
  AOI220     o204(.A0(x08), .A1(ori_ori_n226_), .B0(ori_ori_n146_), .B1(x08), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n200_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n228_), .B(ori_ori_n92_), .Y(ori_ori_n229_));
  NA2        o207(.A(ori_ori_n136_), .B(ori_ori_n93_), .Y(ori_ori_n230_));
  NA2        o208(.A(x12), .B(ori_ori_n103_), .Y(ori_ori_n231_));
  NA4        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .C(ori_ori_n229_), .D(ori_ori_n48_), .Y(ori_ori_n232_));
  INV        o210(.A(ori_ori_n146_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n233_), .B(ori_ori_n55_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n234_), .B(x02), .Y(ori_ori_n235_));
  NO3        o213(.A(ori_ori_n144_), .B(ori_ori_n131_), .C(ori_ori_n51_), .Y(ori_ori_n236_));
  OAI210     o214(.A0(ori_ori_n121_), .A1(ori_ori_n36_), .B0(ori_ori_n90_), .Y(ori_ori_n237_));
  OAI210     o215(.A0(ori_ori_n237_), .A1(ori_ori_n138_), .B0(ori_ori_n236_), .Y(ori_ori_n238_));
  NA3        o216(.A(ori_ori_n238_), .B(ori_ori_n235_), .C(x06), .Y(ori_ori_n239_));
  NA2        o217(.A(x09), .B(x03), .Y(ori_ori_n240_));
  OAI220     o218(.A0(ori_ori_n240_), .A1(ori_ori_n102_), .B0(ori_ori_n153_), .B1(ori_ori_n59_), .Y(ori_ori_n241_));
  NO3        o219(.A(ori_ori_n200_), .B(ori_ori_n101_), .C(x08), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n242_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n244_));
  NO3        o222(.A(ori_ori_n95_), .B(ori_ori_n102_), .C(ori_ori_n38_), .Y(ori_ori_n245_));
  AOI210     o223(.A0(ori_ori_n236_), .A1(ori_ori_n244_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  OAI210     o224(.A0(ori_ori_n243_), .A1(ori_ori_n28_), .B0(ori_ori_n246_), .Y(ori_ori_n247_));
  AO220      o225(.A0(ori_ori_n247_), .A1(x04), .B0(ori_ori_n241_), .B1(x05), .Y(ori_ori_n248_));
  AOI210     o226(.A0(ori_ori_n239_), .A1(ori_ori_n232_), .B0(ori_ori_n248_), .Y(ori_ori_n249_));
  OAI210     o227(.A0(ori_ori_n225_), .A1(x12), .B0(ori_ori_n249_), .Y(ori03));
  OR2        o228(.A(ori_ori_n42_), .B(ori_ori_n164_), .Y(ori_ori_n251_));
  AOI210     o229(.A0(ori_ori_n125_), .A1(ori_ori_n90_), .B0(ori_ori_n251_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n144_), .B(ori_ori_n124_), .Y(ori_ori_n253_));
  NA2        o231(.A(ori_ori_n253_), .B(ori_ori_n147_), .Y(ori_ori_n254_));
  OAI210     o232(.A0(ori_ori_n254_), .A1(ori_ori_n252_), .B0(x05), .Y(ori_ori_n255_));
  AOI210     o233(.A0(ori_ori_n166_), .A1(ori_ori_n71_), .B0(ori_ori_n98_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n256_), .B(ori_ori_n55_), .Y(ori_ori_n257_));
  NA2        o235(.A(ori_ori_n257_), .B(ori_ori_n90_), .Y(ori_ori_n258_));
  AOI210     o236(.A0(ori_ori_n119_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n135_), .B(ori_ori_n107_), .Y(ori_ori_n260_));
  OAI220     o238(.A0(ori_ori_n260_), .A1(ori_ori_n37_), .B0(ori_ori_n122_), .B1(x13), .Y(ori_ori_n261_));
  OAI210     o239(.A0(ori_ori_n261_), .A1(ori_ori_n259_), .B0(x04), .Y(ori_ori_n262_));
  NO3        o240(.A(x12), .B(ori_ori_n76_), .C(ori_ori_n55_), .Y(ori_ori_n263_));
  AOI210     o241(.A0(x13), .A1(ori_ori_n90_), .B0(ori_ori_n119_), .Y(ori_ori_n264_));
  AN2        o242(.A(x12), .B(ori_ori_n107_), .Y(ori_ori_n265_));
  NO3        o243(.A(ori_ori_n265_), .B(ori_ori_n264_), .C(ori_ori_n263_), .Y(ori_ori_n266_));
  NA4        o244(.A(ori_ori_n266_), .B(ori_ori_n262_), .C(ori_ori_n258_), .D(ori_ori_n255_), .Y(ori04));
  NO2        o245(.A(ori_ori_n79_), .B(ori_ori_n39_), .Y(ori_ori_n268_));
  XO2        o246(.A(ori_ori_n268_), .B(ori_ori_n182_), .Y(ori05));
  OAI210     o247(.A0(ori_ori_n23_), .A1(x03), .B0(ori_ori_n90_), .Y(ori_ori_n270_));
  OAI210     o248(.A0(ori_ori_n26_), .A1(ori_ori_n90_), .B0(x07), .Y(ori_ori_n271_));
  INV        o249(.A(ori_ori_n271_), .Y(ori_ori_n272_));
  BUFFER     o250(.A(ori_ori_n175_), .Y(ori_ori_n273_));
  NA2        o251(.A(ori_ori_n176_), .B(ori_ori_n173_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n274_), .B(ori_ori_n273_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n275_), .B(ori_ori_n90_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n33_), .B(ori_ori_n90_), .Y(ori_ori_n277_));
  AOI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n81_), .B0(x07), .Y(ori_ori_n278_));
  AOI220     o256(.A0(ori_ori_n278_), .A1(ori_ori_n276_), .B0(ori_ori_n272_), .B1(ori_ori_n270_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n298_), .B(x08), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n104_), .B(ori_ori_n28_), .Y(ori_ori_n281_));
  INV        o259(.A(ori_ori_n281_), .Y(ori_ori_n282_));
  OR3        o260(.A(ori_ori_n282_), .B(x12), .C(x03), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n283_), .B(x08), .Y(ori_ori_n284_));
  INV        o262(.A(ori_ori_n284_), .Y(ori_ori_n285_));
  NO2        o263(.A(ori_ori_n280_), .B(ori_ori_n285_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n56_), .B(x12), .Y(ori_ori_n287_));
  INV        o265(.A(x14), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n299_), .B(ori_ori_n53_), .Y(ori_ori_n289_));
  NO2        o267(.A(ori_ori_n289_), .B(ori_ori_n288_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n290_), .B(ori_ori_n287_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n95_), .B(ori_ori_n90_), .Y(ori_ori_n292_));
  OAI210     o270(.A0(ori_ori_n300_), .A1(ori_ori_n80_), .B0(ori_ori_n292_), .Y(ori_ori_n293_));
  NO4        o271(.A(ori_ori_n293_), .B(ori_ori_n291_), .C(ori_ori_n286_), .D(ori_ori_n279_), .Y(ori06));
  INV        o272(.A(ori_ori_n166_), .Y(ori_ori_n297_));
  INV        o273(.A(x02), .Y(ori_ori_n298_));
  INV        o274(.A(x01), .Y(ori_ori_n299_));
  INV        o275(.A(x06), .Y(ori_ori_n300_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NO2        m026(.A(x02), .B(x11), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  INV        m029(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(x07), .Y(mai_mai_n53_));
  OAI210     m031(.A0(mai_mai_n53_), .A1(mai_mai_n49_), .B0(mai_mai_n47_), .Y(mai_mai_n54_));
  NOi21      m032(.An(x01), .B(x09), .Y(mai_mai_n55_));
  INV        m033(.A(x00), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n56_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(x09), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m037(.A(x07), .Y(mai_mai_n60_));
  AOI220     m038(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n60_), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n58_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n63_));
  OAI220     m041(.A0(x02), .A1(mai_mai_n62_), .B0(mai_mai_n61_), .B1(mai_mai_n59_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n60_), .B(mai_mai_n48_), .Y(mai_mai_n65_));
  OAI210     m043(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n65_), .Y(mai_mai_n66_));
  AOI220     m044(.A0(mai_mai_n66_), .A1(mai_mai_n58_), .B0(mai_mai_n64_), .B1(mai_mai_n31_), .Y(mai_mai_n67_));
  AOI210     m045(.A0(mai_mai_n67_), .A1(mai_mai_n54_), .B0(x05), .Y(mai_mai_n68_));
  NA2        m046(.A(x09), .B(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x10), .B(x06), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n60_), .B(mai_mai_n41_), .Y(mai_mai_n71_));
  NOi31      m049(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n72_));
  NO2        m050(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n36_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n73_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n76_));
  NO2        m054(.A(x08), .B(x01), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n77_), .A1(mai_mai_n76_), .B0(mai_mai_n35_), .Y(mai_mai_n78_));
  NA2        m056(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n79_));
  INV        m057(.A(mai_mai_n78_), .Y(mai_mai_n80_));
  NO2        m058(.A(x06), .B(x05), .Y(mai_mai_n81_));
  NA2        m059(.A(x11), .B(x00), .Y(mai_mai_n82_));
  NO2        m060(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n83_));
  NOi21      m061(.An(mai_mai_n82_), .B(mai_mai_n83_), .Y(mai_mai_n84_));
  AOI210     m062(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n84_), .Y(mai_mai_n85_));
  NOi21      m063(.An(x01), .B(x10), .Y(mai_mai_n86_));
  NO2        m064(.A(mai_mai_n29_), .B(mai_mai_n56_), .Y(mai_mai_n87_));
  NO3        m065(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(x06), .Y(mai_mai_n88_));
  NA2        m066(.A(mai_mai_n88_), .B(mai_mai_n27_), .Y(mai_mai_n89_));
  OAI210     m067(.A0(mai_mai_n85_), .A1(x07), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n90_), .B(mai_mai_n68_), .Y(mai01));
  INV        m069(.A(x12), .Y(mai_mai_n92_));
  INV        m070(.A(x13), .Y(mai_mai_n93_));
  NA2        m071(.A(x08), .B(mai_mai_n81_), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n86_), .B(mai_mai_n28_), .Y(mai_mai_n95_));
  NO2        m073(.A(x10), .B(x01), .Y(mai_mai_n96_));
  NO2        m074(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n97_));
  AOI210     m075(.A0(mai_mai_n95_), .A1(mai_mai_n94_), .B0(mai_mai_n93_), .Y(mai_mai_n98_));
  NO2        m076(.A(mai_mai_n55_), .B(x05), .Y(mai_mai_n99_));
  NOi21      m077(.An(mai_mai_n99_), .B(mai_mai_n57_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n77_), .B(x13), .Y(mai_mai_n102_));
  NA2        m080(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NA2        m082(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n105_), .B(x05), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(mai_mai_n104_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n35_), .B(mai_mai_n56_), .Y(mai_mai_n108_));
  AOI210     m086(.A0(mai_mai_n56_), .A1(mai_mai_n74_), .B0(mai_mai_n100_), .Y(mai_mai_n109_));
  AOI210     m087(.A0(mai_mai_n109_), .A1(mai_mai_n107_), .B0(mai_mai_n70_), .Y(mai_mai_n110_));
  NA2        m088(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n111_));
  NA2        m089(.A(x10), .B(mai_mai_n56_), .Y(mai_mai_n112_));
  NA2        m090(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n59_), .B(x05), .Y(mai_mai_n115_));
  NO3        m093(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n116_));
  NO3        m094(.A(mai_mai_n116_), .B(mai_mai_n110_), .C(mai_mai_n98_), .Y(mai_mai_n117_));
  OAI210     m095(.A0(mai_mai_n77_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n120_));
  NO2        m098(.A(x09), .B(x05), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(mai_mai_n47_), .Y(mai_mai_n122_));
  AOI210     m100(.A0(mai_mai_n122_), .A1(x01), .B0(x02), .Y(mai_mai_n123_));
  NA2        m101(.A(x09), .B(x00), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n99_), .B(mai_mai_n124_), .Y(mai_mai_n125_));
  AOI210     m103(.A0(x09), .A1(mai_mai_n125_), .B0(mai_mai_n120_), .Y(mai_mai_n126_));
  NO2        m104(.A(mai_mai_n126_), .B(mai_mai_n123_), .Y(mai_mai_n127_));
  NO2        m105(.A(x03), .B(x02), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n78_), .B(mai_mai_n93_), .Y(mai_mai_n129_));
  OR2        m107(.A(mai_mai_n127_), .B(x11), .Y(mai_mai_n130_));
  OAI210     m108(.A0(mai_mai_n117_), .A1(mai_mai_n23_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NAi21      m109(.An(x06), .B(x10), .Y(mai_mai_n132_));
  NOi21      m110(.An(x01), .B(x13), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NO2        m112(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n135_));
  NA2        m113(.A(mai_mai_n93_), .B(x01), .Y(mai_mai_n136_));
  NO2        m114(.A(mai_mai_n136_), .B(x08), .Y(mai_mai_n137_));
  AOI210     m115(.A0(x09), .A1(mai_mai_n135_), .B0(mai_mai_n48_), .Y(mai_mai_n138_));
  NO2        m116(.A(x11), .B(mai_mai_n28_), .Y(mai_mai_n139_));
  OAI210     m117(.A0(mai_mai_n138_), .A1(mai_mai_n133_), .B0(mai_mai_n139_), .Y(mai_mai_n140_));
  NA2        m118(.A(x04), .B(x02), .Y(mai_mai_n141_));
  NA2        m119(.A(x10), .B(x05), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n96_), .B(mai_mai_n31_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(x00), .Y(mai_mai_n144_));
  OAI210     m122(.A0(mai_mai_n361_), .A1(x11), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NAi21      m123(.An(mai_mai_n141_), .B(mai_mai_n145_), .Y(mai_mai_n146_));
  INV        m124(.A(mai_mai_n25_), .Y(mai_mai_n147_));
  NAi21      m125(.An(x13), .B(x00), .Y(mai_mai_n148_));
  AOI210     m126(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n148_), .Y(mai_mai_n149_));
  AOI220     m127(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n35_), .B(mai_mai_n150_), .Y(mai_mai_n151_));
  NO2        m129(.A(mai_mai_n87_), .B(x06), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n152_), .B(mai_mai_n362_), .Y(mai_mai_n154_));
  OAI210     m132(.A0(mai_mai_n154_), .A1(x06), .B0(mai_mai_n147_), .Y(mai_mai_n155_));
  NOi21      m133(.An(x09), .B(x00), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n156_), .B(mai_mai_n47_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n93_), .B(x12), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n159_));
  NO2        m137(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n159_), .B(x12), .Y(mai_mai_n161_));
  NA4        m139(.A(mai_mai_n161_), .B(mai_mai_n155_), .C(mai_mai_n146_), .D(mai_mai_n140_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n131_), .A1(mai_mai_n92_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  NA2        m141(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n164_));
  NA2        m142(.A(mai_mai_n164_), .B(mai_mai_n118_), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n111_), .B(x06), .Y(mai_mai_n166_));
  AOI210     m144(.A0(mai_mai_n363_), .A1(mai_mai_n165_), .B0(mai_mai_n166_), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n167_), .B(x12), .Y(mai_mai_n168_));
  INV        m146(.A(mai_mai_n72_), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n134_), .B(mai_mai_n56_), .Y(mai_mai_n170_));
  NA2        m148(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(x09), .A1(mai_mai_n171_), .B0(mai_mai_n23_), .Y(mai_mai_n173_));
  OAI210     m151(.A0(mai_mai_n168_), .A1(mai_mai_n56_), .B0(mai_mai_n173_), .Y(mai_mai_n174_));
  INV        m152(.A(mai_mai_n120_), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n176_));
  OAI210     m154(.A0(mai_mai_n73_), .A1(mai_mai_n36_), .B0(mai_mai_n103_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n93_), .B(x03), .Y(mai_mai_n178_));
  AOI220     m156(.A0(mai_mai_n178_), .A1(mai_mai_n177_), .B0(mai_mai_n72_), .B1(mai_mai_n176_), .Y(mai_mai_n179_));
  NA2        m157(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n180_));
  INV        m158(.A(mai_mai_n132_), .Y(mai_mai_n181_));
  NOi21      m159(.An(x13), .B(x04), .Y(mai_mai_n182_));
  NO3        m160(.A(mai_mai_n182_), .B(mai_mai_n72_), .C(mai_mai_n156_), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n183_), .B(x05), .Y(mai_mai_n184_));
  AOI220     m162(.A0(mai_mai_n184_), .A1(mai_mai_n180_), .B0(mai_mai_n181_), .B1(mai_mai_n56_), .Y(mai_mai_n185_));
  OAI210     m163(.A0(mai_mai_n179_), .A1(mai_mai_n175_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n83_), .Y(mai_mai_n187_));
  NO2        m165(.A(mai_mai_n187_), .B(x12), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n190_));
  OAI210     m168(.A0(mai_mai_n190_), .A1(mai_mai_n151_), .B0(mai_mai_n149_), .Y(mai_mai_n191_));
  AOI210     m169(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n193_), .B(x03), .Y(mai_mai_n194_));
  OA210      m172(.A0(mai_mai_n194_), .A1(mai_mai_n124_), .B0(mai_mai_n191_), .Y(mai_mai_n195_));
  NA2        m173(.A(x13), .B(mai_mai_n92_), .Y(mai_mai_n196_));
  NA3        m174(.A(mai_mai_n196_), .B(x12), .C(mai_mai_n84_), .Y(mai_mai_n197_));
  OAI210     m175(.A0(mai_mai_n195_), .A1(mai_mai_n189_), .B0(mai_mai_n197_), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n188_), .A1(mai_mai_n186_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  AOI210     m177(.A0(mai_mai_n199_), .A1(mai_mai_n174_), .B0(x07), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n69_), .B(mai_mai_n29_), .Y(mai_mai_n201_));
  INV        m179(.A(mai_mai_n201_), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n203_));
  NO2        m181(.A(x08), .B(x05), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(mai_mai_n192_), .Y(mai_mai_n205_));
  OAI210     m183(.A0(mai_mai_n205_), .A1(x06), .B0(x03), .Y(mai_mai_n206_));
  NO2        m184(.A(x12), .B(x02), .Y(mai_mai_n207_));
  INV        m185(.A(mai_mai_n207_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n208_), .B(mai_mai_n187_), .Y(mai_mai_n209_));
  OA210      m187(.A0(mai_mai_n206_), .A1(mai_mai_n202_), .B0(mai_mai_n209_), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n211_), .B(x01), .Y(mai_mai_n212_));
  NOi21      m190(.An(mai_mai_n77_), .B(mai_mai_n103_), .Y(mai_mai_n213_));
  NA2        m191(.A(mai_mai_n203_), .B(mai_mai_n177_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n93_), .B(x04), .Y(mai_mai_n215_));
  NA2        m193(.A(mai_mai_n215_), .B(mai_mai_n28_), .Y(mai_mai_n216_));
  OAI210     m194(.A0(mai_mai_n216_), .A1(mai_mai_n102_), .B0(mai_mai_n214_), .Y(mai_mai_n217_));
  NO3        m195(.A(mai_mai_n82_), .B(x12), .C(x03), .Y(mai_mai_n218_));
  OAI210     m196(.A0(mai_mai_n217_), .A1(mai_mai_n213_), .B0(mai_mai_n218_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n220_));
  OAI210     m198(.A0(x06), .A1(mai_mai_n86_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n172_), .B(mai_mai_n152_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n189_), .B(mai_mai_n28_), .Y(mai_mai_n223_));
  OAI210     m201(.A0(mai_mai_n222_), .A1(mai_mai_n175_), .B0(mai_mai_n223_), .Y(mai_mai_n224_));
  NA3        m202(.A(mai_mai_n224_), .B(mai_mai_n221_), .C(mai_mai_n219_), .Y(mai_mai_n225_));
  NO3        m203(.A(mai_mai_n225_), .B(mai_mai_n210_), .C(mai_mai_n200_), .Y(mai_mai_n226_));
  OAI210     m204(.A0(mai_mai_n163_), .A1(mai_mai_n60_), .B0(mai_mai_n226_), .Y(mai02));
  BUFFER     m205(.A(mai_mai_n183_), .Y(mai_mai_n228_));
  NA3        m206(.A(x13), .B(x10), .C(mai_mai_n55_), .Y(mai_mai_n229_));
  OAI210     m207(.A0(mai_mai_n228_), .A1(mai_mai_n32_), .B0(mai_mai_n229_), .Y(mai_mai_n230_));
  NA2        m208(.A(mai_mai_n230_), .B(mai_mai_n142_), .Y(mai_mai_n231_));
  INV        m209(.A(mai_mai_n142_), .Y(mai_mai_n232_));
  AOI210     m210(.A0(mai_mai_n101_), .A1(mai_mai_n79_), .B0(mai_mai_n172_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n233_), .B(mai_mai_n93_), .Y(mai_mai_n234_));
  AOI220     m212(.A0(mai_mai_n234_), .A1(mai_mai_n232_), .B0(mai_mai_n129_), .B1(mai_mai_n128_), .Y(mai_mai_n235_));
  AOI210     m213(.A0(mai_mai_n235_), .A1(mai_mai_n231_), .B0(mai_mai_n48_), .Y(mai_mai_n236_));
  AOI220     m214(.A0(mai_mai_n204_), .A1(mai_mai_n57_), .B0(mai_mai_n55_), .B1(mai_mai_n36_), .Y(mai_mai_n237_));
  NOi21      m215(.An(x13), .B(mai_mai_n237_), .Y(mai_mai_n238_));
  AOI210     m216(.A0(mai_mai_n182_), .A1(mai_mai_n73_), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n239_), .B(mai_mai_n120_), .Y(mai_mai_n240_));
  INV        m218(.A(mai_mai_n179_), .Y(mai_mai_n241_));
  NO2        m219(.A(mai_mai_n193_), .B(mai_mai_n47_), .Y(mai_mai_n242_));
  NA2        m220(.A(mai_mai_n242_), .B(mai_mai_n241_), .Y(mai_mai_n243_));
  AN2        m221(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n244_));
  OAI210     m222(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n245_));
  AOI210     m223(.A0(x02), .A1(mai_mai_n118_), .B0(mai_mai_n245_), .Y(mai_mai_n246_));
  OAI210     m224(.A0(mai_mai_n246_), .A1(mai_mai_n244_), .B0(mai_mai_n87_), .Y(mai_mai_n247_));
  NA3        m225(.A(mai_mai_n87_), .B(mai_mai_n77_), .C(mai_mai_n176_), .Y(mai_mai_n248_));
  NA3        m226(.A(mai_mai_n86_), .B(mai_mai_n76_), .C(mai_mai_n42_), .Y(mai_mai_n249_));
  AOI210     m227(.A0(mai_mai_n249_), .A1(mai_mai_n248_), .B0(x04), .Y(mai_mai_n250_));
  INV        m228(.A(mai_mai_n128_), .Y(mai_mai_n251_));
  OAI220     m229(.A0(mai_mai_n205_), .A1(mai_mai_n95_), .B0(mai_mai_n251_), .B1(mai_mai_n113_), .Y(mai_mai_n252_));
  AOI210     m230(.A0(mai_mai_n252_), .A1(x13), .B0(mai_mai_n250_), .Y(mai_mai_n253_));
  NA3        m231(.A(mai_mai_n253_), .B(mai_mai_n247_), .C(mai_mai_n243_), .Y(mai_mai_n254_));
  NO3        m232(.A(mai_mai_n254_), .B(mai_mai_n240_), .C(mai_mai_n236_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n119_), .B(x03), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n148_), .B(mai_mai_n256_), .Y(mai_mai_n257_));
  NA2        m235(.A(mai_mai_n257_), .B(mai_mai_n96_), .Y(mai_mai_n258_));
  OAI220     m236(.A0(mai_mai_n215_), .A1(x09), .B0(mai_mai_n114_), .B1(mai_mai_n28_), .Y(mai_mai_n259_));
  NA2        m237(.A(mai_mai_n259_), .B(mai_mai_n97_), .Y(mai_mai_n260_));
  NA2        m238(.A(mai_mai_n215_), .B(mai_mai_n92_), .Y(mai_mai_n261_));
  NA2        m239(.A(mai_mai_n261_), .B(mai_mai_n113_), .Y(mai_mai_n262_));
  NA4        m240(.A(mai_mai_n262_), .B(mai_mai_n260_), .C(mai_mai_n258_), .D(mai_mai_n48_), .Y(mai_mai_n263_));
  INV        m241(.A(mai_mai_n160_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n137_), .B(mai_mai_n40_), .Y(mai_mai_n265_));
  NA2        m243(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n266_));
  OAI220     m244(.A0(mai_mai_n266_), .A1(mai_mai_n265_), .B0(mai_mai_n264_), .B1(mai_mai_n58_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n267_), .B(x02), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n190_), .Y(mai_mai_n269_));
  NA2        m247(.A(mai_mai_n158_), .B(x04), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n270_), .B(mai_mai_n269_), .Y(mai_mai_n271_));
  NO2        m249(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n272_));
  OAI210     m250(.A0(mai_mai_n272_), .A1(mai_mai_n271_), .B0(mai_mai_n87_), .Y(mai_mai_n273_));
  NO3        m251(.A(mai_mai_n158_), .B(mai_mai_n135_), .C(mai_mai_n51_), .Y(mai_mai_n274_));
  OAI210     m252(.A0(mai_mai_n124_), .A1(mai_mai_n36_), .B0(mai_mai_n92_), .Y(mai_mai_n275_));
  OAI210     m253(.A0(mai_mai_n275_), .A1(mai_mai_n157_), .B0(mai_mai_n274_), .Y(mai_mai_n276_));
  NA4        m254(.A(mai_mai_n276_), .B(mai_mai_n273_), .C(mai_mai_n268_), .D(x06), .Y(mai_mai_n277_));
  NA2        m255(.A(x09), .B(x03), .Y(mai_mai_n278_));
  OAI220     m256(.A0(mai_mai_n278_), .A1(mai_mai_n112_), .B0(mai_mai_n164_), .B1(mai_mai_n63_), .Y(mai_mai_n279_));
  NO2        m257(.A(x08), .B(mai_mai_n41_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n280_), .B(mai_mai_n175_), .Y(mai_mai_n281_));
  NO2        m259(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n282_));
  NA2        m260(.A(mai_mai_n274_), .B(mai_mai_n282_), .Y(mai_mai_n283_));
  OAI210     m261(.A0(mai_mai_n281_), .A1(mai_mai_n28_), .B0(mai_mai_n283_), .Y(mai_mai_n284_));
  AO220      m262(.A0(mai_mai_n284_), .A1(x04), .B0(mai_mai_n279_), .B1(x05), .Y(mai_mai_n285_));
  AOI210     m263(.A0(mai_mai_n277_), .A1(mai_mai_n263_), .B0(mai_mai_n285_), .Y(mai_mai_n286_));
  OAI210     m264(.A0(mai_mai_n255_), .A1(x12), .B0(mai_mai_n286_), .Y(mai03));
  OR2        m265(.A(mai_mai_n42_), .B(mai_mai_n176_), .Y(mai_mai_n288_));
  AOI210     m266(.A0(mai_mai_n129_), .A1(mai_mai_n92_), .B0(mai_mai_n288_), .Y(mai_mai_n289_));
  AO210      m267(.A0(mai_mai_n269_), .A1(mai_mai_n79_), .B0(mai_mai_n270_), .Y(mai_mai_n290_));
  INV        m268(.A(mai_mai_n290_), .Y(mai_mai_n291_));
  OAI210     m269(.A0(mai_mai_n291_), .A1(mai_mai_n289_), .B0(x05), .Y(mai_mai_n292_));
  NA2        m270(.A(mai_mai_n288_), .B(x05), .Y(mai_mai_n293_));
  AOI210     m271(.A0(mai_mai_n118_), .A1(mai_mai_n169_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  AOI210     m272(.A0(mai_mai_n178_), .A1(mai_mai_n74_), .B0(mai_mai_n106_), .Y(mai_mai_n295_));
  OAI220     m273(.A0(mai_mai_n295_), .A1(mai_mai_n58_), .B0(x02), .B1(mai_mai_n237_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n296_), .A1(mai_mai_n294_), .B0(mai_mai_n92_), .Y(mai_mai_n297_));
  NO2        m275(.A(mai_mai_n92_), .B(mai_mai_n122_), .Y(mai_mai_n298_));
  OA210      m276(.A0(mai_mai_n137_), .A1(x12), .B0(mai_mai_n115_), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n300_));
  NA3        m278(.A(mai_mai_n300_), .B(mai_mai_n297_), .C(mai_mai_n292_), .Y(mai04));
  NO2        m279(.A(mai_mai_n80_), .B(mai_mai_n39_), .Y(mai_mai_n302_));
  XO2        m280(.A(mai_mai_n302_), .B(mai_mai_n196_), .Y(mai05));
  INV        m281(.A(mai_mai_n166_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n304_), .B(mai_mai_n25_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n120_), .B(mai_mai_n114_), .C(mai_mai_n31_), .Y(mai_mai_n306_));
  NO2        m284(.A(mai_mai_n306_), .B(mai_mai_n24_), .Y(mai_mai_n307_));
  OAI210     m285(.A0(mai_mai_n307_), .A1(mai_mai_n305_), .B0(mai_mai_n92_), .Y(mai_mai_n308_));
  NA2        m286(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n201_), .B(x03), .Y(mai_mai_n311_));
  OAI220     m289(.A0(mai_mai_n311_), .A1(mai_mai_n310_), .B0(mai_mai_n309_), .B1(mai_mai_n75_), .Y(mai_mai_n312_));
  AOI210     m290(.A0(mai_mai_n312_), .A1(x06), .B0(mai_mai_n365_), .Y(mai_mai_n313_));
  AOI220     m291(.A0(mai_mai_n75_), .A1(mai_mai_n31_), .B0(mai_mai_n51_), .B1(mai_mai_n50_), .Y(mai_mai_n314_));
  NO3        m292(.A(mai_mai_n314_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n315_));
  NO2        m293(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n316_));
  OAI210     m294(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n317_));
  OR3        m295(.A(mai_mai_n317_), .B(mai_mai_n316_), .C(mai_mai_n44_), .Y(mai_mai_n318_));
  INV        m296(.A(mai_mai_n318_), .Y(mai_mai_n319_));
  OAI210     m297(.A0(mai_mai_n319_), .A1(mai_mai_n315_), .B0(mai_mai_n92_), .Y(mai_mai_n320_));
  AOI220     m298(.A0(mai_mai_n364_), .A1(mai_mai_n320_), .B0(mai_mai_n313_), .B1(mai_mai_n308_), .Y(mai_mai_n321_));
  AOI210     m299(.A0(mai_mai_n316_), .A1(mai_mai_n71_), .B0(mai_mai_n119_), .Y(mai_mai_n322_));
  OR2        m300(.A(mai_mai_n322_), .B(x03), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n282_), .B(mai_mai_n60_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n324_), .B(x11), .Y(mai_mai_n325_));
  NO3        m303(.A(mai_mai_n325_), .B(mai_mai_n121_), .C(mai_mai_n28_), .Y(mai_mai_n326_));
  AOI210     m304(.A0(mai_mai_n326_), .A1(mai_mai_n323_), .B0(mai_mai_n47_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n327_), .B(mai_mai_n93_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n270_), .B(mai_mai_n207_), .Y(mai_mai_n329_));
  NOi21      m307(.An(mai_mai_n256_), .B(mai_mai_n115_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n330_), .B(mai_mai_n208_), .Y(mai_mai_n331_));
  OAI210     m309(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n196_), .A1(mai_mai_n47_), .B0(mai_mai_n332_), .Y(mai_mai_n333_));
  NO4        m311(.A(mai_mai_n333_), .B(mai_mai_n331_), .C(mai_mai_n329_), .D(x08), .Y(mai_mai_n334_));
  NO2        m312(.A(mai_mai_n114_), .B(mai_mai_n28_), .Y(mai_mai_n335_));
  NO2        m313(.A(mai_mai_n335_), .B(mai_mai_n212_), .Y(mai_mai_n336_));
  OR3        m314(.A(mai_mai_n336_), .B(x12), .C(x03), .Y(mai_mai_n337_));
  NA3        m315(.A(mai_mai_n264_), .B(mai_mai_n108_), .C(x12), .Y(mai_mai_n338_));
  AO210      m316(.A0(mai_mai_n264_), .A1(mai_mai_n108_), .B0(mai_mai_n196_), .Y(mai_mai_n339_));
  NA4        m317(.A(mai_mai_n339_), .B(mai_mai_n338_), .C(mai_mai_n337_), .D(x08), .Y(mai_mai_n340_));
  INV        m318(.A(mai_mai_n340_), .Y(mai_mai_n341_));
  AOI210     m319(.A0(mai_mai_n334_), .A1(mai_mai_n328_), .B0(mai_mai_n341_), .Y(mai_mai_n342_));
  OAI210     m320(.A0(mai_mai_n324_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n232_), .B(x07), .Y(mai_mai_n344_));
  OAI220     m322(.A0(mai_mai_n344_), .A1(mai_mai_n310_), .B0(mai_mai_n121_), .B1(mai_mai_n43_), .Y(mai_mai_n345_));
  OAI210     m323(.A0(mai_mai_n345_), .A1(mai_mai_n343_), .B0(mai_mai_n153_), .Y(mai_mai_n346_));
  NA3        m324(.A(mai_mai_n336_), .B(mai_mai_n330_), .C(mai_mai_n261_), .Y(mai_mai_n347_));
  INV        m325(.A(x14), .Y(mai_mai_n348_));
  NO3        m326(.A(mai_mai_n256_), .B(mai_mai_n95_), .C(x11), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n349_), .B(mai_mai_n348_), .Y(mai_mai_n350_));
  NA3        m328(.A(mai_mai_n350_), .B(mai_mai_n347_), .C(mai_mai_n346_), .Y(mai_mai_n351_));
  AOI220     m329(.A0(x12), .A1(mai_mai_n60_), .B0(mai_mai_n335_), .B1(mai_mai_n135_), .Y(mai_mai_n352_));
  NOi21      m330(.An(mai_mai_n215_), .B(mai_mai_n125_), .Y(mai_mai_n353_));
  NA2        m331(.A(mai_mai_n220_), .B(mai_mai_n181_), .Y(mai_mai_n354_));
  OAI210     m332(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  OAI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n353_), .B0(mai_mai_n92_), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n352_), .A1(mai_mai_n82_), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  NO4        m335(.A(mai_mai_n357_), .B(mai_mai_n351_), .C(mai_mai_n342_), .D(mai_mai_n321_), .Y(mai06));
  INV        m336(.A(x01), .Y(mai_mai_n361_));
  INV        m337(.A(x05), .Y(mai_mai_n362_));
  INV        m338(.A(x05), .Y(mai_mai_n363_));
  INV        m339(.A(x07), .Y(mai_mai_n364_));
  INV        m340(.A(x07), .Y(mai_mai_n365_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NO2        u030(.A(x09), .B(x07), .Y(men_men_n53_));
  OAI210     u031(.A0(men_men_n53_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n54_));
  NOi21      u032(.An(x01), .B(x09), .Y(men_men_n55_));
  INV        u033(.A(x00), .Y(men_men_n56_));
  NO2        u034(.A(men_men_n51_), .B(men_men_n56_), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n57_), .B(men_men_n55_), .Y(men_men_n58_));
  NA2        u036(.A(x09), .B(men_men_n56_), .Y(men_men_n59_));
  INV        u037(.A(x07), .Y(men_men_n60_));
  INV        u038(.A(men_men_n58_), .Y(men_men_n61_));
  OAI220     u039(.A0(men_men_n23_), .A1(men_men_n61_), .B0(x07), .B1(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n62_), .B(men_men_n31_), .Y(men_men_n63_));
  AOI210     u041(.A0(men_men_n63_), .A1(men_men_n54_), .B0(x05), .Y(men_men_n64_));
  NA2        u042(.A(x10), .B(x09), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n60_), .B(men_men_n23_), .Y(men_men_n66_));
  NA2        u044(.A(x09), .B(x05), .Y(men_men_n67_));
  NA2        u045(.A(x10), .B(x06), .Y(men_men_n68_));
  NA3        u046(.A(men_men_n68_), .B(men_men_n67_), .C(men_men_n28_), .Y(men_men_n69_));
  NO2        u047(.A(men_men_n60_), .B(men_men_n41_), .Y(men_men_n70_));
  OAI210     u048(.A0(men_men_n69_), .A1(men_men_n66_), .B0(x03), .Y(men_men_n71_));
  NOi31      u049(.An(x08), .B(x04), .C(x00), .Y(men_men_n72_));
  NO2        u050(.A(x10), .B(x09), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n402_), .B(men_men_n24_), .Y(men_men_n74_));
  NO2        u052(.A(x09), .B(men_men_n41_), .Y(men_men_n75_));
  OAI210     u053(.A0(men_men_n75_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n76_));
  NO2        u054(.A(men_men_n36_), .B(x00), .Y(men_men_n77_));
  NO2        u055(.A(x08), .B(x01), .Y(men_men_n78_));
  OAI210     u056(.A0(men_men_n78_), .A1(men_men_n77_), .B0(men_men_n35_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n79_), .B(men_men_n74_), .Y(men_men_n80_));
  AN2        u058(.A(men_men_n80_), .B(men_men_n71_), .Y(men_men_n81_));
  INV        u059(.A(men_men_n79_), .Y(men_men_n82_));
  NO2        u060(.A(x06), .B(x05), .Y(men_men_n83_));
  NA2        u061(.A(x11), .B(x00), .Y(men_men_n84_));
  NO2        u062(.A(x11), .B(men_men_n47_), .Y(men_men_n85_));
  NOi21      u063(.An(men_men_n84_), .B(men_men_n85_), .Y(men_men_n86_));
  AOI210     u064(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n86_), .Y(men_men_n87_));
  NOi21      u065(.An(x01), .B(x10), .Y(men_men_n88_));
  NO2        u066(.A(men_men_n29_), .B(men_men_n56_), .Y(men_men_n89_));
  NO3        u067(.A(men_men_n89_), .B(men_men_n88_), .C(x06), .Y(men_men_n90_));
  NA2        u068(.A(men_men_n90_), .B(men_men_n27_), .Y(men_men_n91_));
  OAI210     u069(.A0(men_men_n87_), .A1(x07), .B0(men_men_n91_), .Y(men_men_n92_));
  NO3        u070(.A(men_men_n92_), .B(men_men_n81_), .C(men_men_n64_), .Y(men01));
  INV        u071(.A(x12), .Y(men_men_n94_));
  INV        u072(.A(x13), .Y(men_men_n95_));
  NA2        u073(.A(men_men_n403_), .B(men_men_n65_), .Y(men_men_n96_));
  NA2        u074(.A(x08), .B(x04), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n97_), .B(men_men_n56_), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n98_), .B(men_men_n96_), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n88_), .B(men_men_n28_), .Y(men_men_n100_));
  NO2        u078(.A(x10), .B(x01), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n29_), .B(x00), .Y(men_men_n102_));
  INV        u080(.A(men_men_n102_), .Y(men_men_n103_));
  NA2        u081(.A(x04), .B(men_men_n28_), .Y(men_men_n104_));
  NO3        u082(.A(men_men_n104_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n105_));
  INV        u083(.A(men_men_n105_), .Y(men_men_n106_));
  AOI210     u084(.A0(men_men_n106_), .A1(men_men_n99_), .B0(men_men_n95_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n55_), .B(x05), .Y(men_men_n108_));
  NOi21      u086(.An(men_men_n108_), .B(men_men_n57_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n95_), .B(men_men_n36_), .Y(men_men_n110_));
  NA3        u088(.A(men_men_n110_), .B(x04), .C(x06), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n111_), .B(men_men_n109_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n78_), .B(x13), .Y(men_men_n113_));
  NA2        u091(.A(men_men_n35_), .B(men_men_n56_), .Y(men_men_n114_));
  AOI210     u092(.A0(men_men_n114_), .A1(men_men_n113_), .B0(men_men_n68_), .Y(men_men_n115_));
  NA2        u093(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n116_));
  NA2        u094(.A(x10), .B(men_men_n56_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n51_), .B(x05), .Y(men_men_n119_));
  NA3        u097(.A(men_men_n407_), .B(men_men_n119_), .C(x13), .Y(men_men_n120_));
  NO3        u098(.A(men_men_n114_), .B(men_men_n75_), .C(men_men_n36_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n59_), .B(x05), .Y(men_men_n122_));
  NOi41      u100(.An(men_men_n120_), .B(men_men_n122_), .C(men_men_n121_), .D(men_men_n118_), .Y(men_men_n123_));
  NO3        u101(.A(men_men_n123_), .B(x06), .C(x03), .Y(men_men_n124_));
  NO4        u102(.A(men_men_n124_), .B(men_men_n115_), .C(men_men_n112_), .D(men_men_n107_), .Y(men_men_n125_));
  NA2        u103(.A(x13), .B(men_men_n36_), .Y(men_men_n126_));
  OAI210     u104(.A0(men_men_n78_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO2        u106(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n129_));
  OA210      u107(.A0(x00), .A1(men_men_n73_), .B0(men_men_n129_), .Y(men_men_n130_));
  NO2        u108(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n29_), .B(x06), .Y(men_men_n132_));
  AOI210     u110(.A0(men_men_n132_), .A1(men_men_n49_), .B0(men_men_n131_), .Y(men_men_n133_));
  OA210      u111(.A0(men_men_n133_), .A1(men_men_n130_), .B0(men_men_n128_), .Y(men_men_n134_));
  NO2        u112(.A(x09), .B(x05), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(men_men_n47_), .Y(men_men_n136_));
  AOI210     u114(.A0(men_men_n136_), .A1(men_men_n103_), .B0(men_men_n49_), .Y(men_men_n137_));
  NA2        u115(.A(x09), .B(x00), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n108_), .B(men_men_n138_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n72_), .B(men_men_n51_), .Y(men_men_n140_));
  AOI210     u118(.A0(men_men_n140_), .A1(men_men_n139_), .B0(men_men_n132_), .Y(men_men_n141_));
  NO3        u119(.A(men_men_n141_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n142_));
  NO2        u120(.A(x03), .B(x02), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n79_), .B(men_men_n95_), .Y(men_men_n144_));
  OAI210     u122(.A0(men_men_n144_), .A1(men_men_n109_), .B0(men_men_n143_), .Y(men_men_n145_));
  OA210      u123(.A0(men_men_n142_), .A1(x11), .B0(men_men_n145_), .Y(men_men_n146_));
  OAI210     u124(.A0(men_men_n125_), .A1(men_men_n23_), .B0(men_men_n146_), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n103_), .B(men_men_n40_), .Y(men_men_n148_));
  NAi21      u126(.An(x06), .B(x10), .Y(men_men_n149_));
  NOi21      u127(.An(x01), .B(x13), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n150_), .B(men_men_n149_), .Y(men_men_n151_));
  OR2        u129(.A(men_men_n151_), .B(x08), .Y(men_men_n152_));
  AOI210     u130(.A0(men_men_n152_), .A1(men_men_n148_), .B0(men_men_n41_), .Y(men_men_n153_));
  NO2        u131(.A(men_men_n29_), .B(x03), .Y(men_men_n154_));
  NA2        u132(.A(men_men_n95_), .B(x01), .Y(men_men_n155_));
  NO2        u133(.A(men_men_n155_), .B(x08), .Y(men_men_n156_));
  OAI210     u134(.A0(x05), .A1(men_men_n156_), .B0(men_men_n51_), .Y(men_men_n157_));
  AOI210     u135(.A0(men_men_n157_), .A1(men_men_n154_), .B0(men_men_n48_), .Y(men_men_n158_));
  AOI210     u136(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n159_));
  OAI210     u137(.A0(men_men_n158_), .A1(men_men_n153_), .B0(men_men_n159_), .Y(men_men_n160_));
  NA2        u138(.A(x04), .B(x02), .Y(men_men_n161_));
  NA2        u139(.A(x10), .B(x05), .Y(men_men_n162_));
  NO2        u140(.A(x09), .B(x01), .Y(men_men_n163_));
  NO3        u141(.A(men_men_n163_), .B(men_men_n101_), .C(men_men_n31_), .Y(men_men_n164_));
  NA2        u142(.A(men_men_n164_), .B(x00), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n108_), .B(x08), .Y(men_men_n166_));
  NA3        u144(.A(men_men_n150_), .B(men_men_n149_), .C(men_men_n51_), .Y(men_men_n167_));
  NA2        u145(.A(men_men_n88_), .B(x05), .Y(men_men_n168_));
  OAI210     u146(.A0(men_men_n168_), .A1(men_men_n110_), .B0(men_men_n167_), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n166_), .A1(x06), .B0(men_men_n169_), .Y(men_men_n170_));
  OAI210     u148(.A0(men_men_n170_), .A1(x11), .B0(men_men_n165_), .Y(men_men_n171_));
  NAi21      u149(.An(men_men_n161_), .B(men_men_n171_), .Y(men_men_n172_));
  INV        u150(.A(men_men_n25_), .Y(men_men_n173_));
  NAi21      u151(.An(x13), .B(x00), .Y(men_men_n174_));
  AOI210     u152(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n174_), .Y(men_men_n175_));
  AOI220     u153(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n176_));
  OAI210     u154(.A0(men_men_n162_), .A1(men_men_n35_), .B0(men_men_n176_), .Y(men_men_n177_));
  AN2        u155(.A(men_men_n177_), .B(men_men_n175_), .Y(men_men_n178_));
  NO2        u156(.A(men_men_n174_), .B(men_men_n36_), .Y(men_men_n179_));
  INV        u157(.A(men_men_n179_), .Y(men_men_n180_));
  NO2        u158(.A(men_men_n56_), .B(men_men_n67_), .Y(men_men_n181_));
  OAI210     u159(.A0(men_men_n181_), .A1(men_men_n178_), .B0(men_men_n173_), .Y(men_men_n182_));
  NOi21      u160(.An(x09), .B(x00), .Y(men_men_n183_));
  NO3        u161(.A(men_men_n77_), .B(men_men_n183_), .C(men_men_n47_), .Y(men_men_n184_));
  NA2        u162(.A(men_men_n184_), .B(men_men_n117_), .Y(men_men_n185_));
  NA2        u163(.A(x06), .B(x05), .Y(men_men_n186_));
  OAI210     u164(.A0(men_men_n186_), .A1(men_men_n35_), .B0(men_men_n94_), .Y(men_men_n187_));
  AOI210     u165(.A0(x08), .A1(men_men_n57_), .B0(men_men_n187_), .Y(men_men_n188_));
  NA2        u166(.A(men_men_n188_), .B(men_men_n185_), .Y(men_men_n189_));
  NO2        u167(.A(men_men_n95_), .B(x12), .Y(men_men_n190_));
  AOI210     u168(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n190_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n88_), .B(men_men_n51_), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n193_));
  NA2        u171(.A(men_men_n193_), .B(x02), .Y(men_men_n194_));
  NO2        u172(.A(men_men_n194_), .B(men_men_n192_), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n191_), .A1(men_men_n189_), .B0(men_men_n195_), .Y(men_men_n196_));
  NA4        u174(.A(men_men_n196_), .B(men_men_n182_), .C(men_men_n172_), .D(men_men_n160_), .Y(men_men_n197_));
  AOI210     u175(.A0(men_men_n147_), .A1(men_men_n94_), .B0(men_men_n197_), .Y(men_men_n198_));
  NO2        u176(.A(men_men_n116_), .B(x06), .Y(men_men_n199_));
  AOI210     u177(.A0(x06), .A1(men_men_n69_), .B0(x12), .Y(men_men_n200_));
  INV        u178(.A(men_men_n72_), .Y(men_men_n201_));
  NO2        u179(.A(x05), .B(men_men_n51_), .Y(men_men_n202_));
  OAI210     u180(.A0(men_men_n202_), .A1(men_men_n151_), .B0(men_men_n56_), .Y(men_men_n203_));
  NA2        u181(.A(men_men_n203_), .B(men_men_n201_), .Y(men_men_n204_));
  NO2        u182(.A(men_men_n88_), .B(x06), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n205_), .B(men_men_n41_), .Y(men_men_n206_));
  NA4        u184(.A(men_men_n149_), .B(men_men_n55_), .C(men_men_n36_), .D(x04), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(men_men_n132_), .Y(men_men_n208_));
  OAI210     u186(.A0(men_men_n208_), .A1(men_men_n206_), .B0(x02), .Y(men_men_n209_));
  AOI210     u187(.A0(men_men_n209_), .A1(men_men_n204_), .B0(men_men_n23_), .Y(men_men_n210_));
  OAI210     u188(.A0(men_men_n200_), .A1(men_men_n56_), .B0(men_men_n210_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n51_), .B(x03), .Y(men_men_n212_));
  NA2        u190(.A(men_men_n72_), .B(men_men_n212_), .Y(men_men_n213_));
  INV        u191(.A(men_men_n149_), .Y(men_men_n214_));
  NOi21      u192(.An(x13), .B(x04), .Y(men_men_n215_));
  NO3        u193(.A(men_men_n215_), .B(men_men_n72_), .C(men_men_n183_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n216_), .B(x05), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n214_), .B(men_men_n56_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n213_), .B(men_men_n218_), .Y(men_men_n219_));
  INV        u197(.A(men_men_n85_), .Y(men_men_n220_));
  NA2        u198(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n221_));
  NO2        u199(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n222_));
  OAI210     u200(.A0(men_men_n222_), .A1(men_men_n177_), .B0(men_men_n175_), .Y(men_men_n223_));
  AOI210     u201(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n224_));
  NO2        u202(.A(x06), .B(x00), .Y(men_men_n225_));
  NO3        u203(.A(men_men_n225_), .B(men_men_n224_), .C(men_men_n41_), .Y(men_men_n226_));
  OAI210     u204(.A0(men_men_n97_), .A1(men_men_n138_), .B0(men_men_n68_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n229_));
  INV        u207(.A(x03), .Y(men_men_n230_));
  OA210      u208(.A0(men_men_n230_), .A1(men_men_n228_), .B0(men_men_n223_), .Y(men_men_n231_));
  NA2        u209(.A(x13), .B(men_men_n94_), .Y(men_men_n232_));
  NA3        u210(.A(men_men_n232_), .B(men_men_n187_), .C(men_men_n86_), .Y(men_men_n233_));
  OAI210     u211(.A0(men_men_n231_), .A1(men_men_n221_), .B0(men_men_n233_), .Y(men_men_n234_));
  AOI210     u212(.A0(men_men_n85_), .A1(men_men_n219_), .B0(men_men_n234_), .Y(men_men_n235_));
  AOI210     u213(.A0(men_men_n235_), .A1(men_men_n211_), .B0(x07), .Y(men_men_n236_));
  NA2        u214(.A(men_men_n67_), .B(men_men_n29_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n215_), .B(men_men_n183_), .Y(men_men_n238_));
  AOI210     u216(.A0(men_men_n238_), .A1(men_men_n140_), .B0(men_men_n237_), .Y(men_men_n239_));
  NO2        u217(.A(men_men_n95_), .B(x06), .Y(men_men_n240_));
  INV        u218(.A(men_men_n240_), .Y(men_men_n241_));
  NO2        u219(.A(x08), .B(x05), .Y(men_men_n242_));
  NO2        u220(.A(men_men_n242_), .B(men_men_n224_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n72_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n244_));
  OAI210     u222(.A0(men_men_n243_), .A1(men_men_n241_), .B0(men_men_n244_), .Y(men_men_n245_));
  NO2        u223(.A(x12), .B(x02), .Y(men_men_n246_));
  INV        u224(.A(men_men_n246_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n247_), .B(men_men_n220_), .Y(men_men_n248_));
  OA210      u226(.A0(men_men_n245_), .A1(men_men_n239_), .B0(men_men_n248_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n250_), .B(x01), .Y(men_men_n251_));
  NA2        u229(.A(men_men_n95_), .B(x04), .Y(men_men_n252_));
  NO3        u230(.A(men_men_n84_), .B(x12), .C(x03), .Y(men_men_n253_));
  OAI210     u231(.A0(men_men_n406_), .A1(x10), .B0(men_men_n253_), .Y(men_men_n254_));
  AOI210     u232(.A0(men_men_n192_), .A1(men_men_n186_), .B0(men_men_n97_), .Y(men_men_n255_));
  NOi21      u233(.An(men_men_n237_), .B(men_men_n205_), .Y(men_men_n256_));
  NO2        u234(.A(men_men_n25_), .B(x00), .Y(men_men_n257_));
  OAI210     u235(.A0(men_men_n256_), .A1(men_men_n255_), .B0(men_men_n257_), .Y(men_men_n258_));
  NO2        u236(.A(men_men_n57_), .B(x05), .Y(men_men_n259_));
  NA2        u237(.A(men_men_n258_), .B(men_men_n254_), .Y(men_men_n260_));
  NO3        u238(.A(men_men_n260_), .B(men_men_n249_), .C(men_men_n236_), .Y(men_men_n261_));
  OAI210     u239(.A0(men_men_n198_), .A1(men_men_n60_), .B0(men_men_n261_), .Y(men02));
  NA3        u240(.A(x04), .B(x08), .C(men_men_n55_), .Y(men_men_n263_));
  OAI210     u241(.A0(x01), .A1(men_men_n32_), .B0(men_men_n263_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n264_), .B(men_men_n162_), .Y(men_men_n265_));
  INV        u243(.A(men_men_n162_), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n79_), .A1(men_men_n51_), .B0(men_men_n95_), .Y(men_men_n267_));
  NA2        u245(.A(men_men_n267_), .B(men_men_n266_), .Y(men_men_n268_));
  AOI210     u246(.A0(men_men_n268_), .A1(men_men_n265_), .B0(men_men_n48_), .Y(men_men_n269_));
  NO2        u247(.A(x02), .B(men_men_n132_), .Y(men_men_n270_));
  NAi21      u248(.An(men_men_n217_), .B(men_men_n213_), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n229_), .B(men_men_n47_), .Y(men_men_n272_));
  NA2        u250(.A(men_men_n272_), .B(men_men_n271_), .Y(men_men_n273_));
  OAI210     u251(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n274_));
  OA210      u252(.A0(men_men_n409_), .A1(x08), .B0(men_men_n136_), .Y(men_men_n275_));
  NO2        u253(.A(men_men_n275_), .B(men_men_n274_), .Y(men_men_n276_));
  NA2        u254(.A(men_men_n276_), .B(men_men_n89_), .Y(men_men_n277_));
  NA3        u255(.A(men_men_n89_), .B(men_men_n78_), .C(men_men_n212_), .Y(men_men_n278_));
  NA2        u256(.A(men_men_n88_), .B(men_men_n42_), .Y(men_men_n279_));
  AOI210     u257(.A0(men_men_n279_), .A1(men_men_n278_), .B0(x04), .Y(men_men_n280_));
  INV        u258(.A(men_men_n143_), .Y(men_men_n281_));
  OAI220     u259(.A0(men_men_n243_), .A1(men_men_n100_), .B0(men_men_n281_), .B1(men_men_n118_), .Y(men_men_n282_));
  AOI210     u260(.A0(men_men_n282_), .A1(x13), .B0(men_men_n280_), .Y(men_men_n283_));
  NA3        u261(.A(men_men_n283_), .B(men_men_n277_), .C(men_men_n273_), .Y(men_men_n284_));
  NO3        u262(.A(men_men_n284_), .B(men_men_n270_), .C(men_men_n269_), .Y(men_men_n285_));
  NA2        u263(.A(men_men_n131_), .B(x03), .Y(men_men_n286_));
  OAI210     u264(.A0(men_men_n35_), .A1(men_men_n259_), .B0(men_men_n286_), .Y(men_men_n287_));
  NA2        u265(.A(men_men_n287_), .B(men_men_n101_), .Y(men_men_n288_));
  NA2        u266(.A(men_men_n161_), .B(men_men_n155_), .Y(men_men_n289_));
  AN2        u267(.A(men_men_n289_), .B(men_men_n166_), .Y(men_men_n290_));
  INV        u268(.A(men_men_n55_), .Y(men_men_n291_));
  OAI220     u269(.A0(men_men_n252_), .A1(men_men_n291_), .B0(men_men_n119_), .B1(men_men_n28_), .Y(men_men_n292_));
  OAI210     u270(.A0(men_men_n292_), .A1(men_men_n290_), .B0(men_men_n102_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n252_), .B(men_men_n94_), .Y(men_men_n294_));
  NA2        u272(.A(men_men_n94_), .B(men_men_n41_), .Y(men_men_n295_));
  NA3        u273(.A(men_men_n295_), .B(men_men_n294_), .C(men_men_n118_), .Y(men_men_n296_));
  NA4        u274(.A(men_men_n296_), .B(men_men_n293_), .C(men_men_n288_), .D(men_men_n48_), .Y(men_men_n297_));
  INV        u275(.A(men_men_n193_), .Y(men_men_n298_));
  NA2        u276(.A(men_men_n32_), .B(x05), .Y(men_men_n299_));
  NA2        u277(.A(men_men_n404_), .B(x02), .Y(men_men_n300_));
  NA2        u278(.A(men_men_n190_), .B(x04), .Y(men_men_n301_));
  NO2        u279(.A(men_men_n301_), .B(men_men_n51_), .Y(men_men_n302_));
  NO3        u280(.A(men_men_n176_), .B(x13), .C(men_men_n31_), .Y(men_men_n303_));
  OAI210     u281(.A0(men_men_n303_), .A1(men_men_n302_), .B0(men_men_n89_), .Y(men_men_n304_));
  NO3        u282(.A(men_men_n190_), .B(men_men_n154_), .C(men_men_n52_), .Y(men_men_n305_));
  NA2        u283(.A(x12), .B(men_men_n305_), .Y(men_men_n306_));
  NA4        u284(.A(men_men_n306_), .B(men_men_n304_), .C(men_men_n300_), .D(x06), .Y(men_men_n307_));
  NO3        u285(.A(men_men_n108_), .B(men_men_n117_), .C(men_men_n38_), .Y(men_men_n308_));
  INV        u286(.A(men_men_n308_), .Y(men_men_n309_));
  OAI210     u287(.A0(men_men_n132_), .A1(men_men_n28_), .B0(men_men_n309_), .Y(men_men_n310_));
  AN2        u288(.A(men_men_n310_), .B(x04), .Y(men_men_n311_));
  AOI210     u289(.A0(men_men_n307_), .A1(men_men_n297_), .B0(men_men_n311_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n285_), .A1(x12), .B0(men_men_n312_), .Y(men03));
  OR2        u291(.A(men_men_n42_), .B(men_men_n212_), .Y(men_men_n314_));
  AOI210     u292(.A0(men_men_n144_), .A1(men_men_n94_), .B0(men_men_n314_), .Y(men_men_n315_));
  OAI210     u293(.A0(men_men_n405_), .A1(men_men_n315_), .B0(x05), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n314_), .B(x05), .Y(men_men_n317_));
  AOI210     u295(.A0(men_men_n127_), .A1(men_men_n201_), .B0(men_men_n317_), .Y(men_men_n318_));
  NO2        u296(.A(men_men_n409_), .B(x05), .Y(men_men_n319_));
  OAI210     u297(.A0(men_men_n319_), .A1(men_men_n318_), .B0(men_men_n94_), .Y(men_men_n320_));
  NA2        u298(.A(men_men_n408_), .B(x04), .Y(men_men_n321_));
  NO3        u299(.A(men_men_n295_), .B(men_men_n79_), .C(men_men_n58_), .Y(men_men_n322_));
  AOI210     u300(.A0(men_men_n180_), .A1(men_men_n94_), .B0(men_men_n136_), .Y(men_men_n323_));
  BUFFER     u301(.A(men_men_n122_), .Y(men_men_n324_));
  NO3        u302(.A(men_men_n324_), .B(men_men_n323_), .C(men_men_n322_), .Y(men_men_n325_));
  NA4        u303(.A(men_men_n325_), .B(men_men_n321_), .C(men_men_n320_), .D(men_men_n316_), .Y(men04));
  NO2        u304(.A(men_men_n82_), .B(men_men_n39_), .Y(men_men_n327_));
  XO2        u305(.A(men_men_n327_), .B(men_men_n232_), .Y(men05));
  AOI210     u306(.A0(men_men_n67_), .A1(men_men_n52_), .B0(men_men_n199_), .Y(men_men_n329_));
  AOI210     u307(.A0(men_men_n329_), .A1(men_men_n274_), .B0(men_men_n25_), .Y(men_men_n330_));
  NA3        u308(.A(men_men_n132_), .B(men_men_n119_), .C(men_men_n31_), .Y(men_men_n331_));
  AOI210     u309(.A0(men_men_n214_), .A1(men_men_n56_), .B0(men_men_n83_), .Y(men_men_n332_));
  AOI210     u310(.A0(men_men_n332_), .A1(men_men_n331_), .B0(men_men_n24_), .Y(men_men_n333_));
  OAI210     u311(.A0(men_men_n333_), .A1(men_men_n330_), .B0(men_men_n94_), .Y(men_men_n334_));
  NA2        u312(.A(x11), .B(men_men_n31_), .Y(men_men_n335_));
  NA2        u313(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n336_));
  NA2        u314(.A(men_men_n237_), .B(x03), .Y(men_men_n337_));
  OAI220     u315(.A0(men_men_n337_), .A1(men_men_n336_), .B0(men_men_n335_), .B1(men_men_n76_), .Y(men_men_n338_));
  OAI210     u316(.A0(men_men_n26_), .A1(men_men_n94_), .B0(x07), .Y(men_men_n339_));
  AOI210     u317(.A0(men_men_n338_), .A1(x06), .B0(men_men_n339_), .Y(men_men_n340_));
  AOI220     u318(.A0(men_men_n76_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n341_));
  NO3        u319(.A(men_men_n341_), .B(men_men_n23_), .C(x00), .Y(men_men_n342_));
  NA2        u320(.A(men_men_n65_), .B(x02), .Y(men_men_n343_));
  AOI210     u321(.A0(men_men_n343_), .A1(men_men_n337_), .B0(men_men_n240_), .Y(men_men_n344_));
  OR2        u322(.A(men_men_n344_), .B(men_men_n221_), .Y(men_men_n345_));
  NA2        u323(.A(men_men_n150_), .B(x05), .Y(men_men_n346_));
  NA3        u324(.A(men_men_n346_), .B(men_men_n225_), .C(men_men_n220_), .Y(men_men_n347_));
  NO2        u325(.A(men_men_n23_), .B(x10), .Y(men_men_n348_));
  OAI210     u326(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n349_));
  OR3        u327(.A(men_men_n349_), .B(men_men_n348_), .C(men_men_n44_), .Y(men_men_n350_));
  NA3        u328(.A(men_men_n350_), .B(men_men_n347_), .C(men_men_n345_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n351_), .A1(men_men_n342_), .B0(men_men_n94_), .Y(men_men_n352_));
  NA2        u330(.A(men_men_n33_), .B(men_men_n94_), .Y(men_men_n353_));
  AOI210     u331(.A0(men_men_n353_), .A1(men_men_n85_), .B0(x07), .Y(men_men_n354_));
  AOI220     u332(.A0(men_men_n354_), .A1(men_men_n352_), .B0(men_men_n340_), .B1(men_men_n334_), .Y(men_men_n355_));
  NA3        u333(.A(men_men_n23_), .B(men_men_n60_), .C(men_men_n48_), .Y(men_men_n356_));
  AO210      u334(.A0(men_men_n356_), .A1(men_men_n250_), .B0(men_men_n247_), .Y(men_men_n357_));
  AOI210     u335(.A0(men_men_n348_), .A1(men_men_n70_), .B0(men_men_n131_), .Y(men_men_n358_));
  OR2        u336(.A(men_men_n358_), .B(x03), .Y(men_men_n359_));
  NA2        u337(.A(x05), .B(men_men_n60_), .Y(men_men_n360_));
  NO2        u338(.A(men_men_n360_), .B(x11), .Y(men_men_n361_));
  NO3        u339(.A(men_men_n361_), .B(men_men_n135_), .C(men_men_n28_), .Y(men_men_n362_));
  AOI220     u340(.A0(men_men_n362_), .A1(men_men_n359_), .B0(men_men_n357_), .B1(men_men_n47_), .Y(men_men_n363_));
  NO4        u341(.A(men_men_n295_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n364_));
  OAI210     u342(.A0(men_men_n364_), .A1(men_men_n363_), .B0(men_men_n95_), .Y(men_men_n365_));
  AOI210     u343(.A0(men_men_n301_), .A1(men_men_n104_), .B0(men_men_n246_), .Y(men_men_n366_));
  NOi21      u344(.An(men_men_n286_), .B(men_men_n122_), .Y(men_men_n367_));
  OAI210     u345(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n232_), .A1(men_men_n47_), .B0(men_men_n368_), .Y(men_men_n369_));
  NO3        u347(.A(men_men_n369_), .B(men_men_n366_), .C(x08), .Y(men_men_n370_));
  AOI210     u348(.A0(men_men_n348_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n371_));
  NA2        u349(.A(x09), .B(men_men_n41_), .Y(men_men_n372_));
  OAI210     u350(.A0(men_men_n372_), .A1(men_men_n371_), .B0(men_men_n335_), .Y(men_men_n373_));
  NO2        u351(.A(x13), .B(x12), .Y(men_men_n374_));
  NO2        u352(.A(men_men_n119_), .B(men_men_n28_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n375_), .B(men_men_n251_), .Y(men_men_n376_));
  NA3        u354(.A(men_men_n298_), .B(men_men_n114_), .C(x12), .Y(men_men_n377_));
  AO210      u355(.A0(men_men_n298_), .A1(men_men_n114_), .B0(men_men_n232_), .Y(men_men_n378_));
  NA3        u356(.A(men_men_n378_), .B(men_men_n377_), .C(x08), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n374_), .A1(men_men_n373_), .B0(men_men_n379_), .Y(men_men_n380_));
  AOI210     u358(.A0(men_men_n370_), .A1(men_men_n365_), .B0(men_men_n380_), .Y(men_men_n381_));
  OAI210     u359(.A0(men_men_n360_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n382_));
  NA2        u360(.A(men_men_n266_), .B(x07), .Y(men_men_n383_));
  OAI220     u361(.A0(men_men_n383_), .A1(men_men_n336_), .B0(men_men_n135_), .B1(men_men_n43_), .Y(men_men_n384_));
  OAI210     u362(.A0(men_men_n384_), .A1(men_men_n382_), .B0(men_men_n179_), .Y(men_men_n385_));
  NA3        u363(.A(men_men_n376_), .B(men_men_n367_), .C(men_men_n294_), .Y(men_men_n386_));
  INV        u364(.A(x14), .Y(men_men_n387_));
  NO3        u365(.A(men_men_n286_), .B(men_men_n100_), .C(x11), .Y(men_men_n388_));
  NO3        u366(.A(men_men_n155_), .B(men_men_n70_), .C(men_men_n56_), .Y(men_men_n389_));
  NO3        u367(.A(men_men_n356_), .B(men_men_n295_), .C(men_men_n174_), .Y(men_men_n390_));
  NO4        u368(.A(men_men_n390_), .B(men_men_n389_), .C(men_men_n388_), .D(men_men_n387_), .Y(men_men_n391_));
  NA3        u369(.A(men_men_n391_), .B(men_men_n386_), .C(men_men_n385_), .Y(men_men_n392_));
  AOI220     u370(.A0(men_men_n353_), .A1(men_men_n60_), .B0(men_men_n375_), .B1(men_men_n154_), .Y(men_men_n393_));
  NO3        u371(.A(men_men_n116_), .B(men_men_n24_), .C(x06), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n257_), .A1(men_men_n214_), .B0(men_men_n394_), .Y(men_men_n395_));
  OAI210     u373(.A0(men_men_n44_), .A1(x04), .B0(men_men_n395_), .Y(men_men_n396_));
  NA2        u374(.A(men_men_n396_), .B(men_men_n94_), .Y(men_men_n397_));
  OAI210     u375(.A0(men_men_n393_), .A1(men_men_n84_), .B0(men_men_n397_), .Y(men_men_n398_));
  NO4        u376(.A(men_men_n398_), .B(men_men_n392_), .C(men_men_n381_), .D(men_men_n355_), .Y(men06));
  INV        u377(.A(x07), .Y(men_men_n402_));
  INV        u378(.A(x01), .Y(men_men_n403_));
  INV        u379(.A(men_men_n299_), .Y(men_men_n404_));
  INV        u380(.A(men_men_n301_), .Y(men_men_n405_));
  INV        u381(.A(x02), .Y(men_men_n406_));
  INV        u382(.A(x04), .Y(men_men_n407_));
  INV        u383(.A(men_men_n139_), .Y(men_men_n408_));
  INV        u384(.A(x13), .Y(men_men_n409_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule