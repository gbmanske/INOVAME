library verilog;
use verilog.vl_types.all;
entity Parity_Partes_vlg_vec_tst is
end Parity_Partes_vlg_vec_tst;
