//Benchmark atmr_intb_466_0.0313

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n341_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n396_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n363_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n429_, mai_mai_n430_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n373_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  AOI220     o039(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o040(.A(ori_ori_n59_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n64_), .B(ori_ori_n24_), .Y(ori_ori_n65_));
  OAI220     o043(.A0(ori_ori_n65_), .A1(ori_ori_n63_), .B0(ori_ori_n62_), .B1(ori_ori_n60_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n67_));
  OAI210     o045(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n67_), .Y(ori_ori_n68_));
  AOI220     o046(.A0(ori_ori_n68_), .A1(ori_ori_n59_), .B0(ori_ori_n66_), .B1(ori_ori_n31_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(ori_ori_n69_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n61_), .B(ori_ori_n23_), .Y(ori_ori_n71_));
  NA2        o049(.A(x09), .B(x05), .Y(ori_ori_n72_));
  NA2        o050(.A(x10), .B(x06), .Y(ori_ori_n73_));
  NA2        o051(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n74_), .A1(ori_ori_n71_), .B0(x03), .Y(ori_ori_n76_));
  NOi31      o054(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n77_));
  INV        o055(.A(x07), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n24_), .Y(ori_ori_n79_));
  NO2        o057(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(ori_ori_n36_), .Y(ori_ori_n81_));
  OAI210     o059(.A0(ori_ori_n80_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n82_));
  AOI210     o060(.A0(ori_ori_n81_), .A1(ori_ori_n48_), .B0(ori_ori_n82_), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n84_));
  NO2        o062(.A(x08), .B(x01), .Y(ori_ori_n85_));
  OAI210     o063(.A0(ori_ori_n85_), .A1(ori_ori_n84_), .B0(ori_ori_n35_), .Y(ori_ori_n86_));
  NA2        o064(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n87_));
  NO3        o065(.A(ori_ori_n86_), .B(ori_ori_n83_), .C(ori_ori_n79_), .Y(ori_ori_n88_));
  AN2        o066(.A(ori_ori_n88_), .B(ori_ori_n76_), .Y(ori_ori_n89_));
  INV        o067(.A(ori_ori_n86_), .Y(ori_ori_n90_));
  NA2        o068(.A(x11), .B(x00), .Y(ori_ori_n91_));
  NO2        o069(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n92_));
  NOi21      o070(.An(ori_ori_n91_), .B(ori_ori_n92_), .Y(ori_ori_n93_));
  NOi21      o071(.An(x01), .B(x10), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n94_), .C(x06), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n96_), .B(ori_ori_n27_), .Y(ori_ori_n97_));
  OAI210     o075(.A0(ori_ori_n396_), .A1(x07), .B0(ori_ori_n97_), .Y(ori_ori_n98_));
  NO3        o076(.A(ori_ori_n98_), .B(ori_ori_n89_), .C(ori_ori_n70_), .Y(ori01));
  INV        o077(.A(x12), .Y(ori_ori_n100_));
  INV        o078(.A(x13), .Y(ori_ori_n101_));
  NA2        o079(.A(x08), .B(x04), .Y(ori_ori_n102_));
  NO2        o080(.A(x10), .B(x01), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(ori_ori_n103_), .Y(ori_ori_n105_));
  NA2        o083(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n107_));
  NOi21      o085(.An(ori_ori_n107_), .B(ori_ori_n58_), .Y(ori_ori_n108_));
  INV        o086(.A(x13), .Y(ori_ori_n109_));
  NA2        o087(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n110_));
  NA2        o088(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(x05), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n113_));
  INV        o091(.A(ori_ori_n108_), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n114_), .B(ori_ori_n73_), .Y(ori_ori_n115_));
  NA2        o093(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n116_));
  NA2        o094(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n117_), .B(ori_ori_n116_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n120_));
  NA3        o098(.A(ori_ori_n120_), .B(ori_ori_n119_), .C(x13), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n122_));
  NOi31      o100(.An(ori_ori_n121_), .B(ori_ori_n122_), .C(ori_ori_n118_), .Y(ori_ori_n123_));
  NO3        o101(.A(ori_ori_n123_), .B(x06), .C(x03), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n124_), .B(ori_ori_n115_), .Y(ori_ori_n125_));
  NA2        o103(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n126_));
  OAI210     o104(.A0(ori_ori_n85_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n129_));
  NO2        o107(.A(x09), .B(x05), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(ori_ori_n47_), .Y(ori_ori_n131_));
  AOI210     o109(.A0(ori_ori_n131_), .A1(ori_ori_n105_), .B0(ori_ori_n49_), .Y(ori_ori_n132_));
  NA2        o110(.A(x09), .B(x00), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n107_), .B(ori_ori_n133_), .Y(ori_ori_n134_));
  INV        o112(.A(ori_ori_n132_), .Y(ori_ori_n135_));
  NO2        o113(.A(x03), .B(x02), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n86_), .B(ori_ori_n101_), .Y(ori_ori_n137_));
  OAI210     o115(.A0(ori_ori_n137_), .A1(ori_ori_n108_), .B0(ori_ori_n136_), .Y(ori_ori_n138_));
  OA210      o116(.A0(ori_ori_n135_), .A1(x11), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  OAI210     o117(.A0(ori_ori_n125_), .A1(ori_ori_n23_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n105_), .B(ori_ori_n40_), .Y(ori_ori_n141_));
  NAi21      o119(.An(x06), .B(x10), .Y(ori_ori_n142_));
  NOi21      o120(.An(x01), .B(x13), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(ori_ori_n142_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n141_), .B(ori_ori_n41_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n101_), .B(x01), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n147_), .B(x08), .Y(ori_ori_n148_));
  OAI210     o126(.A0(x05), .A1(ori_ori_n148_), .B0(ori_ori_n51_), .Y(ori_ori_n149_));
  AOI210     o127(.A0(ori_ori_n149_), .A1(ori_ori_n146_), .B0(ori_ori_n48_), .Y(ori_ori_n150_));
  AOI210     o128(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n151_));
  OAI210     o129(.A0(ori_ori_n150_), .A1(ori_ori_n145_), .B0(ori_ori_n151_), .Y(ori_ori_n152_));
  NA2        o130(.A(x10), .B(x05), .Y(ori_ori_n153_));
  NO2        o131(.A(x09), .B(x01), .Y(ori_ori_n154_));
  INV        o132(.A(ori_ori_n25_), .Y(ori_ori_n155_));
  NAi21      o133(.An(x13), .B(x00), .Y(ori_ori_n156_));
  AN2        o134(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n95_), .B(x06), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n156_), .B(ori_ori_n36_), .Y(ori_ori_n159_));
  INV        o137(.A(ori_ori_n159_), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n158_), .B(ori_ori_n157_), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n161_), .B(ori_ori_n155_), .Y(ori_ori_n162_));
  NOi21      o140(.An(x09), .B(x00), .Y(ori_ori_n163_));
  NO3        o141(.A(ori_ori_n84_), .B(ori_ori_n163_), .C(ori_ori_n47_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n164_), .B(ori_ori_n117_), .Y(ori_ori_n165_));
  NA2        o143(.A(x10), .B(x08), .Y(ori_ori_n166_));
  INV        o144(.A(ori_ori_n166_), .Y(ori_ori_n167_));
  NA2        o145(.A(x06), .B(x05), .Y(ori_ori_n168_));
  OAI210     o146(.A0(ori_ori_n168_), .A1(ori_ori_n35_), .B0(ori_ori_n100_), .Y(ori_ori_n169_));
  AOI210     o147(.A0(ori_ori_n167_), .A1(ori_ori_n58_), .B0(ori_ori_n169_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n170_), .B(ori_ori_n165_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n101_), .B(x12), .Y(ori_ori_n172_));
  AOI210     o150(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n172_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n94_), .B(ori_ori_n51_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(x02), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n173_), .B(ori_ori_n171_), .Y(ori_ori_n177_));
  NA3        o155(.A(ori_ori_n177_), .B(ori_ori_n162_), .C(ori_ori_n152_), .Y(ori_ori_n178_));
  AOI210     o156(.A0(ori_ori_n140_), .A1(ori_ori_n100_), .B0(ori_ori_n178_), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n180_), .B(ori_ori_n127_), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n116_), .B(x06), .Y(ori_ori_n183_));
  AOI210     o161(.A0(ori_ori_n182_), .A1(ori_ori_n181_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n184_), .B(x12), .Y(ori_ori_n185_));
  INV        o163(.A(ori_ori_n77_), .Y(ori_ori_n186_));
  NO2        o164(.A(x05), .B(ori_ori_n51_), .Y(ori_ori_n187_));
  OAI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n144_), .B0(ori_ori_n57_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n188_), .B(ori_ori_n186_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n94_), .B(x06), .Y(ori_ori_n190_));
  AOI210     o168(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n191_));
  NO3        o169(.A(ori_ori_n191_), .B(ori_ori_n190_), .C(ori_ori_n41_), .Y(ori_ori_n192_));
  INV        o170(.A(ori_ori_n129_), .Y(ori_ori_n193_));
  OAI210     o171(.A0(ori_ori_n193_), .A1(ori_ori_n192_), .B0(x02), .Y(ori_ori_n194_));
  AOI210     o172(.A0(ori_ori_n194_), .A1(ori_ori_n189_), .B0(ori_ori_n23_), .Y(ori_ori_n195_));
  OAI210     o173(.A0(ori_ori_n185_), .A1(ori_ori_n57_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n129_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n198_));
  OAI210     o176(.A0(ori_ori_n80_), .A1(ori_ori_n36_), .B0(ori_ori_n110_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n101_), .B(x03), .Y(ori_ori_n200_));
  AOI220     o178(.A0(ori_ori_n200_), .A1(ori_ori_n199_), .B0(ori_ori_n77_), .B1(ori_ori_n198_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n202_));
  INV        o180(.A(ori_ori_n142_), .Y(ori_ori_n203_));
  NOi21      o181(.An(x13), .B(x04), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n204_), .B(ori_ori_n77_), .C(ori_ori_n163_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n205_), .B(x05), .Y(ori_ori_n206_));
  AOI220     o184(.A0(ori_ori_n206_), .A1(ori_ori_n202_), .B0(ori_ori_n203_), .B1(ori_ori_n57_), .Y(ori_ori_n207_));
  OAI210     o185(.A0(ori_ori_n201_), .A1(ori_ori_n197_), .B0(ori_ori_n207_), .Y(ori_ori_n208_));
  INV        o186(.A(ori_ori_n92_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n209_), .B(x12), .Y(ori_ori_n210_));
  NA2        o188(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n212_));
  NO2        o190(.A(x06), .B(x00), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n213_), .B(ori_ori_n41_), .Y(ori_ori_n214_));
  INV        o192(.A(ori_ori_n73_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n215_), .B(ori_ori_n214_), .Y(ori_ori_n216_));
  NA2        o194(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n217_), .B(x03), .Y(ori_ori_n218_));
  OR2        o196(.A(ori_ori_n218_), .B(ori_ori_n216_), .Y(ori_ori_n219_));
  NA2        o197(.A(x13), .B(ori_ori_n100_), .Y(ori_ori_n220_));
  NA3        o198(.A(ori_ori_n220_), .B(ori_ori_n169_), .C(ori_ori_n93_), .Y(ori_ori_n221_));
  OAI210     o199(.A0(ori_ori_n219_), .A1(ori_ori_n211_), .B0(ori_ori_n221_), .Y(ori_ori_n222_));
  AOI210     o200(.A0(ori_ori_n210_), .A1(ori_ori_n208_), .B0(ori_ori_n222_), .Y(ori_ori_n223_));
  AOI210     o201(.A0(ori_ori_n223_), .A1(ori_ori_n196_), .B0(x07), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n72_), .B(ori_ori_n29_), .Y(ori_ori_n225_));
  NOi31      o203(.An(ori_ori_n126_), .B(ori_ori_n204_), .C(ori_ori_n163_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(ori_ori_n225_), .Y(ori_ori_n227_));
  NO2        o205(.A(x08), .B(x05), .Y(ori_ori_n228_));
  OAI210     o206(.A0(ori_ori_n77_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n229_));
  INV        o207(.A(ori_ori_n229_), .Y(ori_ori_n230_));
  NO2        o208(.A(x12), .B(x02), .Y(ori_ori_n231_));
  INV        o209(.A(ori_ori_n231_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n232_), .B(ori_ori_n209_), .Y(ori_ori_n233_));
  OA210      o211(.A0(ori_ori_n230_), .A1(ori_ori_n227_), .B0(ori_ori_n233_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n235_), .B(x01), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  AOI210     o215(.A0(ori_ori_n237_), .A1(ori_ori_n121_), .B0(ori_ori_n29_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n101_), .B(x04), .Y(ori_ori_n239_));
  NO2        o217(.A(x02), .B(ori_ori_n109_), .Y(ori_ori_n240_));
  NO3        o218(.A(ori_ori_n91_), .B(x12), .C(x03), .Y(ori_ori_n241_));
  OAI210     o219(.A0(ori_ori_n240_), .A1(ori_ori_n238_), .B0(ori_ori_n241_), .Y(ori_ori_n242_));
  AOI210     o220(.A0(ori_ori_n174_), .A1(ori_ori_n168_), .B0(ori_ori_n102_), .Y(ori_ori_n243_));
  NOi21      o221(.An(ori_ori_n225_), .B(ori_ori_n190_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n245_));
  OAI210     o223(.A0(ori_ori_n244_), .A1(ori_ori_n243_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  NO2        o224(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n247_));
  NO3        o225(.A(ori_ori_n247_), .B(ori_ori_n191_), .C(ori_ori_n158_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n211_), .B(ori_ori_n28_), .Y(ori_ori_n249_));
  OAI210     o227(.A0(ori_ori_n248_), .A1(ori_ori_n197_), .B0(ori_ori_n249_), .Y(ori_ori_n250_));
  NA3        o228(.A(ori_ori_n250_), .B(ori_ori_n246_), .C(ori_ori_n242_), .Y(ori_ori_n251_));
  NO3        o229(.A(ori_ori_n251_), .B(ori_ori_n234_), .C(ori_ori_n224_), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n179_), .A1(ori_ori_n61_), .B0(ori_ori_n252_), .Y(ori02));
  AOI210     o231(.A0(ori_ori_n126_), .A1(ori_ori_n86_), .B0(ori_ori_n119_), .Y(ori_ori_n254_));
  NOi21      o232(.An(ori_ori_n205_), .B(ori_ori_n154_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n101_), .B(ori_ori_n35_), .Y(ori_ori_n256_));
  NA3        o234(.A(ori_ori_n256_), .B(ori_ori_n167_), .C(ori_ori_n56_), .Y(ori_ori_n257_));
  OAI210     o235(.A0(ori_ori_n255_), .A1(ori_ori_n32_), .B0(ori_ori_n257_), .Y(ori_ori_n258_));
  OAI210     o236(.A0(ori_ori_n258_), .A1(ori_ori_n254_), .B0(ori_ori_n153_), .Y(ori_ori_n259_));
  INV        o237(.A(ori_ori_n153_), .Y(ori_ori_n260_));
  INV        o238(.A(ori_ori_n191_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n261_), .B(ori_ori_n101_), .Y(ori_ori_n262_));
  AOI220     o240(.A0(ori_ori_n262_), .A1(ori_ori_n260_), .B0(ori_ori_n137_), .B1(ori_ori_n136_), .Y(ori_ori_n263_));
  AOI210     o241(.A0(ori_ori_n263_), .A1(ori_ori_n259_), .B0(ori_ori_n48_), .Y(ori_ori_n264_));
  NO2        o242(.A(x05), .B(x02), .Y(ori_ori_n265_));
  OAI210     o243(.A0(ori_ori_n181_), .A1(ori_ori_n163_), .B0(ori_ori_n265_), .Y(ori_ori_n266_));
  AOI220     o244(.A0(ori_ori_n228_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n267_));
  NOi21      o245(.An(ori_ori_n256_), .B(ori_ori_n267_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n204_), .A1(ori_ori_n80_), .B0(ori_ori_n268_), .Y(ori_ori_n269_));
  AOI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n266_), .B0(ori_ori_n129_), .Y(ori_ori_n270_));
  NAi21      o248(.An(ori_ori_n206_), .B(ori_ori_n201_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n217_), .B(ori_ori_n47_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n272_), .B(ori_ori_n271_), .Y(ori_ori_n273_));
  AN2        o251(.A(ori_ori_n200_), .B(ori_ori_n199_), .Y(ori_ori_n274_));
  OAI210     o252(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n275_));
  NA2        o253(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n276_));
  BUFFER     o254(.A(ori_ori_n131_), .Y(ori_ori_n277_));
  AOI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n127_), .B0(ori_ori_n275_), .Y(ori_ori_n278_));
  OAI210     o256(.A0(ori_ori_n278_), .A1(ori_ori_n274_), .B0(ori_ori_n95_), .Y(ori_ori_n279_));
  INV        o257(.A(ori_ori_n136_), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n280_), .B(ori_ori_n118_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n281_), .B(x13), .Y(ori_ori_n282_));
  NA3        o260(.A(ori_ori_n282_), .B(ori_ori_n279_), .C(ori_ori_n273_), .Y(ori_ori_n283_));
  NO3        o261(.A(ori_ori_n283_), .B(ori_ori_n270_), .C(ori_ori_n264_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n128_), .B(x03), .Y(ori_ori_n285_));
  INV        o263(.A(ori_ori_n156_), .Y(ori_ori_n286_));
  OAI210     o264(.A0(ori_ori_n51_), .A1(ori_ori_n35_), .B0(ori_ori_n36_), .Y(ori_ori_n287_));
  AOI220     o265(.A0(ori_ori_n287_), .A1(ori_ori_n286_), .B0(ori_ori_n175_), .B1(x08), .Y(ori_ori_n288_));
  OAI210     o266(.A0(ori_ori_n288_), .A1(ori_ori_n247_), .B0(ori_ori_n285_), .Y(ori_ori_n289_));
  NA2        o267(.A(ori_ori_n289_), .B(ori_ori_n103_), .Y(ori_ori_n290_));
  INV        o268(.A(ori_ori_n56_), .Y(ori_ori_n291_));
  OAI220     o269(.A0(ori_ori_n239_), .A1(ori_ori_n291_), .B0(ori_ori_n119_), .B1(ori_ori_n28_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n292_), .B(ori_ori_n104_), .Y(ori_ori_n293_));
  NA2        o271(.A(ori_ori_n239_), .B(ori_ori_n100_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n100_), .B(ori_ori_n41_), .Y(ori_ori_n295_));
  NA3        o273(.A(ori_ori_n295_), .B(ori_ori_n294_), .C(ori_ori_n118_), .Y(ori_ori_n296_));
  NA4        o274(.A(ori_ori_n296_), .B(ori_ori_n293_), .C(ori_ori_n290_), .D(ori_ori_n48_), .Y(ori_ori_n297_));
  INV        o275(.A(ori_ori_n175_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n148_), .B(ori_ori_n40_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n300_));
  OAI220     o278(.A0(ori_ori_n300_), .A1(ori_ori_n299_), .B0(ori_ori_n298_), .B1(ori_ori_n59_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n301_), .B(x02), .Y(ori_ori_n302_));
  INV        o280(.A(ori_ori_n212_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n172_), .B(x04), .Y(ori_ori_n304_));
  NO3        o282(.A(ori_ori_n172_), .B(ori_ori_n146_), .C(ori_ori_n52_), .Y(ori_ori_n305_));
  OAI210     o283(.A0(ori_ori_n133_), .A1(ori_ori_n36_), .B0(ori_ori_n100_), .Y(ori_ori_n306_));
  OAI210     o284(.A0(ori_ori_n306_), .A1(ori_ori_n164_), .B0(ori_ori_n305_), .Y(ori_ori_n307_));
  NA3        o285(.A(ori_ori_n307_), .B(ori_ori_n302_), .C(x06), .Y(ori_ori_n308_));
  NA2        o286(.A(x09), .B(x03), .Y(ori_ori_n309_));
  OAI220     o287(.A0(ori_ori_n309_), .A1(ori_ori_n117_), .B0(ori_ori_n180_), .B1(ori_ori_n64_), .Y(ori_ori_n310_));
  OAI220     o288(.A0(ori_ori_n147_), .A1(x09), .B0(x08), .B1(ori_ori_n41_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n247_), .B(ori_ori_n116_), .C(x08), .Y(ori_ori_n312_));
  AOI210     o290(.A0(ori_ori_n311_), .A1(ori_ori_n197_), .B0(ori_ori_n312_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n314_));
  NO3        o292(.A(ori_ori_n107_), .B(ori_ori_n117_), .C(ori_ori_n38_), .Y(ori_ori_n315_));
  AOI210     o293(.A0(ori_ori_n305_), .A1(ori_ori_n314_), .B0(ori_ori_n315_), .Y(ori_ori_n316_));
  OAI210     o294(.A0(ori_ori_n313_), .A1(ori_ori_n28_), .B0(ori_ori_n316_), .Y(ori_ori_n317_));
  AO220      o295(.A0(ori_ori_n317_), .A1(x04), .B0(ori_ori_n310_), .B1(x05), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n308_), .A1(ori_ori_n297_), .B0(ori_ori_n318_), .Y(ori_ori_n319_));
  OAI210     o297(.A0(ori_ori_n284_), .A1(x12), .B0(ori_ori_n319_), .Y(ori03));
  OR2        o298(.A(ori_ori_n42_), .B(ori_ori_n198_), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n137_), .A1(ori_ori_n100_), .B0(ori_ori_n321_), .Y(ori_ori_n322_));
  AO210      o300(.A0(ori_ori_n303_), .A1(ori_ori_n87_), .B0(ori_ori_n304_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n172_), .B(ori_ori_n136_), .Y(ori_ori_n324_));
  NA3        o302(.A(ori_ori_n324_), .B(ori_ori_n323_), .C(ori_ori_n176_), .Y(ori_ori_n325_));
  OAI210     o303(.A0(ori_ori_n325_), .A1(ori_ori_n322_), .B0(x05), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n321_), .B(x05), .Y(ori_ori_n327_));
  AOI210     o305(.A0(ori_ori_n127_), .A1(ori_ori_n186_), .B0(ori_ori_n327_), .Y(ori_ori_n328_));
  AOI210     o306(.A0(ori_ori_n200_), .A1(ori_ori_n81_), .B0(ori_ori_n112_), .Y(ori_ori_n329_));
  OAI220     o307(.A0(ori_ori_n329_), .A1(ori_ori_n59_), .B0(ori_ori_n276_), .B1(ori_ori_n267_), .Y(ori_ori_n330_));
  OAI210     o308(.A0(ori_ori_n330_), .A1(ori_ori_n328_), .B0(ori_ori_n100_), .Y(ori_ori_n331_));
  AOI210     o309(.A0(ori_ori_n131_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n154_), .B(ori_ori_n122_), .Y(ori_ori_n333_));
  OAI220     o311(.A0(ori_ori_n333_), .A1(ori_ori_n37_), .B0(ori_ori_n134_), .B1(x13), .Y(ori_ori_n334_));
  OAI210     o312(.A0(ori_ori_n334_), .A1(ori_ori_n332_), .B0(x04), .Y(ori_ori_n335_));
  NO3        o313(.A(ori_ori_n295_), .B(ori_ori_n86_), .C(ori_ori_n59_), .Y(ori_ori_n336_));
  AOI210     o314(.A0(ori_ori_n160_), .A1(ori_ori_n100_), .B0(ori_ori_n131_), .Y(ori_ori_n337_));
  OA210      o315(.A0(ori_ori_n148_), .A1(x12), .B0(ori_ori_n122_), .Y(ori_ori_n338_));
  NO3        o316(.A(ori_ori_n338_), .B(ori_ori_n337_), .C(ori_ori_n336_), .Y(ori_ori_n339_));
  NA4        o317(.A(ori_ori_n339_), .B(ori_ori_n335_), .C(ori_ori_n331_), .D(ori_ori_n326_), .Y(ori04));
  NO2        o318(.A(ori_ori_n90_), .B(ori_ori_n39_), .Y(ori_ori_n341_));
  XO2        o319(.A(ori_ori_n341_), .B(ori_ori_n220_), .Y(ori05));
  AOI210     o320(.A0(ori_ori_n72_), .A1(ori_ori_n52_), .B0(ori_ori_n183_), .Y(ori_ori_n343_));
  AOI210     o321(.A0(ori_ori_n343_), .A1(ori_ori_n275_), .B0(ori_ori_n25_), .Y(ori_ori_n344_));
  NA3        o322(.A(ori_ori_n129_), .B(ori_ori_n119_), .C(ori_ori_n31_), .Y(ori_ori_n345_));
  NA2        o323(.A(ori_ori_n203_), .B(ori_ori_n57_), .Y(ori_ori_n346_));
  AOI210     o324(.A0(ori_ori_n346_), .A1(ori_ori_n345_), .B0(ori_ori_n24_), .Y(ori_ori_n347_));
  OAI210     o325(.A0(ori_ori_n347_), .A1(ori_ori_n344_), .B0(ori_ori_n100_), .Y(ori_ori_n348_));
  OAI210     o326(.A0(ori_ori_n26_), .A1(ori_ori_n100_), .B0(x07), .Y(ori_ori_n349_));
  INV        o327(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NO3        o328(.A(x02), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n351_));
  OR2        o329(.A(x02), .B(ori_ori_n211_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n213_), .B(ori_ori_n209_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n353_), .B(ori_ori_n352_), .Y(ori_ori_n354_));
  OAI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n351_), .B0(ori_ori_n100_), .Y(ori_ori_n355_));
  NA2        o333(.A(ori_ori_n33_), .B(ori_ori_n100_), .Y(ori_ori_n356_));
  AOI210     o334(.A0(ori_ori_n356_), .A1(ori_ori_n92_), .B0(x07), .Y(ori_ori_n357_));
  AOI220     o335(.A0(ori_ori_n357_), .A1(ori_ori_n355_), .B0(ori_ori_n350_), .B1(ori_ori_n348_), .Y(ori_ori_n358_));
  NO2        o336(.A(ori_ori_n47_), .B(x02), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n359_), .B(ori_ori_n101_), .Y(ori_ori_n360_));
  AOI210     o338(.A0(ori_ori_n304_), .A1(ori_ori_n106_), .B0(ori_ori_n231_), .Y(ori_ori_n361_));
  NOi21      o339(.An(ori_ori_n285_), .B(ori_ori_n122_), .Y(ori_ori_n362_));
  NO2        o340(.A(ori_ori_n362_), .B(ori_ori_n232_), .Y(ori_ori_n363_));
  OAI210     o341(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n364_));
  AOI210     o342(.A0(ori_ori_n220_), .A1(ori_ori_n47_), .B0(ori_ori_n364_), .Y(ori_ori_n365_));
  NO4        o343(.A(ori_ori_n365_), .B(ori_ori_n363_), .C(ori_ori_n361_), .D(x08), .Y(ori_ori_n366_));
  NA2        o344(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n367_));
  NO2        o345(.A(ori_ori_n367_), .B(x03), .Y(ori_ori_n368_));
  NO2        o346(.A(x13), .B(x12), .Y(ori_ori_n369_));
  NO2        o347(.A(ori_ori_n119_), .B(ori_ori_n28_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n370_), .B(ori_ori_n236_), .Y(ori_ori_n371_));
  OR3        o349(.A(ori_ori_n371_), .B(x12), .C(x03), .Y(ori_ori_n372_));
  NA3        o350(.A(ori_ori_n298_), .B(ori_ori_n113_), .C(x12), .Y(ori_ori_n373_));
  AO210      o351(.A0(ori_ori_n298_), .A1(ori_ori_n113_), .B0(ori_ori_n220_), .Y(ori_ori_n374_));
  NA4        o352(.A(ori_ori_n374_), .B(ori_ori_n373_), .C(ori_ori_n372_), .D(x08), .Y(ori_ori_n375_));
  AOI210     o353(.A0(ori_ori_n369_), .A1(ori_ori_n368_), .B0(ori_ori_n375_), .Y(ori_ori_n376_));
  AOI210     o354(.A0(ori_ori_n366_), .A1(ori_ori_n360_), .B0(ori_ori_n376_), .Y(ori_ori_n377_));
  INV        o355(.A(x03), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n130_), .B(ori_ori_n43_), .Y(ori_ori_n379_));
  OAI210     o357(.A0(ori_ori_n379_), .A1(ori_ori_n378_), .B0(ori_ori_n159_), .Y(ori_ori_n380_));
  NA3        o358(.A(ori_ori_n371_), .B(ori_ori_n362_), .C(ori_ori_n294_), .Y(ori_ori_n381_));
  INV        o359(.A(x14), .Y(ori_ori_n382_));
  NO3        o360(.A(ori_ori_n147_), .B(ori_ori_n75_), .C(ori_ori_n57_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n383_), .B(ori_ori_n382_), .Y(ori_ori_n384_));
  NA3        o362(.A(ori_ori_n384_), .B(ori_ori_n381_), .C(ori_ori_n380_), .Y(ori_ori_n385_));
  NA2        o363(.A(ori_ori_n356_), .B(ori_ori_n61_), .Y(ori_ori_n386_));
  NOi21      o364(.An(ori_ori_n239_), .B(ori_ori_n134_), .Y(ori_ori_n387_));
  NO3        o365(.A(ori_ori_n116_), .B(ori_ori_n24_), .C(x06), .Y(ori_ori_n388_));
  AOI210     o366(.A0(ori_ori_n245_), .A1(ori_ori_n203_), .B0(ori_ori_n388_), .Y(ori_ori_n389_));
  OAI210     o367(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n389_), .Y(ori_ori_n390_));
  OAI210     o368(.A0(ori_ori_n390_), .A1(ori_ori_n387_), .B0(ori_ori_n100_), .Y(ori_ori_n391_));
  OAI210     o369(.A0(ori_ori_n386_), .A1(ori_ori_n91_), .B0(ori_ori_n391_), .Y(ori_ori_n392_));
  NO4        o370(.A(ori_ori_n392_), .B(ori_ori_n385_), .C(ori_ori_n377_), .D(ori_ori_n358_), .Y(ori06));
  INV        o371(.A(ori_ori_n93_), .Y(ori_ori_n396_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NOi21      m029(.An(x01), .B(x09), .Y(mai_mai_n52_));
  INV        m030(.A(x00), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  NO2        m032(.A(mai_mai_n54_), .B(mai_mai_n52_), .Y(mai_mai_n55_));
  NA2        m033(.A(x09), .B(mai_mai_n53_), .Y(mai_mai_n56_));
  INV        m034(.A(x07), .Y(mai_mai_n57_));
  AOI220     m035(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n57_), .Y(mai_mai_n58_));
  INV        m036(.A(mai_mai_n55_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n60_), .B(mai_mai_n24_), .Y(mai_mai_n61_));
  OAI220     m039(.A0(mai_mai_n61_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .B1(mai_mai_n56_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n57_), .B(mai_mai_n48_), .Y(mai_mai_n63_));
  OAI210     m041(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n63_), .Y(mai_mai_n64_));
  AOI220     m042(.A0(mai_mai_n64_), .A1(mai_mai_n55_), .B0(mai_mai_n62_), .B1(mai_mai_n31_), .Y(mai_mai_n65_));
  NO2        m043(.A(mai_mai_n65_), .B(x05), .Y(mai_mai_n66_));
  NO2        m044(.A(mai_mai_n57_), .B(mai_mai_n23_), .Y(mai_mai_n67_));
  NA2        m045(.A(x09), .B(x05), .Y(mai_mai_n68_));
  NA2        m046(.A(x10), .B(x06), .Y(mai_mai_n69_));
  NA3        m047(.A(mai_mai_n69_), .B(mai_mai_n68_), .C(mai_mai_n28_), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n57_), .B(mai_mai_n41_), .Y(mai_mai_n71_));
  OAI210     m049(.A0(mai_mai_n70_), .A1(mai_mai_n67_), .B0(x03), .Y(mai_mai_n72_));
  NOi31      m050(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n73_));
  INV        m051(.A(mai_mai_n24_), .Y(mai_mai_n74_));
  NO2        m052(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n75_), .B(mai_mai_n36_), .Y(mai_mai_n76_));
  OAI210     m054(.A0(mai_mai_n75_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n77_));
  INV        m055(.A(mai_mai_n77_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n79_));
  NO2        m057(.A(x08), .B(x01), .Y(mai_mai_n80_));
  OAI210     m058(.A0(mai_mai_n80_), .A1(mai_mai_n79_), .B0(mai_mai_n35_), .Y(mai_mai_n81_));
  NA2        m059(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n82_));
  NO3        m060(.A(mai_mai_n81_), .B(mai_mai_n78_), .C(mai_mai_n74_), .Y(mai_mai_n83_));
  AN2        m061(.A(mai_mai_n83_), .B(mai_mai_n72_), .Y(mai_mai_n84_));
  INV        m062(.A(mai_mai_n81_), .Y(mai_mai_n85_));
  NO2        m063(.A(x06), .B(x05), .Y(mai_mai_n86_));
  NA2        m064(.A(x11), .B(x00), .Y(mai_mai_n87_));
  NO2        m065(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n88_));
  NOi21      m066(.An(mai_mai_n87_), .B(mai_mai_n88_), .Y(mai_mai_n89_));
  AOI210     m067(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NOi21      m068(.An(x01), .B(x10), .Y(mai_mai_n91_));
  NO2        m069(.A(mai_mai_n29_), .B(mai_mai_n53_), .Y(mai_mai_n92_));
  NO3        m070(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(x06), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n93_), .B(mai_mai_n27_), .Y(mai_mai_n94_));
  OAI210     m072(.A0(mai_mai_n90_), .A1(x07), .B0(mai_mai_n94_), .Y(mai_mai_n95_));
  NO3        m073(.A(mai_mai_n95_), .B(mai_mai_n84_), .C(mai_mai_n66_), .Y(mai01));
  INV        m074(.A(x12), .Y(mai_mai_n97_));
  INV        m075(.A(x13), .Y(mai_mai_n98_));
  NA2        m076(.A(x08), .B(x04), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n91_), .B(mai_mai_n28_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n68_), .Y(mai_mai_n101_));
  NO2        m079(.A(x10), .B(x01), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NA2        m082(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n105_), .B(mai_mai_n36_), .Y(mai_mai_n106_));
  AOI210     m084(.A0(mai_mai_n106_), .A1(mai_mai_n104_), .B0(mai_mai_n101_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(mai_mai_n98_), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n52_), .B(x05), .Y(mai_mai_n109_));
  NOi21      m087(.An(mai_mai_n109_), .B(mai_mai_n54_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n111_));
  NA3        m089(.A(x13), .B(mai_mai_n111_), .C(x06), .Y(mai_mai_n112_));
  INV        m090(.A(mai_mai_n112_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n80_), .B(x13), .Y(mai_mai_n114_));
  NA2        m092(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NA2        m094(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n117_), .B(x05), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n118_), .B(mai_mai_n116_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n35_), .B(mai_mai_n53_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n120_), .B(mai_mai_n98_), .Y(mai_mai_n121_));
  AOI210     m099(.A0(mai_mai_n121_), .A1(mai_mai_n76_), .B0(mai_mai_n110_), .Y(mai_mai_n122_));
  AOI210     m100(.A0(mai_mai_n122_), .A1(mai_mai_n119_), .B0(mai_mai_n69_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n124_));
  NA2        m102(.A(x10), .B(mai_mai_n53_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n127_));
  NO3        m105(.A(mai_mai_n120_), .B(mai_mai_n75_), .C(mai_mai_n36_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n128_), .C(mai_mai_n126_), .Y(mai_mai_n130_));
  NO3        m108(.A(mai_mai_n130_), .B(x06), .C(x03), .Y(mai_mai_n131_));
  NO4        m109(.A(mai_mai_n131_), .B(mai_mai_n123_), .C(mai_mai_n113_), .D(mai_mai_n108_), .Y(mai_mai_n132_));
  NA2        m110(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n133_));
  OAI210     m111(.A0(mai_mai_n80_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n137_));
  AOI210     m115(.A0(mai_mai_n137_), .A1(mai_mai_n49_), .B0(mai_mai_n136_), .Y(mai_mai_n138_));
  AN2        m116(.A(mai_mai_n138_), .B(mai_mai_n135_), .Y(mai_mai_n139_));
  NO2        m117(.A(x09), .B(x05), .Y(mai_mai_n140_));
  NA2        m118(.A(mai_mai_n140_), .B(mai_mai_n47_), .Y(mai_mai_n141_));
  NO2        m119(.A(mai_mai_n104_), .B(mai_mai_n49_), .Y(mai_mai_n142_));
  NA2        m120(.A(x09), .B(x00), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n109_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n73_), .B(mai_mai_n50_), .Y(mai_mai_n145_));
  AOI210     m123(.A0(mai_mai_n145_), .A1(mai_mai_n144_), .B0(mai_mai_n137_), .Y(mai_mai_n146_));
  NO3        m124(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n139_), .Y(mai_mai_n147_));
  NO2        m125(.A(x03), .B(x02), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n81_), .B(mai_mai_n98_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n149_), .A1(mai_mai_n110_), .B0(mai_mai_n148_), .Y(mai_mai_n150_));
  OA210      m128(.A0(mai_mai_n147_), .A1(x11), .B0(mai_mai_n150_), .Y(mai_mai_n151_));
  OAI210     m129(.A0(mai_mai_n132_), .A1(mai_mai_n23_), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  NA2        m130(.A(mai_mai_n104_), .B(mai_mai_n40_), .Y(mai_mai_n153_));
  NAi21      m131(.An(x06), .B(x10), .Y(mai_mai_n154_));
  NOi21      m132(.An(x01), .B(x13), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n154_), .Y(mai_mai_n156_));
  BUFFER     m134(.A(mai_mai_n156_), .Y(mai_mai_n157_));
  AOI210     m135(.A0(mai_mai_n157_), .A1(mai_mai_n153_), .B0(mai_mai_n41_), .Y(mai_mai_n158_));
  NO2        m136(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n98_), .B(x01), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(x08), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n159_), .B(mai_mai_n48_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n163_));
  OAI210     m141(.A0(mai_mai_n162_), .A1(mai_mai_n158_), .B0(mai_mai_n163_), .Y(mai_mai_n164_));
  NA2        m142(.A(x04), .B(x02), .Y(mai_mai_n165_));
  NA2        m143(.A(x10), .B(x05), .Y(mai_mai_n166_));
  NA2        m144(.A(x09), .B(x06), .Y(mai_mai_n167_));
  NO2        m145(.A(x09), .B(x01), .Y(mai_mai_n168_));
  NO3        m146(.A(mai_mai_n168_), .B(mai_mai_n102_), .C(mai_mai_n31_), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n169_), .B(x00), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n109_), .B(x08), .Y(mai_mai_n171_));
  OAI210     m149(.A0(mai_mai_n430_), .A1(x11), .B0(mai_mai_n170_), .Y(mai_mai_n172_));
  NAi21      m150(.An(mai_mai_n165_), .B(mai_mai_n172_), .Y(mai_mai_n173_));
  INV        m151(.A(mai_mai_n25_), .Y(mai_mai_n174_));
  NAi21      m152(.An(x13), .B(x00), .Y(mai_mai_n175_));
  AOI210     m153(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n175_), .Y(mai_mai_n176_));
  AOI220     m154(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n177_));
  OAI210     m155(.A0(mai_mai_n166_), .A1(mai_mai_n35_), .B0(mai_mai_n177_), .Y(mai_mai_n178_));
  AN2        m156(.A(mai_mai_n178_), .B(mai_mai_n176_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n92_), .B(x06), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n175_), .B(mai_mai_n36_), .Y(mai_mai_n181_));
  INV        m159(.A(mai_mai_n181_), .Y(mai_mai_n182_));
  OAI210     m160(.A0(mai_mai_n182_), .A1(mai_mai_n167_), .B0(mai_mai_n69_), .Y(mai_mai_n183_));
  OAI210     m161(.A0(mai_mai_n183_), .A1(mai_mai_n179_), .B0(mai_mai_n174_), .Y(mai_mai_n184_));
  NOi21      m162(.An(x09), .B(x00), .Y(mai_mai_n185_));
  NO3        m163(.A(mai_mai_n79_), .B(mai_mai_n185_), .C(mai_mai_n47_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n186_), .B(mai_mai_n125_), .Y(mai_mai_n187_));
  NA2        m165(.A(mai_mai_n97_), .B(mai_mai_n187_), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n98_), .B(x12), .Y(mai_mai_n189_));
  AOI210     m167(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n189_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n91_), .B(mai_mai_n50_), .Y(mai_mai_n191_));
  NO2        m169(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n192_), .B(x02), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n193_), .B(mai_mai_n191_), .Y(mai_mai_n194_));
  AOI210     m172(.A0(mai_mai_n190_), .A1(mai_mai_n188_), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  NA4        m173(.A(mai_mai_n195_), .B(mai_mai_n184_), .C(mai_mai_n173_), .D(mai_mai_n164_), .Y(mai_mai_n196_));
  AOI210     m174(.A0(mai_mai_n152_), .A1(mai_mai_n97_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  INV        m175(.A(mai_mai_n70_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n198_), .B(mai_mai_n135_), .Y(mai_mai_n199_));
  NA2        m177(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n200_), .B(mai_mai_n134_), .Y(mai_mai_n201_));
  AOI210     m179(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n124_), .B(x06), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n202_), .A1(mai_mai_n201_), .B0(mai_mai_n203_), .Y(mai_mai_n204_));
  AOI210     m182(.A0(mai_mai_n204_), .A1(mai_mai_n199_), .B0(x12), .Y(mai_mai_n205_));
  INV        m183(.A(mai_mai_n73_), .Y(mai_mai_n206_));
  NO2        m184(.A(x05), .B(mai_mai_n50_), .Y(mai_mai_n207_));
  OAI210     m185(.A0(mai_mai_n207_), .A1(mai_mai_n156_), .B0(mai_mai_n53_), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n208_), .B(mai_mai_n206_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n91_), .B(x06), .Y(mai_mai_n210_));
  AOI210     m188(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n211_));
  NA4        m189(.A(mai_mai_n154_), .B(mai_mai_n52_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n212_));
  NA2        m190(.A(mai_mai_n212_), .B(mai_mai_n137_), .Y(mai_mai_n213_));
  NA2        m191(.A(mai_mai_n213_), .B(x02), .Y(mai_mai_n214_));
  AOI210     m192(.A0(mai_mai_n214_), .A1(mai_mai_n209_), .B0(mai_mai_n23_), .Y(mai_mai_n215_));
  OAI210     m193(.A0(mai_mai_n205_), .A1(mai_mai_n53_), .B0(mai_mai_n215_), .Y(mai_mai_n216_));
  INV        m194(.A(mai_mai_n137_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n218_));
  OAI210     m196(.A0(mai_mai_n75_), .A1(mai_mai_n36_), .B0(mai_mai_n115_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n98_), .B(x03), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n221_));
  INV        m199(.A(mai_mai_n154_), .Y(mai_mai_n222_));
  NOi21      m200(.An(x13), .B(x04), .Y(mai_mai_n223_));
  NO3        m201(.A(mai_mai_n223_), .B(mai_mai_n73_), .C(mai_mai_n185_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n224_), .B(x05), .Y(mai_mai_n225_));
  AOI220     m203(.A0(mai_mai_n225_), .A1(mai_mai_n221_), .B0(mai_mai_n222_), .B1(mai_mai_n53_), .Y(mai_mai_n226_));
  INV        m204(.A(mai_mai_n226_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n88_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n228_), .B(x12), .Y(mai_mai_n229_));
  NA2        m207(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n231_));
  OAI210     m209(.A0(mai_mai_n231_), .A1(mai_mai_n178_), .B0(mai_mai_n176_), .Y(mai_mai_n232_));
  AOI210     m210(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n233_));
  NO2        m211(.A(x06), .B(x00), .Y(mai_mai_n234_));
  NO3        m212(.A(mai_mai_n234_), .B(mai_mai_n233_), .C(mai_mai_n41_), .Y(mai_mai_n235_));
  OAI210     m213(.A0(mai_mai_n99_), .A1(mai_mai_n143_), .B0(mai_mai_n69_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n238_), .B(x03), .Y(mai_mai_n239_));
  OA210      m217(.A0(mai_mai_n239_), .A1(mai_mai_n237_), .B0(mai_mai_n232_), .Y(mai_mai_n240_));
  NA2        m218(.A(x13), .B(mai_mai_n97_), .Y(mai_mai_n241_));
  NA3        m219(.A(mai_mai_n241_), .B(x12), .C(mai_mai_n89_), .Y(mai_mai_n242_));
  OAI210     m220(.A0(mai_mai_n240_), .A1(mai_mai_n230_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n229_), .A1(mai_mai_n227_), .B0(mai_mai_n243_), .Y(mai_mai_n244_));
  AOI210     m222(.A0(mai_mai_n244_), .A1(mai_mai_n216_), .B0(x07), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n68_), .B(mai_mai_n29_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n223_), .B(mai_mai_n185_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n247_), .A1(mai_mai_n145_), .B0(mai_mai_n246_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n98_), .B(x06), .Y(mai_mai_n249_));
  INV        m227(.A(mai_mai_n249_), .Y(mai_mai_n250_));
  NO2        m228(.A(x08), .B(x05), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n251_), .B(mai_mai_n233_), .Y(mai_mai_n252_));
  NA2        m230(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n253_));
  OAI210     m231(.A0(mai_mai_n252_), .A1(mai_mai_n250_), .B0(mai_mai_n253_), .Y(mai_mai_n254_));
  NO2        m232(.A(x12), .B(x02), .Y(mai_mai_n255_));
  INV        m233(.A(mai_mai_n255_), .Y(mai_mai_n256_));
  NO2        m234(.A(mai_mai_n256_), .B(mai_mai_n228_), .Y(mai_mai_n257_));
  OA210      m235(.A0(mai_mai_n254_), .A1(mai_mai_n248_), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  NA2        m236(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n259_), .B(x01), .Y(mai_mai_n260_));
  NOi21      m238(.An(mai_mai_n80_), .B(mai_mai_n115_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n261_), .B(mai_mai_n260_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n262_), .B(mai_mai_n29_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n249_), .B(mai_mai_n219_), .Y(mai_mai_n264_));
  NA2        m242(.A(mai_mai_n98_), .B(x04), .Y(mai_mai_n265_));
  NA2        m243(.A(mai_mai_n265_), .B(mai_mai_n28_), .Y(mai_mai_n266_));
  OAI210     m244(.A0(mai_mai_n266_), .A1(mai_mai_n114_), .B0(mai_mai_n264_), .Y(mai_mai_n267_));
  NO3        m245(.A(mai_mai_n87_), .B(x12), .C(x03), .Y(mai_mai_n268_));
  OAI210     m246(.A0(mai_mai_n267_), .A1(mai_mai_n263_), .B0(mai_mai_n268_), .Y(mai_mai_n269_));
  NOi21      m247(.An(mai_mai_n246_), .B(mai_mai_n210_), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n270_), .B(mai_mai_n271_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n54_), .B(x05), .Y(mai_mai_n273_));
  NO3        m251(.A(mai_mai_n273_), .B(mai_mai_n211_), .C(mai_mai_n180_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n230_), .B(mai_mai_n28_), .Y(mai_mai_n275_));
  OAI210     m253(.A0(mai_mai_n274_), .A1(mai_mai_n217_), .B0(mai_mai_n275_), .Y(mai_mai_n276_));
  NA3        m254(.A(mai_mai_n276_), .B(mai_mai_n272_), .C(mai_mai_n269_), .Y(mai_mai_n277_));
  NO3        m255(.A(mai_mai_n277_), .B(mai_mai_n258_), .C(mai_mai_n245_), .Y(mai_mai_n278_));
  OAI210     m256(.A0(mai_mai_n197_), .A1(mai_mai_n57_), .B0(mai_mai_n278_), .Y(mai02));
  AOI210     m257(.A0(mai_mai_n133_), .A1(mai_mai_n81_), .B0(mai_mai_n127_), .Y(mai_mai_n280_));
  NOi21      m258(.An(mai_mai_n224_), .B(mai_mai_n168_), .Y(mai_mai_n281_));
  NO2        m259(.A(mai_mai_n281_), .B(mai_mai_n32_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n282_), .A1(mai_mai_n280_), .B0(mai_mai_n166_), .Y(mai_mai_n283_));
  INV        m261(.A(mai_mai_n166_), .Y(mai_mai_n284_));
  AOI210     m262(.A0(mai_mai_n111_), .A1(mai_mai_n82_), .B0(mai_mai_n211_), .Y(mai_mai_n285_));
  OAI220     m263(.A0(mai_mai_n285_), .A1(mai_mai_n98_), .B0(mai_mai_n81_), .B1(mai_mai_n50_), .Y(mai_mai_n286_));
  AOI220     m264(.A0(mai_mai_n286_), .A1(mai_mai_n284_), .B0(mai_mai_n149_), .B1(mai_mai_n148_), .Y(mai_mai_n287_));
  AOI210     m265(.A0(mai_mai_n287_), .A1(mai_mai_n283_), .B0(mai_mai_n48_), .Y(mai_mai_n288_));
  NO2        m266(.A(x05), .B(x02), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n201_), .A1(mai_mai_n185_), .B0(mai_mai_n289_), .Y(mai_mai_n290_));
  AOI220     m268(.A0(mai_mai_n251_), .A1(mai_mai_n54_), .B0(mai_mai_n52_), .B1(mai_mai_n36_), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n290_), .B(mai_mai_n137_), .Y(mai_mai_n292_));
  NO2        m270(.A(mai_mai_n238_), .B(mai_mai_n47_), .Y(mai_mai_n293_));
  NA2        m271(.A(mai_mai_n293_), .B(mai_mai_n225_), .Y(mai_mai_n294_));
  AN2        m272(.A(mai_mai_n220_), .B(mai_mai_n219_), .Y(mai_mai_n295_));
  OAI210     m273(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n296_));
  NA2        m274(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n297_));
  OA210      m275(.A0(mai_mai_n297_), .A1(x08), .B0(mai_mai_n141_), .Y(mai_mai_n298_));
  AOI210     m276(.A0(mai_mai_n298_), .A1(mai_mai_n134_), .B0(mai_mai_n296_), .Y(mai_mai_n299_));
  OAI210     m277(.A0(mai_mai_n299_), .A1(mai_mai_n295_), .B0(mai_mai_n92_), .Y(mai_mai_n300_));
  NA3        m278(.A(mai_mai_n92_), .B(mai_mai_n80_), .C(mai_mai_n218_), .Y(mai_mai_n301_));
  NA3        m279(.A(mai_mai_n91_), .B(mai_mai_n79_), .C(mai_mai_n42_), .Y(mai_mai_n302_));
  AOI210     m280(.A0(mai_mai_n302_), .A1(mai_mai_n301_), .B0(x04), .Y(mai_mai_n303_));
  INV        m281(.A(mai_mai_n148_), .Y(mai_mai_n304_));
  OAI220     m282(.A0(mai_mai_n252_), .A1(mai_mai_n100_), .B0(mai_mai_n304_), .B1(mai_mai_n126_), .Y(mai_mai_n305_));
  AOI210     m283(.A0(mai_mai_n305_), .A1(x13), .B0(mai_mai_n303_), .Y(mai_mai_n306_));
  NA3        m284(.A(mai_mai_n306_), .B(mai_mai_n300_), .C(mai_mai_n294_), .Y(mai_mai_n307_));
  NO3        m285(.A(mai_mai_n307_), .B(mai_mai_n292_), .C(mai_mai_n288_), .Y(mai_mai_n308_));
  NA2        m286(.A(mai_mai_n136_), .B(x03), .Y(mai_mai_n309_));
  OAI210     m287(.A0(mai_mai_n175_), .A1(mai_mai_n273_), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n310_), .B(mai_mai_n102_), .Y(mai_mai_n311_));
  NA2        m289(.A(mai_mai_n165_), .B(mai_mai_n160_), .Y(mai_mai_n312_));
  AN2        m290(.A(mai_mai_n312_), .B(mai_mai_n171_), .Y(mai_mai_n313_));
  INV        m291(.A(mai_mai_n52_), .Y(mai_mai_n314_));
  OAI220     m292(.A0(mai_mai_n265_), .A1(mai_mai_n314_), .B0(mai_mai_n127_), .B1(mai_mai_n28_), .Y(mai_mai_n315_));
  OAI210     m293(.A0(mai_mai_n315_), .A1(mai_mai_n313_), .B0(mai_mai_n103_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n265_), .B(mai_mai_n97_), .Y(mai_mai_n317_));
  NA2        m295(.A(mai_mai_n97_), .B(mai_mai_n41_), .Y(mai_mai_n318_));
  NA3        m296(.A(mai_mai_n318_), .B(mai_mai_n317_), .C(mai_mai_n126_), .Y(mai_mai_n319_));
  NA4        m297(.A(mai_mai_n319_), .B(mai_mai_n316_), .C(mai_mai_n311_), .D(mai_mai_n48_), .Y(mai_mai_n320_));
  INV        m298(.A(mai_mai_n192_), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n161_), .B(mai_mai_n40_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n323_));
  OAI220     m301(.A0(mai_mai_n323_), .A1(mai_mai_n322_), .B0(mai_mai_n321_), .B1(mai_mai_n55_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n324_), .B(x02), .Y(mai_mai_n325_));
  INV        m303(.A(mai_mai_n231_), .Y(mai_mai_n326_));
  NA2        m304(.A(mai_mai_n189_), .B(x04), .Y(mai_mai_n327_));
  NO2        m305(.A(mai_mai_n327_), .B(mai_mai_n326_), .Y(mai_mai_n328_));
  NO3        m306(.A(mai_mai_n177_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n329_));
  OAI210     m307(.A0(mai_mai_n329_), .A1(mai_mai_n328_), .B0(mai_mai_n92_), .Y(mai_mai_n330_));
  NO3        m308(.A(mai_mai_n189_), .B(mai_mai_n159_), .C(mai_mai_n51_), .Y(mai_mai_n331_));
  OAI210     m309(.A0(mai_mai_n143_), .A1(mai_mai_n36_), .B0(mai_mai_n97_), .Y(mai_mai_n332_));
  OAI210     m310(.A0(mai_mai_n332_), .A1(mai_mai_n186_), .B0(mai_mai_n331_), .Y(mai_mai_n333_));
  NA4        m311(.A(mai_mai_n333_), .B(mai_mai_n330_), .C(mai_mai_n325_), .D(x06), .Y(mai_mai_n334_));
  NA2        m312(.A(x09), .B(x03), .Y(mai_mai_n335_));
  OAI220     m313(.A0(mai_mai_n335_), .A1(mai_mai_n125_), .B0(mai_mai_n200_), .B1(mai_mai_n60_), .Y(mai_mai_n336_));
  NO2        m314(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n331_), .B(mai_mai_n337_), .Y(mai_mai_n338_));
  INV        m316(.A(mai_mai_n338_), .Y(mai_mai_n339_));
  AO220      m317(.A0(mai_mai_n339_), .A1(x04), .B0(mai_mai_n336_), .B1(x05), .Y(mai_mai_n340_));
  AOI210     m318(.A0(mai_mai_n334_), .A1(mai_mai_n320_), .B0(mai_mai_n340_), .Y(mai_mai_n341_));
  OAI210     m319(.A0(mai_mai_n308_), .A1(x12), .B0(mai_mai_n341_), .Y(mai03));
  OR2        m320(.A(mai_mai_n42_), .B(mai_mai_n218_), .Y(mai_mai_n343_));
  AOI210     m321(.A0(mai_mai_n149_), .A1(mai_mai_n97_), .B0(mai_mai_n343_), .Y(mai_mai_n344_));
  AO210      m322(.A0(mai_mai_n326_), .A1(mai_mai_n82_), .B0(mai_mai_n327_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n189_), .B(mai_mai_n148_), .Y(mai_mai_n346_));
  NA3        m324(.A(mai_mai_n346_), .B(mai_mai_n345_), .C(mai_mai_n193_), .Y(mai_mai_n347_));
  OAI210     m325(.A0(mai_mai_n347_), .A1(mai_mai_n344_), .B0(x05), .Y(mai_mai_n348_));
  NA2        m326(.A(mai_mai_n343_), .B(x05), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n134_), .A1(mai_mai_n206_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  AOI210     m328(.A0(mai_mai_n220_), .A1(mai_mai_n76_), .B0(mai_mai_n118_), .Y(mai_mai_n351_));
  OAI220     m329(.A0(mai_mai_n351_), .A1(mai_mai_n55_), .B0(mai_mai_n297_), .B1(mai_mai_n291_), .Y(mai_mai_n352_));
  OAI210     m330(.A0(mai_mai_n352_), .A1(mai_mai_n350_), .B0(mai_mai_n97_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n141_), .A1(mai_mai_n56_), .B0(mai_mai_n38_), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n168_), .B(mai_mai_n129_), .Y(mai_mai_n355_));
  OAI220     m333(.A0(mai_mai_n355_), .A1(mai_mai_n37_), .B0(mai_mai_n144_), .B1(x13), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n356_), .A1(mai_mai_n354_), .B0(x04), .Y(mai_mai_n357_));
  NO3        m335(.A(mai_mai_n318_), .B(mai_mai_n81_), .C(mai_mai_n55_), .Y(mai_mai_n358_));
  AOI210     m336(.A0(mai_mai_n182_), .A1(mai_mai_n97_), .B0(mai_mai_n141_), .Y(mai_mai_n359_));
  OA210      m337(.A0(mai_mai_n161_), .A1(x12), .B0(mai_mai_n129_), .Y(mai_mai_n360_));
  NO3        m338(.A(mai_mai_n360_), .B(mai_mai_n359_), .C(mai_mai_n358_), .Y(mai_mai_n361_));
  NA4        m339(.A(mai_mai_n361_), .B(mai_mai_n357_), .C(mai_mai_n353_), .D(mai_mai_n348_), .Y(mai04));
  NO2        m340(.A(mai_mai_n85_), .B(mai_mai_n39_), .Y(mai_mai_n363_));
  XO2        m341(.A(mai_mai_n363_), .B(mai_mai_n241_), .Y(mai05));
  AOI210     m342(.A0(mai_mai_n68_), .A1(mai_mai_n51_), .B0(mai_mai_n203_), .Y(mai_mai_n365_));
  AOI210     m343(.A0(mai_mai_n365_), .A1(mai_mai_n296_), .B0(mai_mai_n25_), .Y(mai_mai_n366_));
  NO2        m344(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n367_));
  OAI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n366_), .B0(mai_mai_n97_), .Y(mai_mai_n368_));
  NA2        m346(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n369_));
  NA2        m347(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n370_));
  NA2        m348(.A(mai_mai_n246_), .B(x03), .Y(mai_mai_n371_));
  OAI220     m349(.A0(mai_mai_n371_), .A1(mai_mai_n370_), .B0(mai_mai_n369_), .B1(mai_mai_n77_), .Y(mai_mai_n372_));
  OAI210     m350(.A0(mai_mai_n26_), .A1(mai_mai_n97_), .B0(x07), .Y(mai_mai_n373_));
  AOI210     m351(.A0(mai_mai_n372_), .A1(x06), .B0(mai_mai_n373_), .Y(mai_mai_n374_));
  AOI220     m352(.A0(mai_mai_n77_), .A1(mai_mai_n31_), .B0(mai_mai_n51_), .B1(mai_mai_n50_), .Y(mai_mai_n375_));
  NO3        m353(.A(mai_mai_n375_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n376_));
  NO2        m354(.A(mai_mai_n371_), .B(mai_mai_n249_), .Y(mai_mai_n377_));
  OR2        m355(.A(mai_mai_n377_), .B(mai_mai_n230_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n155_), .B(x05), .Y(mai_mai_n379_));
  NA3        m357(.A(mai_mai_n379_), .B(mai_mai_n234_), .C(mai_mai_n228_), .Y(mai_mai_n380_));
  NO2        m358(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n381_));
  OAI210     m359(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n382_));
  OR3        m360(.A(mai_mai_n382_), .B(mai_mai_n381_), .C(mai_mai_n44_), .Y(mai_mai_n383_));
  NA3        m361(.A(mai_mai_n383_), .B(mai_mai_n380_), .C(mai_mai_n378_), .Y(mai_mai_n384_));
  OAI210     m362(.A0(mai_mai_n384_), .A1(mai_mai_n376_), .B0(mai_mai_n97_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n33_), .B(mai_mai_n97_), .Y(mai_mai_n386_));
  AOI210     m364(.A0(mai_mai_n386_), .A1(mai_mai_n88_), .B0(x07), .Y(mai_mai_n387_));
  AOI220     m365(.A0(mai_mai_n387_), .A1(mai_mai_n385_), .B0(mai_mai_n374_), .B1(mai_mai_n368_), .Y(mai_mai_n388_));
  NA3        m366(.A(mai_mai_n23_), .B(mai_mai_n57_), .C(mai_mai_n48_), .Y(mai_mai_n389_));
  OR2        m367(.A(mai_mai_n259_), .B(mai_mai_n256_), .Y(mai_mai_n390_));
  AOI210     m368(.A0(mai_mai_n381_), .A1(mai_mai_n71_), .B0(mai_mai_n136_), .Y(mai_mai_n391_));
  OR2        m369(.A(mai_mai_n391_), .B(x03), .Y(mai_mai_n392_));
  NA2        m370(.A(mai_mai_n337_), .B(mai_mai_n57_), .Y(mai_mai_n393_));
  NO2        m371(.A(mai_mai_n393_), .B(x11), .Y(mai_mai_n394_));
  NO3        m372(.A(mai_mai_n394_), .B(mai_mai_n140_), .C(mai_mai_n28_), .Y(mai_mai_n395_));
  AOI220     m373(.A0(mai_mai_n395_), .A1(mai_mai_n392_), .B0(mai_mai_n390_), .B1(mai_mai_n47_), .Y(mai_mai_n396_));
  NA2        m374(.A(mai_mai_n396_), .B(mai_mai_n98_), .Y(mai_mai_n397_));
  AOI210     m375(.A0(mai_mai_n327_), .A1(mai_mai_n105_), .B0(mai_mai_n255_), .Y(mai_mai_n398_));
  NOi21      m376(.An(mai_mai_n309_), .B(mai_mai_n129_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n399_), .B(mai_mai_n256_), .Y(mai_mai_n400_));
  OAI210     m378(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n401_));
  AOI210     m379(.A0(mai_mai_n241_), .A1(mai_mai_n47_), .B0(mai_mai_n401_), .Y(mai_mai_n402_));
  NO4        m380(.A(mai_mai_n402_), .B(mai_mai_n400_), .C(mai_mai_n398_), .D(x08), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n127_), .B(mai_mai_n28_), .Y(mai_mai_n404_));
  NO2        m382(.A(mai_mai_n404_), .B(mai_mai_n260_), .Y(mai_mai_n405_));
  NA3        m383(.A(mai_mai_n321_), .B(mai_mai_n120_), .C(x12), .Y(mai_mai_n406_));
  AO210      m384(.A0(mai_mai_n321_), .A1(mai_mai_n120_), .B0(mai_mai_n241_), .Y(mai_mai_n407_));
  NA3        m385(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(x08), .Y(mai_mai_n408_));
  INV        m386(.A(mai_mai_n408_), .Y(mai_mai_n409_));
  AOI210     m387(.A0(mai_mai_n403_), .A1(mai_mai_n397_), .B0(mai_mai_n409_), .Y(mai_mai_n410_));
  OAI210     m388(.A0(mai_mai_n393_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n429_), .B(mai_mai_n370_), .Y(mai_mai_n412_));
  OAI210     m390(.A0(mai_mai_n412_), .A1(mai_mai_n411_), .B0(mai_mai_n181_), .Y(mai_mai_n413_));
  NA3        m391(.A(mai_mai_n405_), .B(mai_mai_n399_), .C(mai_mai_n317_), .Y(mai_mai_n414_));
  INV        m392(.A(x14), .Y(mai_mai_n415_));
  NO3        m393(.A(mai_mai_n309_), .B(mai_mai_n100_), .C(x11), .Y(mai_mai_n416_));
  NO3        m394(.A(mai_mai_n160_), .B(mai_mai_n71_), .C(mai_mai_n53_), .Y(mai_mai_n417_));
  NO3        m395(.A(mai_mai_n389_), .B(mai_mai_n318_), .C(mai_mai_n175_), .Y(mai_mai_n418_));
  NO4        m396(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(mai_mai_n416_), .D(mai_mai_n415_), .Y(mai_mai_n419_));
  NA3        m397(.A(mai_mai_n419_), .B(mai_mai_n414_), .C(mai_mai_n413_), .Y(mai_mai_n420_));
  AOI220     m398(.A0(mai_mai_n386_), .A1(mai_mai_n57_), .B0(mai_mai_n404_), .B1(mai_mai_n159_), .Y(mai_mai_n421_));
  NOi21      m399(.An(mai_mai_n265_), .B(mai_mai_n144_), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n423_));
  OAI210     m401(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n97_), .Y(mai_mai_n424_));
  OAI210     m402(.A0(mai_mai_n421_), .A1(mai_mai_n87_), .B0(mai_mai_n424_), .Y(mai_mai_n425_));
  NO4        m403(.A(mai_mai_n425_), .B(mai_mai_n420_), .C(mai_mai_n410_), .D(mai_mai_n388_), .Y(mai06));
  INV        m404(.A(x07), .Y(mai_mai_n429_));
  INV        m405(.A(x01), .Y(mai_mai_n430_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  INV        u039(.A(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  NO2        u042(.A(men_men_n64_), .B(men_men_n62_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  NA3        u050(.A(men_men_n72_), .B(men_men_n71_), .C(men_men_n28_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n73_), .A1(x11), .B0(x03), .Y(men_men_n74_));
  NOi31      u052(.An(x08), .B(x04), .C(x00), .Y(men_men_n75_));
  NO2        u053(.A(x10), .B(x09), .Y(men_men_n76_));
  NO2        u054(.A(men_men_n445_), .B(men_men_n24_), .Y(men_men_n77_));
  NO2        u055(.A(x09), .B(men_men_n41_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n78_), .B(men_men_n36_), .Y(men_men_n79_));
  OAI210     u057(.A0(men_men_n78_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n80_));
  AOI210     u058(.A0(men_men_n79_), .A1(men_men_n48_), .B0(men_men_n80_), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n36_), .B(x00), .Y(men_men_n82_));
  NO2        u060(.A(x08), .B(x01), .Y(men_men_n83_));
  OAI210     u061(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n35_), .Y(men_men_n84_));
  NA2        u062(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n85_));
  NO3        u063(.A(men_men_n84_), .B(men_men_n81_), .C(men_men_n77_), .Y(men_men_n86_));
  AN2        u064(.A(men_men_n86_), .B(men_men_n74_), .Y(men_men_n87_));
  INV        u065(.A(men_men_n84_), .Y(men_men_n88_));
  NA2        u066(.A(x11), .B(x00), .Y(men_men_n89_));
  NO2        u067(.A(x11), .B(men_men_n47_), .Y(men_men_n90_));
  NOi21      u068(.An(men_men_n89_), .B(men_men_n90_), .Y(men_men_n91_));
  NOi21      u069(.An(x01), .B(x10), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n93_));
  NO3        u071(.A(men_men_n93_), .B(men_men_n92_), .C(x06), .Y(men_men_n94_));
  NA2        u072(.A(men_men_n94_), .B(men_men_n27_), .Y(men_men_n95_));
  OAI210     u073(.A0(men_men_n446_), .A1(x07), .B0(men_men_n95_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n87_), .C(men_men_n69_), .Y(men01));
  INV        u075(.A(x12), .Y(men_men_n98_));
  INV        u076(.A(x13), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n449_), .B(men_men_n70_), .Y(men_men_n100_));
  NA2        u078(.A(x08), .B(x04), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n101_), .B(men_men_n57_), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n102_), .B(men_men_n100_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n92_), .B(men_men_n28_), .Y(men_men_n104_));
  NO2        u082(.A(x10), .B(x01), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n29_), .B(x00), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NA2        u085(.A(x04), .B(men_men_n28_), .Y(men_men_n108_));
  NO3        u086(.A(men_men_n108_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n109_));
  NA2        u087(.A(men_men_n109_), .B(men_men_n107_), .Y(men_men_n110_));
  AOI210     u088(.A0(men_men_n110_), .A1(men_men_n103_), .B0(men_men_n99_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n56_), .B(x05), .Y(men_men_n112_));
  NOi21      u090(.An(men_men_n112_), .B(men_men_n58_), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n99_), .B(men_men_n36_), .Y(men_men_n114_));
  NA3        u092(.A(men_men_n114_), .B(men_men_n450_), .C(x06), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n115_), .B(men_men_n113_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n83_), .B(x13), .Y(men_men_n117_));
  NA2        u095(.A(x09), .B(men_men_n35_), .Y(men_men_n118_));
  NA2        u096(.A(x13), .B(men_men_n35_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(x05), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n121_));
  NO2        u099(.A(x00), .B(men_men_n72_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n123_));
  NA2        u101(.A(x10), .B(men_men_n57_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n51_), .B(x05), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n126_), .B(x13), .Y(men_men_n127_));
  NO3        u105(.A(men_men_n121_), .B(men_men_n78_), .C(men_men_n36_), .Y(men_men_n128_));
  NO2        u106(.A(men_men_n60_), .B(x05), .Y(men_men_n129_));
  NOi41      u107(.An(men_men_n127_), .B(men_men_n129_), .C(men_men_n128_), .D(men_men_n125_), .Y(men_men_n130_));
  NO3        u108(.A(men_men_n130_), .B(x06), .C(x03), .Y(men_men_n131_));
  NO4        u109(.A(men_men_n131_), .B(men_men_n122_), .C(men_men_n116_), .D(men_men_n111_), .Y(men_men_n132_));
  NA2        u110(.A(x13), .B(men_men_n36_), .Y(men_men_n133_));
  OAI210     u111(.A0(men_men_n83_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n134_));
  NA2        u112(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NO2        u113(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n136_));
  OA210      u114(.A0(x00), .A1(men_men_n76_), .B0(men_men_n136_), .Y(men_men_n137_));
  NO2        u115(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n29_), .B(x06), .Y(men_men_n139_));
  AOI210     u117(.A0(men_men_n139_), .A1(men_men_n49_), .B0(men_men_n138_), .Y(men_men_n140_));
  OA210      u118(.A0(men_men_n140_), .A1(men_men_n137_), .B0(men_men_n135_), .Y(men_men_n141_));
  NO2        u119(.A(x09), .B(x05), .Y(men_men_n142_));
  NA2        u120(.A(men_men_n142_), .B(men_men_n47_), .Y(men_men_n143_));
  AOI210     u121(.A0(men_men_n143_), .A1(men_men_n107_), .B0(men_men_n49_), .Y(men_men_n144_));
  NA2        u122(.A(x09), .B(x00), .Y(men_men_n145_));
  NA2        u123(.A(men_men_n112_), .B(men_men_n145_), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n75_), .B(men_men_n51_), .Y(men_men_n147_));
  AOI210     u125(.A0(men_men_n147_), .A1(men_men_n146_), .B0(men_men_n139_), .Y(men_men_n148_));
  NO3        u126(.A(men_men_n148_), .B(men_men_n144_), .C(men_men_n141_), .Y(men_men_n149_));
  NO2        u127(.A(x03), .B(x02), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n84_), .B(men_men_n99_), .Y(men_men_n151_));
  OAI210     u129(.A0(men_men_n151_), .A1(men_men_n113_), .B0(men_men_n150_), .Y(men_men_n152_));
  OA210      u130(.A0(men_men_n149_), .A1(x11), .B0(men_men_n152_), .Y(men_men_n153_));
  OAI210     u131(.A0(men_men_n132_), .A1(men_men_n23_), .B0(men_men_n153_), .Y(men_men_n154_));
  NA2        u132(.A(men_men_n107_), .B(men_men_n40_), .Y(men_men_n155_));
  NAi21      u133(.An(x06), .B(x10), .Y(men_men_n156_));
  NOi21      u134(.An(x01), .B(x13), .Y(men_men_n157_));
  NA2        u135(.A(men_men_n157_), .B(men_men_n156_), .Y(men_men_n158_));
  OR2        u136(.A(men_men_n158_), .B(x08), .Y(men_men_n159_));
  AOI210     u137(.A0(men_men_n159_), .A1(men_men_n155_), .B0(men_men_n41_), .Y(men_men_n160_));
  NO2        u138(.A(men_men_n29_), .B(x03), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n99_), .B(x01), .Y(men_men_n162_));
  NO2        u140(.A(men_men_n162_), .B(x08), .Y(men_men_n163_));
  OAI210     u141(.A0(x05), .A1(men_men_n163_), .B0(men_men_n51_), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n161_), .B0(men_men_n48_), .Y(men_men_n165_));
  AOI210     u143(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n166_));
  OAI210     u144(.A0(men_men_n165_), .A1(men_men_n160_), .B0(men_men_n166_), .Y(men_men_n167_));
  NA2        u145(.A(x04), .B(x02), .Y(men_men_n168_));
  NA2        u146(.A(x10), .B(x05), .Y(men_men_n169_));
  NO2        u147(.A(x09), .B(x01), .Y(men_men_n170_));
  NO2        u148(.A(men_men_n105_), .B(men_men_n31_), .Y(men_men_n171_));
  NA2        u149(.A(men_men_n171_), .B(x00), .Y(men_men_n172_));
  NO2        u150(.A(men_men_n112_), .B(x08), .Y(men_men_n173_));
  NA3        u151(.A(men_men_n157_), .B(men_men_n156_), .C(men_men_n51_), .Y(men_men_n174_));
  NA2        u152(.A(men_men_n92_), .B(x05), .Y(men_men_n175_));
  OAI210     u153(.A0(men_men_n175_), .A1(men_men_n114_), .B0(men_men_n174_), .Y(men_men_n176_));
  AOI210     u154(.A0(men_men_n173_), .A1(x06), .B0(men_men_n176_), .Y(men_men_n177_));
  OAI210     u155(.A0(men_men_n177_), .A1(x11), .B0(men_men_n172_), .Y(men_men_n178_));
  NAi21      u156(.An(men_men_n168_), .B(men_men_n178_), .Y(men_men_n179_));
  INV        u157(.A(men_men_n25_), .Y(men_men_n180_));
  NAi21      u158(.An(x13), .B(x00), .Y(men_men_n181_));
  AOI210     u159(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n181_), .Y(men_men_n182_));
  AOI220     u160(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n169_), .A1(men_men_n35_), .B0(men_men_n183_), .Y(men_men_n184_));
  BUFFER     u162(.A(men_men_n182_), .Y(men_men_n185_));
  BUFFER     u163(.A(men_men_n71_), .Y(men_men_n186_));
  NO2        u164(.A(men_men_n181_), .B(men_men_n36_), .Y(men_men_n187_));
  INV        u165(.A(men_men_n187_), .Y(men_men_n188_));
  NO2        u166(.A(men_men_n57_), .B(men_men_n186_), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n185_), .B0(men_men_n180_), .Y(men_men_n190_));
  NOi21      u168(.An(x09), .B(x00), .Y(men_men_n191_));
  NO3        u169(.A(men_men_n82_), .B(men_men_n191_), .C(men_men_n47_), .Y(men_men_n192_));
  NA2        u170(.A(men_men_n192_), .B(men_men_n124_), .Y(men_men_n193_));
  NA2        u171(.A(x06), .B(x05), .Y(men_men_n194_));
  OAI210     u172(.A0(men_men_n194_), .A1(men_men_n35_), .B0(men_men_n98_), .Y(men_men_n195_));
  AOI210     u173(.A0(x10), .A1(men_men_n58_), .B0(men_men_n195_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n196_), .B(men_men_n193_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n99_), .B(x12), .Y(men_men_n198_));
  AOI210     u176(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n198_), .Y(men_men_n199_));
  NA2        u177(.A(men_men_n92_), .B(men_men_n51_), .Y(men_men_n200_));
  NO2        u178(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n201_));
  NA2        u179(.A(men_men_n201_), .B(x02), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n202_), .B(men_men_n200_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n199_), .A1(men_men_n197_), .B0(men_men_n203_), .Y(men_men_n204_));
  NA4        u182(.A(men_men_n204_), .B(men_men_n190_), .C(men_men_n179_), .D(men_men_n167_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n154_), .A1(men_men_n98_), .B0(men_men_n205_), .Y(men_men_n206_));
  INV        u184(.A(men_men_n73_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(men_men_n135_), .Y(men_men_n208_));
  NA2        u186(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n209_), .B(men_men_n134_), .Y(men_men_n210_));
  NO2        u188(.A(men_men_n123_), .B(x06), .Y(men_men_n211_));
  INV        u189(.A(men_men_n211_), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n212_), .A1(men_men_n208_), .B0(x12), .Y(men_men_n213_));
  INV        u191(.A(men_men_n75_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n92_), .B(x06), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n215_), .B(men_men_n41_), .Y(men_men_n216_));
  NA4        u194(.A(men_men_n156_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n139_), .Y(men_men_n218_));
  OAI210     u196(.A0(men_men_n218_), .A1(men_men_n216_), .B0(x02), .Y(men_men_n219_));
  AOI210     u197(.A0(men_men_n219_), .A1(men_men_n57_), .B0(men_men_n23_), .Y(men_men_n220_));
  OAI210     u198(.A0(men_men_n213_), .A1(men_men_n57_), .B0(men_men_n220_), .Y(men_men_n221_));
  INV        u199(.A(men_men_n139_), .Y(men_men_n222_));
  NO2        u200(.A(men_men_n51_), .B(x03), .Y(men_men_n223_));
  OAI210     u201(.A0(men_men_n78_), .A1(men_men_n36_), .B0(men_men_n118_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n99_), .B(x03), .Y(men_men_n225_));
  AOI220     u203(.A0(men_men_n225_), .A1(men_men_n224_), .B0(men_men_n75_), .B1(men_men_n223_), .Y(men_men_n226_));
  INV        u204(.A(men_men_n156_), .Y(men_men_n227_));
  NOi21      u205(.An(x13), .B(x04), .Y(men_men_n228_));
  NO3        u206(.A(men_men_n228_), .B(men_men_n75_), .C(men_men_n191_), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n229_), .B(x05), .Y(men_men_n230_));
  AOI220     u208(.A0(men_men_n230_), .A1(men_men_n448_), .B0(men_men_n227_), .B1(men_men_n57_), .Y(men_men_n231_));
  OAI210     u209(.A0(men_men_n226_), .A1(men_men_n222_), .B0(men_men_n231_), .Y(men_men_n232_));
  INV        u210(.A(men_men_n90_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n233_), .B(x12), .Y(men_men_n234_));
  NA2        u212(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n236_));
  OAI210     u214(.A0(men_men_n236_), .A1(men_men_n184_), .B0(men_men_n182_), .Y(men_men_n237_));
  AOI210     u215(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n238_));
  NA2        u216(.A(men_men_n145_), .B(men_men_n72_), .Y(men_men_n239_));
  INV        u217(.A(men_men_n239_), .Y(men_men_n240_));
  NA2        u218(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n241_));
  NA2        u219(.A(men_men_n241_), .B(x03), .Y(men_men_n242_));
  OA210      u220(.A0(men_men_n242_), .A1(men_men_n240_), .B0(men_men_n237_), .Y(men_men_n243_));
  NA2        u221(.A(x13), .B(men_men_n98_), .Y(men_men_n244_));
  NA3        u222(.A(men_men_n244_), .B(men_men_n195_), .C(men_men_n91_), .Y(men_men_n245_));
  OAI210     u223(.A0(men_men_n243_), .A1(men_men_n235_), .B0(men_men_n245_), .Y(men_men_n246_));
  AOI210     u224(.A0(men_men_n234_), .A1(men_men_n232_), .B0(men_men_n246_), .Y(men_men_n247_));
  AOI210     u225(.A0(men_men_n247_), .A1(men_men_n221_), .B0(x07), .Y(men_men_n248_));
  NA2        u226(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n249_));
  AOI210     u227(.A0(men_men_n133_), .A1(men_men_n147_), .B0(men_men_n249_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n99_), .B(x06), .Y(men_men_n251_));
  INV        u229(.A(men_men_n251_), .Y(men_men_n252_));
  NO2        u230(.A(x08), .B(x05), .Y(men_men_n253_));
  NO2        u231(.A(men_men_n253_), .B(men_men_n238_), .Y(men_men_n254_));
  OAI210     u232(.A0(men_men_n75_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n255_));
  OAI210     u233(.A0(men_men_n254_), .A1(men_men_n252_), .B0(men_men_n255_), .Y(men_men_n256_));
  NO2        u234(.A(x12), .B(x02), .Y(men_men_n257_));
  INV        u235(.A(men_men_n257_), .Y(men_men_n258_));
  NO2        u236(.A(men_men_n258_), .B(men_men_n233_), .Y(men_men_n259_));
  OA210      u237(.A0(men_men_n256_), .A1(men_men_n250_), .B0(men_men_n259_), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n261_));
  NO2        u239(.A(men_men_n261_), .B(x01), .Y(men_men_n262_));
  NOi21      u240(.An(men_men_n83_), .B(men_men_n118_), .Y(men_men_n263_));
  NO2        u241(.A(men_men_n263_), .B(men_men_n262_), .Y(men_men_n264_));
  AOI210     u242(.A0(men_men_n264_), .A1(men_men_n127_), .B0(men_men_n29_), .Y(men_men_n265_));
  NA2        u243(.A(men_men_n251_), .B(men_men_n224_), .Y(men_men_n266_));
  NA2        u244(.A(men_men_n99_), .B(x04), .Y(men_men_n267_));
  NA2        u245(.A(men_men_n267_), .B(men_men_n28_), .Y(men_men_n268_));
  OAI210     u246(.A0(men_men_n268_), .A1(men_men_n117_), .B0(men_men_n266_), .Y(men_men_n269_));
  NO3        u247(.A(men_men_n89_), .B(x12), .C(x03), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n269_), .A1(men_men_n265_), .B0(men_men_n270_), .Y(men_men_n271_));
  AOI210     u249(.A0(men_men_n200_), .A1(men_men_n194_), .B0(men_men_n101_), .Y(men_men_n272_));
  NOi21      u250(.An(men_men_n249_), .B(men_men_n215_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n25_), .B(x00), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n274_), .Y(men_men_n275_));
  NO2        u253(.A(men_men_n58_), .B(x05), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n235_), .B(men_men_n28_), .Y(men_men_n277_));
  NA2        u255(.A(men_men_n222_), .B(men_men_n277_), .Y(men_men_n278_));
  NA3        u256(.A(men_men_n278_), .B(men_men_n275_), .C(men_men_n271_), .Y(men_men_n279_));
  NO3        u257(.A(men_men_n279_), .B(men_men_n260_), .C(men_men_n248_), .Y(men_men_n280_));
  OAI210     u258(.A0(men_men_n206_), .A1(men_men_n61_), .B0(men_men_n280_), .Y(men02));
  NOi21      u259(.An(men_men_n229_), .B(men_men_n170_), .Y(men_men_n282_));
  NO2        u260(.A(men_men_n99_), .B(men_men_n35_), .Y(men_men_n283_));
  NA3        u261(.A(men_men_n283_), .B(x10), .C(men_men_n56_), .Y(men_men_n284_));
  OAI210     u262(.A0(men_men_n282_), .A1(men_men_n32_), .B0(men_men_n284_), .Y(men_men_n285_));
  NA2        u263(.A(men_men_n285_), .B(men_men_n169_), .Y(men_men_n286_));
  INV        u264(.A(men_men_n169_), .Y(men_men_n287_));
  NA2        u265(.A(men_men_n450_), .B(men_men_n85_), .Y(men_men_n288_));
  OAI220     u266(.A0(men_men_n288_), .A1(men_men_n99_), .B0(men_men_n84_), .B1(men_men_n51_), .Y(men_men_n289_));
  AOI220     u267(.A0(men_men_n289_), .A1(men_men_n287_), .B0(men_men_n151_), .B1(men_men_n150_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n290_), .A1(men_men_n286_), .B0(men_men_n48_), .Y(men_men_n291_));
  NO2        u269(.A(x05), .B(x02), .Y(men_men_n292_));
  OAI210     u270(.A0(men_men_n210_), .A1(men_men_n191_), .B0(men_men_n292_), .Y(men_men_n293_));
  AOI220     u271(.A0(men_men_n253_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n294_));
  NOi21      u272(.An(men_men_n283_), .B(men_men_n294_), .Y(men_men_n295_));
  AOI210     u273(.A0(men_men_n228_), .A1(men_men_n78_), .B0(men_men_n295_), .Y(men_men_n296_));
  AOI210     u274(.A0(men_men_n296_), .A1(men_men_n293_), .B0(men_men_n139_), .Y(men_men_n297_));
  NAi21      u275(.An(men_men_n230_), .B(men_men_n226_), .Y(men_men_n298_));
  NO2        u276(.A(men_men_n241_), .B(men_men_n47_), .Y(men_men_n299_));
  NA2        u277(.A(men_men_n299_), .B(men_men_n298_), .Y(men_men_n300_));
  AN2        u278(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n302_));
  NA2        u280(.A(x13), .B(men_men_n28_), .Y(men_men_n303_));
  OA210      u281(.A0(men_men_n303_), .A1(x08), .B0(men_men_n143_), .Y(men_men_n304_));
  AOI210     u282(.A0(men_men_n304_), .A1(men_men_n134_), .B0(men_men_n302_), .Y(men_men_n305_));
  OAI210     u283(.A0(men_men_n305_), .A1(men_men_n301_), .B0(men_men_n93_), .Y(men_men_n306_));
  NA3        u284(.A(men_men_n93_), .B(men_men_n83_), .C(men_men_n223_), .Y(men_men_n307_));
  NA3        u285(.A(men_men_n92_), .B(men_men_n82_), .C(men_men_n42_), .Y(men_men_n308_));
  AOI210     u286(.A0(men_men_n308_), .A1(men_men_n307_), .B0(x04), .Y(men_men_n309_));
  INV        u287(.A(men_men_n150_), .Y(men_men_n310_));
  OAI220     u288(.A0(men_men_n254_), .A1(men_men_n104_), .B0(men_men_n310_), .B1(men_men_n125_), .Y(men_men_n311_));
  AOI210     u289(.A0(men_men_n311_), .A1(x13), .B0(men_men_n309_), .Y(men_men_n312_));
  NA3        u290(.A(men_men_n312_), .B(men_men_n306_), .C(men_men_n300_), .Y(men_men_n313_));
  NO3        u291(.A(men_men_n313_), .B(men_men_n297_), .C(men_men_n291_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n138_), .B(x03), .Y(men_men_n315_));
  INV        u293(.A(men_men_n181_), .Y(men_men_n316_));
  AOI220     u294(.A0(x08), .A1(men_men_n316_), .B0(men_men_n201_), .B1(x08), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n317_), .A1(men_men_n276_), .B0(men_men_n315_), .Y(men_men_n318_));
  NA2        u296(.A(men_men_n318_), .B(men_men_n105_), .Y(men_men_n319_));
  NA2        u297(.A(men_men_n168_), .B(men_men_n162_), .Y(men_men_n320_));
  AN2        u298(.A(men_men_n320_), .B(men_men_n173_), .Y(men_men_n321_));
  NO2        u299(.A(men_men_n126_), .B(men_men_n28_), .Y(men_men_n322_));
  OAI210     u300(.A0(men_men_n322_), .A1(men_men_n321_), .B0(men_men_n106_), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n267_), .B(men_men_n98_), .Y(men_men_n324_));
  NA2        u302(.A(men_men_n98_), .B(men_men_n41_), .Y(men_men_n325_));
  NA3        u303(.A(men_men_n325_), .B(men_men_n324_), .C(men_men_n125_), .Y(men_men_n326_));
  NA4        u304(.A(men_men_n326_), .B(men_men_n323_), .C(men_men_n319_), .D(men_men_n48_), .Y(men_men_n327_));
  INV        u305(.A(men_men_n201_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n32_), .B(x05), .Y(men_men_n329_));
  OAI220     u307(.A0(men_men_n329_), .A1(men_men_n447_), .B0(men_men_n328_), .B1(men_men_n59_), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(x02), .Y(men_men_n331_));
  INV        u309(.A(men_men_n236_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n198_), .B(x04), .Y(men_men_n333_));
  NO2        u311(.A(men_men_n333_), .B(men_men_n332_), .Y(men_men_n334_));
  NO3        u312(.A(men_men_n183_), .B(x13), .C(men_men_n31_), .Y(men_men_n335_));
  OAI210     u313(.A0(men_men_n335_), .A1(men_men_n334_), .B0(men_men_n93_), .Y(men_men_n336_));
  NO3        u314(.A(men_men_n198_), .B(men_men_n161_), .C(men_men_n52_), .Y(men_men_n337_));
  OAI210     u315(.A0(men_men_n145_), .A1(men_men_n36_), .B0(men_men_n98_), .Y(men_men_n338_));
  OAI210     u316(.A0(men_men_n338_), .A1(men_men_n192_), .B0(men_men_n337_), .Y(men_men_n339_));
  NA4        u317(.A(men_men_n339_), .B(men_men_n336_), .C(men_men_n331_), .D(x06), .Y(men_men_n340_));
  NA2        u318(.A(x09), .B(x03), .Y(men_men_n341_));
  OAI220     u319(.A0(men_men_n341_), .A1(men_men_n124_), .B0(men_men_n209_), .B1(men_men_n63_), .Y(men_men_n342_));
  OAI220     u320(.A0(men_men_n162_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n343_));
  NO3        u321(.A(men_men_n276_), .B(men_men_n123_), .C(x08), .Y(men_men_n344_));
  AOI210     u322(.A0(men_men_n343_), .A1(men_men_n222_), .B0(men_men_n344_), .Y(men_men_n345_));
  NO2        u323(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n346_));
  NO3        u324(.A(men_men_n112_), .B(men_men_n124_), .C(men_men_n38_), .Y(men_men_n347_));
  AOI210     u325(.A0(men_men_n337_), .A1(men_men_n346_), .B0(men_men_n347_), .Y(men_men_n348_));
  OAI210     u326(.A0(men_men_n345_), .A1(men_men_n28_), .B0(men_men_n348_), .Y(men_men_n349_));
  AO220      u327(.A0(men_men_n349_), .A1(x04), .B0(men_men_n342_), .B1(x05), .Y(men_men_n350_));
  AOI210     u328(.A0(men_men_n340_), .A1(men_men_n327_), .B0(men_men_n350_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n314_), .A1(x12), .B0(men_men_n351_), .Y(men03));
  OR2        u330(.A(men_men_n42_), .B(men_men_n223_), .Y(men_men_n353_));
  AOI210     u331(.A0(men_men_n151_), .A1(men_men_n98_), .B0(men_men_n353_), .Y(men_men_n354_));
  AO210      u332(.A0(men_men_n332_), .A1(men_men_n85_), .B0(men_men_n333_), .Y(men_men_n355_));
  NA2        u333(.A(men_men_n198_), .B(men_men_n150_), .Y(men_men_n356_));
  NA3        u334(.A(men_men_n356_), .B(men_men_n355_), .C(men_men_n202_), .Y(men_men_n357_));
  OAI210     u335(.A0(men_men_n357_), .A1(men_men_n354_), .B0(x05), .Y(men_men_n358_));
  NA2        u336(.A(men_men_n353_), .B(x05), .Y(men_men_n359_));
  AOI210     u337(.A0(men_men_n134_), .A1(men_men_n214_), .B0(men_men_n359_), .Y(men_men_n360_));
  AOI210     u338(.A0(men_men_n225_), .A1(men_men_n79_), .B0(men_men_n120_), .Y(men_men_n361_));
  OAI220     u339(.A0(men_men_n361_), .A1(men_men_n59_), .B0(men_men_n303_), .B1(men_men_n294_), .Y(men_men_n362_));
  OAI210     u340(.A0(men_men_n362_), .A1(men_men_n360_), .B0(men_men_n98_), .Y(men_men_n363_));
  AOI210     u341(.A0(men_men_n143_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n364_));
  NO2        u342(.A(men_men_n170_), .B(men_men_n129_), .Y(men_men_n365_));
  OAI220     u343(.A0(men_men_n365_), .A1(men_men_n37_), .B0(men_men_n146_), .B1(x13), .Y(men_men_n366_));
  OAI210     u344(.A0(men_men_n366_), .A1(men_men_n364_), .B0(x04), .Y(men_men_n367_));
  NO3        u345(.A(men_men_n325_), .B(men_men_n84_), .C(men_men_n59_), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n188_), .A1(men_men_n98_), .B0(men_men_n143_), .Y(men_men_n369_));
  OA210      u347(.A0(men_men_n163_), .A1(x12), .B0(men_men_n129_), .Y(men_men_n370_));
  NO3        u348(.A(men_men_n370_), .B(men_men_n369_), .C(men_men_n368_), .Y(men_men_n371_));
  NA4        u349(.A(men_men_n371_), .B(men_men_n367_), .C(men_men_n363_), .D(men_men_n358_), .Y(men04));
  NO2        u350(.A(men_men_n88_), .B(men_men_n39_), .Y(men_men_n373_));
  XO2        u351(.A(men_men_n373_), .B(men_men_n244_), .Y(men05));
  NO2        u352(.A(men_men_n302_), .B(men_men_n25_), .Y(men_men_n375_));
  NAi31      u353(.An(men_men_n76_), .B(men_men_n126_), .C(men_men_n31_), .Y(men_men_n376_));
  AOI210     u354(.A0(x05), .A1(men_men_n376_), .B0(men_men_n24_), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n377_), .A1(men_men_n375_), .B0(men_men_n98_), .Y(men_men_n378_));
  NA2        u356(.A(x11), .B(men_men_n31_), .Y(men_men_n379_));
  NA2        u357(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n380_));
  NA2        u358(.A(men_men_n249_), .B(x03), .Y(men_men_n381_));
  OAI220     u359(.A0(men_men_n381_), .A1(men_men_n380_), .B0(men_men_n379_), .B1(men_men_n80_), .Y(men_men_n382_));
  OAI210     u360(.A0(men_men_n26_), .A1(men_men_n98_), .B0(x07), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n382_), .A1(x06), .B0(men_men_n383_), .Y(men_men_n384_));
  NA2        u362(.A(men_men_n80_), .B(men_men_n31_), .Y(men_men_n385_));
  NO3        u363(.A(men_men_n385_), .B(men_men_n23_), .C(x00), .Y(men_men_n386_));
  NA2        u364(.A(men_men_n70_), .B(x02), .Y(men_men_n387_));
  AOI210     u365(.A0(men_men_n387_), .A1(men_men_n381_), .B0(men_men_n251_), .Y(men_men_n388_));
  OR2        u366(.A(men_men_n388_), .B(men_men_n235_), .Y(men_men_n389_));
  NO2        u367(.A(men_men_n23_), .B(x10), .Y(men_men_n390_));
  OAI210     u368(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n391_));
  OR3        u369(.A(men_men_n391_), .B(men_men_n390_), .C(men_men_n44_), .Y(men_men_n392_));
  NA2        u370(.A(men_men_n392_), .B(men_men_n389_), .Y(men_men_n393_));
  OAI210     u371(.A0(men_men_n393_), .A1(men_men_n386_), .B0(men_men_n98_), .Y(men_men_n394_));
  NA2        u372(.A(men_men_n33_), .B(men_men_n98_), .Y(men_men_n395_));
  AOI210     u373(.A0(men_men_n395_), .A1(men_men_n90_), .B0(x07), .Y(men_men_n396_));
  AOI220     u374(.A0(men_men_n396_), .A1(men_men_n394_), .B0(men_men_n384_), .B1(men_men_n378_), .Y(men_men_n397_));
  NA3        u375(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n398_));
  AO210      u376(.A0(men_men_n398_), .A1(men_men_n261_), .B0(men_men_n258_), .Y(men_men_n399_));
  AOI210     u377(.A0(men_men_n390_), .A1(x07), .B0(men_men_n138_), .Y(men_men_n400_));
  OR2        u378(.A(men_men_n400_), .B(x03), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n346_), .B(men_men_n61_), .Y(men_men_n402_));
  NO2        u380(.A(men_men_n402_), .B(x11), .Y(men_men_n403_));
  NO3        u381(.A(men_men_n403_), .B(men_men_n142_), .C(men_men_n28_), .Y(men_men_n404_));
  AOI220     u382(.A0(men_men_n404_), .A1(men_men_n401_), .B0(men_men_n399_), .B1(men_men_n47_), .Y(men_men_n405_));
  NO4        u383(.A(men_men_n325_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n406_));
  OAI210     u384(.A0(men_men_n406_), .A1(men_men_n405_), .B0(men_men_n99_), .Y(men_men_n407_));
  AOI210     u385(.A0(men_men_n333_), .A1(men_men_n108_), .B0(men_men_n257_), .Y(men_men_n408_));
  NOi21      u386(.An(men_men_n315_), .B(men_men_n129_), .Y(men_men_n409_));
  NO2        u387(.A(men_men_n409_), .B(men_men_n258_), .Y(men_men_n410_));
  OAI210     u388(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n411_));
  AOI210     u389(.A0(men_men_n244_), .A1(men_men_n47_), .B0(men_men_n411_), .Y(men_men_n412_));
  NO4        u390(.A(men_men_n412_), .B(men_men_n410_), .C(men_men_n408_), .D(x08), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n390_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n414_));
  OAI220     u392(.A0(x05), .A1(men_men_n414_), .B0(men_men_n379_), .B1(men_men_n66_), .Y(men_men_n415_));
  NO2        u393(.A(x13), .B(x12), .Y(men_men_n416_));
  NO2        u394(.A(men_men_n126_), .B(men_men_n28_), .Y(men_men_n417_));
  NO2        u395(.A(men_men_n417_), .B(men_men_n262_), .Y(men_men_n418_));
  OR3        u396(.A(men_men_n418_), .B(x12), .C(x03), .Y(men_men_n419_));
  NA3        u397(.A(men_men_n328_), .B(men_men_n121_), .C(x12), .Y(men_men_n420_));
  AO210      u398(.A0(men_men_n328_), .A1(men_men_n121_), .B0(men_men_n244_), .Y(men_men_n421_));
  NA4        u399(.A(men_men_n421_), .B(men_men_n420_), .C(men_men_n419_), .D(x08), .Y(men_men_n422_));
  AOI210     u400(.A0(men_men_n416_), .A1(men_men_n415_), .B0(men_men_n422_), .Y(men_men_n423_));
  AOI210     u401(.A0(men_men_n413_), .A1(men_men_n407_), .B0(men_men_n423_), .Y(men_men_n424_));
  OAI210     u402(.A0(men_men_n402_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n425_));
  NA2        u403(.A(men_men_n287_), .B(x07), .Y(men_men_n426_));
  OAI220     u404(.A0(men_men_n426_), .A1(men_men_n380_), .B0(men_men_n142_), .B1(men_men_n43_), .Y(men_men_n427_));
  OAI210     u405(.A0(men_men_n427_), .A1(men_men_n425_), .B0(men_men_n187_), .Y(men_men_n428_));
  NA3        u406(.A(men_men_n418_), .B(men_men_n409_), .C(men_men_n324_), .Y(men_men_n429_));
  INV        u407(.A(x14), .Y(men_men_n430_));
  NO3        u408(.A(men_men_n315_), .B(men_men_n104_), .C(x11), .Y(men_men_n431_));
  NO3        u409(.A(men_men_n398_), .B(men_men_n325_), .C(men_men_n181_), .Y(men_men_n432_));
  NO3        u410(.A(men_men_n432_), .B(men_men_n431_), .C(men_men_n430_), .Y(men_men_n433_));
  NA3        u411(.A(men_men_n433_), .B(men_men_n429_), .C(men_men_n428_), .Y(men_men_n434_));
  AOI220     u412(.A0(men_men_n395_), .A1(men_men_n61_), .B0(men_men_n417_), .B1(men_men_n161_), .Y(men_men_n435_));
  NOi21      u413(.An(men_men_n267_), .B(men_men_n146_), .Y(men_men_n436_));
  NO3        u414(.A(men_men_n123_), .B(men_men_n24_), .C(x06), .Y(men_men_n437_));
  AOI210     u415(.A0(men_men_n274_), .A1(men_men_n227_), .B0(men_men_n437_), .Y(men_men_n438_));
  OAI210     u416(.A0(men_men_n44_), .A1(x04), .B0(men_men_n438_), .Y(men_men_n439_));
  OAI210     u417(.A0(men_men_n439_), .A1(men_men_n436_), .B0(men_men_n98_), .Y(men_men_n440_));
  OAI210     u418(.A0(men_men_n435_), .A1(men_men_n89_), .B0(men_men_n440_), .Y(men_men_n441_));
  NO4        u419(.A(men_men_n441_), .B(men_men_n434_), .C(men_men_n424_), .D(men_men_n397_), .Y(men06));
  INV        u420(.A(x07), .Y(men_men_n445_));
  INV        u421(.A(men_men_n91_), .Y(men_men_n446_));
  INV        u422(.A(men_men_n40_), .Y(men_men_n447_));
  INV        u423(.A(x06), .Y(men_men_n448_));
  INV        u424(.A(x01), .Y(men_men_n449_));
  INV        u425(.A(x02), .Y(men_men_n450_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule