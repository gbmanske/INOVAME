//Benchmark atmr_max1024_476_0.5

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n475_, men_men_n476_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  INV        o003(.A(ori_ori_n19_), .Y(ori_ori_n20_));
  NA2        o004(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n21_));
  INV        o005(.A(x5), .Y(ori_ori_n22_));
  INV        o006(.A(ori_ori_n21_), .Y(ori_ori_n23_));
  NO2        o007(.A(x4), .B(x3), .Y(ori_ori_n24_));
  INV        o008(.A(ori_ori_n24_), .Y(ori_ori_n25_));
  NOi21      o009(.An(ori_ori_n20_), .B(ori_ori_n23_), .Y(ori00));
  NO2        o010(.A(x1), .B(x0), .Y(ori_ori_n27_));
  INV        o011(.A(x6), .Y(ori_ori_n28_));
  NA2        o012(.A(x4), .B(x3), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n20_), .B(ori_ori_n29_), .Y(ori_ori_n30_));
  NO2        o014(.A(x2), .B(x0), .Y(ori_ori_n31_));
  INV        o015(.A(x3), .Y(ori_ori_n32_));
  NO2        o016(.A(ori_ori_n32_), .B(ori_ori_n18_), .Y(ori_ori_n33_));
  INV        o017(.A(ori_ori_n33_), .Y(ori_ori_n34_));
  INV        o018(.A(x4), .Y(ori_ori_n35_));
  INV        o019(.A(ori_ori_n27_), .Y(ori_ori_n36_));
  INV        o020(.A(x2), .Y(ori_ori_n37_));
  NO2        o021(.A(ori_ori_n37_), .B(ori_ori_n17_), .Y(ori_ori_n38_));
  NA2        o022(.A(ori_ori_n32_), .B(ori_ori_n18_), .Y(ori_ori_n39_));
  NA2        o023(.A(ori_ori_n39_), .B(ori_ori_n38_), .Y(ori_ori_n40_));
  OAI210     o024(.A0(ori_ori_n36_), .A1(ori_ori_n25_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO3        o025(.A(ori_ori_n41_), .B(ori_ori_n31_), .C(ori_ori_n30_), .Y(ori01));
  NA2        o026(.A(ori_ori_n32_), .B(x1), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(x5), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n33_), .A1(ori_ori_n22_), .B0(ori_ori_n37_), .Y(ori_ori_n45_));
  NA2        o029(.A(ori_ori_n39_), .B(ori_ori_n45_), .Y(ori_ori_n46_));
  INV        o030(.A(ori_ori_n46_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(x4), .Y(ori_ori_n48_));
  NA2        o032(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n49_));
  OAI210     o033(.A0(ori_ori_n49_), .A1(ori_ori_n39_), .B0(x0), .Y(ori_ori_n50_));
  INV        o034(.A(x6), .Y(ori_ori_n51_));
  NAi21      o035(.An(x4), .B(x3), .Y(ori_ori_n52_));
  NO2        o036(.A(x4), .B(x2), .Y(ori_ori_n53_));
  NO2        o037(.A(ori_ori_n52_), .B(ori_ori_n18_), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n50_), .Y(ori_ori_n55_));
  NA2        o039(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NO2        o040(.A(ori_ori_n56_), .B(ori_ori_n22_), .Y(ori_ori_n57_));
  AOI210     o041(.A0(ori_ori_n39_), .A1(ori_ori_n22_), .B0(ori_ori_n37_), .Y(ori_ori_n58_));
  NA2        o042(.A(ori_ori_n34_), .B(ori_ori_n35_), .Y(ori_ori_n59_));
  NO2        o043(.A(ori_ori_n59_), .B(ori_ori_n58_), .Y(ori_ori_n60_));
  NA2        o044(.A(x4), .B(ori_ori_n32_), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n35_), .B(ori_ori_n37_), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n61_), .B(x1), .Y(ori_ori_n63_));
  NA2        o047(.A(ori_ori_n37_), .B(x1), .Y(ori_ori_n64_));
  NO3        o048(.A(x0), .B(ori_ori_n63_), .C(ori_ori_n60_), .Y(ori_ori_n65_));
  AO210      o049(.A0(ori_ori_n55_), .A1(ori_ori_n48_), .B0(ori_ori_n65_), .Y(ori02));
  NO2        o050(.A(x4), .B(x1), .Y(ori_ori_n67_));
  NO2        o051(.A(x5), .B(ori_ori_n35_), .Y(ori_ori_n68_));
  NAi21      o052(.An(x0), .B(x4), .Y(ori_ori_n69_));
  NO2        o053(.A(ori_ori_n53_), .B(ori_ori_n62_), .Y(ori_ori_n70_));
  INV        o054(.A(x0), .Y(ori_ori_n71_));
  NO2        o055(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n72_));
  NO2        o056(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n73_));
  NA2        o057(.A(ori_ori_n22_), .B(ori_ori_n18_), .Y(ori_ori_n74_));
  NA2        o058(.A(ori_ori_n22_), .B(ori_ori_n17_), .Y(ori_ori_n75_));
  NA3        o059(.A(ori_ori_n75_), .B(ori_ori_n74_), .C(ori_ori_n21_), .Y(ori_ori_n76_));
  AN2        o060(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  NA2        o061(.A(x2), .B(x0), .Y(ori_ori_n78_));
  BUFFER     o062(.A(ori_ori_n67_), .Y(ori_ori_n79_));
  NOi21      o063(.An(ori_ori_n79_), .B(ori_ori_n78_), .Y(ori_ori_n80_));
  NO3        o064(.A(ori_ori_n80_), .B(ori_ori_n77_), .C(ori_ori_n73_), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(ori_ori_n32_), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n76_), .B(ori_ori_n49_), .Y(ori_ori_n83_));
  INV        o067(.A(ori_ori_n68_), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n64_), .B(ori_ori_n84_), .Y(ori_ori_n85_));
  NA2        o069(.A(ori_ori_n79_), .B(ori_ori_n31_), .Y(ori_ori_n86_));
  OAI210     o070(.A0(ori_ori_n75_), .A1(ori_ori_n70_), .B0(ori_ori_n86_), .Y(ori_ori_n87_));
  NO3        o071(.A(ori_ori_n87_), .B(ori_ori_n85_), .C(ori_ori_n83_), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n88_), .B(x3), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n89_), .B(ori_ori_n82_), .Y(ori03));
  NO2        o074(.A(x0), .B(x6), .Y(ori_ori_n91_));
  NOi21      o075(.An(ori_ori_n53_), .B(ori_ori_n91_), .Y(ori_ori_n92_));
  INV        o076(.A(ori_ori_n92_), .Y(ori_ori_n93_));
  OR2        o077(.A(ori_ori_n93_), .B(x5), .Y(ori_ori_n94_));
  NA2        o078(.A(ori_ori_n72_), .B(ori_ori_n57_), .Y(ori_ori_n95_));
  NA2        o079(.A(ori_ori_n51_), .B(x4), .Y(ori_ori_n96_));
  INV        o080(.A(ori_ori_n96_), .Y(ori_ori_n97_));
  OAI210     o081(.A0(ori_ori_n44_), .A1(ori_ori_n97_), .B0(x2), .Y(ori_ori_n98_));
  NA3        o082(.A(ori_ori_n98_), .B(ori_ori_n95_), .C(ori_ori_n94_), .Y(ori_ori_n99_));
  INV        o083(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n32_), .B(ori_ori_n17_), .Y(ori_ori_n101_));
  INV        o085(.A(ori_ori_n33_), .Y(ori_ori_n102_));
  NO2        o086(.A(ori_ori_n102_), .B(ori_ori_n84_), .Y(ori_ori_n103_));
  NO2        o087(.A(x4), .B(x2), .Y(ori_ori_n104_));
  NA2        o088(.A(ori_ori_n18_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  AOI220     o089(.A0(ori_ori_n17_), .A1(x3), .B0(ori_ori_n18_), .B1(ori_ori_n24_), .Y(ori_ori_n106_));
  AOI210     o090(.A0(ori_ori_n106_), .A1(ori_ori_n105_), .B0(ori_ori_n22_), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n107_), .B(ori_ori_n103_), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n100_), .B(ori_ori_n108_), .Y(ori04));
  INV        o093(.A(x2), .Y(ori_ori_n110_));
  OAI210     o094(.A0(ori_ori_n101_), .A1(ori_ori_n110_), .B0(ori_ori_n28_), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n37_), .B(x0), .Y(ori_ori_n112_));
  NA2        o096(.A(x6), .B(ori_ori_n112_), .Y(ori_ori_n113_));
  NA2        o097(.A(ori_ori_n113_), .B(ori_ori_n111_), .Y(ori_ori_n114_));
  INV        o098(.A(ori_ori_n114_), .Y(ori_ori_n115_));
  NA3        o099(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n116_));
  INV        o100(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NA2        o101(.A(ori_ori_n117_), .B(x6), .Y(ori_ori_n118_));
  INV        o102(.A(ori_ori_n69_), .Y(ori_ori_n119_));
  NO2        o103(.A(x2), .B(ori_ori_n119_), .Y(ori_ori_n120_));
  AOI210     o104(.A0(ori_ori_n120_), .A1(ori_ori_n25_), .B0(ori_ori_n22_), .Y(ori_ori_n121_));
  NA2        o105(.A(ori_ori_n121_), .B(ori_ori_n28_), .Y(ori_ori_n122_));
  NA2        o106(.A(ori_ori_n122_), .B(ori_ori_n118_), .Y(ori_ori_n123_));
  AOI210     o107(.A0(ori_ori_n115_), .A1(ori_ori_n22_), .B0(ori_ori_n123_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  NAi21      m004(.An(mai_mai_n20_), .B(mai_mai_n19_), .Y(mai_mai_n21_));
  NA2        m005(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n22_));
  INV        m006(.A(x5), .Y(mai_mai_n23_));
  NA2        m007(.A(x7), .B(x6), .Y(mai_mai_n24_));
  NA2        m008(.A(x4), .B(x2), .Y(mai_mai_n25_));
  NO3        m009(.A(mai_mai_n25_), .B(mai_mai_n24_), .C(mai_mai_n23_), .Y(mai_mai_n26_));
  NO2        m010(.A(mai_mai_n26_), .B(mai_mai_n22_), .Y(mai_mai_n27_));
  NO2        m011(.A(x4), .B(x3), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OA210      m013(.A0(mai_mai_n29_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n30_));
  NOi31      m014(.An(mai_mai_n21_), .B(mai_mai_n30_), .C(mai_mai_n27_), .Y(mai00));
  NO2        m015(.A(x1), .B(x0), .Y(mai_mai_n32_));
  INV        m016(.A(x6), .Y(mai_mai_n33_));
  NO2        m017(.A(mai_mai_n33_), .B(mai_mai_n23_), .Y(mai_mai_n34_));
  NA2        m018(.A(mai_mai_n34_), .B(mai_mai_n32_), .Y(mai_mai_n35_));
  NA2        m019(.A(x4), .B(x3), .Y(mai_mai_n36_));
  AOI210     m020(.A0(mai_mai_n35_), .A1(mai_mai_n21_), .B0(mai_mai_n36_), .Y(mai_mai_n37_));
  NO2        m021(.A(x2), .B(x0), .Y(mai_mai_n38_));
  INV        m022(.A(x3), .Y(mai_mai_n39_));
  NO2        m023(.A(mai_mai_n39_), .B(mai_mai_n18_), .Y(mai_mai_n40_));
  INV        m024(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(mai_mai_n34_), .B(x4), .Y(mai_mai_n42_));
  OAI210     m026(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n38_), .Y(mai_mai_n43_));
  INV        m027(.A(x4), .Y(mai_mai_n44_));
  NO2        m028(.A(mai_mai_n44_), .B(mai_mai_n17_), .Y(mai_mai_n45_));
  NA2        m029(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n20_), .B0(mai_mai_n43_), .Y(mai_mai_n47_));
  NA2        m031(.A(x7), .B(mai_mai_n34_), .Y(mai_mai_n48_));
  AOI220     m032(.A0(mai_mai_n48_), .A1(mai_mai_n32_), .B0(mai_mai_n20_), .B1(mai_mai_n19_), .Y(mai_mai_n49_));
  INV        m033(.A(x2), .Y(mai_mai_n50_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n39_), .B(mai_mai_n18_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  OAI210     m037(.A0(mai_mai_n49_), .A1(mai_mai_n29_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  NO3        m038(.A(mai_mai_n54_), .B(mai_mai_n47_), .C(mai_mai_n37_), .Y(mai01));
  NA2        m039(.A(x8), .B(x7), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n39_), .B(x1), .Y(mai_mai_n57_));
  INV        m041(.A(x9), .Y(mai_mai_n58_));
  NO2        m042(.A(mai_mai_n33_), .B(mai_mai_n57_), .Y(mai_mai_n59_));
  NO2        m043(.A(x7), .B(x6), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n61_));
  NO2        m045(.A(x8), .B(x2), .Y(mai_mai_n62_));
  OA210      m046(.A0(mai_mai_n62_), .A1(mai_mai_n61_), .B0(mai_mai_n60_), .Y(mai_mai_n63_));
  OAI210     m047(.A0(mai_mai_n40_), .A1(mai_mai_n23_), .B0(mai_mai_n50_), .Y(mai_mai_n64_));
  OAI210     m048(.A0(mai_mai_n52_), .A1(mai_mai_n20_), .B0(mai_mai_n64_), .Y(mai_mai_n65_));
  NAi31      m049(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(mai_mai_n65_), .B(mai_mai_n63_), .Y(mai_mai_n67_));
  OAI210     m051(.A0(mai_mai_n67_), .A1(mai_mai_n59_), .B0(x4), .Y(mai_mai_n68_));
  NA2        m052(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n69_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n70_));
  NA2        m054(.A(x5), .B(x3), .Y(mai_mai_n71_));
  NO2        m055(.A(x8), .B(x6), .Y(mai_mai_n72_));
  NO2        m056(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n73_));
  NAi21      m057(.An(x4), .B(x3), .Y(mai_mai_n74_));
  INV        m058(.A(mai_mai_n74_), .Y(mai_mai_n75_));
  NO2        m059(.A(mai_mai_n75_), .B(mai_mai_n20_), .Y(mai_mai_n76_));
  NO2        m060(.A(x4), .B(x2), .Y(mai_mai_n77_));
  NO2        m061(.A(mai_mai_n77_), .B(x3), .Y(mai_mai_n78_));
  NO3        m062(.A(mai_mai_n78_), .B(mai_mai_n76_), .C(mai_mai_n18_), .Y(mai_mai_n79_));
  NO3        m063(.A(mai_mai_n79_), .B(mai_mai_n73_), .C(mai_mai_n70_), .Y(mai_mai_n80_));
  NO3        m064(.A(x7), .B(mai_mai_n39_), .C(x1), .Y(mai_mai_n81_));
  INV        m065(.A(x4), .Y(mai_mai_n82_));
  NA2        m066(.A(mai_mai_n81_), .B(mai_mai_n82_), .Y(mai_mai_n83_));
  NA2        m067(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(mai_mai_n23_), .Y(mai_mai_n85_));
  INV        m069(.A(x8), .Y(mai_mai_n86_));
  NO2        m070(.A(x2), .B(mai_mai_n85_), .Y(mai_mai_n87_));
  NO2        m071(.A(mai_mai_n87_), .B(mai_mai_n24_), .Y(mai_mai_n88_));
  AOI210     m072(.A0(mai_mai_n52_), .A1(mai_mai_n23_), .B0(mai_mai_n50_), .Y(mai_mai_n89_));
  OAI210     m073(.A0(mai_mai_n41_), .A1(mai_mai_n34_), .B0(mai_mai_n44_), .Y(mai_mai_n90_));
  NO3        m074(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(mai_mai_n88_), .Y(mai_mai_n91_));
  NA2        m075(.A(x4), .B(mai_mai_n39_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n44_), .B(mai_mai_n50_), .Y(mai_mai_n93_));
  OAI210     m077(.A0(mai_mai_n93_), .A1(mai_mai_n39_), .B0(mai_mai_n18_), .Y(mai_mai_n94_));
  AOI210     m078(.A0(mai_mai_n92_), .A1(mai_mai_n48_), .B0(mai_mai_n94_), .Y(mai_mai_n95_));
  NO2        m079(.A(x3), .B(x2), .Y(mai_mai_n96_));
  NA2        m080(.A(mai_mai_n96_), .B(mai_mai_n23_), .Y(mai_mai_n97_));
  INV        m081(.A(mai_mai_n97_), .Y(mai_mai_n98_));
  NA2        m082(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n99_));
  OAI210     m083(.A0(mai_mai_n99_), .A1(mai_mai_n36_), .B0(mai_mai_n17_), .Y(mai_mai_n100_));
  NO4        m084(.A(mai_mai_n100_), .B(mai_mai_n98_), .C(mai_mai_n95_), .D(mai_mai_n91_), .Y(mai_mai_n101_));
  AO220      m085(.A0(mai_mai_n101_), .A1(mai_mai_n83_), .B0(mai_mai_n80_), .B1(mai_mai_n68_), .Y(mai02));
  NO2        m086(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n103_));
  NA2        m087(.A(mai_mai_n39_), .B(x0), .Y(mai_mai_n104_));
  OAI210     m088(.A0(x4), .A1(x0), .B0(mai_mai_n104_), .Y(mai_mai_n105_));
  AOI220     m089(.A0(mai_mai_n105_), .A1(x1), .B0(mai_mai_n103_), .B1(x4), .Y(mai_mai_n106_));
  NO3        m090(.A(mai_mai_n106_), .B(x7), .C(x5), .Y(mai_mai_n107_));
  NA2        m091(.A(x9), .B(x2), .Y(mai_mai_n108_));
  OR2        m092(.A(x8), .B(x0), .Y(mai_mai_n109_));
  INV        m093(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NAi21      m094(.An(x2), .B(x8), .Y(mai_mai_n111_));
  NO2        m095(.A(x4), .B(x1), .Y(mai_mai_n112_));
  NA3        m096(.A(mai_mai_n112_), .B(x2), .C(mai_mai_n56_), .Y(mai_mai_n113_));
  NOi21      m097(.An(x0), .B(x1), .Y(mai_mai_n114_));
  NOi21      m098(.An(x0), .B(x4), .Y(mai_mai_n115_));
  INV        m099(.A(x8), .Y(mai_mai_n116_));
  NA2        m100(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  AOI210     m101(.A0(mai_mai_n117_), .A1(mai_mai_n113_), .B0(mai_mai_n71_), .Y(mai_mai_n118_));
  NO2        m102(.A(x5), .B(mai_mai_n44_), .Y(mai_mai_n119_));
  NA2        m103(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n120_));
  AOI210     m104(.A0(mai_mai_n120_), .A1(mai_mai_n99_), .B0(mai_mai_n104_), .Y(mai_mai_n121_));
  OAI210     m105(.A0(mai_mai_n121_), .A1(mai_mai_n32_), .B0(mai_mai_n119_), .Y(mai_mai_n122_));
  NAi21      m106(.An(x0), .B(x4), .Y(mai_mai_n123_));
  NO2        m107(.A(mai_mai_n123_), .B(x1), .Y(mai_mai_n124_));
  NO2        m108(.A(x7), .B(x0), .Y(mai_mai_n125_));
  NO2        m109(.A(mai_mai_n77_), .B(mai_mai_n93_), .Y(mai_mai_n126_));
  NO2        m110(.A(mai_mai_n126_), .B(x3), .Y(mai_mai_n127_));
  OAI210     m111(.A0(mai_mai_n125_), .A1(mai_mai_n124_), .B0(mai_mai_n127_), .Y(mai_mai_n128_));
  NO2        m112(.A(x7), .B(mai_mai_n39_), .Y(mai_mai_n129_));
  NA2        m113(.A(x5), .B(x0), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n131_));
  NA2        m115(.A(mai_mai_n131_), .B(mai_mai_n129_), .Y(mai_mai_n132_));
  NA4        m116(.A(mai_mai_n132_), .B(mai_mai_n128_), .C(mai_mai_n122_), .D(mai_mai_n33_), .Y(mai_mai_n133_));
  NO3        m117(.A(mai_mai_n133_), .B(mai_mai_n118_), .C(mai_mai_n107_), .Y(mai_mai_n134_));
  NO3        m118(.A(mai_mai_n71_), .B(mai_mai_n69_), .C(mai_mai_n22_), .Y(mai_mai_n135_));
  AOI220     m119(.A0(mai_mai_n114_), .A1(x4), .B0(mai_mai_n61_), .B1(mai_mai_n17_), .Y(mai_mai_n136_));
  NO2        m120(.A(mai_mai_n136_), .B(mai_mai_n56_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n92_), .B(x5), .Y(mai_mai_n138_));
  NO2        m122(.A(x9), .B(x7), .Y(mai_mai_n139_));
  NOi21      m123(.An(x8), .B(x0), .Y(mai_mai_n140_));
  INV        m124(.A(x7), .Y(mai_mai_n141_));
  AOI220     m125(.A0(x1), .A1(mai_mai_n331_), .B0(mai_mai_n103_), .B1(x7), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n23_), .B(x4), .Y(mai_mai_n143_));
  NO2        m127(.A(mai_mai_n143_), .B(mai_mai_n115_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n144_), .B(mai_mai_n142_), .Y(mai_mai_n145_));
  NA2        m129(.A(x5), .B(x1), .Y(mai_mai_n146_));
  INV        m130(.A(mai_mai_n146_), .Y(mai_mai_n147_));
  AOI210     m131(.A0(mai_mai_n147_), .A1(mai_mai_n115_), .B0(mai_mai_n33_), .Y(mai_mai_n148_));
  NAi21      m132(.An(x2), .B(x7), .Y(mai_mai_n149_));
  NAi31      m133(.An(mai_mai_n71_), .B(x7), .C(mai_mai_n32_), .Y(mai_mai_n150_));
  NA2        m134(.A(mai_mai_n150_), .B(mai_mai_n148_), .Y(mai_mai_n151_));
  NO4        m135(.A(mai_mai_n151_), .B(mai_mai_n145_), .C(mai_mai_n137_), .D(mai_mai_n135_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n152_), .B(mai_mai_n134_), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n130_), .B(mai_mai_n126_), .Y(mai_mai_n154_));
  NA2        m138(.A(mai_mai_n23_), .B(mai_mai_n18_), .Y(mai_mai_n155_));
  NA2        m139(.A(mai_mai_n23_), .B(mai_mai_n17_), .Y(mai_mai_n156_));
  NA3        m140(.A(mai_mai_n156_), .B(mai_mai_n155_), .C(mai_mai_n22_), .Y(mai_mai_n157_));
  AN2        m141(.A(mai_mai_n157_), .B(mai_mai_n131_), .Y(mai_mai_n158_));
  NA2        m142(.A(x8), .B(x0), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n114_), .B(x4), .Y(mai_mai_n160_));
  NA2        m144(.A(mai_mai_n160_), .B(x5), .Y(mai_mai_n161_));
  AOI210     m145(.A0(mai_mai_n159_), .A1(mai_mai_n120_), .B0(mai_mai_n161_), .Y(mai_mai_n162_));
  NA2        m146(.A(x2), .B(x0), .Y(mai_mai_n163_));
  NA2        m147(.A(x4), .B(x1), .Y(mai_mai_n164_));
  NAi21      m148(.An(mai_mai_n112_), .B(mai_mai_n164_), .Y(mai_mai_n165_));
  NOi31      m149(.An(mai_mai_n165_), .B(mai_mai_n143_), .C(mai_mai_n163_), .Y(mai_mai_n166_));
  NO4        m150(.A(mai_mai_n166_), .B(mai_mai_n162_), .C(mai_mai_n158_), .D(mai_mai_n154_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n167_), .B(mai_mai_n39_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n157_), .B(mai_mai_n69_), .Y(mai_mai_n169_));
  INV        m153(.A(mai_mai_n119_), .Y(mai_mai_n170_));
  NO3        m154(.A(mai_mai_n324_), .B(mai_mai_n170_), .C(x7), .Y(mai_mai_n171_));
  NA3        m155(.A(mai_mai_n165_), .B(mai_mai_n170_), .C(mai_mai_n38_), .Y(mai_mai_n172_));
  OAI210     m156(.A0(mai_mai_n156_), .A1(mai_mai_n126_), .B0(mai_mai_n172_), .Y(mai_mai_n173_));
  NO3        m157(.A(mai_mai_n173_), .B(mai_mai_n171_), .C(mai_mai_n169_), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n174_), .B(x3), .Y(mai_mai_n175_));
  NO3        m159(.A(mai_mai_n175_), .B(mai_mai_n168_), .C(mai_mai_n153_), .Y(mai03));
  NO2        m160(.A(mai_mai_n44_), .B(x3), .Y(mai_mai_n177_));
  NO2        m161(.A(x6), .B(mai_mai_n23_), .Y(mai_mai_n178_));
  NA2        m162(.A(x6), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  NA2        m163(.A(x6), .B(mai_mai_n23_), .Y(mai_mai_n180_));
  NA2        m164(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NA2        m166(.A(mai_mai_n180_), .B(mai_mai_n74_), .Y(mai_mai_n183_));
  AOI210     m167(.A0(mai_mai_n23_), .A1(x3), .B0(mai_mai_n163_), .Y(mai_mai_n184_));
  AOI210     m168(.A0(mai_mai_n184_), .A1(mai_mai_n183_), .B0(mai_mai_n182_), .Y(mai_mai_n185_));
  NO2        m169(.A(x5), .B(x1), .Y(mai_mai_n186_));
  NA2        m170(.A(mai_mai_n186_), .B(mai_mai_n17_), .Y(mai_mai_n187_));
  NO2        m171(.A(mai_mai_n181_), .B(mai_mai_n155_), .Y(mai_mai_n188_));
  NA2        m172(.A(mai_mai_n325_), .B(mai_mai_n44_), .Y(mai_mai_n189_));
  NA3        m173(.A(mai_mai_n189_), .B(mai_mai_n185_), .C(mai_mai_n179_), .Y(mai_mai_n190_));
  NA2        m174(.A(mai_mai_n39_), .B(mai_mai_n50_), .Y(mai_mai_n191_));
  NA2        m175(.A(mai_mai_n131_), .B(mai_mai_n85_), .Y(mai_mai_n192_));
  NA2        m176(.A(x6), .B(mai_mai_n44_), .Y(mai_mai_n193_));
  NA2        m177(.A(mai_mai_n178_), .B(mai_mai_n124_), .Y(mai_mai_n194_));
  NA2        m178(.A(mai_mai_n119_), .B(x6), .Y(mai_mai_n195_));
  OAI210     m179(.A0(mai_mai_n86_), .A1(mai_mai_n33_), .B0(mai_mai_n61_), .Y(mai_mai_n196_));
  NA3        m180(.A(mai_mai_n196_), .B(mai_mai_n195_), .C(mai_mai_n194_), .Y(mai_mai_n197_));
  NA2        m181(.A(mai_mai_n197_), .B(x2), .Y(mai_mai_n198_));
  NA3        m182(.A(mai_mai_n198_), .B(mai_mai_n192_), .C(x7), .Y(mai_mai_n199_));
  AOI210     m183(.A0(mai_mai_n190_), .A1(x8), .B0(mai_mai_n199_), .Y(mai_mai_n200_));
  NA3        m184(.A(mai_mai_n23_), .B(x3), .C(x2), .Y(mai_mai_n201_));
  INV        m185(.A(mai_mai_n201_), .Y(mai_mai_n202_));
  NA2        m186(.A(mai_mai_n202_), .B(mai_mai_n112_), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n181_), .B(x6), .Y(mai_mai_n204_));
  NA2        m188(.A(mai_mai_n203_), .B(mai_mai_n141_), .Y(mai_mai_n205_));
  NA2        m189(.A(mai_mai_n178_), .B(mai_mai_n330_), .Y(mai_mai_n206_));
  NO2        m190(.A(mai_mai_n130_), .B(mai_mai_n18_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n44_), .B(mai_mai_n207_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n206_), .Y(mai_mai_n209_));
  NA2        m193(.A(mai_mai_n58_), .B(x2), .Y(mai_mai_n210_));
  INV        m194(.A(mai_mai_n206_), .Y(mai_mai_n211_));
  NO3        m195(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n212_));
  NA2        m196(.A(x6), .B(x2), .Y(mai_mai_n213_));
  NA2        m197(.A(mai_mai_n50_), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  OAI220     m198(.A0(mai_mai_n214_), .A1(mai_mai_n39_), .B0(mai_mai_n160_), .B1(mai_mai_n42_), .Y(mai_mai_n215_));
  OAI210     m199(.A0(mai_mai_n215_), .A1(mai_mai_n211_), .B0(mai_mai_n209_), .Y(mai_mai_n216_));
  NA2        m200(.A(x4), .B(x0), .Y(mai_mai_n217_));
  NA2        m201(.A(mai_mai_n138_), .B(mai_mai_n38_), .Y(mai_mai_n218_));
  AOI210     m202(.A0(mai_mai_n218_), .A1(mai_mai_n216_), .B0(x8), .Y(mai_mai_n219_));
  NA2        m203(.A(x4), .B(mai_mai_n20_), .Y(mai_mai_n220_));
  NO2        m204(.A(mai_mai_n220_), .B(mai_mai_n191_), .Y(mai_mai_n221_));
  NO3        m205(.A(mai_mai_n221_), .B(mai_mai_n219_), .C(mai_mai_n205_), .Y(mai_mai_n222_));
  INV        m206(.A(x1), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n204_), .B(x2), .Y(mai_mai_n224_));
  NA2        m208(.A(x6), .B(mai_mai_n40_), .Y(mai_mai_n225_));
  AOI210     m209(.A0(mai_mai_n225_), .A1(mai_mai_n224_), .B0(mai_mai_n170_), .Y(mai_mai_n226_));
  NA3        m210(.A(mai_mai_n213_), .B(mai_mai_n186_), .C(mai_mai_n36_), .Y(mai_mai_n227_));
  NA2        m211(.A(x3), .B(x2), .Y(mai_mai_n228_));
  AOI220     m212(.A0(mai_mai_n228_), .A1(mai_mai_n191_), .B0(mai_mai_n146_), .B1(mai_mai_n227_), .Y(mai_mai_n229_));
  NA2        m213(.A(x0), .B(mai_mai_n75_), .Y(mai_mai_n230_));
  NO2        m214(.A(mai_mai_n230_), .B(mai_mai_n23_), .Y(mai_mai_n231_));
  NA3        m215(.A(mai_mai_n33_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n232_));
  NA2        m216(.A(mai_mai_n213_), .B(mai_mai_n232_), .Y(mai_mai_n233_));
  INV        m217(.A(mai_mai_n188_), .Y(mai_mai_n234_));
  NA2        m218(.A(mai_mai_n33_), .B(mai_mai_n39_), .Y(mai_mai_n235_));
  OR2        m219(.A(mai_mai_n235_), .B(mai_mai_n217_), .Y(mai_mai_n236_));
  OAI220     m220(.A0(mai_mai_n236_), .A1(mai_mai_n146_), .B0(mai_mai_n193_), .B1(mai_mai_n234_), .Y(mai_mai_n237_));
  AO210      m221(.A0(mai_mai_n233_), .A1(mai_mai_n138_), .B0(mai_mai_n237_), .Y(mai_mai_n238_));
  NO4        m222(.A(mai_mai_n238_), .B(mai_mai_n231_), .C(mai_mai_n229_), .D(mai_mai_n226_), .Y(mai_mai_n239_));
  OAI210     m223(.A0(mai_mai_n222_), .A1(mai_mai_n200_), .B0(mai_mai_n239_), .Y(mai04));
  NA3        m224(.A(x1), .B(mai_mai_n212_), .C(mai_mai_n78_), .Y(mai_mai_n241_));
  NO2        m225(.A(mai_mai_n210_), .B(mai_mai_n84_), .Y(mai_mai_n242_));
  NO2        m226(.A(mai_mai_n242_), .B(mai_mai_n33_), .Y(mai_mai_n243_));
  NA2        m227(.A(mai_mai_n327_), .B(mai_mai_n86_), .Y(mai_mai_n244_));
  NA2        m228(.A(mai_mai_n244_), .B(mai_mai_n243_), .Y(mai_mai_n245_));
  NA2        m229(.A(mai_mai_n245_), .B(x6), .Y(mai_mai_n246_));
  NOi21      m230(.An(mai_mai_n140_), .B(mai_mai_n120_), .Y(mai_mai_n247_));
  OAI210     m231(.A0(mai_mai_n210_), .A1(mai_mai_n232_), .B0(mai_mai_n235_), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n247_), .B(mai_mai_n248_), .Y(mai_mai_n249_));
  NA2        m233(.A(mai_mai_n326_), .B(mai_mai_n249_), .Y(mai_mai_n250_));
  AOI210     m234(.A0(mai_mai_n250_), .A1(x4), .B0(x7), .Y(mai_mai_n251_));
  NOi21      m235(.An(x4), .B(x0), .Y(mai_mai_n252_));
  NO2        m236(.A(x0), .B(mai_mai_n108_), .Y(mai_mai_n253_));
  NA2        m237(.A(mai_mai_n253_), .B(x8), .Y(mai_mai_n254_));
  NO2        m238(.A(mai_mai_n254_), .B(x3), .Y(mai_mai_n255_));
  NO2        m239(.A(mai_mai_n86_), .B(x4), .Y(mai_mai_n256_));
  NA2        m240(.A(mai_mai_n256_), .B(mai_mai_n40_), .Y(mai_mai_n257_));
  NO2        m241(.A(mai_mai_n25_), .B(mai_mai_n22_), .Y(mai_mai_n258_));
  INV        m242(.A(mai_mai_n258_), .Y(mai_mai_n259_));
  NA3        m243(.A(mai_mai_n259_), .B(mai_mai_n257_), .C(x6), .Y(mai_mai_n260_));
  NO2        m244(.A(mai_mai_n140_), .B(mai_mai_n74_), .Y(mai_mai_n261_));
  NO2        m245(.A(mai_mai_n32_), .B(x2), .Y(mai_mai_n262_));
  OAI210     m246(.A0(mai_mai_n329_), .A1(mai_mai_n58_), .B0(mai_mai_n74_), .Y(mai_mai_n263_));
  OAI220     m247(.A0(mai_mai_n263_), .A1(x6), .B0(mai_mai_n260_), .B1(mai_mai_n255_), .Y(mai_mai_n264_));
  INV        m248(.A(mai_mai_n236_), .Y(mai_mai_n265_));
  AOI210     m249(.A0(mai_mai_n265_), .A1(mai_mai_n18_), .B0(mai_mai_n141_), .Y(mai_mai_n266_));
  AO220      m250(.A0(mai_mai_n266_), .A1(mai_mai_n264_), .B0(mai_mai_n251_), .B1(mai_mai_n246_), .Y(mai_mai_n267_));
  NA2        m251(.A(mai_mai_n262_), .B(x6), .Y(mai_mai_n268_));
  NA2        m252(.A(mai_mai_n77_), .B(mai_mai_n268_), .Y(mai_mai_n269_));
  NA3        m253(.A(mai_mai_n269_), .B(mai_mai_n267_), .C(mai_mai_n241_), .Y(mai_mai_n270_));
  NA2        m254(.A(mai_mai_n177_), .B(mai_mai_n141_), .Y(mai_mai_n271_));
  AO210      m255(.A0(mai_mai_n103_), .A1(x4), .B0(mai_mai_n139_), .Y(mai_mai_n272_));
  NA2        m256(.A(x3), .B(x0), .Y(mai_mai_n273_));
  NO2        m257(.A(mai_mai_n273_), .B(x2), .Y(mai_mai_n274_));
  AOI210     m258(.A0(mai_mai_n272_), .A1(mai_mai_n110_), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  AOI210     m259(.A0(mai_mai_n275_), .A1(mai_mai_n271_), .B0(mai_mai_n23_), .Y(mai_mai_n276_));
  NO2        m260(.A(x3), .B(mai_mai_n23_), .Y(mai_mai_n277_));
  AOI210     m261(.A0(mai_mai_n111_), .A1(mai_mai_n109_), .B0(mai_mai_n38_), .Y(mai_mai_n278_));
  NOi21      m262(.An(mai_mai_n278_), .B(mai_mai_n164_), .Y(mai_mai_n279_));
  OAI210     m263(.A0(mai_mai_n279_), .A1(mai_mai_n277_), .B0(mai_mai_n139_), .Y(mai_mai_n280_));
  NAi31      m264(.An(mai_mai_n46_), .B(mai_mai_n223_), .C(x5), .Y(mai_mai_n281_));
  NA2        m265(.A(mai_mai_n281_), .B(mai_mai_n280_), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n282_), .A1(mai_mai_n276_), .B0(x6), .Y(mai_mai_n283_));
  NA2        m267(.A(mai_mai_n177_), .B(mai_mai_n141_), .Y(mai_mai_n284_));
  INV        m268(.A(x1), .Y(mai_mai_n285_));
  OAI210     m269(.A0(mai_mai_n284_), .A1(x8), .B0(mai_mai_n285_), .Y(mai_mai_n286_));
  NAi31      m270(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n287_));
  OAI210     m271(.A0(mai_mai_n287_), .A1(x4), .B0(mai_mai_n149_), .Y(mai_mai_n288_));
  NA2        m272(.A(mai_mai_n288_), .B(x9), .Y(mai_mai_n289_));
  NA2        m273(.A(mai_mai_n261_), .B(mai_mai_n141_), .Y(mai_mai_n290_));
  NA4        m274(.A(mai_mai_n290_), .B(x1), .C(mai_mai_n289_), .D(mai_mai_n46_), .Y(mai_mai_n291_));
  NA2        m275(.A(mai_mai_n286_), .B(mai_mai_n291_), .Y(mai_mai_n292_));
  NOi31      m276(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n293_));
  AOI210     m277(.A0(mai_mai_n115_), .A1(x3), .B0(mai_mai_n252_), .Y(mai_mai_n294_));
  NO2        m278(.A(mai_mai_n56_), .B(mai_mai_n114_), .Y(mai_mai_n295_));
  OAI210     m279(.A0(mai_mai_n295_), .A1(x3), .B0(mai_mai_n294_), .Y(mai_mai_n296_));
  NO3        m280(.A(mai_mai_n296_), .B(x9), .C(x2), .Y(mai_mai_n297_));
  INV        m281(.A(mai_mai_n297_), .Y(mai_mai_n298_));
  AOI210     m282(.A0(mai_mai_n298_), .A1(mai_mai_n292_), .B0(mai_mai_n23_), .Y(mai_mai_n299_));
  AOI220     m283(.A0(x1), .A1(mai_mai_n328_), .B0(mai_mai_n323_), .B1(mai_mai_n278_), .Y(mai_mai_n300_));
  NO2        m284(.A(mai_mai_n300_), .B(mai_mai_n96_), .Y(mai_mai_n301_));
  NO3        m285(.A(mai_mai_n210_), .B(mai_mai_n159_), .C(mai_mai_n36_), .Y(mai_mai_n302_));
  OAI210     m286(.A0(mai_mai_n302_), .A1(mai_mai_n301_), .B0(x7), .Y(mai_mai_n303_));
  NA2        m287(.A(x9), .B(x7), .Y(mai_mai_n304_));
  NA3        m288(.A(mai_mai_n304_), .B(mai_mai_n331_), .C(mai_mai_n124_), .Y(mai_mai_n305_));
  NA2        m289(.A(mai_mai_n305_), .B(mai_mai_n303_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n306_), .A1(mai_mai_n299_), .B0(mai_mai_n33_), .Y(mai_mai_n307_));
  NA2        m291(.A(x3), .B(x7), .Y(mai_mai_n308_));
  NO2        m292(.A(mai_mai_n146_), .B(mai_mai_n125_), .Y(mai_mai_n309_));
  NA2        m293(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  AOI210     m294(.A0(mai_mai_n310_), .A1(mai_mai_n150_), .B0(mai_mai_n25_), .Y(mai_mai_n311_));
  NA2        m295(.A(x0), .B(mai_mai_n287_), .Y(mai_mai_n312_));
  NA2        m296(.A(mai_mai_n312_), .B(x5), .Y(mai_mai_n313_));
  INV        m297(.A(mai_mai_n66_), .Y(mai_mai_n314_));
  NO3        m298(.A(mai_mai_n293_), .B(x3), .C(mai_mai_n50_), .Y(mai_mai_n315_));
  AOI210     m299(.A0(mai_mai_n315_), .A1(x1), .B0(mai_mai_n314_), .Y(mai_mai_n316_));
  AOI210     m300(.A0(mai_mai_n316_), .A1(mai_mai_n313_), .B0(mai_mai_n193_), .Y(mai_mai_n317_));
  NO2        m301(.A(mai_mai_n317_), .B(mai_mai_n311_), .Y(mai_mai_n318_));
  NA3        m302(.A(mai_mai_n318_), .B(mai_mai_n307_), .C(mai_mai_n283_), .Y(mai_mai_n319_));
  AOI210     m303(.A0(mai_mai_n270_), .A1(mai_mai_n23_), .B0(mai_mai_n319_), .Y(mai05));
  INV        m304(.A(x4), .Y(mai_mai_n323_));
  INV        m305(.A(mai_mai_n32_), .Y(mai_mai_n324_));
  INV        m306(.A(mai_mai_n187_), .Y(mai_mai_n325_));
  INV        m307(.A(mai_mai_n72_), .Y(mai_mai_n326_));
  INV        m308(.A(mai_mai_n228_), .Y(mai_mai_n327_));
  INV        m309(.A(x2), .Y(mai_mai_n328_));
  INV        m310(.A(x0), .Y(mai_mai_n329_));
  INV        m311(.A(x3), .Y(mai_mai_n330_));
  INV        m312(.A(x2), .Y(mai_mai_n331_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO3        u012(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  NOi21      u016(.An(men_men_n23_), .B(men_men_n30_), .Y(men00));
  NO2        u017(.A(x1), .B(x0), .Y(men_men_n34_));
  INV        u018(.A(x6), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA2        u020(.A(men_men_n36_), .B(men_men_n34_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n23_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NA2        u027(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u028(.A(x4), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n45_), .B(men_men_n17_), .Y(men_men_n46_));
  NA2        u030(.A(men_men_n46_), .B(x2), .Y(men_men_n47_));
  INV        u031(.A(men_men_n44_), .Y(men_men_n48_));
  AOI210     u032(.A0(men_men_n475_), .A1(men_men_n34_), .B0(men_men_n22_), .Y(men_men_n49_));
  INV        u033(.A(x2), .Y(men_men_n50_));
  NO2        u034(.A(men_men_n50_), .B(men_men_n17_), .Y(men_men_n51_));
  INV        u035(.A(men_men_n51_), .Y(men_men_n52_));
  OAI210     u036(.A0(men_men_n49_), .A1(men_men_n32_), .B0(men_men_n52_), .Y(men_men_n53_));
  NO3        u037(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n39_), .Y(men01));
  NA2        u038(.A(x8), .B(x7), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n41_), .B(x1), .Y(men_men_n56_));
  INV        u040(.A(x9), .Y(men_men_n57_));
  NO2        u041(.A(men_men_n57_), .B(men_men_n35_), .Y(men_men_n58_));
  INV        u042(.A(men_men_n58_), .Y(men_men_n59_));
  NO2        u043(.A(men_men_n59_), .B(men_men_n55_), .Y(men_men_n60_));
  NO2        u044(.A(x7), .B(x6), .Y(men_men_n61_));
  NO2        u045(.A(men_men_n56_), .B(x5), .Y(men_men_n62_));
  NO2        u046(.A(x8), .B(x2), .Y(men_men_n63_));
  INV        u047(.A(men_men_n63_), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n64_), .B(x1), .Y(men_men_n65_));
  OA210      u049(.A0(men_men_n65_), .A1(men_men_n62_), .B0(men_men_n61_), .Y(men_men_n66_));
  NA2        u050(.A(men_men_n25_), .B(men_men_n50_), .Y(men_men_n67_));
  INV        u051(.A(men_men_n67_), .Y(men_men_n68_));
  NAi31      u052(.An(x1), .B(x9), .C(x5), .Y(men_men_n69_));
  OAI220     u053(.A0(men_men_n69_), .A1(men_men_n41_), .B0(men_men_n68_), .B1(men_men_n66_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n70_), .A1(men_men_n60_), .B0(x4), .Y(men_men_n71_));
  NA2        u055(.A(men_men_n45_), .B(x2), .Y(men_men_n72_));
  INV        u056(.A(x0), .Y(men_men_n73_));
  NA2        u057(.A(x5), .B(x3), .Y(men_men_n74_));
  NO2        u058(.A(x8), .B(x6), .Y(men_men_n75_));
  NO3        u059(.A(men_men_n75_), .B(men_men_n61_), .C(men_men_n50_), .Y(men_men_n76_));
  NAi21      u060(.An(x4), .B(x3), .Y(men_men_n77_));
  INV        u061(.A(men_men_n77_), .Y(men_men_n78_));
  NO2        u062(.A(x4), .B(x2), .Y(men_men_n79_));
  NO2        u063(.A(men_men_n79_), .B(x3), .Y(men_men_n80_));
  NO3        u064(.A(men_men_n80_), .B(men_men_n21_), .C(men_men_n18_), .Y(men_men_n81_));
  NO3        u065(.A(men_men_n81_), .B(men_men_n76_), .C(men_men_n73_), .Y(men_men_n82_));
  NO3        u066(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .Y(men_men_n83_));
  NA2        u067(.A(men_men_n57_), .B(men_men_n45_), .Y(men_men_n84_));
  INV        u068(.A(men_men_n84_), .Y(men_men_n85_));
  OAI210     u069(.A0(men_men_n83_), .A1(men_men_n62_), .B0(men_men_n85_), .Y(men_men_n86_));
  NA2        u070(.A(x3), .B(men_men_n18_), .Y(men_men_n87_));
  NO2        u071(.A(men_men_n87_), .B(men_men_n25_), .Y(men_men_n88_));
  INV        u072(.A(x8), .Y(men_men_n89_));
  NA2        u073(.A(x2), .B(x1), .Y(men_men_n90_));
  NO2        u074(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n88_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n26_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n25_), .B(men_men_n50_), .Y(men_men_n94_));
  NO3        u078(.A(x4), .B(men_men_n94_), .C(men_men_n93_), .Y(men_men_n95_));
  NA2        u079(.A(x4), .B(men_men_n41_), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n45_), .B(men_men_n50_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n97_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n98_));
  AOI210     u082(.A0(men_men_n96_), .A1(men_men_n475_), .B0(men_men_n98_), .Y(men_men_n99_));
  NO2        u083(.A(x3), .B(x2), .Y(men_men_n100_));
  NA2        u084(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n101_));
  AOI210     u085(.A0(x8), .A1(x6), .B0(men_men_n101_), .Y(men_men_n102_));
  NA2        u086(.A(men_men_n50_), .B(x1), .Y(men_men_n103_));
  OAI210     u087(.A0(men_men_n103_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n104_));
  NO4        u088(.A(men_men_n104_), .B(men_men_n102_), .C(men_men_n99_), .D(men_men_n95_), .Y(men_men_n105_));
  AO220      u089(.A0(men_men_n105_), .A1(men_men_n86_), .B0(men_men_n82_), .B1(men_men_n71_), .Y(men02));
  NO2        u090(.A(x3), .B(men_men_n50_), .Y(men_men_n107_));
  NO2        u091(.A(x8), .B(men_men_n18_), .Y(men_men_n108_));
  NA2        u092(.A(men_men_n50_), .B(men_men_n17_), .Y(men_men_n109_));
  NA2        u093(.A(men_men_n41_), .B(x0), .Y(men_men_n110_));
  OAI210     u094(.A0(men_men_n84_), .A1(men_men_n109_), .B0(men_men_n110_), .Y(men_men_n111_));
  AOI220     u095(.A0(men_men_n111_), .A1(men_men_n108_), .B0(men_men_n107_), .B1(x4), .Y(men_men_n112_));
  NO3        u096(.A(men_men_n112_), .B(x7), .C(x5), .Y(men_men_n113_));
  NA2        u097(.A(x9), .B(x2), .Y(men_men_n114_));
  OR2        u098(.A(x8), .B(x0), .Y(men_men_n115_));
  INV        u099(.A(men_men_n115_), .Y(men_men_n116_));
  NAi21      u100(.An(x2), .B(x8), .Y(men_men_n117_));
  INV        u101(.A(men_men_n117_), .Y(men_men_n118_));
  OAI210     u102(.A0(men_men_n114_), .A1(x7), .B0(men_men_n116_), .Y(men_men_n119_));
  NO2        u103(.A(x4), .B(x1), .Y(men_men_n120_));
  NA3        u104(.A(men_men_n120_), .B(men_men_n119_), .C(men_men_n55_), .Y(men_men_n121_));
  NOi21      u105(.An(x0), .B(x1), .Y(men_men_n122_));
  NO3        u106(.A(x9), .B(x8), .C(x7), .Y(men_men_n123_));
  NOi21      u107(.An(x0), .B(x4), .Y(men_men_n124_));
  NAi21      u108(.An(x8), .B(x7), .Y(men_men_n125_));
  NO2        u109(.A(men_men_n125_), .B(men_men_n57_), .Y(men_men_n126_));
  AOI220     u110(.A0(men_men_n126_), .A1(men_men_n124_), .B0(men_men_n123_), .B1(men_men_n122_), .Y(men_men_n127_));
  AOI210     u111(.A0(men_men_n127_), .A1(men_men_n121_), .B0(men_men_n74_), .Y(men_men_n128_));
  NO2        u112(.A(x5), .B(men_men_n45_), .Y(men_men_n129_));
  NA2        u113(.A(x2), .B(men_men_n18_), .Y(men_men_n130_));
  INV        u114(.A(men_men_n110_), .Y(men_men_n131_));
  OAI210     u115(.A0(men_men_n131_), .A1(men_men_n34_), .B0(men_men_n129_), .Y(men_men_n132_));
  NAi21      u116(.An(x0), .B(x4), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n133_), .B(x1), .Y(men_men_n134_));
  NO2        u118(.A(x7), .B(x0), .Y(men_men_n135_));
  NO2        u119(.A(men_men_n79_), .B(men_men_n97_), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x3), .Y(men_men_n137_));
  OAI210     u121(.A0(men_men_n135_), .A1(men_men_n134_), .B0(men_men_n137_), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n139_));
  NA2        u123(.A(x5), .B(x0), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n45_), .B(x2), .Y(men_men_n141_));
  NA3        u125(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n139_), .Y(men_men_n142_));
  NA4        u126(.A(men_men_n142_), .B(men_men_n138_), .C(men_men_n132_), .D(men_men_n35_), .Y(men_men_n143_));
  NO3        u127(.A(men_men_n143_), .B(men_men_n128_), .C(men_men_n113_), .Y(men_men_n144_));
  NO3        u128(.A(men_men_n74_), .B(men_men_n72_), .C(men_men_n24_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n146_));
  AOI220     u130(.A0(men_men_n122_), .A1(men_men_n146_), .B0(men_men_n62_), .B1(men_men_n17_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n147_), .B(men_men_n55_), .C(men_men_n57_), .Y(men_men_n148_));
  NA2        u132(.A(x7), .B(x3), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n96_), .B(x5), .Y(men_men_n150_));
  NO2        u134(.A(x9), .B(x7), .Y(men_men_n151_));
  NOi21      u135(.An(x8), .B(x0), .Y(men_men_n152_));
  OA210      u136(.A0(men_men_n151_), .A1(x1), .B0(men_men_n152_), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n41_), .B(x2), .Y(men_men_n154_));
  INV        u138(.A(x7), .Y(men_men_n155_));
  NA2        u139(.A(men_men_n155_), .B(men_men_n18_), .Y(men_men_n156_));
  AOI220     u140(.A0(men_men_n156_), .A1(men_men_n154_), .B0(men_men_n107_), .B1(men_men_n36_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n25_), .B(x4), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n158_), .B(men_men_n124_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n159_), .B(men_men_n157_), .Y(men_men_n160_));
  AOI210     u144(.A0(men_men_n153_), .A1(men_men_n150_), .B0(men_men_n160_), .Y(men_men_n161_));
  OAI210     u145(.A0(men_men_n149_), .A1(men_men_n47_), .B0(men_men_n161_), .Y(men_men_n162_));
  NA2        u146(.A(x5), .B(x1), .Y(men_men_n163_));
  INV        u147(.A(men_men_n163_), .Y(men_men_n164_));
  AOI210     u148(.A0(men_men_n164_), .A1(men_men_n124_), .B0(men_men_n35_), .Y(men_men_n165_));
  NO2        u149(.A(men_men_n57_), .B(men_men_n89_), .Y(men_men_n166_));
  NAi21      u150(.An(x2), .B(x7), .Y(men_men_n167_));
  NO3        u151(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n45_), .Y(men_men_n168_));
  NA2        u152(.A(men_men_n168_), .B(men_men_n62_), .Y(men_men_n169_));
  NAi31      u153(.An(men_men_n74_), .B(men_men_n36_), .C(men_men_n34_), .Y(men_men_n170_));
  NA3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n165_), .Y(men_men_n171_));
  NO4        u155(.A(men_men_n171_), .B(men_men_n162_), .C(men_men_n148_), .D(men_men_n145_), .Y(men_men_n172_));
  NO2        u156(.A(men_men_n172_), .B(men_men_n144_), .Y(men_men_n173_));
  NA2        u157(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n174_));
  NA2        u158(.A(x8), .B(x0), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n155_), .B(men_men_n25_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n122_), .B(x4), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n177_), .B(men_men_n176_), .Y(men_men_n178_));
  AOI210     u162(.A0(men_men_n175_), .A1(men_men_n130_), .B0(men_men_n178_), .Y(men_men_n179_));
  NA2        u163(.A(x2), .B(x0), .Y(men_men_n180_));
  NA2        u164(.A(x4), .B(x1), .Y(men_men_n181_));
  INV        u165(.A(men_men_n179_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n182_), .B(men_men_n41_), .Y(men_men_n183_));
  INV        u167(.A(men_men_n129_), .Y(men_men_n184_));
  NO2        u168(.A(men_men_n103_), .B(men_men_n17_), .Y(men_men_n185_));
  AOI210     u169(.A0(men_men_n34_), .A1(men_men_n89_), .B0(men_men_n185_), .Y(men_men_n186_));
  NO3        u170(.A(men_men_n186_), .B(men_men_n184_), .C(x7), .Y(men_men_n187_));
  NA3        u171(.A(x4), .B(men_men_n184_), .C(men_men_n40_), .Y(men_men_n188_));
  INV        u172(.A(men_men_n188_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n189_), .B(men_men_n187_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(x3), .Y(men_men_n191_));
  NO3        u175(.A(men_men_n191_), .B(men_men_n183_), .C(men_men_n173_), .Y(men03));
  NO2        u176(.A(men_men_n45_), .B(x3), .Y(men_men_n193_));
  NO2        u177(.A(men_men_n50_), .B(x1), .Y(men_men_n194_));
  OAI210     u178(.A0(men_men_n194_), .A1(men_men_n25_), .B0(men_men_n58_), .Y(men_men_n195_));
  OAI220     u179(.A0(men_men_n195_), .A1(men_men_n17_), .B0(x6), .B1(men_men_n103_), .Y(men_men_n196_));
  NA2        u180(.A(men_men_n196_), .B(men_men_n193_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n74_), .B(x6), .Y(men_men_n198_));
  NA2        u182(.A(x6), .B(men_men_n25_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n199_), .B(x4), .Y(men_men_n200_));
  NO2        u184(.A(men_men_n18_), .B(x0), .Y(men_men_n201_));
  AO220      u185(.A0(men_men_n201_), .A1(men_men_n200_), .B0(men_men_n198_), .B1(men_men_n51_), .Y(men_men_n202_));
  NA2        u186(.A(men_men_n202_), .B(men_men_n57_), .Y(men_men_n203_));
  NA2        u187(.A(x3), .B(men_men_n17_), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n204_), .B(men_men_n199_), .Y(men_men_n205_));
  NA2        u189(.A(x9), .B(men_men_n50_), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n206_), .B(x4), .Y(men_men_n207_));
  NA2        u191(.A(men_men_n199_), .B(men_men_n77_), .Y(men_men_n208_));
  AOI210     u192(.A0(men_men_n25_), .A1(x3), .B0(men_men_n180_), .Y(men_men_n209_));
  AOI220     u193(.A0(men_men_n209_), .A1(men_men_n208_), .B0(men_men_n207_), .B1(men_men_n205_), .Y(men_men_n210_));
  NO3        u194(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n211_));
  NO2        u195(.A(x5), .B(x1), .Y(men_men_n212_));
  AOI220     u196(.A0(men_men_n212_), .A1(men_men_n17_), .B0(men_men_n100_), .B1(x5), .Y(men_men_n213_));
  NO2        u197(.A(men_men_n204_), .B(men_men_n174_), .Y(men_men_n214_));
  NO3        u198(.A(x3), .B(x2), .C(x1), .Y(men_men_n215_));
  NO2        u199(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n216_));
  OAI210     u200(.A0(men_men_n213_), .A1(men_men_n59_), .B0(men_men_n216_), .Y(men_men_n217_));
  AOI220     u201(.A0(men_men_n217_), .A1(men_men_n45_), .B0(men_men_n211_), .B1(men_men_n129_), .Y(men_men_n218_));
  NA4        u202(.A(men_men_n218_), .B(men_men_n210_), .C(men_men_n203_), .D(men_men_n197_), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n45_), .B(men_men_n41_), .Y(men_men_n220_));
  NA2        u204(.A(men_men_n220_), .B(men_men_n19_), .Y(men_men_n221_));
  NO2        u205(.A(x3), .B(men_men_n17_), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n222_), .B(x6), .Y(men_men_n223_));
  NOi21      u207(.An(men_men_n79_), .B(men_men_n223_), .Y(men_men_n224_));
  NA2        u208(.A(men_men_n57_), .B(men_men_n89_), .Y(men_men_n225_));
  NA3        u209(.A(men_men_n225_), .B(men_men_n222_), .C(x6), .Y(men_men_n226_));
  AOI210     u210(.A0(men_men_n226_), .A1(men_men_n224_), .B0(men_men_n155_), .Y(men_men_n227_));
  AO210      u211(.A0(men_men_n227_), .A1(men_men_n221_), .B0(men_men_n176_), .Y(men_men_n228_));
  NA2        u212(.A(men_men_n41_), .B(men_men_n50_), .Y(men_men_n229_));
  OAI210     u213(.A0(men_men_n229_), .A1(men_men_n25_), .B0(x5), .Y(men_men_n230_));
  NO3        u214(.A(men_men_n181_), .B(men_men_n57_), .C(x6), .Y(men_men_n231_));
  NA2        u215(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  NA2        u216(.A(x6), .B(men_men_n45_), .Y(men_men_n233_));
  OAI210     u217(.A0(men_men_n116_), .A1(men_men_n75_), .B0(x4), .Y(men_men_n234_));
  AOI210     u218(.A0(men_men_n234_), .A1(men_men_n233_), .B0(men_men_n74_), .Y(men_men_n235_));
  NO2        u219(.A(men_men_n57_), .B(x6), .Y(men_men_n236_));
  NO2        u220(.A(men_men_n163_), .B(men_men_n41_), .Y(men_men_n237_));
  OAI210     u221(.A0(men_men_n237_), .A1(men_men_n214_), .B0(men_men_n236_), .Y(men_men_n238_));
  NA3        u222(.A(men_men_n204_), .B(men_men_n129_), .C(x6), .Y(men_men_n239_));
  NA2        u223(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  OAI210     u224(.A0(men_men_n240_), .A1(men_men_n235_), .B0(x2), .Y(men_men_n241_));
  NA3        u225(.A(men_men_n241_), .B(men_men_n232_), .C(men_men_n228_), .Y(men_men_n242_));
  AOI210     u226(.A0(men_men_n219_), .A1(x8), .B0(men_men_n242_), .Y(men_men_n243_));
  NO2        u227(.A(men_men_n89_), .B(x3), .Y(men_men_n244_));
  NA2        u228(.A(men_men_n244_), .B(men_men_n200_), .Y(men_men_n245_));
  NO3        u229(.A(men_men_n87_), .B(men_men_n75_), .C(men_men_n25_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n223_), .A1(men_men_n158_), .B0(men_men_n246_), .Y(men_men_n247_));
  AOI210     u231(.A0(men_men_n247_), .A1(men_men_n245_), .B0(x2), .Y(men_men_n248_));
  NO2        u232(.A(x4), .B(men_men_n50_), .Y(men_men_n249_));
  AOI220     u233(.A0(men_men_n200_), .A1(men_men_n185_), .B0(men_men_n249_), .B1(men_men_n62_), .Y(men_men_n250_));
  NA2        u234(.A(men_men_n57_), .B(x6), .Y(men_men_n251_));
  NA3        u235(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n252_));
  AOI210     u236(.A0(men_men_n252_), .A1(men_men_n140_), .B0(men_men_n251_), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n254_));
  NO2        u238(.A(men_men_n254_), .B(men_men_n25_), .Y(men_men_n255_));
  OAI210     u239(.A0(men_men_n255_), .A1(men_men_n253_), .B0(men_men_n120_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n204_), .B(x6), .Y(men_men_n257_));
  NO2        u241(.A(men_men_n204_), .B(x6), .Y(men_men_n258_));
  NAi21      u242(.An(men_men_n166_), .B(men_men_n258_), .Y(men_men_n259_));
  NA3        u243(.A(men_men_n259_), .B(men_men_n257_), .C(men_men_n146_), .Y(men_men_n260_));
  NA4        u244(.A(men_men_n260_), .B(men_men_n256_), .C(men_men_n250_), .D(men_men_n155_), .Y(men_men_n261_));
  NA2        u245(.A(x5), .B(men_men_n222_), .Y(men_men_n262_));
  NO2        u246(.A(x9), .B(x6), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n140_), .B(men_men_n18_), .Y(men_men_n264_));
  NAi21      u248(.An(men_men_n264_), .B(men_men_n252_), .Y(men_men_n265_));
  NAi21      u249(.An(x1), .B(x4), .Y(men_men_n266_));
  AOI210     u250(.A0(x3), .A1(x2), .B0(men_men_n45_), .Y(men_men_n267_));
  OAI210     u251(.A0(men_men_n140_), .A1(x3), .B0(men_men_n267_), .Y(men_men_n268_));
  AOI220     u252(.A0(men_men_n268_), .A1(men_men_n266_), .B0(men_men_n265_), .B1(men_men_n263_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n269_), .B(men_men_n262_), .Y(men_men_n270_));
  NA2        u254(.A(men_men_n57_), .B(x2), .Y(men_men_n271_));
  NO2        u255(.A(men_men_n271_), .B(men_men_n262_), .Y(men_men_n272_));
  NO3        u256(.A(x9), .B(x6), .C(x0), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n103_), .B(men_men_n25_), .Y(men_men_n274_));
  NA2        u258(.A(x6), .B(x2), .Y(men_men_n275_));
  NO2        u259(.A(men_men_n275_), .B(men_men_n174_), .Y(men_men_n276_));
  AOI210     u260(.A0(men_men_n274_), .A1(men_men_n273_), .B0(men_men_n276_), .Y(men_men_n277_));
  OAI210     u261(.A0(men_men_n277_), .A1(men_men_n41_), .B0(men_men_n476_), .Y(men_men_n278_));
  OAI210     u262(.A0(men_men_n278_), .A1(men_men_n272_), .B0(men_men_n270_), .Y(men_men_n279_));
  NA2        u263(.A(x9), .B(men_men_n41_), .Y(men_men_n280_));
  NO2        u264(.A(men_men_n280_), .B(men_men_n199_), .Y(men_men_n281_));
  OR3        u265(.A(men_men_n281_), .B(men_men_n198_), .C(men_men_n150_), .Y(men_men_n282_));
  NA2        u266(.A(x4), .B(x0), .Y(men_men_n283_));
  NO3        u267(.A(men_men_n69_), .B(men_men_n283_), .C(x6), .Y(men_men_n284_));
  AOI210     u268(.A0(men_men_n282_), .A1(men_men_n40_), .B0(men_men_n284_), .Y(men_men_n285_));
  AOI210     u269(.A0(men_men_n285_), .A1(men_men_n279_), .B0(x8), .Y(men_men_n286_));
  INV        u270(.A(men_men_n251_), .Y(men_men_n287_));
  OAI210     u271(.A0(men_men_n264_), .A1(men_men_n212_), .B0(men_men_n287_), .Y(men_men_n288_));
  INV        u272(.A(men_men_n175_), .Y(men_men_n289_));
  OAI210     u273(.A0(men_men_n289_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n290_), .A1(men_men_n288_), .B0(men_men_n229_), .Y(men_men_n291_));
  NO4        u275(.A(men_men_n291_), .B(men_men_n286_), .C(men_men_n261_), .D(men_men_n248_), .Y(men_men_n292_));
  NO2        u276(.A(men_men_n166_), .B(x1), .Y(men_men_n293_));
  NO3        u277(.A(men_men_n293_), .B(x3), .C(men_men_n35_), .Y(men_men_n294_));
  NA2        u278(.A(men_men_n294_), .B(x2), .Y(men_men_n295_));
  OAI210     u279(.A0(men_men_n289_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n296_));
  AOI210     u280(.A0(men_men_n296_), .A1(men_men_n295_), .B0(men_men_n184_), .Y(men_men_n297_));
  NOi21      u281(.An(men_men_n275_), .B(men_men_n17_), .Y(men_men_n298_));
  NA3        u282(.A(men_men_n298_), .B(men_men_n212_), .C(men_men_n38_), .Y(men_men_n299_));
  AOI210     u283(.A0(men_men_n35_), .A1(men_men_n50_), .B0(x0), .Y(men_men_n300_));
  NA3        u284(.A(men_men_n300_), .B(men_men_n164_), .C(men_men_n32_), .Y(men_men_n301_));
  NA2        u285(.A(x3), .B(x2), .Y(men_men_n302_));
  AOI220     u286(.A0(men_men_n302_), .A1(men_men_n229_), .B0(men_men_n301_), .B1(men_men_n299_), .Y(men_men_n303_));
  NAi21      u287(.An(x4), .B(x0), .Y(men_men_n304_));
  NO3        u288(.A(men_men_n304_), .B(men_men_n42_), .C(x2), .Y(men_men_n305_));
  OAI210     u289(.A0(x6), .A1(men_men_n18_), .B0(men_men_n305_), .Y(men_men_n306_));
  OAI220     u290(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n307_));
  NO2        u291(.A(x9), .B(x8), .Y(men_men_n308_));
  NA3        u292(.A(men_men_n308_), .B(men_men_n35_), .C(men_men_n50_), .Y(men_men_n309_));
  OAI210     u293(.A0(men_men_n300_), .A1(men_men_n298_), .B0(men_men_n309_), .Y(men_men_n310_));
  AOI220     u294(.A0(men_men_n310_), .A1(men_men_n78_), .B0(men_men_n307_), .B1(men_men_n31_), .Y(men_men_n311_));
  AOI210     u295(.A0(men_men_n311_), .A1(men_men_n306_), .B0(men_men_n25_), .Y(men_men_n312_));
  NA3        u296(.A(men_men_n35_), .B(x1), .C(men_men_n17_), .Y(men_men_n313_));
  NO2        u297(.A(men_men_n300_), .B(men_men_n298_), .Y(men_men_n314_));
  INV        u298(.A(men_men_n214_), .Y(men_men_n315_));
  NA2        u299(.A(men_men_n35_), .B(men_men_n41_), .Y(men_men_n316_));
  OR2        u300(.A(men_men_n316_), .B(men_men_n283_), .Y(men_men_n317_));
  OAI220     u301(.A0(men_men_n317_), .A1(men_men_n163_), .B0(men_men_n233_), .B1(men_men_n315_), .Y(men_men_n318_));
  AO210      u302(.A0(men_men_n314_), .A1(men_men_n150_), .B0(men_men_n318_), .Y(men_men_n319_));
  NO4        u303(.A(men_men_n319_), .B(men_men_n312_), .C(men_men_n303_), .D(men_men_n297_), .Y(men_men_n320_));
  OAI210     u304(.A0(men_men_n292_), .A1(men_men_n243_), .B0(men_men_n320_), .Y(men04));
  OAI210     u305(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n322_));
  NA3        u306(.A(men_men_n322_), .B(men_men_n273_), .C(men_men_n80_), .Y(men_men_n323_));
  NO2        u307(.A(x2), .B(x1), .Y(men_men_n324_));
  OAI210     u308(.A0(men_men_n254_), .A1(men_men_n324_), .B0(men_men_n35_), .Y(men_men_n325_));
  NO2        u309(.A(men_men_n324_), .B(men_men_n304_), .Y(men_men_n326_));
  AOI210     u310(.A0(men_men_n57_), .A1(x4), .B0(men_men_n109_), .Y(men_men_n327_));
  OAI210     u311(.A0(men_men_n327_), .A1(men_men_n326_), .B0(men_men_n244_), .Y(men_men_n328_));
  NO2        u312(.A(men_men_n271_), .B(men_men_n87_), .Y(men_men_n329_));
  NO2        u313(.A(men_men_n329_), .B(men_men_n35_), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n302_), .B(men_men_n201_), .Y(men_men_n331_));
  NA2        u315(.A(x9), .B(x0), .Y(men_men_n332_));
  AOI210     u316(.A0(men_men_n87_), .A1(men_men_n72_), .B0(men_men_n332_), .Y(men_men_n333_));
  OAI210     u317(.A0(men_men_n333_), .A1(men_men_n331_), .B0(men_men_n89_), .Y(men_men_n334_));
  NA3        u318(.A(men_men_n334_), .B(men_men_n330_), .C(men_men_n328_), .Y(men_men_n335_));
  NA2        u319(.A(men_men_n335_), .B(men_men_n325_), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n206_), .B(men_men_n110_), .Y(men_men_n337_));
  NO3        u321(.A(men_men_n251_), .B(men_men_n117_), .C(men_men_n18_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n338_), .B(men_men_n337_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n115_), .A1(men_men_n103_), .B0(men_men_n175_), .Y(men_men_n340_));
  NA3        u324(.A(men_men_n340_), .B(x6), .C(x3), .Y(men_men_n341_));
  NOi21      u325(.An(men_men_n152_), .B(men_men_n130_), .Y(men_men_n342_));
  AOI210     u326(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n343_));
  OAI220     u327(.A0(men_men_n343_), .A1(men_men_n316_), .B0(men_men_n271_), .B1(men_men_n313_), .Y(men_men_n344_));
  AOI210     u328(.A0(men_men_n342_), .A1(men_men_n58_), .B0(men_men_n344_), .Y(men_men_n345_));
  NA2        u329(.A(x2), .B(men_men_n17_), .Y(men_men_n346_));
  OAI210     u330(.A0(men_men_n103_), .A1(men_men_n17_), .B0(men_men_n346_), .Y(men_men_n347_));
  AOI220     u331(.A0(men_men_n347_), .A1(men_men_n75_), .B0(men_men_n329_), .B1(men_men_n89_), .Y(men_men_n348_));
  NA4        u332(.A(men_men_n348_), .B(men_men_n345_), .C(men_men_n341_), .D(men_men_n339_), .Y(men_men_n349_));
  OAI210     u333(.A0(men_men_n108_), .A1(x3), .B0(men_men_n305_), .Y(men_men_n350_));
  NA3        u334(.A(men_men_n225_), .B(men_men_n211_), .C(men_men_n79_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n351_), .B(men_men_n350_), .C(men_men_n155_), .Y(men_men_n352_));
  AOI210     u336(.A0(men_men_n349_), .A1(x4), .B0(men_men_n352_), .Y(men_men_n353_));
  NA3        u337(.A(men_men_n326_), .B(men_men_n206_), .C(men_men_n89_), .Y(men_men_n354_));
  NOi21      u338(.An(x4), .B(x0), .Y(men_men_n355_));
  XO2        u339(.A(x4), .B(x0), .Y(men_men_n356_));
  OAI210     u340(.A0(men_men_n356_), .A1(men_men_n114_), .B0(men_men_n266_), .Y(men_men_n357_));
  AOI220     u341(.A0(men_men_n357_), .A1(x8), .B0(men_men_n355_), .B1(men_men_n90_), .Y(men_men_n358_));
  AOI210     u342(.A0(men_men_n358_), .A1(men_men_n354_), .B0(x3), .Y(men_men_n359_));
  INV        u343(.A(men_men_n90_), .Y(men_men_n360_));
  NO2        u344(.A(men_men_n89_), .B(x4), .Y(men_men_n361_));
  AOI220     u345(.A0(men_men_n361_), .A1(men_men_n42_), .B0(men_men_n124_), .B1(men_men_n360_), .Y(men_men_n362_));
  NO3        u346(.A(men_men_n356_), .B(men_men_n166_), .C(x2), .Y(men_men_n363_));
  NO3        u347(.A(men_men_n225_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n364_));
  NO2        u348(.A(men_men_n364_), .B(men_men_n363_), .Y(men_men_n365_));
  NA4        u349(.A(men_men_n365_), .B(men_men_n362_), .C(men_men_n221_), .D(x6), .Y(men_men_n366_));
  OAI220     u350(.A0(men_men_n304_), .A1(men_men_n87_), .B0(men_men_n180_), .B1(men_men_n89_), .Y(men_men_n367_));
  NO2        u351(.A(men_men_n41_), .B(x0), .Y(men_men_n368_));
  OR2        u352(.A(men_men_n361_), .B(men_men_n368_), .Y(men_men_n369_));
  NO2        u353(.A(men_men_n152_), .B(men_men_n103_), .Y(men_men_n370_));
  AOI220     u354(.A0(men_men_n370_), .A1(men_men_n369_), .B0(men_men_n367_), .B1(men_men_n56_), .Y(men_men_n371_));
  NO2        u355(.A(men_men_n152_), .B(men_men_n77_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n34_), .B(x2), .Y(men_men_n373_));
  NOi21      u357(.An(men_men_n120_), .B(men_men_n27_), .Y(men_men_n374_));
  AOI210     u358(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n374_), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n371_), .A1(men_men_n57_), .B0(men_men_n375_), .Y(men_men_n376_));
  OAI220     u360(.A0(men_men_n376_), .A1(x6), .B0(men_men_n366_), .B1(men_men_n359_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n58_), .A1(men_men_n45_), .B0(men_men_n40_), .Y(men_men_n378_));
  OAI210     u362(.A0(men_men_n378_), .A1(men_men_n89_), .B0(men_men_n317_), .Y(men_men_n379_));
  AOI210     u363(.A0(men_men_n379_), .A1(men_men_n18_), .B0(men_men_n155_), .Y(men_men_n380_));
  AO220      u364(.A0(men_men_n380_), .A1(men_men_n377_), .B0(men_men_n353_), .B1(men_men_n336_), .Y(men_men_n381_));
  NA2        u365(.A(men_men_n373_), .B(x6), .Y(men_men_n382_));
  AOI210     u366(.A0(x6), .A1(x1), .B0(men_men_n154_), .Y(men_men_n383_));
  NA2        u367(.A(men_men_n361_), .B(x0), .Y(men_men_n384_));
  NO2        u368(.A(men_men_n384_), .B(men_men_n383_), .Y(men_men_n385_));
  AOI220     u369(.A0(men_men_n385_), .A1(men_men_n382_), .B0(men_men_n215_), .B1(men_men_n46_), .Y(men_men_n386_));
  NA3        u370(.A(men_men_n386_), .B(men_men_n381_), .C(men_men_n323_), .Y(men_men_n387_));
  AOI210     u371(.A0(men_men_n194_), .A1(x8), .B0(men_men_n108_), .Y(men_men_n388_));
  NA2        u372(.A(men_men_n388_), .B(men_men_n346_), .Y(men_men_n389_));
  NA3        u373(.A(men_men_n389_), .B(men_men_n193_), .C(men_men_n155_), .Y(men_men_n390_));
  OAI210     u374(.A0(men_men_n28_), .A1(x1), .B0(men_men_n229_), .Y(men_men_n391_));
  AO220      u375(.A0(men_men_n391_), .A1(men_men_n151_), .B0(men_men_n107_), .B1(x4), .Y(men_men_n392_));
  NA3        u376(.A(x7), .B(x3), .C(x0), .Y(men_men_n393_));
  NA2        u377(.A(men_men_n220_), .B(x0), .Y(men_men_n394_));
  NO2        u378(.A(men_men_n394_), .B(men_men_n206_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n392_), .A1(men_men_n116_), .B0(men_men_n395_), .Y(men_men_n396_));
  AOI210     u380(.A0(men_men_n396_), .A1(men_men_n390_), .B0(men_men_n25_), .Y(men_men_n397_));
  NA3        u381(.A(men_men_n118_), .B(men_men_n220_), .C(x0), .Y(men_men_n398_));
  OAI210     u382(.A0(men_men_n193_), .A1(men_men_n63_), .B0(men_men_n201_), .Y(men_men_n399_));
  NA3        u383(.A(men_men_n194_), .B(men_men_n222_), .C(x8), .Y(men_men_n400_));
  AOI210     u384(.A0(men_men_n400_), .A1(men_men_n399_), .B0(men_men_n25_), .Y(men_men_n401_));
  AOI210     u385(.A0(men_men_n117_), .A1(men_men_n115_), .B0(men_men_n40_), .Y(men_men_n402_));
  NOi31      u386(.An(men_men_n402_), .B(men_men_n368_), .C(men_men_n181_), .Y(men_men_n403_));
  OAI210     u387(.A0(men_men_n403_), .A1(men_men_n401_), .B0(men_men_n151_), .Y(men_men_n404_));
  NAi31      u388(.An(men_men_n47_), .B(men_men_n293_), .C(men_men_n176_), .Y(men_men_n405_));
  NA3        u389(.A(men_men_n405_), .B(men_men_n404_), .C(men_men_n398_), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n406_), .A1(men_men_n397_), .B0(x6), .Y(men_men_n407_));
  OAI210     u391(.A0(men_men_n166_), .A1(men_men_n45_), .B0(men_men_n135_), .Y(men_men_n408_));
  NA3        u392(.A(men_men_n51_), .B(men_men_n36_), .C(men_men_n31_), .Y(men_men_n409_));
  AOI220     u393(.A0(men_men_n409_), .A1(men_men_n408_), .B0(men_men_n38_), .B1(men_men_n32_), .Y(men_men_n410_));
  NO2        u394(.A(men_men_n155_), .B(x0), .Y(men_men_n411_));
  NA2        u395(.A(men_men_n193_), .B(men_men_n155_), .Y(men_men_n412_));
  AOI210     u396(.A0(men_men_n126_), .A1(men_men_n249_), .B0(x1), .Y(men_men_n413_));
  OAI210     u397(.A0(men_men_n412_), .A1(x8), .B0(men_men_n413_), .Y(men_men_n414_));
  NAi31      u398(.An(x2), .B(x8), .C(x0), .Y(men_men_n415_));
  OAI210     u399(.A0(men_men_n415_), .A1(x4), .B0(men_men_n167_), .Y(men_men_n416_));
  NA3        u400(.A(men_men_n416_), .B(men_men_n149_), .C(x9), .Y(men_men_n417_));
  NO4        u401(.A(men_men_n125_), .B(men_men_n304_), .C(x9), .D(x2), .Y(men_men_n418_));
  NOi21      u402(.An(men_men_n123_), .B(men_men_n180_), .Y(men_men_n419_));
  NO3        u403(.A(men_men_n419_), .B(men_men_n418_), .C(men_men_n18_), .Y(men_men_n420_));
  NO3        u404(.A(x9), .B(men_men_n155_), .C(x0), .Y(men_men_n421_));
  AOI220     u405(.A0(men_men_n421_), .A1(men_men_n244_), .B0(men_men_n372_), .B1(men_men_n155_), .Y(men_men_n422_));
  NA4        u406(.A(men_men_n422_), .B(men_men_n420_), .C(men_men_n417_), .D(men_men_n47_), .Y(men_men_n423_));
  OAI210     u407(.A0(men_men_n414_), .A1(men_men_n410_), .B0(men_men_n423_), .Y(men_men_n424_));
  NOi31      u408(.An(men_men_n411_), .B(men_men_n32_), .C(x8), .Y(men_men_n425_));
  AOI210     u409(.A0(men_men_n36_), .A1(x9), .B0(men_men_n133_), .Y(men_men_n426_));
  NO3        u410(.A(men_men_n426_), .B(men_men_n123_), .C(men_men_n41_), .Y(men_men_n427_));
  NOi31      u411(.An(x1), .B(x8), .C(x7), .Y(men_men_n428_));
  AOI220     u412(.A0(men_men_n428_), .A1(men_men_n355_), .B0(men_men_n124_), .B1(x3), .Y(men_men_n429_));
  AOI210     u413(.A0(men_men_n266_), .A1(men_men_n55_), .B0(men_men_n122_), .Y(men_men_n430_));
  OAI210     u414(.A0(men_men_n430_), .A1(x3), .B0(men_men_n429_), .Y(men_men_n431_));
  NO3        u415(.A(men_men_n431_), .B(men_men_n427_), .C(x2), .Y(men_men_n432_));
  OAI220     u416(.A0(men_men_n356_), .A1(men_men_n308_), .B0(men_men_n304_), .B1(men_men_n41_), .Y(men_men_n433_));
  AOI210     u417(.A0(x9), .A1(men_men_n45_), .B0(men_men_n393_), .Y(men_men_n434_));
  AOI220     u418(.A0(men_men_n434_), .A1(men_men_n89_), .B0(men_men_n433_), .B1(men_men_n155_), .Y(men_men_n435_));
  NO2        u419(.A(men_men_n435_), .B(men_men_n50_), .Y(men_men_n436_));
  NO3        u420(.A(men_men_n436_), .B(men_men_n432_), .C(men_men_n425_), .Y(men_men_n437_));
  AOI210     u421(.A0(men_men_n437_), .A1(men_men_n424_), .B0(men_men_n25_), .Y(men_men_n438_));
  NA4        u422(.A(men_men_n31_), .B(men_men_n89_), .C(x2), .D(men_men_n17_), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n57_), .B(x4), .C(x1), .Y(men_men_n440_));
  NO3        u424(.A(men_men_n63_), .B(men_men_n18_), .C(x0), .Y(men_men_n441_));
  AOI220     u425(.A0(men_men_n441_), .A1(men_men_n267_), .B0(men_men_n440_), .B1(men_men_n402_), .Y(men_men_n442_));
  NO2        u426(.A(men_men_n442_), .B(men_men_n100_), .Y(men_men_n443_));
  NO3        u427(.A(men_men_n271_), .B(men_men_n175_), .C(men_men_n38_), .Y(men_men_n444_));
  OAI210     u428(.A0(men_men_n444_), .A1(men_men_n443_), .B0(x7), .Y(men_men_n445_));
  NA2        u429(.A(men_men_n225_), .B(x7), .Y(men_men_n446_));
  NA3        u430(.A(men_men_n446_), .B(men_men_n154_), .C(men_men_n134_), .Y(men_men_n447_));
  NA3        u431(.A(men_men_n447_), .B(men_men_n445_), .C(men_men_n439_), .Y(men_men_n448_));
  OAI210     u432(.A0(men_men_n448_), .A1(men_men_n438_), .B0(men_men_n35_), .Y(men_men_n449_));
  NO2        u433(.A(men_men_n421_), .B(men_men_n201_), .Y(men_men_n450_));
  NO4        u434(.A(men_men_n450_), .B(men_men_n74_), .C(x4), .D(men_men_n50_), .Y(men_men_n451_));
  NA2        u435(.A(men_men_n254_), .B(men_men_n21_), .Y(men_men_n452_));
  NO2        u436(.A(men_men_n163_), .B(men_men_n135_), .Y(men_men_n453_));
  NA2        u437(.A(men_men_n453_), .B(men_men_n452_), .Y(men_men_n454_));
  AOI210     u438(.A0(men_men_n454_), .A1(men_men_n170_), .B0(men_men_n28_), .Y(men_men_n455_));
  AOI220     u439(.A0(men_men_n368_), .A1(men_men_n89_), .B0(men_men_n152_), .B1(men_men_n194_), .Y(men_men_n456_));
  NA3        u440(.A(men_men_n456_), .B(men_men_n415_), .C(men_men_n87_), .Y(men_men_n457_));
  NA2        u441(.A(men_men_n457_), .B(men_men_n176_), .Y(men_men_n458_));
  OAI220     u442(.A0(men_men_n280_), .A1(men_men_n64_), .B0(men_men_n163_), .B1(men_men_n41_), .Y(men_men_n459_));
  NA2        u443(.A(x3), .B(men_men_n50_), .Y(men_men_n460_));
  AOI210     u444(.A0(men_men_n167_), .A1(men_men_n27_), .B0(men_men_n69_), .Y(men_men_n461_));
  OAI210     u445(.A0(men_men_n151_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n462_));
  NO3        u446(.A(men_men_n428_), .B(x3), .C(men_men_n50_), .Y(men_men_n463_));
  AOI210     u447(.A0(men_men_n463_), .A1(men_men_n462_), .B0(men_men_n461_), .Y(men_men_n464_));
  OAI210     u448(.A0(men_men_n156_), .A1(men_men_n460_), .B0(men_men_n464_), .Y(men_men_n465_));
  AOI220     u449(.A0(men_men_n465_), .A1(x0), .B0(men_men_n459_), .B1(men_men_n135_), .Y(men_men_n466_));
  AOI210     u450(.A0(men_men_n466_), .A1(men_men_n458_), .B0(men_men_n233_), .Y(men_men_n467_));
  NA2        u451(.A(x9), .B(x5), .Y(men_men_n468_));
  NO4        u452(.A(men_men_n103_), .B(men_men_n468_), .C(men_men_n55_), .D(men_men_n32_), .Y(men_men_n469_));
  NO4        u453(.A(men_men_n469_), .B(men_men_n467_), .C(men_men_n455_), .D(men_men_n451_), .Y(men_men_n470_));
  NA3        u454(.A(men_men_n470_), .B(men_men_n449_), .C(men_men_n407_), .Y(men_men_n471_));
  AOI210     u455(.A0(men_men_n387_), .A1(men_men_n25_), .B0(men_men_n471_), .Y(men05));
  INV        u456(.A(men_men_n36_), .Y(men_men_n475_));
  INV        u457(.A(x4), .Y(men_men_n476_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule