library verilog;
use verilog.vl_types.all;
entity spi_slave_ex_vlg_vec_tst is
end spi_slave_ex_vlg_vec_tst;
