// Benchmark "top" written by ABC on Fri Jun 21 17:49:22 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n142_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1078_, new_new_n1079_,
    new_new_n1080_, new_new_n1081_, new_new_n1082_, new_new_n1083_,
    new_new_n1084_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA2        g0042(.A(i_1_), .B(i_10_), .Y(new_new_n65_));
  NO2        g0043(.A(new_new_n65_), .B(i_6_), .Y(new_new_n66_));
  NAi21      g0044(.An(new_new_n66_), .B(new_new_n61_), .Y(new_new_n67_));
  NA2        g0045(.A(new_new_n50_), .B(i_2_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  INV        g0053(.A(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n67_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(new_new_n79_), .B(new_new_n58_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  NO3        g0060(.A(new_new_n82_), .B(new_new_n81_), .C(new_new_n63_), .Y(new_new_n83_));
  INV        g0061(.A(i_6_), .Y(new_new_n84_));
  OR4        g0062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n85_));
  INV        g0063(.A(new_new_n85_), .Y(new_new_n86_));
  NO2        g0064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  NO2        g0065(.A(new_new_n86_), .B(new_new_n87_), .Y(new_new_n88_));
  OAI210     g0066(.A0(new_new_n83_), .A1(new_new_n80_), .B0(new_new_n88_), .Y(new_new_n89_));
  NAi21      g0067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g0068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g0069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n63_), .Y(new_new_n92_));
  NA2        g0070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  NO3        g0071(.A(new_new_n93_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n94_));
  NO2        g0072(.A(new_new_n94_), .B(new_new_n92_), .Y(new_new_n95_));
  AOI210     g0073(.A0(new_new_n95_), .A1(new_new_n89_), .B0(new_new_n78_), .Y(new_new_n96_));
  AN3        g0074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n97_));
  NAi21      g0075(.An(i_6_), .B(i_11_), .Y(new_new_n98_));
  NO2        g0076(.A(i_5_), .B(i_8_), .Y(new_new_n99_));
  NOi21      g0077(.An(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  AOI220     g0078(.A0(new_new_n100_), .A1(new_new_n62_), .B0(new_new_n97_), .B1(new_new_n32_), .Y(new_new_n101_));
  INV        g0079(.A(i_7_), .Y(new_new_n102_));
  NA2        g0080(.A(new_new_n46_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g0081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g0082(.A(new_new_n104_), .B(new_new_n84_), .Y(new_new_n105_));
  NA2        g0083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  INV        g0084(.A(new_new_n106_), .Y(new_new_n107_));
  NA3        g0085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n103_), .Y(new_new_n108_));
  NAi21      g0086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g0087(.A(new_new_n109_), .B(new_new_n90_), .C(new_new_n53_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g0089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g0090(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n113_));
  NO2        g0091(.A(i_8_), .B(new_new_n102_), .Y(new_new_n114_));
  NO3        g0092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g0093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g0094(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g0096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g0097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g0098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NAi41      g0099(.An(new_new_n110_), .B(new_new_n121_), .C(new_new_n108_), .D(new_new_n101_), .Y(new_new_n122_));
  NOi21      g0100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g0103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g0105(.A(new_new_n127_), .B(new_new_n46_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n129_));
  NAi21      g0107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n130_), .B(new_new_n62_), .Y(new_new_n131_));
  NOi31      g0109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g0110(.A(i_1_), .B(new_new_n84_), .Y(new_new_n133_));
  NO2        g0111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g0113(.A0(new_new_n135_), .A1(new_new_n47_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g0114(.A0(new_new_n136_), .A1(new_new_n109_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g0115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n96_), .Y(new_new_n138_));
  NA3        g0116(.A(new_new_n138_), .B(new_new_n77_), .C(new_new_n56_), .Y(men2));
  NO2        g0117(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n140_));
  INV        g0118(.A(i_6_), .Y(new_new_n141_));
  NA2        g0119(.A(new_new_n141_), .B(new_new_n140_), .Y(new_new_n142_));
  NA4        g0120(.A(new_new_n142_), .B(new_new_n75_), .C(new_new_n68_), .D(new_new_n30_), .Y(men0));
  AN2        g0121(.A(i_8_), .B(i_7_), .Y(new_new_n144_));
  NA2        g0122(.A(new_new_n144_), .B(i_6_), .Y(new_new_n145_));
  NO2        g0123(.A(i_12_), .B(i_13_), .Y(new_new_n146_));
  NAi21      g0124(.An(i_5_), .B(i_11_), .Y(new_new_n147_));
  NOi21      g0125(.An(new_new_n146_), .B(new_new_n147_), .Y(new_new_n148_));
  NO2        g0126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NA2        g0127(.A(i_2_), .B(i_3_), .Y(new_new_n150_));
  NO2        g0128(.A(new_new_n150_), .B(i_4_), .Y(new_new_n151_));
  NA3        g0129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  OR2        g0130(.A(new_new_n152_), .B(new_new_n25_), .Y(new_new_n153_));
  AN2        g0131(.A(new_new_n146_), .B(new_new_n81_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n154_), .B(new_new_n27_), .Y(new_new_n155_));
  NA2        g0133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  NO2        g0134(.A(new_new_n71_), .B(new_new_n46_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n36_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n156_), .C(new_new_n155_), .Y(new_new_n159_));
  OR2        g0137(.A(i_0_), .B(i_1_), .Y(new_new_n160_));
  NO3        g0138(.A(new_new_n160_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n161_));
  NAi32      g0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n162_));
  NAi21      g0140(.An(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NOi21      g0141(.An(i_4_), .B(i_10_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n39_), .Y(new_new_n165_));
  NO2        g0143(.A(i_3_), .B(i_5_), .Y(new_new_n166_));
  NO3        g0144(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n167_));
  NA2        g0145(.A(new_new_n167_), .B(new_new_n166_), .Y(new_new_n168_));
  OAI210     g0146(.A0(new_new_n168_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n169_));
  NO2        g0147(.A(new_new_n169_), .B(new_new_n159_), .Y(new_new_n170_));
  AOI210     g0148(.A0(new_new_n170_), .A1(new_new_n153_), .B0(new_new_n145_), .Y(new_new_n171_));
  NA3        g0149(.A(new_new_n71_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n172_));
  NA2        g0150(.A(i_3_), .B(new_new_n48_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_4_), .B(i_9_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_11_), .B(i_13_), .Y(new_new_n175_));
  NA2        g0153(.A(new_new_n175_), .B(new_new_n174_), .Y(new_new_n176_));
  OR2        g0154(.A(new_new_n176_), .B(new_new_n173_), .Y(new_new_n177_));
  NO2        g0155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g0156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n81_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n172_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n71_), .B(new_new_n63_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n183_), .B(new_new_n46_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n36_), .B(i_5_), .Y(new_new_n185_));
  NAi31      g0163(.An(new_new_n185_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n186_));
  NA2        g0164(.A(i_3_), .B(i_5_), .Y(new_new_n187_));
  OR2        g0165(.A(new_new_n187_), .B(new_new_n176_), .Y(new_new_n188_));
  AOI210     g0166(.A0(new_new_n188_), .A1(new_new_n186_), .B0(new_new_n184_), .Y(new_new_n189_));
  NO2        g0167(.A(new_new_n71_), .B(i_5_), .Y(new_new_n190_));
  NO2        g0168(.A(i_13_), .B(i_10_), .Y(new_new_n191_));
  NA3        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n44_), .Y(new_new_n192_));
  NO2        g0170(.A(i_2_), .B(i_1_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_3_), .Y(new_new_n194_));
  NAi21      g0172(.An(i_4_), .B(i_12_), .Y(new_new_n195_));
  NO4        g0173(.A(new_new_n195_), .B(new_new_n194_), .C(new_new_n192_), .D(new_new_n25_), .Y(new_new_n196_));
  NO3        g0174(.A(new_new_n196_), .B(new_new_n189_), .C(new_new_n182_), .Y(new_new_n197_));
  INV        g0175(.A(i_8_), .Y(new_new_n198_));
  NO2        g0176(.A(new_new_n198_), .B(i_7_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(i_6_), .Y(new_new_n200_));
  NO3        g0178(.A(i_3_), .B(new_new_n84_), .C(new_new_n48_), .Y(new_new_n201_));
  NA2        g0179(.A(new_new_n201_), .B(new_new_n114_), .Y(new_new_n202_));
  NO3        g0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n205_));
  OAI210     g0183(.A0(new_new_n97_), .A1(i_12_), .B0(new_new_n205_), .Y(new_new_n206_));
  AOI210     g0184(.A0(new_new_n206_), .A1(new_new_n204_), .B0(new_new_n202_), .Y(new_new_n207_));
  NO2        g0185(.A(i_3_), .B(i_8_), .Y(new_new_n208_));
  NO3        g0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(new_new_n208_), .C(new_new_n39_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n104_), .B(new_new_n58_), .Y(new_new_n211_));
  NO2        g0189(.A(i_13_), .B(i_9_), .Y(new_new_n212_));
  NAi21      g0190(.An(i_12_), .B(i_3_), .Y(new_new_n213_));
  OR2        g0191(.A(new_new_n213_), .B(i_8_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n44_), .B(i_5_), .Y(new_new_n215_));
  NO3        g0193(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n216_));
  NA3        g0194(.A(new_new_n216_), .B(new_new_n215_), .C(i_10_), .Y(new_new_n217_));
  OAI220     g0195(.A0(new_new_n217_), .A1(new_new_n214_), .B0(new_new_n104_), .B1(new_new_n210_), .Y(new_new_n218_));
  AOI210     g0196(.A0(new_new_n218_), .A1(i_7_), .B0(new_new_n207_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n219_), .A1(i_4_), .B0(new_new_n200_), .B1(new_new_n197_), .Y(new_new_n220_));
  NAi21      g0198(.An(i_12_), .B(i_7_), .Y(new_new_n221_));
  NA3        g0199(.A(i_13_), .B(new_new_n198_), .C(i_10_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n223_));
  NA2        g0201(.A(i_0_), .B(i_5_), .Y(new_new_n224_));
  NA2        g0202(.A(new_new_n224_), .B(new_new_n105_), .Y(new_new_n225_));
  OAI220     g0203(.A0(new_new_n225_), .A1(new_new_n194_), .B0(new_new_n184_), .B1(new_new_n135_), .Y(new_new_n226_));
  NAi31      g0204(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n36_), .B(i_13_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n230_));
  NA3        g0208(.A(new_new_n230_), .B(new_new_n229_), .C(new_new_n228_), .Y(new_new_n231_));
  INV        g0209(.A(i_13_), .Y(new_new_n232_));
  NO2        g0210(.A(i_12_), .B(new_new_n232_), .Y(new_new_n233_));
  NA3        g0211(.A(new_new_n233_), .B(new_new_n203_), .C(new_new_n201_), .Y(new_new_n234_));
  OAI210     g0212(.A0(new_new_n231_), .A1(new_new_n227_), .B0(new_new_n234_), .Y(new_new_n235_));
  AOI220     g0213(.A0(new_new_n235_), .A1(new_new_n144_), .B0(new_new_n226_), .B1(new_new_n223_), .Y(new_new_n236_));
  NO2        g0214(.A(i_12_), .B(new_new_n37_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n187_), .B(i_4_), .Y(new_new_n238_));
  NA2        g0216(.A(new_new_n238_), .B(new_new_n237_), .Y(new_new_n239_));
  OR2        g0217(.A(i_8_), .B(i_7_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n240_), .B(new_new_n84_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n53_), .B(i_1_), .Y(new_new_n242_));
  NA2        g0220(.A(new_new_n242_), .B(new_new_n241_), .Y(new_new_n243_));
  INV        g0221(.A(i_12_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n44_), .B(new_new_n244_), .Y(new_new_n245_));
  NO3        g0223(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n246_));
  NA2        g0224(.A(i_2_), .B(i_1_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n243_), .B(new_new_n239_), .Y(new_new_n248_));
  NO3        g0226(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n249_));
  NAi21      g0227(.An(i_4_), .B(i_3_), .Y(new_new_n250_));
  NO2        g0228(.A(new_new_n250_), .B(new_new_n73_), .Y(new_new_n251_));
  NO2        g0229(.A(i_0_), .B(i_6_), .Y(new_new_n252_));
  NOi41      g0230(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n253_), .B(new_new_n252_), .Y(new_new_n254_));
  NO2        g0232(.A(new_new_n247_), .B(new_new_n187_), .Y(new_new_n255_));
  INV        g0233(.A(new_new_n248_), .Y(new_new_n256_));
  NO2        g0234(.A(i_11_), .B(new_new_n232_), .Y(new_new_n257_));
  NOi21      g0235(.An(i_1_), .B(i_6_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n244_), .B(i_9_), .Y(new_new_n259_));
  OR4        g0237(.A(new_new_n259_), .B(i_3_), .C(new_new_n258_), .D(new_new_n190_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n71_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NA3        g0244(.A(new_new_n266_), .B(new_new_n263_), .C(new_new_n64_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n267_), .B(new_new_n260_), .Y(new_new_n268_));
  NA3        g0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n269_));
  INV        g0247(.A(new_new_n145_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n244_), .B(i_13_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n73_), .Y(new_new_n272_));
  AOI220     g0250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n268_), .B1(new_new_n257_), .Y(new_new_n273_));
  NO2        g0251(.A(new_new_n240_), .B(new_new_n37_), .Y(new_new_n274_));
  NA2        g0252(.A(i_12_), .B(i_6_), .Y(new_new_n275_));
  OR2        g0253(.A(i_13_), .B(i_9_), .Y(new_new_n276_));
  NO3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n48_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n250_), .B(i_2_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n277_), .C(new_new_n44_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n257_), .B(i_9_), .Y(new_new_n280_));
  OAI210     g0258(.A0(new_new_n71_), .A1(new_new_n280_), .B0(new_new_n279_), .Y(new_new_n281_));
  NA2        g0259(.A(new_new_n157_), .B(new_new_n63_), .Y(new_new_n282_));
  NO3        g0260(.A(i_11_), .B(new_new_n232_), .C(new_new_n25_), .Y(new_new_n283_));
  NO2        g0261(.A(i_6_), .B(new_new_n48_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(i_7_), .C(new_new_n283_), .Y(new_new_n285_));
  NA3        g0263(.A(new_new_n1084_), .B(new_new_n274_), .C(new_new_n233_), .Y(new_new_n286_));
  AOI210     g0264(.A0(new_new_n286_), .A1(new_new_n285_), .B0(new_new_n282_), .Y(new_new_n287_));
  AOI210     g0265(.A0(new_new_n281_), .A1(new_new_n274_), .B0(new_new_n287_), .Y(new_new_n288_));
  NA4        g0266(.A(new_new_n288_), .B(new_new_n273_), .C(new_new_n256_), .D(new_new_n236_), .Y(new_new_n289_));
  NO3        g0267(.A(i_12_), .B(new_new_n232_), .C(new_new_n37_), .Y(new_new_n290_));
  INV        g0268(.A(new_new_n290_), .Y(new_new_n291_));
  NOi21      g0269(.An(new_new_n166_), .B(new_new_n84_), .Y(new_new_n292_));
  NO3        g0270(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n201_), .B0(new_new_n292_), .B1(new_new_n242_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(i_7_), .Y(new_new_n295_));
  NO3        g0273(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n247_), .B(i_0_), .Y(new_new_n297_));
  AOI220     g0275(.A0(new_new_n297_), .A1(new_new_n199_), .B0(new_new_n296_), .B1(new_new_n144_), .Y(new_new_n298_));
  NA2        g0276(.A(new_new_n284_), .B(new_new_n26_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(new_new_n298_), .Y(new_new_n300_));
  NA2        g0278(.A(i_0_), .B(i_1_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n301_), .B(i_2_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n59_), .B(i_6_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n302_), .C(new_new_n166_), .Y(new_new_n304_));
  OAI210     g0282(.A0(new_new_n168_), .A1(new_new_n145_), .B0(new_new_n304_), .Y(new_new_n305_));
  NO3        g0283(.A(new_new_n305_), .B(new_new_n300_), .C(new_new_n295_), .Y(new_new_n306_));
  NO2        g0284(.A(i_3_), .B(i_10_), .Y(new_new_n307_));
  NA3        g0285(.A(new_new_n307_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n308_));
  NO2        g0286(.A(i_2_), .B(new_new_n102_), .Y(new_new_n309_));
  NOi21      g0287(.An(new_new_n224_), .B(new_new_n104_), .Y(new_new_n310_));
  NA3        g0288(.A(new_new_n310_), .B(new_new_n36_), .C(new_new_n309_), .Y(new_new_n311_));
  AN2        g0289(.A(i_3_), .B(i_10_), .Y(new_new_n312_));
  NA4        g0290(.A(new_new_n312_), .B(new_new_n203_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n313_));
  NO2        g0291(.A(i_5_), .B(new_new_n37_), .Y(new_new_n314_));
  NO2        g0292(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n315_));
  OR2        g0293(.A(new_new_n311_), .B(new_new_n308_), .Y(new_new_n316_));
  OAI220     g0294(.A0(new_new_n316_), .A1(i_6_), .B0(new_new_n306_), .B1(new_new_n291_), .Y(new_new_n317_));
  NO4        g0295(.A(new_new_n317_), .B(new_new_n289_), .C(new_new_n220_), .D(new_new_n171_), .Y(new_new_n318_));
  NO3        g0296(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n319_));
  NO3        g0297(.A(i_6_), .B(new_new_n198_), .C(i_7_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n320_), .B(new_new_n203_), .Y(new_new_n321_));
  AOI210     g0299(.A0(new_new_n321_), .A1(new_new_n247_), .B0(new_new_n173_), .Y(new_new_n322_));
  NO2        g0300(.A(i_2_), .B(i_3_), .Y(new_new_n323_));
  OR2        g0301(.A(i_0_), .B(i_5_), .Y(new_new_n324_));
  NA2        g0302(.A(new_new_n224_), .B(new_new_n324_), .Y(new_new_n325_));
  NA3        g0303(.A(new_new_n325_), .B(new_new_n241_), .C(new_new_n323_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n297_), .B(new_new_n292_), .C(new_new_n114_), .Y(new_new_n327_));
  NO2        g0305(.A(i_8_), .B(i_6_), .Y(new_new_n328_));
  NO2        g0306(.A(new_new_n160_), .B(new_new_n46_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n329_), .B(new_new_n328_), .C(new_new_n166_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n330_), .B(new_new_n327_), .C(new_new_n326_), .Y(new_new_n331_));
  OAI210     g0309(.A0(new_new_n331_), .A1(new_new_n322_), .B0(i_4_), .Y(new_new_n332_));
  NO2        g0310(.A(i_12_), .B(i_10_), .Y(new_new_n333_));
  NOi21      g0311(.An(i_5_), .B(i_0_), .Y(new_new_n334_));
  AOI210     g0312(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n102_), .Y(new_new_n335_));
  NO4        g0313(.A(new_new_n335_), .B(i_4_), .C(new_new_n334_), .D(new_new_n130_), .Y(new_new_n336_));
  NA4        g0314(.A(new_new_n82_), .B(new_new_n36_), .C(new_new_n84_), .D(i_8_), .Y(new_new_n337_));
  NA2        g0315(.A(new_new_n336_), .B(new_new_n333_), .Y(new_new_n338_));
  NO2        g0316(.A(i_6_), .B(i_8_), .Y(new_new_n339_));
  AN2        g0317(.A(i_0_), .B(new_new_n339_), .Y(new_new_n340_));
  NO2        g0318(.A(i_1_), .B(i_7_), .Y(new_new_n341_));
  NA3        g0319(.A(new_new_n340_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n342_));
  NA3        g0320(.A(new_new_n342_), .B(new_new_n338_), .C(new_new_n332_), .Y(new_new_n343_));
  NO2        g0321(.A(i_8_), .B(new_new_n325_), .Y(new_new_n344_));
  NOi21      g0322(.An(new_new_n156_), .B(new_new_n105_), .Y(new_new_n345_));
  NO2        g0323(.A(new_new_n345_), .B(new_new_n126_), .Y(new_new_n346_));
  OAI210     g0324(.A0(new_new_n346_), .A1(new_new_n344_), .B0(i_3_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n301_), .B(new_new_n79_), .Y(new_new_n348_));
  NA2        g0326(.A(new_new_n348_), .B(new_new_n134_), .Y(new_new_n349_));
  NO2        g0327(.A(new_new_n93_), .B(new_new_n198_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n310_), .B(new_new_n350_), .C(new_new_n63_), .Y(new_new_n351_));
  AOI210     g0329(.A0(new_new_n351_), .A1(new_new_n349_), .B0(i_3_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n198_), .B(i_9_), .Y(new_new_n353_));
  NA2        g0331(.A(new_new_n353_), .B(new_new_n211_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n354_), .B(new_new_n46_), .Y(new_new_n355_));
  NO3        g0333(.A(new_new_n355_), .B(new_new_n352_), .C(new_new_n300_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n356_), .A1(new_new_n347_), .B0(new_new_n165_), .Y(new_new_n357_));
  AOI210     g0335(.A0(new_new_n343_), .A1(new_new_n319_), .B0(new_new_n357_), .Y(new_new_n358_));
  NOi32      g0336(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n359_));
  INV        g0337(.A(new_new_n359_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_0_), .B(i_6_), .Y(new_new_n361_));
  NAi21      g0339(.An(i_1_), .B(i_5_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n361_), .Y(new_new_n363_));
  NA2        g0341(.A(new_new_n363_), .B(new_new_n25_), .Y(new_new_n364_));
  OAI210     g0342(.A0(new_new_n364_), .A1(new_new_n162_), .B0(new_new_n254_), .Y(new_new_n365_));
  NAi41      g0343(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n366_));
  OAI220     g0344(.A0(new_new_n366_), .A1(new_new_n362_), .B0(new_new_n227_), .B1(new_new_n162_), .Y(new_new_n367_));
  AOI210     g0345(.A0(new_new_n366_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n368_));
  NOi32      g0346(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n369_));
  NA2        g0347(.A(new_new_n369_), .B(new_new_n46_), .Y(new_new_n370_));
  NO2        g0348(.A(new_new_n370_), .B(i_0_), .Y(new_new_n371_));
  OR3        g0349(.A(new_new_n371_), .B(new_new_n368_), .C(new_new_n367_), .Y(new_new_n372_));
  NO2        g0350(.A(i_1_), .B(new_new_n102_), .Y(new_new_n373_));
  NAi21      g0351(.An(i_3_), .B(i_4_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n374_), .B(i_9_), .Y(new_new_n375_));
  AN2        g0353(.A(i_6_), .B(i_7_), .Y(new_new_n376_));
  OAI210     g0354(.A0(new_new_n376_), .A1(new_new_n373_), .B0(new_new_n375_), .Y(new_new_n377_));
  NA2        g0355(.A(i_2_), .B(i_7_), .Y(new_new_n378_));
  NO2        g0356(.A(new_new_n374_), .B(i_10_), .Y(new_new_n379_));
  NA3        g0357(.A(new_new_n379_), .B(new_new_n378_), .C(new_new_n252_), .Y(new_new_n380_));
  AOI210     g0358(.A0(new_new_n380_), .A1(new_new_n377_), .B0(new_new_n190_), .Y(new_new_n381_));
  AOI210     g0359(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n382_));
  OAI210     g0360(.A0(new_new_n382_), .A1(new_new_n193_), .B0(new_new_n379_), .Y(new_new_n383_));
  AOI220     g0361(.A0(new_new_n379_), .A1(new_new_n341_), .B0(new_new_n246_), .B1(new_new_n193_), .Y(new_new_n384_));
  AOI210     g0362(.A0(new_new_n384_), .A1(new_new_n383_), .B0(i_5_), .Y(new_new_n385_));
  NO4        g0363(.A(new_new_n385_), .B(new_new_n381_), .C(new_new_n372_), .D(new_new_n365_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n386_), .B(new_new_n360_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n388_));
  AN2        g0366(.A(i_12_), .B(i_5_), .Y(new_new_n389_));
  NO2        g0367(.A(i_4_), .B(new_new_n26_), .Y(new_new_n390_));
  NA2        g0368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  NO2        g0369(.A(i_11_), .B(i_6_), .Y(new_new_n392_));
  NA3        g0370(.A(new_new_n392_), .B(new_new_n329_), .C(new_new_n232_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n393_), .B(new_new_n391_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n250_), .B(i_5_), .Y(new_new_n395_));
  NO2        g0373(.A(i_5_), .B(i_10_), .Y(new_new_n396_));
  AOI220     g0374(.A0(new_new_n396_), .A1(new_new_n278_), .B0(new_new_n395_), .B1(new_new_n203_), .Y(new_new_n397_));
  NA2        g0375(.A(new_new_n146_), .B(new_new_n45_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n397_), .Y(new_new_n399_));
  OAI210     g0377(.A0(new_new_n399_), .A1(new_new_n394_), .B0(new_new_n388_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n152_), .B(new_new_n84_), .Y(new_new_n402_));
  OAI210     g0380(.A0(new_new_n402_), .A1(new_new_n394_), .B0(new_new_n401_), .Y(new_new_n403_));
  NO2        g0381(.A(i_11_), .B(i_12_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n396_), .B(new_new_n244_), .Y(new_new_n405_));
  NA3        g0383(.A(new_new_n114_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n406_), .B(new_new_n227_), .Y(new_new_n407_));
  NAi21      g0385(.An(i_13_), .B(i_0_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n407_), .B(i_0_), .Y(new_new_n409_));
  NA3        g0387(.A(new_new_n409_), .B(new_new_n403_), .C(new_new_n400_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n44_), .B(new_new_n232_), .Y(new_new_n411_));
  NO3        g0389(.A(i_1_), .B(i_12_), .C(new_new_n84_), .Y(new_new_n412_));
  NO2        g0390(.A(i_0_), .B(i_11_), .Y(new_new_n413_));
  AN2        g0391(.A(i_1_), .B(i_6_), .Y(new_new_n414_));
  NOi21      g0392(.An(i_2_), .B(i_12_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n415_), .B(new_new_n414_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n416_), .B(new_new_n1079_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n144_), .B(i_9_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n418_), .B(i_4_), .Y(new_new_n419_));
  NA2        g0397(.A(new_new_n417_), .B(new_new_n419_), .Y(new_new_n420_));
  NAi21      g0398(.An(i_9_), .B(i_4_), .Y(new_new_n421_));
  OR2        g0399(.A(i_13_), .B(i_10_), .Y(new_new_n422_));
  NO3        g0400(.A(new_new_n422_), .B(new_new_n119_), .C(new_new_n421_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n176_), .B(new_new_n125_), .Y(new_new_n424_));
  OR2        g0402(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n290_), .B(new_new_n426_), .Y(new_new_n427_));
  INV        g0405(.A(new_new_n216_), .Y(new_new_n428_));
  OAI220     g0406(.A0(new_new_n428_), .A1(new_new_n425_), .B0(new_new_n427_), .B1(new_new_n345_), .Y(new_new_n429_));
  INV        g0407(.A(new_new_n429_), .Y(new_new_n430_));
  AOI210     g0408(.A0(new_new_n430_), .A1(new_new_n420_), .B0(new_new_n26_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n327_), .B(new_new_n326_), .Y(new_new_n432_));
  AOI220     g0410(.A0(new_new_n303_), .A1(new_new_n293_), .B0(new_new_n297_), .B1(i_7_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n433_), .B(new_new_n173_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n187_), .B(new_new_n84_), .Y(new_new_n435_));
  AOI220     g0413(.A0(new_new_n435_), .A1(new_new_n302_), .B0(new_new_n1084_), .B1(new_new_n216_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(i_7_), .Y(new_new_n437_));
  NO3        g0415(.A(new_new_n437_), .B(new_new_n434_), .C(new_new_n432_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n201_), .B(new_new_n97_), .Y(new_new_n439_));
  NA3        g0417(.A(new_new_n329_), .B(new_new_n166_), .C(new_new_n84_), .Y(new_new_n440_));
  AOI210     g0418(.A0(new_new_n440_), .A1(new_new_n439_), .B0(i_8_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n198_), .B(i_10_), .Y(new_new_n442_));
  NA3        g0420(.A(new_new_n263_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n303_), .B(new_new_n242_), .Y(new_new_n444_));
  OAI220     g0422(.A0(new_new_n444_), .A1(new_new_n187_), .B0(new_new_n443_), .B1(new_new_n442_), .Y(new_new_n445_));
  NO2        g0423(.A(i_3_), .B(new_new_n48_), .Y(new_new_n446_));
  NA3        g0424(.A(new_new_n341_), .B(new_new_n340_), .C(new_new_n446_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n320_), .B(new_new_n325_), .Y(new_new_n448_));
  OAI210     g0426(.A0(new_new_n448_), .A1(new_new_n194_), .B0(new_new_n447_), .Y(new_new_n449_));
  NO3        g0427(.A(new_new_n449_), .B(new_new_n445_), .C(new_new_n441_), .Y(new_new_n450_));
  AOI210     g0428(.A0(new_new_n450_), .A1(new_new_n438_), .B0(new_new_n280_), .Y(new_new_n451_));
  NO4        g0429(.A(new_new_n451_), .B(new_new_n431_), .C(new_new_n410_), .D(new_new_n387_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n63_), .B(i_4_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n71_), .B(i_13_), .Y(new_new_n454_));
  NA3        g0432(.A(new_new_n454_), .B(new_new_n453_), .C(i_2_), .Y(new_new_n455_));
  NO2        g0433(.A(i_10_), .B(i_9_), .Y(new_new_n456_));
  NAi21      g0434(.An(i_12_), .B(i_8_), .Y(new_new_n457_));
  NO2        g0435(.A(new_new_n457_), .B(i_3_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n458_), .B(new_new_n456_), .Y(new_new_n459_));
  NO2        g0437(.A(new_new_n46_), .B(i_4_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n460_), .B(new_new_n105_), .Y(new_new_n461_));
  OAI220     g0439(.A0(new_new_n461_), .A1(new_new_n210_), .B0(new_new_n459_), .B1(new_new_n455_), .Y(new_new_n462_));
  NA2        g0440(.A(new_new_n315_), .B(i_0_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n464_));
  NA2        g0442(.A(new_new_n275_), .B(new_new_n98_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n465_), .B(new_new_n464_), .Y(new_new_n466_));
  NA2        g0444(.A(i_8_), .B(i_9_), .Y(new_new_n467_));
  AOI210     g0445(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n468_));
  OR2        g0446(.A(new_new_n468_), .B(new_new_n467_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n290_), .B(new_new_n211_), .Y(new_new_n470_));
  OAI220     g0448(.A0(new_new_n470_), .A1(new_new_n469_), .B0(new_new_n466_), .B1(new_new_n463_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n257_), .B(new_new_n314_), .Y(new_new_n472_));
  NO3        g0450(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n473_));
  INV        g0451(.A(new_new_n473_), .Y(new_new_n474_));
  NA3        g0452(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n475_));
  NA4        g0453(.A(new_new_n147_), .B(new_new_n117_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n476_));
  OAI220     g0454(.A0(new_new_n476_), .A1(new_new_n475_), .B0(new_new_n474_), .B1(new_new_n472_), .Y(new_new_n477_));
  NO3        g0455(.A(new_new_n477_), .B(new_new_n471_), .C(new_new_n462_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n302_), .B(new_new_n109_), .Y(new_new_n479_));
  OR2        g0457(.A(new_new_n479_), .B(i_8_), .Y(new_new_n480_));
  OA210      g0458(.A0(new_new_n354_), .A1(new_new_n102_), .B0(new_new_n304_), .Y(new_new_n481_));
  OA220      g0459(.A0(new_new_n481_), .A1(new_new_n165_), .B0(new_new_n480_), .B1(new_new_n239_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n97_), .B(i_13_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n435_), .B(new_new_n388_), .Y(new_new_n484_));
  NO2        g0462(.A(i_2_), .B(i_13_), .Y(new_new_n485_));
  NA3        g0463(.A(new_new_n485_), .B(new_new_n164_), .C(new_new_n100_), .Y(new_new_n486_));
  OAI220     g0464(.A0(new_new_n486_), .A1(new_new_n244_), .B0(new_new_n484_), .B1(new_new_n483_), .Y(new_new_n487_));
  NO3        g0465(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n488_));
  NO2        g0466(.A(i_6_), .B(i_7_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n71_), .B(i_3_), .Y(new_new_n491_));
  NOi21      g0469(.An(i_2_), .B(i_7_), .Y(new_new_n492_));
  NAi31      g0470(.An(i_11_), .B(new_new_n492_), .C(new_new_n491_), .Y(new_new_n493_));
  NO2        g0471(.A(new_new_n422_), .B(i_6_), .Y(new_new_n494_));
  NA3        g0472(.A(new_new_n494_), .B(new_new_n453_), .C(new_new_n73_), .Y(new_new_n495_));
  NO2        g0473(.A(new_new_n495_), .B(new_new_n493_), .Y(new_new_n496_));
  NO2        g0474(.A(i_3_), .B(new_new_n198_), .Y(new_new_n497_));
  NO2        g0475(.A(i_6_), .B(i_10_), .Y(new_new_n498_));
  NA3        g0476(.A(new_new_n253_), .B(new_new_n175_), .C(new_new_n134_), .Y(new_new_n499_));
  NA2        g0477(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n160_), .B(i_3_), .Y(new_new_n501_));
  NAi31      g0479(.An(new_new_n500_), .B(new_new_n501_), .C(new_new_n233_), .Y(new_new_n502_));
  NA3        g0480(.A(new_new_n401_), .B(new_new_n183_), .C(new_new_n151_), .Y(new_new_n503_));
  NA3        g0481(.A(new_new_n503_), .B(new_new_n502_), .C(new_new_n499_), .Y(new_new_n504_));
  NO3        g0482(.A(new_new_n504_), .B(new_new_n496_), .C(new_new_n487_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n464_), .B(new_new_n389_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n473_), .B(new_new_n396_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n507_), .B(new_new_n231_), .Y(new_new_n508_));
  NAi21      g0486(.An(new_new_n222_), .B(new_new_n404_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n341_), .B(new_new_n224_), .Y(new_new_n510_));
  NO2        g0488(.A(new_new_n26_), .B(i_5_), .Y(new_new_n511_));
  NO2        g0489(.A(i_0_), .B(new_new_n84_), .Y(new_new_n512_));
  NA3        g0490(.A(new_new_n512_), .B(new_new_n511_), .C(new_new_n144_), .Y(new_new_n513_));
  OAI220     g0491(.A0(new_new_n38_), .A1(new_new_n513_), .B0(new_new_n510_), .B1(new_new_n509_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n27_), .B(i_10_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n319_), .B(new_new_n246_), .Y(new_new_n516_));
  OAI220     g0494(.A0(new_new_n516_), .A1(new_new_n443_), .B0(new_new_n515_), .B1(new_new_n483_), .Y(new_new_n517_));
  NA4        g0495(.A(new_new_n312_), .B(new_new_n230_), .C(new_new_n71_), .D(new_new_n244_), .Y(new_new_n518_));
  NO2        g0496(.A(new_new_n518_), .B(new_new_n490_), .Y(new_new_n519_));
  NO4        g0497(.A(new_new_n519_), .B(new_new_n517_), .C(new_new_n514_), .D(new_new_n508_), .Y(new_new_n520_));
  NA4        g0498(.A(new_new_n520_), .B(new_new_n505_), .C(new_new_n482_), .D(new_new_n478_), .Y(new_new_n521_));
  NA3        g0499(.A(new_new_n312_), .B(new_new_n180_), .C(new_new_n178_), .Y(new_new_n522_));
  OAI210     g0500(.A0(new_new_n308_), .A1(new_new_n185_), .B0(new_new_n522_), .Y(new_new_n523_));
  AN2        g0501(.A(new_new_n293_), .B(new_new_n241_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n524_), .B(new_new_n523_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n319_), .B(new_new_n167_), .Y(new_new_n526_));
  OAI210     g0504(.A0(new_new_n526_), .A1(new_new_n239_), .B0(new_new_n313_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n527_), .B(new_new_n328_), .Y(new_new_n528_));
  NA4        g0506(.A(new_new_n454_), .B(new_new_n453_), .C(new_new_n208_), .D(i_2_), .Y(new_new_n529_));
  INV        g0507(.A(new_new_n529_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n389_), .B(new_new_n232_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n359_), .B(new_new_n71_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n376_), .B(new_new_n369_), .Y(new_new_n533_));
  AO210      g0511(.A0(new_new_n532_), .A1(new_new_n531_), .B0(new_new_n533_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n36_), .B(i_8_), .Y(new_new_n535_));
  INV        g0513(.A(new_new_n423_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n536_), .B(new_new_n534_), .Y(new_new_n537_));
  AOI210     g0515(.A0(new_new_n530_), .A1(new_new_n209_), .B0(new_new_n537_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n539_));
  OAI210     g0517(.A0(i_8_), .A1(new_new_n539_), .B0(new_new_n136_), .Y(new_new_n540_));
  AOI210     g0518(.A0(new_new_n199_), .A1(i_9_), .B0(new_new_n274_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n541_), .B(new_new_n204_), .Y(new_new_n542_));
  AOI220     g0520(.A0(i_6_), .A1(new_new_n542_), .B0(new_new_n540_), .B1(new_new_n424_), .Y(new_new_n543_));
  NA4        g0521(.A(new_new_n543_), .B(new_new_n538_), .C(new_new_n528_), .D(new_new_n525_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n395_), .B(new_new_n302_), .Y(new_new_n545_));
  OAI210     g0523(.A0(new_new_n391_), .A1(new_new_n172_), .B0(new_new_n545_), .Y(new_new_n546_));
  NO2        g0524(.A(i_12_), .B(new_new_n198_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n498_), .B(new_new_n178_), .C(new_new_n27_), .Y(new_new_n548_));
  NO3        g0526(.A(new_new_n548_), .B(i_13_), .C(new_new_n479_), .Y(new_new_n549_));
  NOi21      g0527(.An(new_new_n320_), .B(new_new_n38_), .Y(new_new_n550_));
  OAI210     g0528(.A0(new_new_n550_), .A1(new_new_n549_), .B0(new_new_n546_), .Y(new_new_n551_));
  NO2        g0529(.A(i_8_), .B(i_7_), .Y(new_new_n552_));
  OAI210     g0530(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n553_), .B(new_new_n230_), .Y(new_new_n554_));
  AOI220     g0532(.A0(new_new_n329_), .A1(new_new_n39_), .B0(new_new_n242_), .B1(new_new_n212_), .Y(new_new_n555_));
  OAI220     g0533(.A0(new_new_n555_), .A1(i_4_), .B0(new_new_n554_), .B1(new_new_n250_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n44_), .B(i_10_), .Y(new_new_n557_));
  NO2        g0535(.A(new_new_n557_), .B(i_6_), .Y(new_new_n558_));
  NA3        g0536(.A(new_new_n558_), .B(new_new_n556_), .C(new_new_n552_), .Y(new_new_n559_));
  AOI220     g0537(.A0(new_new_n435_), .A1(new_new_n329_), .B0(new_new_n255_), .B1(new_new_n252_), .Y(new_new_n560_));
  OAI220     g0538(.A0(new_new_n560_), .A1(new_new_n271_), .B0(new_new_n483_), .B1(new_new_n135_), .Y(new_new_n561_));
  NA2        g0539(.A(new_new_n561_), .B(new_new_n274_), .Y(new_new_n562_));
  NOi31      g0540(.An(new_new_n297_), .B(new_new_n308_), .C(new_new_n185_), .Y(new_new_n563_));
  NA3        g0541(.A(new_new_n312_), .B(new_new_n178_), .C(new_new_n97_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n228_), .B(new_new_n44_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n160_), .B(i_5_), .Y(new_new_n566_));
  NA3        g0544(.A(new_new_n566_), .B(new_new_n411_), .C(new_new_n323_), .Y(new_new_n567_));
  OAI210     g0545(.A0(new_new_n567_), .A1(new_new_n565_), .B0(new_new_n564_), .Y(new_new_n568_));
  OAI210     g0546(.A0(new_new_n568_), .A1(new_new_n563_), .B0(new_new_n473_), .Y(new_new_n569_));
  NA4        g0547(.A(new_new_n569_), .B(new_new_n562_), .C(new_new_n559_), .D(new_new_n551_), .Y(new_new_n570_));
  NA3        g0548(.A(new_new_n224_), .B(new_new_n69_), .C(new_new_n44_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n290_), .B(new_new_n82_), .Y(new_new_n572_));
  AOI210     g0550(.A0(new_new_n571_), .A1(new_new_n349_), .B0(new_new_n572_), .Y(new_new_n573_));
  NA2        g0551(.A(new_new_n303_), .B(new_new_n293_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n574_), .B(new_new_n177_), .Y(new_new_n575_));
  NA2        g0553(.A(new_new_n230_), .B(new_new_n229_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n456_), .B(new_new_n228_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n576_), .B(new_new_n577_), .Y(new_new_n578_));
  NA2        g0556(.A(i_0_), .B(new_new_n48_), .Y(new_new_n579_));
  NA3        g0557(.A(new_new_n547_), .B(new_new_n283_), .C(new_new_n579_), .Y(new_new_n580_));
  INV        g0558(.A(new_new_n580_), .Y(new_new_n581_));
  NO4        g0559(.A(new_new_n581_), .B(new_new_n578_), .C(new_new_n575_), .D(new_new_n573_), .Y(new_new_n582_));
  NO4        g0560(.A(new_new_n258_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n583_));
  NO3        g0561(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n240_), .B(new_new_n36_), .Y(new_new_n585_));
  AN2        g0563(.A(new_new_n585_), .B(new_new_n584_), .Y(new_new_n586_));
  OA210      g0564(.A0(new_new_n586_), .A1(new_new_n583_), .B0(new_new_n359_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n422_), .B(i_1_), .Y(new_new_n588_));
  NOi31      g0566(.An(new_new_n588_), .B(new_new_n465_), .C(new_new_n71_), .Y(new_new_n589_));
  AN3        g0567(.A(new_new_n589_), .B(new_new_n419_), .C(i_2_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n433_), .B(new_new_n181_), .Y(new_new_n591_));
  NO3        g0569(.A(new_new_n591_), .B(new_new_n590_), .C(new_new_n587_), .Y(new_new_n592_));
  NOi21      g0570(.An(i_10_), .B(i_6_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n84_), .B(new_new_n25_), .Y(new_new_n594_));
  AOI220     g0572(.A0(new_new_n290_), .A1(new_new_n594_), .B0(new_new_n283_), .B1(new_new_n593_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n595_), .B(new_new_n463_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n597_));
  NA2        g0575(.A(new_new_n320_), .B(new_new_n167_), .Y(new_new_n598_));
  AOI220     g0576(.A0(new_new_n598_), .A1(new_new_n444_), .B0(new_new_n188_), .B1(new_new_n186_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n203_), .B(new_new_n37_), .Y(new_new_n600_));
  NOi31      g0578(.An(new_new_n148_), .B(new_new_n600_), .C(new_new_n337_), .Y(new_new_n601_));
  NO3        g0579(.A(new_new_n601_), .B(new_new_n599_), .C(new_new_n596_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n532_), .B(new_new_n384_), .Y(new_new_n603_));
  INV        g0581(.A(new_new_n323_), .Y(new_new_n604_));
  NO2        g0582(.A(i_12_), .B(new_new_n84_), .Y(new_new_n605_));
  NA3        g0583(.A(new_new_n392_), .B(new_new_n290_), .C(new_new_n224_), .Y(new_new_n606_));
  NO2        g0584(.A(new_new_n606_), .B(new_new_n604_), .Y(new_new_n607_));
  NA2        g0585(.A(new_new_n178_), .B(i_0_), .Y(new_new_n608_));
  NO3        g0586(.A(new_new_n608_), .B(new_new_n1081_), .C(new_new_n308_), .Y(new_new_n609_));
  OR2        g0587(.A(i_2_), .B(i_5_), .Y(new_new_n610_));
  OR2        g0588(.A(new_new_n610_), .B(new_new_n414_), .Y(new_new_n611_));
  NO2        g0589(.A(new_new_n252_), .B(new_new_n203_), .Y(new_new_n612_));
  AOI210     g0590(.A0(new_new_n612_), .A1(new_new_n611_), .B0(new_new_n509_), .Y(new_new_n613_));
  NO4        g0591(.A(new_new_n613_), .B(new_new_n609_), .C(new_new_n607_), .D(new_new_n603_), .Y(new_new_n614_));
  NA4        g0592(.A(new_new_n614_), .B(new_new_n602_), .C(new_new_n592_), .D(new_new_n582_), .Y(new_new_n615_));
  NO4        g0593(.A(new_new_n615_), .B(new_new_n570_), .C(new_new_n544_), .D(new_new_n521_), .Y(new_new_n616_));
  NA4        g0594(.A(new_new_n616_), .B(new_new_n452_), .C(new_new_n358_), .D(new_new_n318_), .Y(men7));
  NO2        g0595(.A(new_new_n93_), .B(new_new_n54_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n109_), .B(new_new_n90_), .Y(new_new_n619_));
  NA2        g0597(.A(new_new_n390_), .B(new_new_n619_), .Y(new_new_n620_));
  NA2        g0598(.A(new_new_n498_), .B(new_new_n82_), .Y(new_new_n621_));
  NA2        g0599(.A(i_11_), .B(new_new_n198_), .Y(new_new_n622_));
  INV        g0600(.A(new_new_n620_), .Y(new_new_n623_));
  NA3        g0601(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n244_), .B(i_4_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n625_), .B(i_8_), .Y(new_new_n626_));
  AOI210     g0604(.A0(new_new_n626_), .A1(new_new_n106_), .B0(new_new_n624_), .Y(new_new_n627_));
  NA2        g0605(.A(i_2_), .B(new_new_n84_), .Y(new_new_n628_));
  OAI210     g0606(.A0(new_new_n87_), .A1(new_new_n208_), .B0(new_new_n209_), .Y(new_new_n629_));
  NO2        g0607(.A(i_7_), .B(new_new_n37_), .Y(new_new_n630_));
  NA2        g0608(.A(i_4_), .B(i_8_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n312_), .B(new_new_n630_), .Y(new_new_n632_));
  OAI220     g0610(.A0(new_new_n632_), .A1(new_new_n628_), .B0(new_new_n629_), .B1(i_13_), .Y(new_new_n633_));
  NO4        g0611(.A(new_new_n633_), .B(new_new_n627_), .C(new_new_n623_), .D(new_new_n618_), .Y(new_new_n634_));
  AOI210     g0612(.A0(new_new_n130_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n635_));
  AOI210     g0613(.A0(new_new_n635_), .A1(new_new_n244_), .B0(new_new_n164_), .Y(new_new_n636_));
  OR2        g0614(.A(i_6_), .B(i_10_), .Y(new_new_n637_));
  NO2        g0615(.A(new_new_n637_), .B(new_new_n23_), .Y(new_new_n638_));
  OR3        g0616(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n639_));
  NO3        g0617(.A(new_new_n639_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n640_));
  INV        g0618(.A(new_new_n205_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n640_), .B(new_new_n638_), .Y(new_new_n642_));
  OA220      g0620(.A0(new_new_n642_), .A1(new_new_n604_), .B0(new_new_n636_), .B1(new_new_n276_), .Y(new_new_n643_));
  AOI210     g0621(.A0(new_new_n643_), .A1(new_new_n634_), .B0(new_new_n63_), .Y(new_new_n644_));
  NOi21      g0622(.An(i_11_), .B(i_7_), .Y(new_new_n645_));
  AO210      g0623(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n647_), .B(new_new_n212_), .Y(new_new_n648_));
  NA3        g0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n649_));
  NAi21      g0627(.An(new_new_n649_), .B(i_11_), .Y(new_new_n650_));
  AOI210     g0628(.A0(new_new_n650_), .A1(new_new_n648_), .B0(new_new_n63_), .Y(new_new_n651_));
  NA2        g0629(.A(new_new_n86_), .B(new_new_n63_), .Y(new_new_n652_));
  AO210      g0630(.A0(new_new_n652_), .A1(new_new_n384_), .B0(new_new_n40_), .Y(new_new_n653_));
  NO3        g0631(.A(new_new_n265_), .B(new_new_n213_), .C(new_new_n622_), .Y(new_new_n654_));
  OAI210     g0632(.A0(new_new_n654_), .A1(new_new_n233_), .B0(new_new_n63_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n415_), .B(new_new_n31_), .Y(new_new_n656_));
  OR2        g0634(.A(new_new_n213_), .B(new_new_n109_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(new_new_n656_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n63_), .B(i_9_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n659_), .B(i_4_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n660_), .B(new_new_n658_), .Y(new_new_n661_));
  NO2        g0639(.A(i_1_), .B(i_12_), .Y(new_new_n662_));
  NA3        g0640(.A(new_new_n662_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n663_));
  NA4        g0641(.A(new_new_n663_), .B(new_new_n661_), .C(new_new_n655_), .D(new_new_n653_), .Y(new_new_n664_));
  OAI210     g0642(.A0(new_new_n664_), .A1(new_new_n651_), .B0(i_6_), .Y(new_new_n665_));
  OAI210     g0643(.A0(new_new_n649_), .A1(new_new_n109_), .B0(new_new_n475_), .Y(new_new_n666_));
  NA2        g0644(.A(new_new_n666_), .B(new_new_n605_), .Y(new_new_n667_));
  NO2        g0645(.A(i_6_), .B(i_11_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n667_), .B(new_new_n466_), .Y(new_new_n669_));
  NO4        g0647(.A(new_new_n221_), .B(new_new_n130_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n670_));
  NA2        g0648(.A(new_new_n670_), .B(new_new_n659_), .Y(new_new_n671_));
  NO3        g0649(.A(new_new_n637_), .B(new_new_n240_), .C(new_new_n23_), .Y(new_new_n672_));
  AOI210     g0650(.A0(i_1_), .A1(new_new_n266_), .B0(new_new_n672_), .Y(new_new_n673_));
  OAI210     g0651(.A0(new_new_n673_), .A1(new_new_n44_), .B0(new_new_n671_), .Y(new_new_n674_));
  NA3        g0652(.A(new_new_n552_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n140_), .B(i_9_), .Y(new_new_n676_));
  NA3        g0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n46_), .B(i_1_), .Y(new_new_n678_));
  NA3        g0656(.A(new_new_n678_), .B(new_new_n275_), .C(new_new_n44_), .Y(new_new_n679_));
  OAI220     g0657(.A0(new_new_n679_), .A1(new_new_n677_), .B0(new_new_n676_), .B1(new_new_n1078_), .Y(new_new_n680_));
  NA3        g0658(.A(new_new_n659_), .B(new_new_n323_), .C(i_6_), .Y(new_new_n681_));
  NAi21      g0659(.An(new_new_n675_), .B(new_new_n92_), .Y(new_new_n682_));
  NA2        g0660(.A(new_new_n678_), .B(new_new_n275_), .Y(new_new_n683_));
  NO2        g0661(.A(i_11_), .B(new_new_n37_), .Y(new_new_n684_));
  NA2        g0662(.A(new_new_n684_), .B(new_new_n24_), .Y(new_new_n685_));
  OAI210     g0663(.A0(new_new_n685_), .A1(new_new_n683_), .B0(new_new_n682_), .Y(new_new_n686_));
  OR2        g0664(.A(new_new_n686_), .B(new_new_n680_), .Y(new_new_n687_));
  NO3        g0665(.A(new_new_n687_), .B(new_new_n674_), .C(new_new_n669_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n244_), .B(new_new_n102_), .Y(new_new_n689_));
  NO2        g0667(.A(new_new_n689_), .B(new_new_n645_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n421_), .B(new_new_n84_), .Y(new_new_n691_));
  NA2        g0669(.A(i_3_), .B(new_new_n198_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n692_), .B(new_new_n116_), .Y(new_new_n693_));
  AN2        g0671(.A(new_new_n693_), .B(new_new_n558_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n240_), .B(new_new_n44_), .Y(new_new_n695_));
  NO3        g0673(.A(new_new_n695_), .B(new_new_n315_), .C(new_new_n245_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n697_), .B(i_6_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n84_), .B(i_9_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n699_), .B(new_new_n63_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n700_), .B(new_new_n662_), .Y(new_new_n701_));
  NO4        g0679(.A(new_new_n701_), .B(new_new_n698_), .C(new_new_n696_), .D(i_4_), .Y(new_new_n702_));
  NA2        g0680(.A(i_1_), .B(i_3_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n467_), .B(new_new_n93_), .Y(new_new_n704_));
  AOI210     g0682(.A0(new_new_n695_), .A1(new_new_n593_), .B0(new_new_n704_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n703_), .Y(new_new_n706_));
  NO3        g0684(.A(new_new_n706_), .B(new_new_n702_), .C(new_new_n694_), .Y(new_new_n707_));
  NA3        g0685(.A(new_new_n707_), .B(new_new_n688_), .C(new_new_n665_), .Y(new_new_n708_));
  NO3        g0686(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n709_));
  NOi21      g0687(.An(new_new_n709_), .B(i_10_), .Y(new_new_n710_));
  OA210      g0688(.A0(new_new_n710_), .A1(new_new_n253_), .B0(new_new_n84_), .Y(new_new_n711_));
  NA2        g0689(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n712_));
  NA3        g0690(.A(new_new_n498_), .B(new_new_n535_), .C(new_new_n46_), .Y(new_new_n713_));
  NO3        g0691(.A(new_new_n492_), .B(new_new_n631_), .C(new_new_n84_), .Y(new_new_n714_));
  NA2        g0692(.A(new_new_n714_), .B(new_new_n25_), .Y(new_new_n715_));
  NA3        g0693(.A(new_new_n715_), .B(new_new_n713_), .C(new_new_n712_), .Y(new_new_n716_));
  OAI210     g0694(.A0(new_new_n716_), .A1(new_new_n711_), .B0(i_1_), .Y(new_new_n717_));
  INV        g0695(.A(i_1_), .Y(new_new_n718_));
  NO2        g0696(.A(new_new_n374_), .B(i_2_), .Y(new_new_n719_));
  AOI210     g0697(.A0(new_new_n681_), .A1(new_new_n717_), .B0(i_13_), .Y(new_new_n720_));
  OR2        g0698(.A(i_11_), .B(i_7_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n107_), .B(new_new_n140_), .Y(new_new_n722_));
  AOI220     g0700(.A0(new_new_n485_), .A1(new_new_n164_), .B0(new_new_n460_), .B1(new_new_n140_), .Y(new_new_n723_));
  OAI210     g0701(.A0(new_new_n723_), .A1(new_new_n44_), .B0(new_new_n722_), .Y(new_new_n724_));
  NO2        g0702(.A(new_new_n492_), .B(new_new_n24_), .Y(new_new_n725_));
  AOI220     g0703(.A0(new_new_n725_), .A1(new_new_n691_), .B0(new_new_n253_), .B1(new_new_n133_), .Y(new_new_n726_));
  NO2        g0704(.A(new_new_n726_), .B(new_new_n40_), .Y(new_new_n727_));
  AOI210     g0705(.A0(new_new_n724_), .A1(new_new_n339_), .B0(new_new_n727_), .Y(new_new_n728_));
  AOI220     g0706(.A0(i_7_), .A1(new_new_n70_), .B0(new_new_n392_), .B1(new_new_n678_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n729_), .B(new_new_n250_), .Y(new_new_n730_));
  AOI210     g0708(.A0(new_new_n457_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n731_));
  NOi31      g0709(.An(new_new_n731_), .B(new_new_n621_), .C(new_new_n44_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n129_), .B(i_13_), .Y(new_new_n733_));
  NO2        g0711(.A(new_new_n677_), .B(new_new_n116_), .Y(new_new_n734_));
  INV        g0712(.A(new_new_n734_), .Y(new_new_n735_));
  OAI220     g0713(.A0(new_new_n735_), .A1(new_new_n69_), .B0(new_new_n733_), .B1(new_new_n718_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n102_), .Y(new_new_n737_));
  NA2        g0715(.A(new_new_n26_), .B(new_new_n198_), .Y(new_new_n738_));
  INV        g0716(.A(i_7_), .Y(new_new_n739_));
  INV        g0717(.A(new_new_n737_), .Y(new_new_n740_));
  AOI220     g0718(.A0(new_new_n392_), .A1(new_new_n678_), .B0(new_new_n92_), .B1(new_new_n103_), .Y(new_new_n741_));
  OAI220     g0719(.A0(new_new_n741_), .A1(new_new_n626_), .B0(new_new_n740_), .B1(new_new_n641_), .Y(new_new_n742_));
  NO4        g0720(.A(new_new_n742_), .B(new_new_n736_), .C(new_new_n732_), .D(new_new_n730_), .Y(new_new_n743_));
  OR2        g0721(.A(i_11_), .B(i_6_), .Y(new_new_n744_));
  NO2        g0722(.A(new_new_n735_), .B(new_new_n744_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n668_), .B(i_13_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n103_), .B(new_new_n738_), .Y(new_new_n747_));
  NAi21      g0725(.An(i_11_), .B(i_12_), .Y(new_new_n748_));
  NO3        g0726(.A(new_new_n748_), .B(i_13_), .C(new_new_n84_), .Y(new_new_n749_));
  NO3        g0727(.A(new_new_n492_), .B(new_new_n605_), .C(new_new_n631_), .Y(new_new_n750_));
  AOI220     g0728(.A0(new_new_n750_), .A1(new_new_n319_), .B0(new_new_n749_), .B1(new_new_n747_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n751_), .B(new_new_n746_), .Y(new_new_n752_));
  OAI210     g0730(.A0(new_new_n752_), .A1(new_new_n745_), .B0(new_new_n63_), .Y(new_new_n753_));
  NO2        g0731(.A(i_2_), .B(i_12_), .Y(new_new_n754_));
  OAI210     g0732(.A0(new_new_n635_), .A1(new_new_n373_), .B0(new_new_n754_), .Y(new_new_n755_));
  NA2        g0733(.A(i_8_), .B(new_new_n25_), .Y(new_new_n756_));
  NO3        g0734(.A(new_new_n756_), .B(new_new_n390_), .C(new_new_n625_), .Y(new_new_n757_));
  OAI210     g0735(.A0(new_new_n757_), .A1(new_new_n375_), .B0(new_new_n373_), .Y(new_new_n758_));
  NO2        g0736(.A(new_new_n130_), .B(i_2_), .Y(new_new_n759_));
  NA2        g0737(.A(new_new_n759_), .B(new_new_n662_), .Y(new_new_n760_));
  NA3        g0738(.A(new_new_n760_), .B(new_new_n758_), .C(new_new_n755_), .Y(new_new_n761_));
  NA3        g0739(.A(new_new_n761_), .B(new_new_n45_), .C(new_new_n232_), .Y(new_new_n762_));
  NA4        g0740(.A(new_new_n762_), .B(new_new_n753_), .C(new_new_n743_), .D(new_new_n728_), .Y(new_new_n763_));
  OR4        g0741(.A(new_new_n763_), .B(new_new_n720_), .C(new_new_n708_), .D(new_new_n644_), .Y(men5));
  AOI210     g0742(.A0(new_new_n690_), .A1(new_new_n278_), .B0(new_new_n424_), .Y(new_new_n765_));
  AO210      g0743(.A0(new_new_n24_), .A1(i_10_), .B0(new_new_n257_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n754_), .C(new_new_n109_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n767_), .B(new_new_n765_), .Y(new_new_n768_));
  NO3        g0746(.A(i_11_), .B(new_new_n244_), .C(i_13_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n770_));
  NA2        g0748(.A(i_12_), .B(i_8_), .Y(new_new_n771_));
  INV        g0749(.A(new_new_n456_), .Y(new_new_n772_));
  AOI220     g0750(.A0(new_new_n323_), .A1(new_new_n597_), .B0(i_12_), .B1(new_new_n770_), .Y(new_new_n773_));
  INV        g0751(.A(new_new_n773_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n774_), .B(new_new_n768_), .Y(new_new_n775_));
  INV        g0753(.A(new_new_n175_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n253_), .Y(new_new_n777_));
  OAI210     g0755(.A0(new_new_n719_), .A1(new_new_n458_), .B0(new_new_n112_), .Y(new_new_n778_));
  AOI210     g0756(.A0(new_new_n778_), .A1(new_new_n777_), .B0(new_new_n776_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n467_), .B(new_new_n26_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n780_), .B(new_new_n426_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n781_), .B(i_2_), .Y(new_new_n782_));
  INV        g0760(.A(new_new_n782_), .Y(new_new_n783_));
  AOI210     g0761(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n422_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n784_), .A1(new_new_n783_), .B0(new_new_n779_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n195_), .B(new_new_n127_), .Y(new_new_n786_));
  OAI210     g0764(.A0(new_new_n786_), .A1(new_new_n770_), .B0(i_2_), .Y(new_new_n787_));
  INV        g0765(.A(new_new_n176_), .Y(new_new_n788_));
  NO3        g0766(.A(new_new_n646_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n789_));
  AOI210     g0767(.A0(new_new_n788_), .A1(new_new_n87_), .B0(new_new_n789_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n790_), .A1(new_new_n787_), .B0(new_new_n198_), .Y(new_new_n791_));
  OA210      g0769(.A0(new_new_n647_), .A1(new_new_n128_), .B0(i_13_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n205_), .B(new_new_n208_), .Y(new_new_n793_));
  INV        g0771(.A(new_new_n154_), .Y(new_new_n794_));
  AOI210     g0772(.A0(new_new_n794_), .A1(new_new_n793_), .B0(new_new_n378_), .Y(new_new_n795_));
  AOI210     g0773(.A0(new_new_n213_), .A1(new_new_n150_), .B0(new_new_n535_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n796_), .B(new_new_n426_), .Y(new_new_n797_));
  NA3        g0775(.A(new_new_n312_), .B(new_new_n126_), .C(new_new_n42_), .Y(new_new_n798_));
  OAI210     g0776(.A0(new_new_n798_), .A1(new_new_n46_), .B0(new_new_n797_), .Y(new_new_n799_));
  NO4        g0777(.A(new_new_n799_), .B(new_new_n795_), .C(new_new_n792_), .D(new_new_n791_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n62_), .B(i_12_), .Y(new_new_n801_));
  NO2        g0779(.A(new_new_n801_), .B(new_new_n128_), .Y(new_new_n802_));
  NO2        g0780(.A(new_new_n802_), .B(new_new_n622_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n803_), .B(new_new_n36_), .Y(new_new_n804_));
  NA4        g0782(.A(new_new_n804_), .B(new_new_n800_), .C(new_new_n785_), .D(new_new_n775_), .Y(men6));
  NA2        g0783(.A(new_new_n25_), .B(new_new_n759_), .Y(new_new_n806_));
  NA4        g0784(.A(new_new_n396_), .B(new_new_n497_), .C(new_new_n69_), .D(new_new_n102_), .Y(new_new_n807_));
  INV        g0785(.A(new_new_n807_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n227_), .B(new_new_n500_), .Y(new_new_n809_));
  NO2        g0787(.A(i_11_), .B(i_9_), .Y(new_new_n810_));
  NO2        g0788(.A(new_new_n808_), .B(new_new_n334_), .Y(new_new_n811_));
  AO210      g0789(.A0(new_new_n811_), .A1(new_new_n806_), .B0(i_12_), .Y(new_new_n812_));
  NA2        g0790(.A(new_new_n379_), .B(new_new_n341_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n605_), .B(new_new_n63_), .Y(new_new_n814_));
  NA2        g0792(.A(new_new_n710_), .B(new_new_n69_), .Y(new_new_n815_));
  NA4        g0793(.A(new_new_n652_), .B(new_new_n815_), .C(new_new_n814_), .D(new_new_n813_), .Y(new_new_n816_));
  INV        g0794(.A(new_new_n202_), .Y(new_new_n817_));
  AOI220     g0795(.A0(new_new_n817_), .A1(new_new_n810_), .B0(new_new_n816_), .B1(new_new_n71_), .Y(new_new_n818_));
  INV        g0796(.A(new_new_n333_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n73_), .B(new_new_n133_), .Y(new_new_n820_));
  INV        g0798(.A(new_new_n126_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n821_), .B(new_new_n46_), .Y(new_new_n822_));
  AOI210     g0800(.A0(new_new_n822_), .A1(new_new_n820_), .B0(new_new_n819_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n1083_), .B(new_new_n801_), .Y(new_new_n824_));
  AOI210     g0802(.A0(new_new_n824_), .A1(new_new_n533_), .B0(new_new_n190_), .Y(new_new_n825_));
  NO2        g0803(.A(new_new_n32_), .B(i_11_), .Y(new_new_n826_));
  NA3        g0804(.A(new_new_n826_), .B(new_new_n489_), .C(new_new_n396_), .Y(new_new_n827_));
  OAI210     g0805(.A0(new_new_n709_), .A1(new_new_n585_), .B0(new_new_n584_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n828_), .B(new_new_n827_), .Y(new_new_n829_));
  OR3        g0807(.A(new_new_n829_), .B(new_new_n825_), .C(new_new_n823_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n721_), .B(i_2_), .Y(new_new_n831_));
  NA2        g0809(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n832_));
  OAI210     g0810(.A0(new_new_n832_), .A1(new_new_n414_), .B0(new_new_n364_), .Y(new_new_n833_));
  NA2        g0811(.A(new_new_n833_), .B(new_new_n831_), .Y(new_new_n834_));
  NA3        g0812(.A(new_new_n353_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n835_));
  BUFFER     g0813(.A(new_new_n458_), .Y(new_new_n836_));
  NA3        g0814(.A(new_new_n836_), .B(new_new_n149_), .C(new_new_n68_), .Y(new_new_n837_));
  AO210      g0815(.A0(new_new_n507_), .A1(new_new_n772_), .B0(new_new_n36_), .Y(new_new_n838_));
  NA4        g0816(.A(new_new_n838_), .B(new_new_n837_), .C(new_new_n835_), .D(new_new_n834_), .Y(new_new_n839_));
  OAI210     g0817(.A0(i_6_), .A1(i_11_), .B0(new_new_n85_), .Y(new_new_n840_));
  AOI220     g0818(.A0(new_new_n840_), .A1(new_new_n584_), .B0(new_new_n809_), .B1(new_new_n739_), .Y(new_new_n841_));
  NA3        g0819(.A(new_new_n378_), .B(new_new_n246_), .C(new_new_n149_), .Y(new_new_n842_));
  NA3        g0820(.A(new_new_n842_), .B(new_new_n841_), .C(new_new_n629_), .Y(new_new_n843_));
  AO210      g0821(.A0(new_new_n535_), .A1(new_new_n46_), .B0(new_new_n86_), .Y(new_new_n844_));
  NA3        g0822(.A(new_new_n844_), .B(new_new_n498_), .C(new_new_n224_), .Y(new_new_n845_));
  INV        g0823(.A(new_new_n583_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n637_), .B(new_new_n103_), .Y(new_new_n847_));
  OAI210     g0825(.A0(new_new_n847_), .A1(new_new_n113_), .B0(new_new_n413_), .Y(new_new_n848_));
  INV        g0826(.A(new_new_n611_), .Y(new_new_n849_));
  NA3        g0827(.A(new_new_n849_), .B(new_new_n333_), .C(i_7_), .Y(new_new_n850_));
  NA4        g0828(.A(new_new_n850_), .B(new_new_n848_), .C(new_new_n846_), .D(new_new_n845_), .Y(new_new_n851_));
  NO4        g0829(.A(new_new_n851_), .B(new_new_n843_), .C(new_new_n839_), .D(new_new_n830_), .Y(new_new_n852_));
  NA4        g0830(.A(new_new_n852_), .B(new_new_n818_), .C(new_new_n812_), .D(new_new_n386_), .Y(men3));
  NA2        g0831(.A(i_6_), .B(i_7_), .Y(new_new_n854_));
  NO2        g0832(.A(new_new_n854_), .B(i_0_), .Y(new_new_n855_));
  NO2        g0833(.A(i_11_), .B(new_new_n244_), .Y(new_new_n856_));
  OAI210     g0834(.A0(new_new_n855_), .A1(new_new_n297_), .B0(new_new_n856_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n857_), .B(new_new_n198_), .Y(new_new_n858_));
  NO3        g0836(.A(new_new_n463_), .B(new_new_n90_), .C(new_new_n44_), .Y(new_new_n859_));
  OA210      g0837(.A0(new_new_n859_), .A1(new_new_n858_), .B0(new_new_n178_), .Y(new_new_n860_));
  NA3        g0838(.A(new_new_n842_), .B(new_new_n629_), .C(new_new_n377_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n861_), .B(new_new_n39_), .Y(new_new_n862_));
  NOi21      g0840(.An(new_new_n97_), .B(new_new_n781_), .Y(new_new_n863_));
  NO3        g0841(.A(new_new_n657_), .B(new_new_n467_), .C(new_new_n133_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n415_), .B(new_new_n45_), .Y(new_new_n865_));
  AN2        g0843(.A(new_new_n465_), .B(new_new_n55_), .Y(new_new_n866_));
  NO3        g0844(.A(new_new_n866_), .B(new_new_n864_), .C(new_new_n863_), .Y(new_new_n867_));
  AOI210     g0845(.A0(new_new_n867_), .A1(new_new_n862_), .B0(new_new_n48_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n731_), .B(new_new_n699_), .Y(new_new_n869_));
  NA2        g0847(.A(i_0_), .B(new_new_n446_), .Y(new_new_n870_));
  NO2        g0848(.A(new_new_n870_), .B(new_new_n869_), .Y(new_new_n871_));
  NOi21      g0849(.An(i_5_), .B(i_9_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n872_), .B(new_new_n454_), .Y(new_new_n873_));
  INV        g0851(.A(new_new_n714_), .Y(new_new_n874_));
  NO3        g0852(.A(new_new_n418_), .B(new_new_n275_), .C(new_new_n71_), .Y(new_new_n875_));
  NO2        g0853(.A(new_new_n179_), .B(new_new_n150_), .Y(new_new_n876_));
  AOI210     g0854(.A0(new_new_n876_), .A1(new_new_n252_), .B0(new_new_n875_), .Y(new_new_n877_));
  OAI220     g0855(.A0(new_new_n877_), .A1(new_new_n185_), .B0(new_new_n874_), .B1(new_new_n873_), .Y(new_new_n878_));
  NO4        g0856(.A(new_new_n878_), .B(new_new_n871_), .C(new_new_n868_), .D(new_new_n860_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n190_), .B(new_new_n24_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n697_), .B(new_new_n619_), .Y(new_new_n881_));
  NO2        g0859(.A(new_new_n881_), .B(new_new_n880_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n319_), .B(new_new_n131_), .Y(new_new_n883_));
  NAi21      g0861(.An(new_new_n165_), .B(new_new_n446_), .Y(new_new_n884_));
  OAI220     g0862(.A0(new_new_n884_), .A1(i_2_), .B0(new_new_n883_), .B1(new_new_n405_), .Y(new_new_n885_));
  NO2        g0863(.A(new_new_n885_), .B(new_new_n882_), .Y(new_new_n886_));
  NO2        g0864(.A(new_new_n396_), .B(new_new_n301_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n887_), .B(new_new_n734_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n594_), .B(i_0_), .Y(new_new_n889_));
  NO3        g0867(.A(new_new_n889_), .B(new_new_n391_), .C(new_new_n87_), .Y(new_new_n890_));
  NO4        g0868(.A(new_new_n610_), .B(new_new_n221_), .C(new_new_n422_), .D(new_new_n414_), .Y(new_new_n891_));
  AOI210     g0869(.A0(new_new_n891_), .A1(i_11_), .B0(new_new_n890_), .Y(new_new_n892_));
  AN2        g0870(.A(new_new_n97_), .B(new_new_n251_), .Y(new_new_n893_));
  NA2        g0871(.A(new_new_n769_), .B(new_new_n334_), .Y(new_new_n894_));
  AOI210     g0872(.A0(new_new_n498_), .A1(new_new_n87_), .B0(new_new_n58_), .Y(new_new_n895_));
  OAI220     g0873(.A0(new_new_n895_), .A1(new_new_n894_), .B0(new_new_n685_), .B1(new_new_n554_), .Y(new_new_n896_));
  NO2        g0874(.A(new_new_n259_), .B(new_new_n156_), .Y(new_new_n897_));
  NA2        g0875(.A(i_0_), .B(i_10_), .Y(new_new_n898_));
  INV        g0876(.A(new_new_n557_), .Y(new_new_n899_));
  NO4        g0877(.A(new_new_n116_), .B(new_new_n58_), .C(new_new_n692_), .D(i_5_), .Y(new_new_n900_));
  AO220      g0878(.A0(new_new_n900_), .A1(new_new_n899_), .B0(new_new_n897_), .B1(i_6_), .Y(new_new_n901_));
  AOI220     g0879(.A0(i_0_), .A1(new_new_n99_), .B0(new_new_n190_), .B1(new_new_n82_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n588_), .B(i_4_), .Y(new_new_n903_));
  NA2        g0881(.A(new_new_n193_), .B(new_new_n208_), .Y(new_new_n904_));
  OAI220     g0882(.A0(new_new_n904_), .A1(new_new_n894_), .B0(new_new_n903_), .B1(new_new_n902_), .Y(new_new_n905_));
  NO4        g0883(.A(new_new_n905_), .B(new_new_n901_), .C(new_new_n896_), .D(new_new_n893_), .Y(new_new_n906_));
  NA4        g0884(.A(new_new_n906_), .B(new_new_n892_), .C(new_new_n888_), .D(new_new_n886_), .Y(new_new_n907_));
  NA2        g0885(.A(i_11_), .B(i_9_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n48_), .B(i_7_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n908_), .B(new_new_n71_), .Y(new_new_n910_));
  NO2        g0888(.A(new_new_n179_), .B(i_0_), .Y(new_new_n911_));
  INV        g0889(.A(new_new_n911_), .Y(new_new_n912_));
  NA2        g0890(.A(new_new_n489_), .B(new_new_n238_), .Y(new_new_n913_));
  INV        g0891(.A(new_new_n412_), .Y(new_new_n914_));
  OAI220     g0892(.A0(new_new_n914_), .A1(new_new_n873_), .B0(new_new_n913_), .B1(new_new_n912_), .Y(new_new_n915_));
  INV        g0893(.A(new_new_n915_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n684_), .B(new_new_n123_), .Y(new_new_n917_));
  NO2        g0895(.A(i_6_), .B(new_new_n917_), .Y(new_new_n918_));
  AOI210     g0896(.A0(new_new_n457_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n919_));
  NA2        g0897(.A(new_new_n175_), .B(new_new_n104_), .Y(new_new_n920_));
  NOi32      g0898(.An(new_new_n919_), .Bn(new_new_n193_), .C(new_new_n920_), .Y(new_new_n921_));
  AOI210     g0899(.A0(new_new_n630_), .A1(new_new_n334_), .B0(new_new_n251_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n922_), .B(new_new_n865_), .Y(new_new_n923_));
  NO3        g0901(.A(new_new_n923_), .B(new_new_n921_), .C(new_new_n918_), .Y(new_new_n924_));
  NOi21      g0902(.An(i_7_), .B(i_5_), .Y(new_new_n925_));
  NOi31      g0903(.An(new_new_n925_), .B(i_0_), .C(new_new_n748_), .Y(new_new_n926_));
  NA3        g0904(.A(new_new_n926_), .B(new_new_n390_), .C(i_6_), .Y(new_new_n927_));
  OA210      g0905(.A0(new_new_n920_), .A1(new_new_n533_), .B0(new_new_n927_), .Y(new_new_n928_));
  NO3        g0906(.A(new_new_n408_), .B(new_new_n366_), .C(new_new_n362_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n269_), .B(new_new_n324_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n748_), .B(new_new_n264_), .Y(new_new_n931_));
  AOI210     g0909(.A0(new_new_n931_), .A1(new_new_n930_), .B0(new_new_n929_), .Y(new_new_n932_));
  NA4        g0910(.A(new_new_n932_), .B(new_new_n928_), .C(new_new_n924_), .D(new_new_n916_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n880_), .B(new_new_n247_), .Y(new_new_n934_));
  AN2        g0912(.A(new_new_n339_), .B(new_new_n334_), .Y(new_new_n935_));
  AN2        g0913(.A(new_new_n935_), .B(new_new_n876_), .Y(new_new_n936_));
  OAI210     g0914(.A0(new_new_n936_), .A1(new_new_n934_), .B0(i_10_), .Y(new_new_n937_));
  OA210      g0915(.A0(new_new_n489_), .A1(new_new_n230_), .B0(new_new_n488_), .Y(new_new_n938_));
  NA2        g0916(.A(i_10_), .B(new_new_n910_), .Y(new_new_n939_));
  NA3        g0917(.A(new_new_n488_), .B(new_new_n415_), .C(new_new_n45_), .Y(new_new_n940_));
  OAI210     g0918(.A0(new_new_n884_), .A1(i_7_), .B0(new_new_n940_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n262_), .B(new_new_n46_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n942_), .B(new_new_n192_), .Y(new_new_n943_));
  AOI220     g0921(.A0(new_new_n943_), .A1(new_new_n489_), .B0(new_new_n941_), .B1(new_new_n71_), .Y(new_new_n944_));
  NA3        g0922(.A(new_new_n832_), .B(new_new_n388_), .C(i_6_), .Y(new_new_n945_));
  NA2        g0923(.A(new_new_n93_), .B(new_new_n44_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n73_), .B(new_new_n771_), .Y(new_new_n947_));
  AOI220     g0925(.A0(new_new_n947_), .A1(new_new_n946_), .B0(new_new_n178_), .B1(new_new_n619_), .Y(new_new_n948_));
  AOI210     g0926(.A0(new_new_n948_), .A1(new_new_n945_), .B0(new_new_n47_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n610_), .B(new_new_n361_), .C(new_new_n24_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n725_), .A1(new_new_n566_), .B0(new_new_n950_), .Y(new_new_n951_));
  NAi21      g0929(.An(i_9_), .B(i_5_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n952_), .B(new_new_n408_), .Y(new_new_n953_));
  NO2        g0931(.A(new_new_n624_), .B(new_new_n106_), .Y(new_new_n954_));
  AOI220     g0932(.A0(new_new_n954_), .A1(i_0_), .B0(new_new_n953_), .B1(new_new_n647_), .Y(new_new_n955_));
  OAI220     g0933(.A0(new_new_n955_), .A1(new_new_n84_), .B0(new_new_n951_), .B1(new_new_n176_), .Y(new_new_n956_));
  NO3        g0934(.A(new_new_n956_), .B(new_new_n949_), .C(new_new_n537_), .Y(new_new_n957_));
  NA4        g0935(.A(new_new_n957_), .B(new_new_n944_), .C(new_new_n939_), .D(new_new_n937_), .Y(new_new_n958_));
  NO3        g0936(.A(new_new_n958_), .B(new_new_n933_), .C(new_new_n907_), .Y(new_new_n959_));
  NO2        g0937(.A(i_0_), .B(new_new_n748_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n71_), .B(new_new_n44_), .Y(new_new_n961_));
  NA2        g0939(.A(new_new_n898_), .B(new_new_n961_), .Y(new_new_n962_));
  NO3        g0940(.A(new_new_n106_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n963_));
  AO220      g0941(.A0(new_new_n963_), .A1(new_new_n962_), .B0(new_new_n960_), .B1(new_new_n178_), .Y(new_new_n964_));
  AOI210     g0942(.A0(new_new_n814_), .A1(new_new_n712_), .B0(new_new_n920_), .Y(new_new_n965_));
  AOI210     g0943(.A0(new_new_n964_), .A1(new_new_n350_), .B0(new_new_n965_), .Y(new_new_n966_));
  NA2        g0944(.A(new_new_n759_), .B(new_new_n148_), .Y(new_new_n967_));
  INV        g0945(.A(new_new_n967_), .Y(new_new_n968_));
  NA3        g0946(.A(new_new_n968_), .B(new_new_n699_), .C(new_new_n71_), .Y(new_new_n969_));
  NO2        g0947(.A(new_new_n828_), .B(new_new_n408_), .Y(new_new_n970_));
  NA3        g0948(.A(new_new_n855_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n856_), .B(i_9_), .Y(new_new_n972_));
  AOI210     g0950(.A0(new_new_n971_), .A1(new_new_n513_), .B0(new_new_n972_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n252_), .B(new_new_n237_), .Y(new_new_n974_));
  AOI210     g0952(.A0(new_new_n974_), .A1(new_new_n889_), .B0(new_new_n156_), .Y(new_new_n975_));
  NO3        g0953(.A(new_new_n975_), .B(new_new_n973_), .C(new_new_n970_), .Y(new_new_n976_));
  NA3        g0954(.A(new_new_n976_), .B(new_new_n969_), .C(new_new_n966_), .Y(new_new_n977_));
  NA2        g0955(.A(new_new_n935_), .B(new_new_n378_), .Y(new_new_n978_));
  AOI210     g0956(.A0(new_new_n308_), .A1(new_new_n165_), .B0(new_new_n978_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n39_), .B(new_new_n44_), .Y(new_new_n980_));
  NA2        g0958(.A(new_new_n909_), .B(new_new_n501_), .Y(new_new_n981_));
  AOI210     g0959(.A0(new_new_n980_), .A1(new_new_n165_), .B0(new_new_n981_), .Y(new_new_n982_));
  NO2        g0960(.A(new_new_n982_), .B(new_new_n979_), .Y(new_new_n983_));
  NO3        g0961(.A(new_new_n898_), .B(new_new_n872_), .C(new_new_n195_), .Y(new_new_n984_));
  AOI220     g0962(.A0(new_new_n984_), .A1(i_11_), .B0(new_new_n589_), .B1(new_new_n73_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n215_), .B(new_new_n389_), .C(i_0_), .Y(new_new_n986_));
  OAI210     g0964(.A0(new_new_n986_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n987_));
  INV        g0965(.A(new_new_n224_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n1082_), .B(new_new_n641_), .Y(new_new_n989_));
  NA3        g0967(.A(new_new_n989_), .B(new_new_n1080_), .C(new_new_n988_), .Y(new_new_n990_));
  NA4        g0968(.A(new_new_n990_), .B(new_new_n987_), .C(new_new_n985_), .D(new_new_n983_), .Y(new_new_n991_));
  NO2        g0969(.A(new_new_n250_), .B(new_new_n93_), .Y(new_new_n992_));
  AOI210     g0970(.A0(new_new_n992_), .A1(new_new_n960_), .B0(new_new_n110_), .Y(new_new_n993_));
  AOI220     g0971(.A0(new_new_n925_), .A1(new_new_n501_), .B0(new_new_n855_), .B1(new_new_n166_), .Y(new_new_n994_));
  NA2        g0972(.A(new_new_n353_), .B(new_new_n180_), .Y(new_new_n995_));
  OA220      g0973(.A0(new_new_n995_), .A1(new_new_n994_), .B0(new_new_n993_), .B1(i_5_), .Y(new_new_n996_));
  AOI210     g0974(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n997_));
  NA2        g0975(.A(new_new_n997_), .B(new_new_n938_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n638_), .B(new_new_n190_), .C(new_new_n82_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n999_), .B(new_new_n564_), .Y(new_new_n1000_));
  NO3        g0978(.A(new_new_n865_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n1001_));
  NA3        g0979(.A(new_new_n506_), .B(new_new_n499_), .C(new_new_n486_), .Y(new_new_n1002_));
  NO3        g0980(.A(new_new_n1002_), .B(new_new_n1001_), .C(new_new_n1000_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n396_), .B(new_new_n175_), .C(new_new_n174_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n909_), .B(new_new_n297_), .C(new_new_n237_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n1005_), .B(new_new_n1004_), .Y(new_new_n1006_));
  NA3        g0984(.A(new_new_n396_), .B(new_new_n340_), .C(new_new_n228_), .Y(new_new_n1007_));
  INV        g0985(.A(new_new_n1007_), .Y(new_new_n1008_));
  NOi31      g0986(.An(new_new_n395_), .B(new_new_n961_), .C(new_new_n247_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n908_), .B(new_new_n224_), .C(new_new_n195_), .Y(new_new_n1010_));
  NO4        g0988(.A(new_new_n1010_), .B(new_new_n1009_), .C(new_new_n1008_), .D(new_new_n1006_), .Y(new_new_n1011_));
  NA4        g0989(.A(new_new_n1011_), .B(new_new_n1003_), .C(new_new_n998_), .D(new_new_n996_), .Y(new_new_n1012_));
  INV        g0990(.A(new_new_n640_), .Y(new_new_n1013_));
  NO3        g0991(.A(new_new_n1013_), .B(new_new_n579_), .C(i_3_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n1014_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n312_), .B(i_5_), .C(new_new_n198_), .Y(new_new_n1016_));
  NAi31      g0994(.An(new_new_n249_), .B(new_new_n1016_), .C(new_new_n250_), .Y(new_new_n1017_));
  NO4        g0995(.A(new_new_n247_), .B(new_new_n215_), .C(i_0_), .D(i_12_), .Y(new_new_n1018_));
  AOI220     g0996(.A0(new_new_n1018_), .A1(new_new_n1017_), .B0(new_new_n808_), .B1(new_new_n180_), .Y(new_new_n1019_));
  AN2        g0997(.A(new_new_n898_), .B(new_new_n156_), .Y(new_new_n1020_));
  NO4        g0998(.A(new_new_n1020_), .B(i_12_), .C(new_new_n675_), .D(new_new_n133_), .Y(new_new_n1021_));
  NA2        g0999(.A(new_new_n1021_), .B(new_new_n224_), .Y(new_new_n1022_));
  NA3        g1000(.A(new_new_n99_), .B(new_new_n593_), .C(i_11_), .Y(new_new_n1023_));
  NA2        g1001(.A(new_new_n925_), .B(new_new_n485_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n64_), .B(new_new_n102_), .Y(new_new_n1025_));
  OAI220     g1003(.A0(new_new_n1025_), .A1(new_new_n1016_), .B0(new_new_n1024_), .B1(new_new_n700_), .Y(new_new_n1026_));
  NA2        g1004(.A(new_new_n1026_), .B(new_new_n911_), .Y(new_new_n1027_));
  NA4        g1005(.A(new_new_n1027_), .B(new_new_n1022_), .C(new_new_n1019_), .D(new_new_n1015_), .Y(new_new_n1028_));
  NO4        g1006(.A(new_new_n1028_), .B(new_new_n1012_), .C(new_new_n991_), .D(new_new_n977_), .Y(new_new_n1029_));
  OAI210     g1007(.A0(new_new_n831_), .A1(new_new_n826_), .B0(new_new_n37_), .Y(new_new_n1030_));
  NA3        g1008(.A(new_new_n919_), .B(new_new_n373_), .C(i_5_), .Y(new_new_n1031_));
  NA3        g1009(.A(new_new_n1031_), .B(new_new_n1030_), .C(new_new_n636_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n1032_), .B(new_new_n212_), .Y(new_new_n1033_));
  AN2        g1011(.A(new_new_n721_), .B(new_new_n374_), .Y(new_new_n1034_));
  NA2        g1012(.A(new_new_n191_), .B(new_new_n193_), .Y(new_new_n1035_));
  AO210      g1013(.A0(new_new_n1034_), .A1(new_new_n33_), .B0(new_new_n1035_), .Y(new_new_n1036_));
  NA2        g1014(.A(new_new_n638_), .B(new_new_n323_), .Y(new_new_n1037_));
  NAi31      g1015(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1038_));
  NA3        g1016(.A(new_new_n1038_), .B(new_new_n1037_), .C(new_new_n1036_), .Y(new_new_n1039_));
  NO2        g1017(.A(new_new_n475_), .B(new_new_n275_), .Y(new_new_n1040_));
  NO4        g1018(.A(new_new_n240_), .B(new_new_n147_), .C(new_new_n703_), .D(new_new_n37_), .Y(new_new_n1041_));
  NO3        g1019(.A(new_new_n1041_), .B(new_new_n1040_), .C(new_new_n891_), .Y(new_new_n1042_));
  NA2        g1020(.A(new_new_n1023_), .B(new_new_n1042_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n1039_), .A1(new_new_n48_), .B0(new_new_n1043_), .Y(new_new_n1044_));
  AOI210     g1022(.A0(new_new_n1044_), .A1(new_new_n1033_), .B0(new_new_n71_), .Y(new_new_n1045_));
  NO2        g1023(.A(new_new_n586_), .B(new_new_n385_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n1046_), .B(new_new_n776_), .Y(new_new_n1047_));
  OAI210     g1025(.A0(new_new_n78_), .A1(new_new_n54_), .B0(new_new_n109_), .Y(new_new_n1048_));
  NA2        g1026(.A(new_new_n1048_), .B(new_new_n74_), .Y(new_new_n1049_));
  AOI210     g1027(.A0(new_new_n997_), .A1(new_new_n909_), .B0(new_new_n926_), .Y(new_new_n1050_));
  AOI210     g1028(.A0(new_new_n1050_), .A1(new_new_n1049_), .B0(new_new_n703_), .Y(new_new_n1051_));
  NA2        g1029(.A(new_new_n269_), .B(new_new_n57_), .Y(new_new_n1052_));
  AOI220     g1030(.A0(new_new_n1052_), .A1(new_new_n74_), .B0(new_new_n348_), .B1(new_new_n261_), .Y(new_new_n1053_));
  NO2        g1031(.A(new_new_n1053_), .B(new_new_n244_), .Y(new_new_n1054_));
  NA3        g1032(.A(new_new_n97_), .B(new_new_n314_), .C(new_new_n31_), .Y(new_new_n1055_));
  INV        g1033(.A(new_new_n1055_), .Y(new_new_n1056_));
  NO3        g1034(.A(new_new_n1056_), .B(new_new_n1054_), .C(new_new_n1051_), .Y(new_new_n1057_));
  OAI210     g1035(.A0(new_new_n277_), .A1(new_new_n161_), .B0(new_new_n87_), .Y(new_new_n1058_));
  NA3        g1036(.A(new_new_n780_), .B(new_new_n297_), .C(new_new_n78_), .Y(new_new_n1059_));
  AOI210     g1037(.A0(new_new_n1059_), .A1(new_new_n1058_), .B0(i_11_), .Y(new_new_n1060_));
  NA2        g1038(.A(new_new_n631_), .B(new_new_n221_), .Y(new_new_n1061_));
  OAI210     g1039(.A0(new_new_n1061_), .A1(new_new_n919_), .B0(new_new_n212_), .Y(new_new_n1062_));
  NA2        g1040(.A(new_new_n167_), .B(i_5_), .Y(new_new_n1063_));
  AOI210     g1041(.A0(new_new_n1062_), .A1(new_new_n793_), .B0(new_new_n1063_), .Y(new_new_n1064_));
  NO3        g1042(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1065_));
  OAI210     g1043(.A0(new_new_n930_), .A1(new_new_n314_), .B0(new_new_n1065_), .Y(new_new_n1066_));
  NO2        g1044(.A(new_new_n1066_), .B(new_new_n748_), .Y(new_new_n1067_));
  NO4        g1045(.A(new_new_n952_), .B(i_11_), .C(i_3_), .D(new_new_n258_), .Y(new_new_n1068_));
  NO2        g1046(.A(new_new_n1068_), .B(new_new_n583_), .Y(new_new_n1069_));
  INV        g1047(.A(new_new_n367_), .Y(new_new_n1070_));
  AOI210     g1048(.A0(new_new_n1070_), .A1(new_new_n1069_), .B0(new_new_n40_), .Y(new_new_n1071_));
  NO4        g1049(.A(new_new_n1071_), .B(new_new_n1067_), .C(new_new_n1064_), .D(new_new_n1060_), .Y(new_new_n1072_));
  OAI210     g1050(.A0(new_new_n1057_), .A1(i_4_), .B0(new_new_n1072_), .Y(new_new_n1073_));
  NO3        g1051(.A(new_new_n1073_), .B(new_new_n1047_), .C(new_new_n1045_), .Y(new_new_n1074_));
  NA4        g1052(.A(new_new_n1074_), .B(new_new_n1029_), .C(new_new_n959_), .D(new_new_n879_), .Y(men4));
  INV        g1053(.A(i_2_), .Y(new_new_n1078_));
  INV        g1054(.A(i_5_), .Y(new_new_n1079_));
  INV        g1055(.A(i_3_), .Y(new_new_n1080_));
  INV        g1056(.A(i_6_), .Y(new_new_n1081_));
  INV        g1057(.A(i_6_), .Y(new_new_n1082_));
  INV        g1058(.A(i_9_), .Y(new_new_n1083_));
  INV        g1059(.A(i_5_), .Y(new_new_n1084_));
endmodule


