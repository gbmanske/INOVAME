//Benchmark atmr_misex3_1774_0.125

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1482_, men_men_n1483_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o000(.A(b), .B(a), .Y(ori_ori_n29_));
  NA2        o001(.A(e), .B(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi32      o002(.An(i), .Bn(g), .C(h), .Y(ori_ori_n31_));
  AN2        o003(.A(m), .B(l), .Y(ori_ori_n32_));
  NOi32      o004(.An(j), .Bn(g), .C(k), .Y(ori_ori_n33_));
  NA2        o005(.A(ori_ori_n33_), .B(ori_ori_n32_), .Y(ori_ori_n34_));
  INV        o006(.A(h), .Y(ori_ori_n35_));
  NAi21      o007(.An(j), .B(l), .Y(ori_ori_n36_));
  INV        o008(.A(i), .Y(ori_ori_n37_));
  AN2        o009(.A(h), .B(g), .Y(ori_ori_n38_));
  NA2        o010(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n39_));
  NAi21      o011(.An(n), .B(m), .Y(ori_ori_n40_));
  NOi32      o012(.An(k), .Bn(h), .C(l), .Y(ori_ori_n41_));
  NOi32      o013(.An(k), .Bn(h), .C(g), .Y(ori_ori_n42_));
  INV        o014(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o015(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o016(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o017(.A(ori_ori_n45_), .B(ori_ori_n30_), .Y(ori_ori_n46_));
  INV        o018(.A(c), .Y(ori_ori_n47_));
  NA2        o019(.A(e), .B(b), .Y(ori_ori_n48_));
  INV        o020(.A(ori_ori_n48_), .Y(ori_ori_n49_));
  INV        o021(.A(d), .Y(ori_ori_n50_));
  NAi21      o022(.An(i), .B(h), .Y(ori_ori_n51_));
  NA2        o023(.A(g), .B(f), .Y(ori_ori_n52_));
  NAi31      o024(.An(l), .B(m), .C(k), .Y(ori_ori_n53_));
  NAi21      o025(.An(e), .B(h), .Y(ori_ori_n54_));
  INV        o026(.A(m), .Y(ori_ori_n55_));
  NOi21      o027(.An(k), .B(l), .Y(ori_ori_n56_));
  NA2        o028(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  AN4        o029(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n58_));
  NOi21      o030(.An(h), .B(f), .Y(ori_ori_n59_));
  NA2        o031(.A(ori_ori_n59_), .B(ori_ori_n58_), .Y(ori_ori_n60_));
  NAi32      o032(.An(m), .Bn(k), .C(j), .Y(ori_ori_n61_));
  OR2        o033(.A(ori_ori_n60_), .B(ori_ori_n57_), .Y(ori_ori_n62_));
  INV        o034(.A(ori_ori_n62_), .Y(ori_ori_n63_));
  INV        o035(.A(n), .Y(ori_ori_n64_));
  NOi32      o036(.An(e), .Bn(b), .C(d), .Y(ori_ori_n65_));
  NA2        o037(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  INV        o038(.A(j), .Y(ori_ori_n67_));
  AN3        o039(.A(m), .B(k), .C(i), .Y(ori_ori_n68_));
  NA3        o040(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(g), .Y(ori_ori_n69_));
  NO2        o041(.A(ori_ori_n69_), .B(f), .Y(ori_ori_n70_));
  NAi32      o042(.An(g), .Bn(f), .C(h), .Y(ori_ori_n71_));
  NAi31      o043(.An(j), .B(m), .C(l), .Y(ori_ori_n72_));
  NO2        o044(.A(ori_ori_n72_), .B(ori_ori_n71_), .Y(ori_ori_n73_));
  NA2        o045(.A(m), .B(l), .Y(ori_ori_n74_));
  NOi32      o046(.An(m), .Bn(l), .C(i), .Y(ori_ori_n75_));
  NOi21      o047(.An(g), .B(i), .Y(ori_ori_n76_));
  AOI220     o048(.A0(m), .A1(ori_ori_n76_), .B0(ori_ori_n75_), .B1(g), .Y(ori_ori_n77_));
  NO2        o049(.A(ori_ori_n73_), .B(ori_ori_n70_), .Y(ori_ori_n78_));
  NAi41      o050(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n79_));
  AN2        o051(.A(e), .B(b), .Y(ori_ori_n80_));
  NOi31      o052(.An(c), .B(h), .C(f), .Y(ori_ori_n81_));
  NA2        o053(.A(ori_ori_n81_), .B(ori_ori_n80_), .Y(ori_ori_n82_));
  NO2        o054(.A(ori_ori_n82_), .B(ori_ori_n79_), .Y(ori_ori_n83_));
  NOi21      o055(.An(i), .B(h), .Y(ori_ori_n84_));
  INV        o056(.A(a), .Y(ori_ori_n85_));
  NA2        o057(.A(ori_ori_n80_), .B(ori_ori_n85_), .Y(ori_ori_n86_));
  INV        o058(.A(l), .Y(ori_ori_n87_));
  NOi21      o059(.An(m), .B(n), .Y(ori_ori_n88_));
  AN2        o060(.A(k), .B(h), .Y(ori_ori_n89_));
  INV        o061(.A(b), .Y(ori_ori_n90_));
  NA2        o062(.A(l), .B(j), .Y(ori_ori_n91_));
  INV        o063(.A(ori_ori_n83_), .Y(ori_ori_n92_));
  OAI210     o064(.A0(ori_ori_n78_), .A1(ori_ori_n66_), .B0(ori_ori_n92_), .Y(ori_ori_n93_));
  NOi31      o065(.An(k), .B(m), .C(j), .Y(ori_ori_n94_));
  NA3        o066(.A(ori_ori_n94_), .B(ori_ori_n59_), .C(ori_ori_n58_), .Y(ori_ori_n95_));
  NOi31      o067(.An(k), .B(m), .C(i), .Y(ori_ori_n96_));
  INV        o068(.A(ori_ori_n95_), .Y(ori_ori_n97_));
  NOi32      o069(.An(f), .Bn(b), .C(e), .Y(ori_ori_n98_));
  NAi21      o070(.An(g), .B(h), .Y(ori_ori_n99_));
  NAi21      o071(.An(m), .B(n), .Y(ori_ori_n100_));
  NAi21      o072(.An(j), .B(k), .Y(ori_ori_n101_));
  NO3        o073(.A(ori_ori_n101_), .B(ori_ori_n100_), .C(ori_ori_n99_), .Y(ori_ori_n102_));
  NAi31      o074(.An(j), .B(k), .C(h), .Y(ori_ori_n103_));
  NA2        o075(.A(ori_ori_n102_), .B(ori_ori_n98_), .Y(ori_ori_n104_));
  INV        o076(.A(ori_ori_n100_), .Y(ori_ori_n105_));
  AN2        o077(.A(k), .B(j), .Y(ori_ori_n106_));
  NAi21      o078(.An(c), .B(b), .Y(ori_ori_n107_));
  NA2        o079(.A(f), .B(d), .Y(ori_ori_n108_));
  NO4        o080(.A(ori_ori_n108_), .B(ori_ori_n107_), .C(ori_ori_n106_), .D(ori_ori_n99_), .Y(ori_ori_n109_));
  NAi31      o081(.An(f), .B(e), .C(b), .Y(ori_ori_n110_));
  NA2        o082(.A(ori_ori_n109_), .B(ori_ori_n105_), .Y(ori_ori_n111_));
  NA2        o083(.A(d), .B(b), .Y(ori_ori_n112_));
  NAi21      o084(.An(e), .B(f), .Y(ori_ori_n113_));
  NA2        o085(.A(b), .B(a), .Y(ori_ori_n114_));
  NAi21      o086(.An(e), .B(g), .Y(ori_ori_n115_));
  NAi21      o087(.An(c), .B(d), .Y(ori_ori_n116_));
  NAi31      o088(.An(l), .B(k), .C(h), .Y(ori_ori_n117_));
  NAi31      o089(.An(ori_ori_n97_), .B(ori_ori_n111_), .C(ori_ori_n104_), .Y(ori_ori_n118_));
  NAi31      o090(.An(e), .B(f), .C(b), .Y(ori_ori_n119_));
  NOi21      o091(.An(h), .B(i), .Y(ori_ori_n120_));
  NOi21      o092(.An(k), .B(m), .Y(ori_ori_n121_));
  NA3        o093(.A(ori_ori_n121_), .B(ori_ori_n120_), .C(n), .Y(ori_ori_n122_));
  NOi21      o094(.An(h), .B(g), .Y(ori_ori_n123_));
  NOi32      o095(.An(n), .Bn(k), .C(m), .Y(ori_ori_n124_));
  NAi31      o096(.An(d), .B(f), .C(c), .Y(ori_ori_n125_));
  NAi31      o097(.An(e), .B(f), .C(c), .Y(ori_ori_n126_));
  NA2        o098(.A(ori_ori_n126_), .B(ori_ori_n125_), .Y(ori_ori_n127_));
  NA2        o099(.A(j), .B(h), .Y(ori_ori_n128_));
  OR3        o100(.A(n), .B(m), .C(k), .Y(ori_ori_n129_));
  NO2        o101(.A(ori_ori_n129_), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  NAi32      o102(.An(m), .Bn(k), .C(n), .Y(ori_ori_n131_));
  NA2        o103(.A(ori_ori_n130_), .B(ori_ori_n127_), .Y(ori_ori_n132_));
  NO2        o104(.A(n), .B(m), .Y(ori_ori_n133_));
  NA2        o105(.A(ori_ori_n133_), .B(ori_ori_n41_), .Y(ori_ori_n134_));
  NAi21      o106(.An(f), .B(e), .Y(ori_ori_n135_));
  NA2        o107(.A(d), .B(c), .Y(ori_ori_n136_));
  NO2        o108(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n137_));
  NOi21      o109(.An(ori_ori_n137_), .B(ori_ori_n134_), .Y(ori_ori_n138_));
  NAi31      o110(.An(m), .B(n), .C(b), .Y(ori_ori_n139_));
  NA2        o111(.A(k), .B(i), .Y(ori_ori_n140_));
  NAi21      o112(.An(h), .B(f), .Y(ori_ori_n141_));
  NO2        o113(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n142_));
  NO2        o114(.A(ori_ori_n139_), .B(ori_ori_n116_), .Y(ori_ori_n143_));
  NA2        o115(.A(ori_ori_n143_), .B(ori_ori_n142_), .Y(ori_ori_n144_));
  NOi32      o116(.An(f), .Bn(c), .C(d), .Y(ori_ori_n145_));
  NOi32      o117(.An(f), .Bn(c), .C(e), .Y(ori_ori_n146_));
  NO2        o118(.A(ori_ori_n146_), .B(ori_ori_n145_), .Y(ori_ori_n147_));
  NO3        o119(.A(n), .B(m), .C(j), .Y(ori_ori_n148_));
  NA2        o120(.A(ori_ori_n148_), .B(ori_ori_n89_), .Y(ori_ori_n149_));
  AO210      o121(.A0(ori_ori_n149_), .A1(ori_ori_n134_), .B0(ori_ori_n147_), .Y(ori_ori_n150_));
  NAi41      o122(.An(ori_ori_n138_), .B(ori_ori_n150_), .C(ori_ori_n144_), .D(ori_ori_n132_), .Y(ori_ori_n151_));
  OR2        o123(.A(ori_ori_n151_), .B(ori_ori_n118_), .Y(ori_ori_n152_));
  NO4        o124(.A(ori_ori_n152_), .B(ori_ori_n93_), .C(ori_ori_n63_), .D(ori_ori_n46_), .Y(ori_ori_n153_));
  NA3        o125(.A(m), .B(ori_ori_n87_), .C(j), .Y(ori_ori_n154_));
  NAi31      o126(.An(n), .B(h), .C(g), .Y(ori_ori_n155_));
  NO2        o127(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NOi32      o128(.An(m), .Bn(k), .C(l), .Y(ori_ori_n157_));
  NA3        o129(.A(ori_ori_n157_), .B(ori_ori_n67_), .C(g), .Y(ori_ori_n158_));
  NOi21      o130(.An(k), .B(j), .Y(ori_ori_n159_));
  NA4        o131(.A(ori_ori_n159_), .B(ori_ori_n88_), .C(i), .D(g), .Y(ori_ori_n160_));
  INV        o132(.A(ori_ori_n156_), .Y(ori_ori_n161_));
  NAi41      o133(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n162_));
  INV        o134(.A(ori_ori_n162_), .Y(ori_ori_n163_));
  INV        o135(.A(f), .Y(ori_ori_n164_));
  INV        o136(.A(g), .Y(ori_ori_n165_));
  NOi31      o137(.An(i), .B(j), .C(h), .Y(ori_ori_n166_));
  NOi21      o138(.An(l), .B(m), .Y(ori_ori_n167_));
  NA2        o139(.A(ori_ori_n167_), .B(ori_ori_n166_), .Y(ori_ori_n168_));
  NO3        o140(.A(ori_ori_n168_), .B(ori_ori_n165_), .C(ori_ori_n164_), .Y(ori_ori_n169_));
  NA2        o141(.A(ori_ori_n169_), .B(ori_ori_n163_), .Y(ori_ori_n170_));
  OAI210     o142(.A0(ori_ori_n161_), .A1(ori_ori_n30_), .B0(ori_ori_n170_), .Y(ori_ori_n171_));
  NOi21      o143(.An(n), .B(m), .Y(ori_ori_n172_));
  OR2        o144(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n173_));
  NAi21      o145(.An(j), .B(h), .Y(ori_ori_n174_));
  XN2        o146(.A(i), .B(h), .Y(ori_ori_n175_));
  NA2        o147(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  NOi31      o148(.An(k), .B(n), .C(m), .Y(ori_ori_n177_));
  NOi31      o149(.An(ori_ori_n177_), .B(ori_ori_n136_), .C(ori_ori_n135_), .Y(ori_ori_n178_));
  NA2        o150(.A(ori_ori_n178_), .B(ori_ori_n176_), .Y(ori_ori_n179_));
  NAi31      o151(.An(f), .B(e), .C(c), .Y(ori_ori_n180_));
  NA3        o152(.A(e), .B(c), .C(b), .Y(ori_ori_n181_));
  NAi32      o153(.An(m), .Bn(i), .C(k), .Y(ori_ori_n182_));
  INV        o154(.A(k), .Y(ori_ori_n183_));
  NAi21      o155(.An(n), .B(a), .Y(ori_ori_n184_));
  NO2        o156(.A(ori_ori_n184_), .B(ori_ori_n112_), .Y(ori_ori_n185_));
  NAi41      o157(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n186_));
  AN2        o158(.A(ori_ori_n179_), .B(ori_ori_n173_), .Y(ori_ori_n187_));
  OR2        o159(.A(h), .B(g), .Y(ori_ori_n188_));
  NO2        o160(.A(ori_ori_n188_), .B(ori_ori_n79_), .Y(ori_ori_n189_));
  NA2        o161(.A(ori_ori_n189_), .B(ori_ori_n98_), .Y(ori_ori_n190_));
  NAi41      o162(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n191_));
  NO2        o163(.A(ori_ori_n191_), .B(ori_ori_n164_), .Y(ori_ori_n192_));
  NA2        o164(.A(ori_ori_n121_), .B(ori_ori_n84_), .Y(ori_ori_n193_));
  NO2        o165(.A(n), .B(a), .Y(ori_ori_n194_));
  NAi31      o166(.An(ori_ori_n186_), .B(ori_ori_n194_), .C(ori_ori_n80_), .Y(ori_ori_n195_));
  NAi21      o167(.An(h), .B(i), .Y(ori_ori_n196_));
  NA2        o168(.A(ori_ori_n133_), .B(k), .Y(ori_ori_n197_));
  NO2        o169(.A(ori_ori_n197_), .B(ori_ori_n196_), .Y(ori_ori_n198_));
  NA2        o170(.A(ori_ori_n198_), .B(ori_ori_n145_), .Y(ori_ori_n199_));
  NA3        o171(.A(ori_ori_n199_), .B(ori_ori_n195_), .C(ori_ori_n190_), .Y(ori_ori_n200_));
  NOi21      o172(.An(g), .B(e), .Y(ori_ori_n201_));
  NOi31      o173(.An(ori_ori_n187_), .B(ori_ori_n200_), .C(ori_ori_n171_), .Y(ori_ori_n202_));
  INV        o174(.A(ori_ori_n156_), .Y(ori_ori_n203_));
  NO2        o175(.A(ori_ori_n203_), .B(ori_ori_n86_), .Y(ori_ori_n204_));
  NA3        o176(.A(ori_ori_n50_), .B(c), .C(b), .Y(ori_ori_n205_));
  NO2        o177(.A(ori_ori_n193_), .B(f), .Y(ori_ori_n206_));
  NAi31      o178(.An(g), .B(k), .C(h), .Y(ori_ori_n207_));
  NA3        o179(.A(ori_ori_n121_), .B(ori_ori_n120_), .C(ori_ori_n64_), .Y(ori_ori_n208_));
  NO2        o180(.A(ori_ori_n208_), .B(ori_ori_n147_), .Y(ori_ori_n209_));
  NA3        o181(.A(e), .B(c), .C(b), .Y(ori_ori_n210_));
  NAi32      o182(.An(j), .Bn(h), .C(i), .Y(ori_ori_n211_));
  NAi21      o183(.An(m), .B(l), .Y(ori_ori_n212_));
  NA2        o184(.A(h), .B(g), .Y(ori_ori_n213_));
  INV        o185(.A(ori_ori_n110_), .Y(ori_ori_n214_));
  NO2        o186(.A(ori_ori_n82_), .B(ori_ori_n79_), .Y(ori_ori_n215_));
  NAi32      o187(.An(n), .Bn(m), .C(l), .Y(ori_ori_n216_));
  NO2        o188(.A(ori_ori_n216_), .B(ori_ori_n211_), .Y(ori_ori_n217_));
  NA2        o189(.A(ori_ori_n217_), .B(ori_ori_n137_), .Y(ori_ori_n218_));
  INV        o190(.A(ori_ori_n218_), .Y(ori_ori_n219_));
  NO3        o191(.A(ori_ori_n219_), .B(ori_ori_n209_), .C(ori_ori_n204_), .Y(ori_ori_n220_));
  NA2        o192(.A(ori_ori_n198_), .B(ori_ori_n146_), .Y(ori_ori_n221_));
  NAi21      o193(.An(m), .B(k), .Y(ori_ori_n222_));
  NO2        o194(.A(ori_ori_n175_), .B(ori_ori_n222_), .Y(ori_ori_n223_));
  NAi41      o195(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n224_));
  NO2        o196(.A(ori_ori_n224_), .B(ori_ori_n115_), .Y(ori_ori_n225_));
  NA2        o197(.A(ori_ori_n225_), .B(ori_ori_n223_), .Y(ori_ori_n226_));
  NA2        o198(.A(e), .B(c), .Y(ori_ori_n227_));
  NO3        o199(.A(ori_ori_n227_), .B(n), .C(d), .Y(ori_ori_n228_));
  NOi21      o200(.An(f), .B(h), .Y(ori_ori_n229_));
  NA2        o201(.A(ori_ori_n229_), .B(k), .Y(ori_ori_n230_));
  NO2        o202(.A(ori_ori_n230_), .B(ori_ori_n165_), .Y(ori_ori_n231_));
  NAi31      o203(.An(d), .B(e), .C(b), .Y(ori_ori_n232_));
  NO2        o204(.A(ori_ori_n100_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NA2        o205(.A(ori_ori_n233_), .B(ori_ori_n231_), .Y(ori_ori_n234_));
  NA3        o206(.A(ori_ori_n234_), .B(ori_ori_n226_), .C(ori_ori_n221_), .Y(ori_ori_n235_));
  NO4        o207(.A(ori_ori_n224_), .B(ori_ori_n61_), .C(ori_ori_n54_), .D(ori_ori_n165_), .Y(ori_ori_n236_));
  NA2        o208(.A(ori_ori_n194_), .B(ori_ori_n80_), .Y(ori_ori_n237_));
  OR2        o209(.A(ori_ori_n237_), .B(ori_ori_n158_), .Y(ori_ori_n238_));
  NOi31      o210(.An(l), .B(n), .C(m), .Y(ori_ori_n239_));
  NA2        o211(.A(ori_ori_n239_), .B(ori_ori_n166_), .Y(ori_ori_n240_));
  NO2        o212(.A(ori_ori_n240_), .B(ori_ori_n147_), .Y(ori_ori_n241_));
  NAi32      o213(.An(ori_ori_n241_), .Bn(ori_ori_n236_), .C(ori_ori_n238_), .Y(ori_ori_n242_));
  NAi32      o214(.An(m), .Bn(j), .C(k), .Y(ori_ori_n243_));
  NAi41      o215(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n244_));
  NA2        o216(.A(ori_ori_n162_), .B(ori_ori_n244_), .Y(ori_ori_n245_));
  NOi31      o217(.An(j), .B(m), .C(k), .Y(ori_ori_n246_));
  NO2        o218(.A(ori_ori_n94_), .B(ori_ori_n246_), .Y(ori_ori_n247_));
  AN3        o219(.A(h), .B(g), .C(f), .Y(ori_ori_n248_));
  NAi31      o220(.An(ori_ori_n247_), .B(ori_ori_n248_), .C(ori_ori_n245_), .Y(ori_ori_n249_));
  NOi32      o221(.An(m), .Bn(j), .C(l), .Y(ori_ori_n250_));
  NO2        o222(.A(ori_ori_n212_), .B(ori_ori_n211_), .Y(ori_ori_n251_));
  NO2        o223(.A(ori_ori_n168_), .B(g), .Y(ori_ori_n252_));
  INV        o224(.A(ori_ori_n119_), .Y(ori_ori_n253_));
  AOI220     o225(.A0(ori_ori_n253_), .A1(ori_ori_n252_), .B0(ori_ori_n192_), .B1(ori_ori_n251_), .Y(ori_ori_n254_));
  NA2        o226(.A(ori_ori_n254_), .B(ori_ori_n249_), .Y(ori_ori_n255_));
  NA3        o227(.A(h), .B(g), .C(f), .Y(ori_ori_n256_));
  NO2        o228(.A(ori_ori_n256_), .B(ori_ori_n57_), .Y(ori_ori_n257_));
  NA2        o229(.A(ori_ori_n244_), .B(ori_ori_n162_), .Y(ori_ori_n258_));
  NA2        o230(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  NOi32      o231(.An(j), .Bn(g), .C(i), .Y(ori_ori_n260_));
  NOi32      o232(.An(e), .Bn(b), .C(a), .Y(ori_ori_n261_));
  AN2        o233(.A(l), .B(j), .Y(ori_ori_n262_));
  NO2        o234(.A(ori_ori_n222_), .B(ori_ori_n262_), .Y(ori_ori_n263_));
  NO3        o235(.A(ori_ori_n224_), .B(ori_ori_n54_), .C(ori_ori_n165_), .Y(ori_ori_n264_));
  NA2        o236(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n265_));
  NAi41      o237(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n266_));
  NA2        o238(.A(ori_ori_n42_), .B(ori_ori_n88_), .Y(ori_ori_n267_));
  NA2        o239(.A(ori_ori_n265_), .B(ori_ori_n259_), .Y(ori_ori_n268_));
  NO4        o240(.A(ori_ori_n268_), .B(ori_ori_n255_), .C(ori_ori_n242_), .D(ori_ori_n235_), .Y(ori_ori_n269_));
  NA4        o241(.A(ori_ori_n269_), .B(ori_ori_n220_), .C(ori_ori_n202_), .D(ori_ori_n153_), .Y(ori10));
  NA3        o242(.A(m), .B(k), .C(i), .Y(ori_ori_n271_));
  NOi21      o243(.An(e), .B(f), .Y(ori_ori_n272_));
  NO3        o244(.A(ori_ori_n116_), .B(n), .C(ori_ori_n85_), .Y(ori_ori_n273_));
  NAi31      o245(.An(b), .B(f), .C(c), .Y(ori_ori_n274_));
  INV        o246(.A(ori_ori_n274_), .Y(ori_ori_n275_));
  NOi32      o247(.An(k), .Bn(h), .C(j), .Y(ori_ori_n276_));
  NA2        o248(.A(ori_ori_n276_), .B(ori_ori_n172_), .Y(ori_ori_n277_));
  NA2        o249(.A(ori_ori_n122_), .B(ori_ori_n277_), .Y(ori_ori_n278_));
  NA2        o250(.A(ori_ori_n278_), .B(ori_ori_n275_), .Y(ori_ori_n279_));
  AN2        o251(.A(j), .B(h), .Y(ori_ori_n280_));
  NO3        o252(.A(n), .B(m), .C(k), .Y(ori_ori_n281_));
  NA2        o253(.A(ori_ori_n281_), .B(ori_ori_n280_), .Y(ori_ori_n282_));
  NO3        o254(.A(ori_ori_n282_), .B(ori_ori_n116_), .C(ori_ori_n164_), .Y(ori_ori_n283_));
  OR2        o255(.A(m), .B(k), .Y(ori_ori_n284_));
  NO2        o256(.A(ori_ori_n128_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  NA4        o257(.A(n), .B(f), .C(c), .D(ori_ori_n90_), .Y(ori_ori_n286_));
  NOi21      o258(.An(ori_ori_n285_), .B(ori_ori_n286_), .Y(ori_ori_n287_));
  NOi32      o259(.An(d), .Bn(a), .C(c), .Y(ori_ori_n288_));
  NA2        o260(.A(ori_ori_n288_), .B(ori_ori_n135_), .Y(ori_ori_n289_));
  NO2        o261(.A(ori_ori_n287_), .B(ori_ori_n283_), .Y(ori_ori_n290_));
  NOi32      o262(.An(f), .Bn(d), .C(c), .Y(ori_ori_n291_));
  NA2        o263(.A(ori_ori_n290_), .B(ori_ori_n279_), .Y(ori_ori_n292_));
  NO2        o264(.A(ori_ori_n50_), .B(ori_ori_n90_), .Y(ori_ori_n293_));
  NA2        o265(.A(ori_ori_n194_), .B(ori_ori_n293_), .Y(ori_ori_n294_));
  INV        o266(.A(e), .Y(ori_ori_n295_));
  NA2        o267(.A(ori_ori_n38_), .B(e), .Y(ori_ori_n296_));
  OAI220     o268(.A0(ori_ori_n296_), .A1(ori_ori_n154_), .B0(ori_ori_n158_), .B1(ori_ori_n295_), .Y(ori_ori_n297_));
  NO2        o269(.A(ori_ori_n69_), .B(ori_ori_n295_), .Y(ori_ori_n298_));
  NO2        o270(.A(ori_ori_n77_), .B(ori_ori_n295_), .Y(ori_ori_n299_));
  NO3        o271(.A(ori_ori_n299_), .B(ori_ori_n298_), .C(ori_ori_n297_), .Y(ori_ori_n300_));
  NOi21      o272(.An(g), .B(h), .Y(ori_ori_n301_));
  NA3        o273(.A(m), .B(ori_ori_n301_), .C(e), .Y(ori_ori_n302_));
  AN3        o274(.A(h), .B(g), .C(e), .Y(ori_ori_n303_));
  NA2        o275(.A(ori_ori_n303_), .B(ori_ori_n75_), .Y(ori_ori_n304_));
  AN2        o276(.A(ori_ori_n304_), .B(ori_ori_n302_), .Y(ori_ori_n305_));
  AOI210     o277(.A0(ori_ori_n305_), .A1(ori_ori_n300_), .B0(ori_ori_n294_), .Y(ori_ori_n306_));
  NAi31      o278(.An(b), .B(c), .C(a), .Y(ori_ori_n307_));
  NO2        o279(.A(ori_ori_n307_), .B(n), .Y(ori_ori_n308_));
  NA2        o280(.A(ori_ori_n42_), .B(m), .Y(ori_ori_n309_));
  NO2        o281(.A(ori_ori_n309_), .B(ori_ori_n113_), .Y(ori_ori_n310_));
  NA2        o282(.A(ori_ori_n310_), .B(ori_ori_n308_), .Y(ori_ori_n311_));
  INV        o283(.A(ori_ori_n311_), .Y(ori_ori_n312_));
  NO3        o284(.A(ori_ori_n312_), .B(ori_ori_n306_), .C(ori_ori_n292_), .Y(ori_ori_n313_));
  NA2        o285(.A(i), .B(g), .Y(ori_ori_n314_));
  NOi21      o286(.An(d), .B(c), .Y(ori_ori_n315_));
  NA3        o287(.A(i), .B(g), .C(f), .Y(ori_ori_n316_));
  OR2        o288(.A(ori_ori_n316_), .B(ori_ori_n53_), .Y(ori_ori_n317_));
  OR2        o289(.A(n), .B(m), .Y(ori_ori_n318_));
  NO2        o290(.A(ori_ori_n318_), .B(ori_ori_n117_), .Y(ori_ori_n319_));
  NO2        o291(.A(ori_ori_n136_), .B(ori_ori_n113_), .Y(ori_ori_n320_));
  OAI210     o292(.A0(ori_ori_n319_), .A1(ori_ori_n130_), .B0(ori_ori_n320_), .Y(ori_ori_n321_));
  INV        o293(.A(ori_ori_n267_), .Y(ori_ori_n322_));
  NA3        o294(.A(ori_ori_n322_), .B(ori_ori_n261_), .C(d), .Y(ori_ori_n323_));
  NO2        o295(.A(ori_ori_n307_), .B(ori_ori_n40_), .Y(ori_ori_n324_));
  NO2        o296(.A(ori_ori_n52_), .B(ori_ori_n87_), .Y(ori_ori_n325_));
  NAi21      o297(.An(k), .B(j), .Y(ori_ori_n326_));
  NA2        o298(.A(ori_ori_n196_), .B(ori_ori_n326_), .Y(ori_ori_n327_));
  NA3        o299(.A(ori_ori_n327_), .B(ori_ori_n325_), .C(ori_ori_n324_), .Y(ori_ori_n328_));
  NAi21      o300(.An(e), .B(d), .Y(ori_ori_n329_));
  INV        o301(.A(ori_ori_n329_), .Y(ori_ori_n330_));
  NO2        o302(.A(ori_ori_n197_), .B(ori_ori_n164_), .Y(ori_ori_n331_));
  NA3        o303(.A(ori_ori_n331_), .B(ori_ori_n330_), .C(ori_ori_n176_), .Y(ori_ori_n332_));
  NA4        o304(.A(ori_ori_n332_), .B(ori_ori_n328_), .C(ori_ori_n323_), .D(ori_ori_n321_), .Y(ori_ori_n333_));
  NO2        o305(.A(ori_ori_n240_), .B(ori_ori_n164_), .Y(ori_ori_n334_));
  NA2        o306(.A(ori_ori_n334_), .B(ori_ori_n330_), .Y(ori_ori_n335_));
  NOi31      o307(.An(n), .B(m), .C(k), .Y(ori_ori_n336_));
  AOI220     o308(.A0(ori_ori_n336_), .A1(ori_ori_n280_), .B0(ori_ori_n172_), .B1(ori_ori_n41_), .Y(ori_ori_n337_));
  NAi31      o309(.An(g), .B(f), .C(c), .Y(ori_ori_n338_));
  OR3        o310(.A(ori_ori_n338_), .B(ori_ori_n337_), .C(e), .Y(ori_ori_n339_));
  NA3        o311(.A(ori_ori_n339_), .B(ori_ori_n335_), .C(ori_ori_n218_), .Y(ori_ori_n340_));
  NO2        o312(.A(ori_ori_n340_), .B(ori_ori_n333_), .Y(ori_ori_n341_));
  NOi32      o313(.An(c), .Bn(a), .C(b), .Y(ori_ori_n342_));
  NA2        o314(.A(ori_ori_n342_), .B(ori_ori_n88_), .Y(ori_ori_n343_));
  INV        o315(.A(ori_ori_n207_), .Y(ori_ori_n344_));
  NO2        o316(.A(ori_ori_n99_), .B(ori_ori_n36_), .Y(ori_ori_n345_));
  NO2        o317(.A(ori_ori_n52_), .B(e), .Y(ori_ori_n346_));
  AOI220     o318(.A0(ori_ori_n56_), .A1(ori_ori_n346_), .B0(ori_ori_n345_), .B1(f), .Y(ori_ori_n347_));
  NO2        o319(.A(ori_ori_n347_), .B(ori_ori_n343_), .Y(ori_ori_n348_));
  NOi21      o320(.An(a), .B(b), .Y(ori_ori_n349_));
  INV        o321(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NO2        o322(.A(ori_ori_n203_), .B(ori_ori_n350_), .Y(ori_ori_n351_));
  NA2        o323(.A(l), .B(k), .Y(ori_ori_n352_));
  INV        o324(.A(ori_ori_n95_), .Y(ori_ori_n353_));
  NO3        o325(.A(ori_ori_n353_), .B(ori_ori_n351_), .C(ori_ori_n348_), .Y(ori_ori_n354_));
  NO2        o326(.A(ori_ori_n141_), .B(ori_ori_n47_), .Y(ori_ori_n355_));
  NAi31      o327(.An(j), .B(l), .C(i), .Y(ori_ori_n356_));
  OAI210     o328(.A0(ori_ori_n356_), .A1(ori_ori_n100_), .B0(ori_ori_n79_), .Y(ori_ori_n357_));
  NA2        o329(.A(ori_ori_n357_), .B(ori_ori_n355_), .Y(ori_ori_n358_));
  NO2        o330(.A(ori_ori_n289_), .B(ori_ori_n267_), .Y(ori_ori_n359_));
  NO3        o331(.A(ori_ori_n359_), .B(ori_ori_n138_), .C(ori_ori_n215_), .Y(ori_ori_n360_));
  NA3        o332(.A(ori_ori_n360_), .B(ori_ori_n358_), .C(ori_ori_n187_), .Y(ori_ori_n361_));
  OAI210     o333(.A0(ori_ori_n96_), .A1(ori_ori_n94_), .B0(n), .Y(ori_ori_n362_));
  XO2        o334(.A(i), .B(h), .Y(ori_ori_n363_));
  NA3        o335(.A(ori_ori_n363_), .B(ori_ori_n121_), .C(n), .Y(ori_ori_n364_));
  NA3        o336(.A(ori_ori_n364_), .B(ori_ori_n337_), .C(ori_ori_n277_), .Y(ori_ori_n365_));
  NOi32      o337(.An(ori_ori_n365_), .Bn(ori_ori_n346_), .C(ori_ori_n205_), .Y(ori_ori_n366_));
  NAi31      o338(.An(c), .B(f), .C(d), .Y(ori_ori_n367_));
  NO2        o339(.A(ori_ori_n149_), .B(ori_ori_n367_), .Y(ori_ori_n368_));
  BUFFER     o340(.A(ori_ori_n62_), .Y(ori_ori_n369_));
  NA2        o341(.A(ori_ori_n177_), .B(ori_ori_n84_), .Y(ori_ori_n370_));
  AOI210     o342(.A0(ori_ori_n370_), .A1(ori_ori_n134_), .B0(ori_ori_n367_), .Y(ori_ori_n371_));
  INV        o343(.A(ori_ori_n371_), .Y(ori_ori_n372_));
  NA3        o344(.A(ori_ori_n33_), .B(ori_ori_n32_), .C(f), .Y(ori_ori_n373_));
  NA2        o345(.A(ori_ori_n372_), .B(ori_ori_n369_), .Y(ori_ori_n374_));
  NO3        o346(.A(ori_ori_n374_), .B(ori_ori_n366_), .C(ori_ori_n361_), .Y(ori_ori_n375_));
  NA4        o347(.A(ori_ori_n375_), .B(ori_ori_n354_), .C(ori_ori_n341_), .D(ori_ori_n313_), .Y(ori11));
  NA2        o348(.A(j), .B(g), .Y(ori_ori_n377_));
  NAi31      o349(.An(i), .B(m), .C(l), .Y(ori_ori_n378_));
  NA3        o350(.A(m), .B(k), .C(j), .Y(ori_ori_n379_));
  NOi32      o351(.An(e), .Bn(b), .C(f), .Y(ori_ori_n380_));
  NA2        o352(.A(ori_ori_n38_), .B(j), .Y(ori_ori_n381_));
  NAi31      o353(.An(d), .B(e), .C(a), .Y(ori_ori_n382_));
  NO2        o354(.A(ori_ori_n382_), .B(n), .Y(ori_ori_n383_));
  NA2        o355(.A(j), .B(i), .Y(ori_ori_n384_));
  NAi31      o356(.An(n), .B(m), .C(k), .Y(ori_ori_n385_));
  NO3        o357(.A(ori_ori_n385_), .B(ori_ori_n384_), .C(ori_ori_n87_), .Y(ori_ori_n386_));
  NO4        o358(.A(n), .B(d), .C(ori_ori_n90_), .D(a), .Y(ori_ori_n387_));
  OR2        o359(.A(n), .B(c), .Y(ori_ori_n388_));
  NO2        o360(.A(ori_ori_n388_), .B(ori_ori_n114_), .Y(ori_ori_n389_));
  NO2        o361(.A(ori_ori_n207_), .B(ori_ori_n40_), .Y(ori_ori_n390_));
  NA2        o362(.A(ori_ori_n106_), .B(ori_ori_n31_), .Y(ori_ori_n391_));
  OAI220     o363(.A0(ori_ori_n391_), .A1(m), .B0(ori_ori_n381_), .B1(ori_ori_n182_), .Y(ori_ori_n392_));
  NOi41      o364(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n393_));
  NAi32      o365(.An(e), .Bn(b), .C(c), .Y(ori_ori_n394_));
  OR2        o366(.A(ori_ori_n394_), .B(ori_ori_n64_), .Y(ori_ori_n395_));
  AN2        o367(.A(ori_ori_n244_), .B(ori_ori_n224_), .Y(ori_ori_n396_));
  NA2        o368(.A(ori_ori_n396_), .B(ori_ori_n395_), .Y(ori_ori_n397_));
  OA210      o369(.A0(ori_ori_n397_), .A1(ori_ori_n393_), .B0(ori_ori_n392_), .Y(ori_ori_n398_));
  NAi31      o370(.An(d), .B(c), .C(a), .Y(ori_ori_n399_));
  NO2        o371(.A(ori_ori_n399_), .B(n), .Y(ori_ori_n400_));
  NAi32      o372(.An(d), .Bn(a), .C(b), .Y(ori_ori_n401_));
  NO3        o373(.A(ori_ori_n131_), .B(ori_ori_n128_), .C(g), .Y(ori_ori_n402_));
  NA2        o374(.A(ori_ori_n402_), .B(ori_ori_n49_), .Y(ori_ori_n403_));
  INV        o375(.A(ori_ori_n403_), .Y(ori_ori_n404_));
  AN3        o376(.A(j), .B(h), .C(g), .Y(ori_ori_n405_));
  NO2        o377(.A(ori_ori_n112_), .B(c), .Y(ori_ori_n406_));
  NA3        o378(.A(ori_ori_n406_), .B(ori_ori_n405_), .C(ori_ori_n336_), .Y(ori_ori_n407_));
  NA3        o379(.A(f), .B(d), .C(b), .Y(ori_ori_n408_));
  NO4        o380(.A(ori_ori_n408_), .B(ori_ori_n131_), .C(ori_ori_n128_), .D(g), .Y(ori_ori_n409_));
  INV        o381(.A(ori_ori_n407_), .Y(ori_ori_n410_));
  NO3        o382(.A(ori_ori_n410_), .B(ori_ori_n404_), .C(ori_ori_n398_), .Y(ori_ori_n411_));
  INV        o383(.A(k), .Y(ori_ori_n412_));
  NAi41      o384(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n413_));
  OAI210     o385(.A0(ori_ori_n382_), .A1(n), .B0(ori_ori_n413_), .Y(ori_ori_n414_));
  NAi31      o386(.An(h), .B(g), .C(f), .Y(ori_ori_n415_));
  NAi31      o387(.An(f), .B(h), .C(g), .Y(ori_ori_n416_));
  NOi32      o388(.An(d), .Bn(a), .C(e), .Y(ori_ori_n417_));
  NO2        o389(.A(n), .B(c), .Y(ori_ori_n418_));
  NOi32      o390(.An(e), .Bn(a), .C(d), .Y(ori_ori_n419_));
  AOI210     o391(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n419_), .Y(ori_ori_n420_));
  NA3        o392(.A(ori_ori_n367_), .B(ori_ori_n126_), .C(ori_ori_n125_), .Y(ori_ori_n421_));
  NA2        o393(.A(ori_ori_n338_), .B(ori_ori_n180_), .Y(ori_ori_n422_));
  NA3        o394(.A(ori_ori_n393_), .B(ori_ori_n246_), .C(ori_ori_n38_), .Y(ori_ori_n423_));
  NOi32      o395(.An(e), .Bn(c), .C(f), .Y(ori_ori_n424_));
  INV        o396(.A(ori_ori_n162_), .Y(ori_ori_n425_));
  AOI220     o397(.A0(ori_ori_n425_), .A1(ori_ori_n285_), .B0(ori_ori_n424_), .B1(ori_ori_n130_), .Y(ori_ori_n426_));
  NA3        o398(.A(ori_ori_n426_), .B(ori_ori_n423_), .C(ori_ori_n132_), .Y(ori_ori_n427_));
  NOi31      o399(.An(m), .B(n), .C(k), .Y(ori_ori_n428_));
  NA2        o400(.A(j), .B(ori_ori_n428_), .Y(ori_ori_n429_));
  AOI210     o401(.A0(ori_ori_n289_), .A1(ori_ori_n266_), .B0(ori_ori_n213_), .Y(ori_ori_n430_));
  NAi21      o402(.An(ori_ori_n429_), .B(ori_ori_n430_), .Y(ori_ori_n431_));
  INV        o403(.A(ori_ori_n431_), .Y(ori_ori_n432_));
  NA2        o404(.A(ori_ori_n84_), .B(ori_ori_n32_), .Y(ori_ori_n433_));
  INV        o405(.A(ori_ori_n261_), .Y(ori_ori_n434_));
  NO2        o406(.A(ori_ori_n434_), .B(n), .Y(ori_ori_n435_));
  NAi31      o407(.An(ori_ori_n433_), .B(ori_ori_n435_), .C(g), .Y(ori_ori_n436_));
  NO2        o408(.A(ori_ori_n381_), .B(ori_ori_n131_), .Y(ori_ori_n437_));
  NA3        o409(.A(ori_ori_n394_), .B(ori_ori_n205_), .C(ori_ori_n110_), .Y(ori_ori_n438_));
  NA2        o410(.A(ori_ori_n363_), .B(ori_ori_n121_), .Y(ori_ori_n439_));
  NO3        o411(.A(ori_ori_n286_), .B(ori_ori_n439_), .C(ori_ori_n67_), .Y(ori_ori_n440_));
  AOI210     o412(.A0(ori_ori_n438_), .A1(ori_ori_n437_), .B0(ori_ori_n440_), .Y(ori_ori_n441_));
  AN3        o413(.A(f), .B(d), .C(b), .Y(ori_ori_n442_));
  NAi31      o414(.An(m), .B(n), .C(k), .Y(ori_ori_n443_));
  INV        o415(.A(ori_ori_n195_), .Y(ori_ori_n444_));
  NA2        o416(.A(ori_ori_n444_), .B(j), .Y(ori_ori_n445_));
  NA3        o417(.A(ori_ori_n445_), .B(ori_ori_n441_), .C(ori_ori_n436_), .Y(ori_ori_n446_));
  NO3        o418(.A(ori_ori_n446_), .B(ori_ori_n432_), .C(ori_ori_n427_), .Y(ori_ori_n447_));
  NA2        o419(.A(ori_ori_n273_), .B(ori_ori_n123_), .Y(ori_ori_n448_));
  NAi31      o420(.An(g), .B(h), .C(f), .Y(ori_ori_n449_));
  OA210      o421(.A0(ori_ori_n382_), .A1(n), .B0(ori_ori_n413_), .Y(ori_ori_n450_));
  NO2        o422(.A(ori_ori_n448_), .B(ori_ori_n379_), .Y(ori_ori_n451_));
  NO3        o423(.A(g), .B(ori_ori_n164_), .C(ori_ori_n47_), .Y(ori_ori_n452_));
  NO2        o424(.A(ori_ori_n370_), .B(ori_ori_n67_), .Y(ori_ori_n453_));
  OAI210     o425(.A0(ori_ori_n453_), .A1(ori_ori_n285_), .B0(ori_ori_n452_), .Y(ori_ori_n454_));
  NA2        o426(.A(h), .B(ori_ori_n33_), .Y(ori_ori_n455_));
  NO2        o427(.A(ori_ori_n455_), .B(ori_ori_n343_), .Y(ori_ori_n456_));
  AOI210     o428(.A0(ori_ori_n401_), .A1(ori_ori_n307_), .B0(ori_ori_n40_), .Y(ori_ori_n457_));
  AOI210     o429(.A0(ori_ori_n924_), .A1(ori_ori_n457_), .B0(ori_ori_n456_), .Y(ori_ori_n458_));
  NA2        o430(.A(ori_ori_n458_), .B(ori_ori_n454_), .Y(ori_ori_n459_));
  NA2        o431(.A(ori_ori_n233_), .B(ori_ori_n106_), .Y(ori_ori_n460_));
  INV        o432(.A(ori_ori_n100_), .Y(ori_ori_n461_));
  NA2        o433(.A(ori_ori_n461_), .B(ori_ori_n380_), .Y(ori_ori_n462_));
  OR2        o434(.A(ori_ori_n462_), .B(ori_ori_n391_), .Y(ori_ori_n463_));
  OAI210     o435(.A0(ori_ori_n460_), .A1(ori_ori_n51_), .B0(ori_ori_n463_), .Y(ori_ori_n464_));
  NO2        o436(.A(ori_ori_n291_), .B(ori_ori_n146_), .Y(ori_ori_n465_));
  NA2        o437(.A(ori_ori_n465_), .B(ori_ori_n180_), .Y(ori_ori_n466_));
  NA3        o438(.A(ori_ori_n466_), .B(ori_ori_n198_), .C(j), .Y(ori_ori_n467_));
  NO3        o439(.A(ori_ori_n338_), .B(ori_ori_n128_), .C(i), .Y(ori_ori_n468_));
  NA2        o440(.A(ori_ori_n342_), .B(ori_ori_n64_), .Y(ori_ori_n469_));
  NO4        o441(.A(ori_ori_n379_), .B(ori_ori_n469_), .C(ori_ori_n99_), .D(ori_ori_n164_), .Y(ori_ori_n470_));
  INV        o442(.A(ori_ori_n470_), .Y(ori_ori_n471_));
  NA3        o443(.A(ori_ori_n471_), .B(ori_ori_n467_), .C(ori_ori_n290_), .Y(ori_ori_n472_));
  NO4        o444(.A(ori_ori_n472_), .B(ori_ori_n464_), .C(ori_ori_n459_), .D(ori_ori_n451_), .Y(ori_ori_n473_));
  NA3        o445(.A(ori_ori_n473_), .B(ori_ori_n447_), .C(ori_ori_n411_), .Y(ori08));
  NO2        o446(.A(k), .B(h), .Y(ori_ori_n475_));
  AO210      o447(.A0(ori_ori_n196_), .A1(ori_ori_n326_), .B0(ori_ori_n475_), .Y(ori_ori_n476_));
  NO2        o448(.A(ori_ori_n476_), .B(ori_ori_n212_), .Y(ori_ori_n477_));
  NA2        o449(.A(ori_ori_n424_), .B(ori_ori_n64_), .Y(ori_ori_n478_));
  NA2        o450(.A(ori_ori_n478_), .B(ori_ori_n338_), .Y(ori_ori_n479_));
  NA2        o451(.A(ori_ori_n479_), .B(ori_ori_n477_), .Y(ori_ori_n480_));
  NA2        o452(.A(ori_ori_n64_), .B(ori_ori_n85_), .Y(ori_ori_n481_));
  NO2        o453(.A(ori_ori_n481_), .B(ori_ori_n48_), .Y(ori_ori_n482_));
  NO3        o454(.A(ori_ori_n271_), .B(j), .C(ori_ori_n165_), .Y(ori_ori_n483_));
  NA2        o455(.A(ori_ori_n408_), .B(ori_ori_n181_), .Y(ori_ori_n484_));
  NA2        o456(.A(ori_ori_n483_), .B(ori_ori_n482_), .Y(ori_ori_n485_));
  AOI210     o457(.A0(ori_ori_n408_), .A1(ori_ori_n119_), .B0(ori_ori_n64_), .Y(ori_ori_n486_));
  NA4        o458(.A(ori_ori_n167_), .B(ori_ori_n106_), .C(ori_ori_n37_), .D(h), .Y(ori_ori_n487_));
  AN2        o459(.A(l), .B(k), .Y(ori_ori_n488_));
  NA3        o460(.A(ori_ori_n488_), .B(ori_ori_n84_), .C(ori_ori_n55_), .Y(ori_ori_n489_));
  OAI210     o461(.A0(ori_ori_n487_), .A1(g), .B0(ori_ori_n489_), .Y(ori_ori_n490_));
  NA2        o462(.A(ori_ori_n490_), .B(ori_ori_n486_), .Y(ori_ori_n491_));
  NA4        o463(.A(ori_ori_n491_), .B(ori_ori_n485_), .C(ori_ori_n480_), .D(ori_ori_n254_), .Y(ori_ori_n492_));
  NO4        o464(.A(ori_ori_n128_), .B(ori_ori_n284_), .C(ori_ori_n87_), .D(g), .Y(ori_ori_n493_));
  NA2        o465(.A(ori_ori_n493_), .B(ori_ori_n484_), .Y(ori_ori_n494_));
  INV        o466(.A(ori_ori_n34_), .Y(ori_ori_n495_));
  NA2        o467(.A(ori_ori_n425_), .B(ori_ori_n251_), .Y(ori_ori_n496_));
  NA2        o468(.A(ori_ori_n496_), .B(ori_ori_n494_), .Y(ori_ori_n497_));
  NO3        o469(.A(ori_ori_n222_), .B(ori_ori_n99_), .C(ori_ori_n36_), .Y(ori_ori_n498_));
  NAi21      o470(.An(ori_ori_n498_), .B(ori_ori_n489_), .Y(ori_ori_n499_));
  NA2        o471(.A(ori_ori_n499_), .B(ori_ori_n58_), .Y(ori_ori_n500_));
  INV        o472(.A(ori_ori_n500_), .Y(ori_ori_n501_));
  NA3        o473(.A(ori_ori_n466_), .B(ori_ori_n239_), .C(ori_ori_n276_), .Y(ori_ori_n502_));
  NA3        o474(.A(m), .B(l), .C(k), .Y(ori_ori_n503_));
  NA3        o475(.A(ori_ori_n88_), .B(k), .C(ori_ori_n67_), .Y(ori_ori_n504_));
  INV        o476(.A(ori_ori_n502_), .Y(ori_ori_n505_));
  NO4        o477(.A(ori_ori_n505_), .B(ori_ori_n501_), .C(ori_ori_n497_), .D(ori_ori_n492_), .Y(ori_ori_n506_));
  NA2        o478(.A(ori_ori_n425_), .B(ori_ori_n285_), .Y(ori_ori_n507_));
  INV        o479(.A(ori_ori_n359_), .Y(ori_ori_n508_));
  NA3        o480(.A(ori_ori_n508_), .B(ori_ori_n507_), .C(ori_ori_n195_), .Y(ori_ori_n509_));
  NA2        o481(.A(ori_ori_n488_), .B(ori_ori_n55_), .Y(ori_ori_n510_));
  NOi21      o482(.An(h), .B(j), .Y(ori_ori_n511_));
  NA2        o483(.A(ori_ori_n511_), .B(f), .Y(ori_ori_n512_));
  NO2        o484(.A(ori_ori_n923_), .B(ori_ori_n510_), .Y(ori_ori_n513_));
  AOI210     o485(.A0(ori_ori_n509_), .A1(l), .B0(ori_ori_n513_), .Y(ori_ori_n514_));
  INV        o486(.A(j), .Y(ori_ori_n515_));
  NO3        o487(.A(ori_ori_n212_), .B(ori_ori_n515_), .C(ori_ori_n35_), .Y(ori_ori_n516_));
  AOI210     o488(.A0(ori_ori_n380_), .A1(n), .B0(ori_ori_n393_), .Y(ori_ori_n517_));
  NA2        o489(.A(ori_ori_n517_), .B(ori_ori_n396_), .Y(ori_ori_n518_));
  AN3        o490(.A(ori_ori_n518_), .B(ori_ori_n516_), .C(ori_ori_n76_), .Y(ori_ori_n519_));
  NA2        o491(.A(ori_ori_n422_), .B(ori_ori_n217_), .Y(ori_ori_n520_));
  NAi31      o492(.An(ori_ori_n420_), .B(ori_ori_n73_), .C(ori_ori_n64_), .Y(ori_ori_n521_));
  NA2        o493(.A(ori_ori_n521_), .B(ori_ori_n520_), .Y(ori_ori_n522_));
  NO2        o494(.A(ori_ori_n212_), .B(ori_ori_n103_), .Y(ori_ori_n523_));
  AOI220     o495(.A0(ori_ori_n523_), .A1(ori_ori_n425_), .B0(ori_ori_n498_), .B1(ori_ori_n486_), .Y(ori_ori_n524_));
  NO2        o496(.A(ori_ori_n503_), .B(ori_ori_n71_), .Y(ori_ori_n525_));
  NA2        o497(.A(ori_ori_n525_), .B(ori_ori_n414_), .Y(ori_ori_n526_));
  NO2        o498(.A(ori_ori_n415_), .B(ori_ori_n91_), .Y(ori_ori_n527_));
  NA2        o499(.A(ori_ori_n527_), .B(ori_ori_n457_), .Y(ori_ori_n528_));
  NA3        o500(.A(ori_ori_n528_), .B(ori_ori_n526_), .C(ori_ori_n524_), .Y(ori_ori_n529_));
  OR3        o501(.A(ori_ori_n529_), .B(ori_ori_n522_), .C(ori_ori_n519_), .Y(ori_ori_n530_));
  NA3        o502(.A(ori_ori_n517_), .B(ori_ori_n396_), .C(ori_ori_n395_), .Y(ori_ori_n531_));
  NA4        o503(.A(ori_ori_n531_), .B(ori_ori_n167_), .C(ori_ori_n326_), .D(ori_ori_n31_), .Y(ori_ori_n532_));
  NO4        o504(.A(ori_ori_n352_), .B(ori_ori_n314_), .C(j), .D(f), .Y(ori_ori_n533_));
  NO2        o505(.A(ori_ori_n72_), .B(ori_ori_n39_), .Y(ori_ori_n534_));
  NA2        o506(.A(ori_ori_n534_), .B(ori_ori_n435_), .Y(ori_ori_n535_));
  NA2        o507(.A(ori_ori_n535_), .B(ori_ori_n532_), .Y(ori_ori_n536_));
  NO2        o508(.A(ori_ori_n450_), .B(ori_ori_n55_), .Y(ori_ori_n537_));
  AOI210     o509(.A0(ori_ori_n533_), .A1(ori_ori_n537_), .B0(ori_ori_n241_), .Y(ori_ori_n538_));
  OAI210     o510(.A0(ori_ori_n503_), .A1(ori_ori_n449_), .B0(ori_ori_n373_), .Y(ori_ori_n539_));
  NA3        o511(.A(ori_ori_n194_), .B(ori_ori_n50_), .C(b), .Y(ori_ori_n540_));
  AOI220     o512(.A0(ori_ori_n418_), .A1(ori_ori_n29_), .B0(ori_ori_n342_), .B1(ori_ori_n64_), .Y(ori_ori_n541_));
  NA2        o513(.A(ori_ori_n541_), .B(ori_ori_n540_), .Y(ori_ori_n542_));
  NA2        o514(.A(ori_ori_n542_), .B(ori_ori_n539_), .Y(ori_ori_n543_));
  NA2        o515(.A(ori_ori_n543_), .B(ori_ori_n538_), .Y(ori_ori_n544_));
  NO3        o516(.A(ori_ori_n544_), .B(ori_ori_n536_), .C(ori_ori_n530_), .Y(ori_ori_n545_));
  NO3        o517(.A(ori_ori_n247_), .B(ori_ori_n213_), .C(ori_ori_n87_), .Y(ori_ori_n546_));
  NA2        o518(.A(ori_ori_n546_), .B(ori_ori_n518_), .Y(ori_ori_n547_));
  NO3        o519(.A(ori_ori_n377_), .B(ori_ori_n74_), .C(h), .Y(ori_ori_n548_));
  NA2        o520(.A(ori_ori_n548_), .B(ori_ori_n482_), .Y(ori_ori_n549_));
  NA2        o521(.A(ori_ori_n549_), .B(ori_ori_n547_), .Y(ori_ori_n550_));
  OR2        o522(.A(ori_ori_n449_), .B(ori_ori_n72_), .Y(ori_ori_n551_));
  NOi31      o523(.An(b), .B(d), .C(a), .Y(ori_ori_n552_));
  NO2        o524(.A(ori_ori_n552_), .B(ori_ori_n417_), .Y(ori_ori_n553_));
  NO2        o525(.A(ori_ori_n553_), .B(n), .Y(ori_ori_n554_));
  BUFFER     o526(.A(ori_ori_n541_), .Y(ori_ori_n555_));
  NO2        o527(.A(ori_ori_n555_), .B(ori_ori_n551_), .Y(ori_ori_n556_));
  NO2        o528(.A(ori_ori_n394_), .B(ori_ori_n64_), .Y(ori_ori_n557_));
  NO2        o529(.A(ori_ori_n487_), .B(ori_ori_n286_), .Y(ori_ori_n558_));
  NO2        o530(.A(ori_ori_n465_), .B(n), .Y(ori_ori_n559_));
  BUFFER     o531(.A(ori_ori_n523_), .Y(ori_ori_n560_));
  AOI220     o532(.A0(ori_ori_n560_), .A1(ori_ori_n452_), .B0(ori_ori_n559_), .B1(ori_ori_n477_), .Y(ori_ori_n561_));
  NO2        o533(.A(ori_ori_n227_), .B(ori_ori_n184_), .Y(ori_ori_n562_));
  NA2        o534(.A(ori_ori_n73_), .B(ori_ori_n562_), .Y(ori_ori_n563_));
  INV        o535(.A(ori_ori_n563_), .Y(ori_ori_n564_));
  NAi21      o536(.An(ori_ori_n564_), .B(ori_ori_n561_), .Y(ori_ori_n565_));
  NO4        o537(.A(ori_ori_n565_), .B(ori_ori_n558_), .C(ori_ori_n556_), .D(ori_ori_n550_), .Y(ori_ori_n566_));
  NA4        o538(.A(ori_ori_n566_), .B(ori_ori_n545_), .C(ori_ori_n514_), .D(ori_ori_n506_), .Y(ori09));
  NA2        o539(.A(f), .B(e), .Y(ori_ori_n568_));
  NA2        o540(.A(ori_ori_n319_), .B(e), .Y(ori_ori_n569_));
  NO2        o541(.A(ori_ori_n569_), .B(ori_ori_n367_), .Y(ori_ori_n570_));
  INV        o542(.A(ori_ori_n570_), .Y(ori_ori_n571_));
  NA3        o543(.A(m), .B(l), .C(i), .Y(ori_ori_n572_));
  OAI220     o544(.A0(ori_ori_n415_), .A1(ori_ori_n572_), .B0(ori_ori_n256_), .B1(ori_ori_n378_), .Y(ori_ori_n573_));
  NA4        o545(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(g), .D(f), .Y(ori_ori_n574_));
  AN2        o546(.A(ori_ori_n573_), .B(ori_ori_n554_), .Y(ori_ori_n575_));
  INV        o547(.A(ori_ori_n244_), .Y(ori_ori_n576_));
  NO2        o548(.A(ori_ori_n96_), .B(ori_ori_n94_), .Y(ori_ori_n577_));
  NOi31      o549(.An(k), .B(m), .C(l), .Y(ori_ori_n578_));
  NO2        o550(.A(ori_ori_n246_), .B(ori_ori_n578_), .Y(ori_ori_n579_));
  AOI210     o551(.A0(ori_ori_n579_), .A1(ori_ori_n577_), .B0(ori_ori_n416_), .Y(ori_ori_n580_));
  NA2        o552(.A(ori_ori_n540_), .B(ori_ori_n237_), .Y(ori_ori_n581_));
  NA2        o553(.A(ori_ori_n248_), .B(ori_ori_n250_), .Y(ori_ori_n582_));
  OAI210     o554(.A0(ori_ori_n158_), .A1(ori_ori_n164_), .B0(ori_ori_n582_), .Y(ori_ori_n583_));
  AOI220     o555(.A0(ori_ori_n583_), .A1(ori_ori_n581_), .B0(ori_ori_n580_), .B1(ori_ori_n576_), .Y(ori_ori_n584_));
  NA2        o556(.A(ori_ori_n476_), .B(ori_ori_n103_), .Y(ori_ori_n585_));
  NA3        o557(.A(ori_ori_n585_), .B(ori_ori_n143_), .C(e), .Y(ori_ori_n586_));
  NA4        o558(.A(ori_ori_n586_), .B(ori_ori_n584_), .C(ori_ori_n426_), .D(ori_ori_n62_), .Y(ori_ori_n587_));
  NA2        o559(.A(f), .B(m), .Y(ori_ori_n588_));
  NO2        o560(.A(ori_ori_n588_), .B(ori_ori_n43_), .Y(ori_ori_n589_));
  NA2        o561(.A(ori_ori_n589_), .B(ori_ori_n389_), .Y(ori_ori_n590_));
  AN2        o562(.A(f), .B(d), .Y(ori_ori_n591_));
  NA3        o563(.A(ori_ori_n349_), .B(ori_ori_n591_), .C(ori_ori_n64_), .Y(ori_ori_n592_));
  NO3        o564(.A(ori_ori_n592_), .B(ori_ori_n55_), .C(ori_ori_n165_), .Y(ori_ori_n593_));
  NA2        o565(.A(j), .B(ori_ori_n593_), .Y(ori_ori_n594_));
  NA2        o566(.A(ori_ori_n594_), .B(ori_ori_n590_), .Y(ori_ori_n595_));
  NO3        o567(.A(ori_ori_n100_), .B(ori_ori_n232_), .C(ori_ori_n117_), .Y(ori_ori_n596_));
  NO2        o568(.A(ori_ori_n443_), .B(ori_ori_n232_), .Y(ori_ori_n597_));
  INV        o569(.A(ori_ori_n596_), .Y(ori_ori_n598_));
  NA3        o570(.A(ori_ori_n121_), .B(ori_ori_n84_), .C(g), .Y(ori_ori_n599_));
  OAI220     o571(.A0(ori_ori_n592_), .A1(ori_ori_n309_), .B0(ori_ori_n244_), .B1(ori_ori_n599_), .Y(ori_ori_n600_));
  NOi31      o572(.An(ori_ori_n173_), .B(ori_ori_n600_), .C(ori_ori_n215_), .Y(ori_ori_n601_));
  NA2        o573(.A(c), .B(ori_ori_n90_), .Y(ori_ori_n602_));
  NO2        o574(.A(ori_ori_n602_), .B(ori_ori_n295_), .Y(ori_ori_n603_));
  NA3        o575(.A(ori_ori_n603_), .B(ori_ori_n365_), .C(f), .Y(ori_ori_n604_));
  OR2        o576(.A(ori_ori_n449_), .B(ori_ori_n385_), .Y(ori_ori_n605_));
  INV        o577(.A(ori_ori_n605_), .Y(ori_ori_n606_));
  NA2        o578(.A(ori_ori_n553_), .B(ori_ori_n86_), .Y(ori_ori_n607_));
  NA2        o579(.A(ori_ori_n607_), .B(ori_ori_n606_), .Y(ori_ori_n608_));
  NA4        o580(.A(ori_ori_n608_), .B(ori_ori_n604_), .C(ori_ori_n601_), .D(ori_ori_n598_), .Y(ori_ori_n609_));
  NO4        o581(.A(ori_ori_n609_), .B(ori_ori_n595_), .C(ori_ori_n587_), .D(ori_ori_n575_), .Y(ori_ori_n610_));
  NO2        o582(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n611_));
  NO2        o583(.A(ori_ori_n180_), .B(ori_ori_n174_), .Y(ori_ori_n612_));
  AOI220     o584(.A0(ori_ori_n612_), .A1(ori_ori_n177_), .B0(ori_ori_n214_), .B1(ori_ori_n611_), .Y(ori_ori_n613_));
  NO2        o585(.A(ori_ori_n309_), .B(ori_ori_n568_), .Y(ori_ori_n614_));
  NA2        o586(.A(ori_ori_n614_), .B(ori_ori_n400_), .Y(ori_ori_n615_));
  NA2        o587(.A(ori_ori_n615_), .B(ori_ori_n613_), .Y(ori_ori_n616_));
  NA2        o588(.A(e), .B(d), .Y(ori_ori_n617_));
  OAI220     o589(.A0(ori_ori_n617_), .A1(c), .B0(ori_ori_n227_), .B1(d), .Y(ori_ori_n618_));
  NA3        o590(.A(ori_ori_n618_), .B(ori_ori_n331_), .C(ori_ori_n363_), .Y(ori_ori_n619_));
  AOI210     o591(.A0(ori_ori_n370_), .A1(ori_ori_n134_), .B0(ori_ori_n180_), .Y(ori_ori_n620_));
  AOI210     o592(.A0(ori_ori_n425_), .A1(ori_ori_n251_), .B0(ori_ori_n620_), .Y(ori_ori_n621_));
  NA3        o593(.A(ori_ori_n124_), .B(ori_ori_n65_), .C(ori_ori_n31_), .Y(ori_ori_n622_));
  NA3        o594(.A(ori_ori_n622_), .B(ori_ori_n621_), .C(ori_ori_n619_), .Y(ori_ori_n623_));
  NO2        o595(.A(ori_ori_n623_), .B(ori_ori_n616_), .Y(ori_ori_n624_));
  OR2        o596(.A(ori_ori_n478_), .B(ori_ori_n168_), .Y(ori_ori_n625_));
  OAI210     o597(.A0(ori_ori_n213_), .A1(j), .B0(ori_ori_n51_), .Y(ori_ori_n626_));
  NA2        o598(.A(ori_ori_n626_), .B(ori_ori_n597_), .Y(ori_ori_n627_));
  OAI210     o599(.A0(ori_ori_n569_), .A1(ori_ori_n125_), .B0(ori_ori_n627_), .Y(ori_ori_n628_));
  AN2        o600(.A(ori_ori_n581_), .B(ori_ori_n573_), .Y(ori_ori_n629_));
  NO2        o601(.A(ori_ori_n629_), .B(ori_ori_n628_), .Y(ori_ori_n630_));
  AN2        o602(.A(ori_ori_n130_), .B(f), .Y(ori_ori_n631_));
  OAI210     o603(.A0(ori_ori_n631_), .A1(ori_ori_n334_), .B0(ori_ori_n618_), .Y(ori_ori_n632_));
  AN3        o604(.A(ori_ori_n632_), .B(ori_ori_n630_), .C(ori_ori_n625_), .Y(ori_ori_n633_));
  NA4        o605(.A(ori_ori_n633_), .B(ori_ori_n624_), .C(ori_ori_n610_), .D(ori_ori_n571_), .Y(ori12));
  NO2        o606(.A(ori_ori_n329_), .B(c), .Y(ori_ori_n635_));
  NO4        o607(.A(ori_ori_n318_), .B(ori_ori_n196_), .C(ori_ori_n412_), .D(ori_ori_n165_), .Y(ori_ori_n636_));
  NA2        o608(.A(ori_ori_n636_), .B(ori_ori_n635_), .Y(ori_ori_n637_));
  NO2        o609(.A(ori_ori_n329_), .B(ori_ori_n90_), .Y(ori_ori_n638_));
  NO2        o610(.A(ori_ori_n449_), .B(ori_ori_n271_), .Y(ori_ori_n639_));
  NA2        o611(.A(ori_ori_n639_), .B(ori_ori_n387_), .Y(ori_ori_n640_));
  NA2        o612(.A(ori_ori_n640_), .B(ori_ori_n637_), .Y(ori_ori_n641_));
  AOI210     o613(.A0(ori_ori_n182_), .A1(ori_ori_n243_), .B0(ori_ori_n155_), .Y(ori_ori_n642_));
  OR2        o614(.A(ori_ori_n642_), .B(ori_ori_n636_), .Y(ori_ori_n643_));
  AOI210     o615(.A0(ori_ori_n240_), .A1(ori_ori_n282_), .B0(ori_ori_n165_), .Y(ori_ori_n644_));
  OAI210     o616(.A0(ori_ori_n644_), .A1(ori_ori_n643_), .B0(ori_ori_n291_), .Y(ori_ori_n645_));
  NO2        o617(.A(ori_ori_n415_), .B(ori_ori_n572_), .Y(ori_ori_n646_));
  NO2        o618(.A(ori_ori_n116_), .B(ori_ori_n184_), .Y(ori_ori_n647_));
  INV        o619(.A(ori_ori_n645_), .Y(ori_ori_n648_));
  OR2        o620(.A(ori_ori_n228_), .B(ori_ori_n638_), .Y(ori_ori_n649_));
  NA2        o621(.A(ori_ori_n649_), .B(ori_ori_n257_), .Y(ori_ori_n650_));
  NO3        o622(.A(ori_ori_n100_), .B(ori_ori_n117_), .C(ori_ori_n165_), .Y(ori_ori_n651_));
  NA2        o623(.A(ori_ori_n651_), .B(ori_ori_n380_), .Y(ori_ori_n652_));
  NA4        o624(.A(ori_ori_n319_), .B(ori_ori_n315_), .C(ori_ori_n135_), .D(g), .Y(ori_ori_n653_));
  NA3        o625(.A(ori_ori_n653_), .B(ori_ori_n652_), .C(ori_ori_n650_), .Y(ori_ori_n654_));
  NO3        o626(.A(ori_ori_n654_), .B(ori_ori_n648_), .C(ori_ori_n641_), .Y(ori_ori_n655_));
  NA2        o627(.A(ori_ori_n394_), .B(ori_ori_n110_), .Y(ori_ori_n656_));
  NOi21      o628(.An(ori_ori_n31_), .B(ori_ori_n443_), .Y(ori_ori_n657_));
  NA2        o629(.A(ori_ori_n657_), .B(ori_ori_n656_), .Y(ori_ori_n658_));
  OAI210     o630(.A0(ori_ori_n195_), .A1(ori_ori_n37_), .B0(ori_ori_n658_), .Y(ori_ori_n659_));
  INV        o631(.A(ori_ori_n226_), .Y(ori_ori_n660_));
  NO2        o632(.A(ori_ori_n362_), .B(ori_ori_n213_), .Y(ori_ori_n661_));
  INV        o633(.A(ori_ori_n661_), .Y(ori_ori_n662_));
  NO2        o634(.A(ori_ori_n662_), .B(ori_ori_n110_), .Y(ori_ori_n663_));
  INV        o635(.A(ori_ori_n265_), .Y(ori_ori_n664_));
  NO4        o636(.A(ori_ori_n664_), .B(ori_ori_n663_), .C(ori_ori_n660_), .D(ori_ori_n659_), .Y(ori_ori_n665_));
  NA2        o637(.A(ori_ori_n251_), .B(g), .Y(ori_ori_n666_));
  NA2        o638(.A(ori_ori_n123_), .B(i), .Y(ori_ori_n667_));
  NA2        o639(.A(ori_ori_n38_), .B(i), .Y(ori_ori_n668_));
  NO2        o640(.A(ori_ori_n668_), .B(ori_ori_n154_), .Y(ori_ori_n669_));
  INV        o641(.A(ori_ori_n669_), .Y(ori_ori_n670_));
  NO2        o642(.A(ori_ori_n110_), .B(ori_ori_n64_), .Y(ori_ori_n671_));
  OR2        o643(.A(ori_ori_n671_), .B(ori_ori_n393_), .Y(ori_ori_n672_));
  INV        o644(.A(ori_ori_n672_), .Y(ori_ori_n673_));
  OAI220     o645(.A0(ori_ori_n673_), .A1(ori_ori_n666_), .B0(ori_ori_n670_), .B1(ori_ori_n237_), .Y(ori_ori_n674_));
  NA2        o646(.A(ori_ori_n574_), .B(ori_ori_n317_), .Y(ori_ori_n675_));
  NO2        o647(.A(ori_ori_n271_), .B(ori_ori_n71_), .Y(ori_ori_n676_));
  NA2        o648(.A(ori_ori_n676_), .B(ori_ori_n185_), .Y(ori_ori_n677_));
  NO2        o649(.A(ori_ori_n337_), .B(ori_ori_n165_), .Y(ori_ori_n678_));
  AOI220     o650(.A0(ori_ori_n678_), .A1(ori_ori_n275_), .B0(ori_ori_n649_), .B1(ori_ori_n169_), .Y(ori_ori_n679_));
  AOI220     o651(.A0(ori_ori_n639_), .A1(ori_ori_n647_), .B0(ori_ori_n414_), .B1(ori_ori_n70_), .Y(ori_ori_n680_));
  NA3        o652(.A(ori_ori_n680_), .B(ori_ori_n679_), .C(ori_ori_n677_), .Y(ori_ori_n681_));
  OAI210     o653(.A0(ori_ori_n675_), .A1(ori_ori_n646_), .B0(ori_ori_n387_), .Y(ori_ori_n682_));
  NA2        o654(.A(ori_ori_n437_), .B(ori_ori_n380_), .Y(ori_ori_n683_));
  NA2        o655(.A(ori_ori_n683_), .B(ori_ori_n682_), .Y(ori_ori_n684_));
  NO3        o656(.A(ori_ori_n684_), .B(ori_ori_n681_), .C(ori_ori_n674_), .Y(ori_ori_n685_));
  NAi31      o657(.An(ori_ori_n107_), .B(ori_ori_n303_), .C(n), .Y(ori_ori_n686_));
  NO3        o658(.A(ori_ori_n94_), .B(ori_ori_n246_), .C(ori_ori_n578_), .Y(ori_ori_n687_));
  NO2        o659(.A(ori_ori_n687_), .B(ori_ori_n686_), .Y(ori_ori_n688_));
  NO3        o660(.A(h), .B(ori_ori_n107_), .C(ori_ori_n295_), .Y(ori_ori_n689_));
  AOI210     o661(.A0(ori_ori_n689_), .A1(ori_ori_n357_), .B0(ori_ori_n688_), .Y(ori_ori_n690_));
  INV        o662(.A(ori_ori_n690_), .Y(ori_ori_n691_));
  NA2        o663(.A(ori_ori_n180_), .B(ori_ori_n126_), .Y(ori_ori_n692_));
  NO3        o664(.A(ori_ori_n217_), .B(ori_ori_n319_), .C(ori_ori_n130_), .Y(ori_ori_n693_));
  NOi31      o665(.An(ori_ori_n692_), .B(ori_ori_n693_), .C(ori_ori_n165_), .Y(ori_ori_n694_));
  NAi21      o666(.An(ori_ori_n394_), .B(ori_ori_n678_), .Y(ori_ori_n695_));
  INV        o667(.A(ori_ori_n695_), .Y(ori_ori_n696_));
  NA2        o668(.A(ori_ori_n642_), .B(ori_ori_n635_), .Y(ori_ori_n697_));
  OAI220     o669(.A0(ori_ori_n639_), .A1(ori_ori_n646_), .B0(ori_ori_n389_), .B1(ori_ori_n308_), .Y(ori_ori_n698_));
  NA3        o670(.A(ori_ori_n698_), .B(ori_ori_n697_), .C(ori_ori_n423_), .Y(ori_ori_n699_));
  OAI210     o671(.A0(ori_ori_n642_), .A1(ori_ori_n636_), .B0(ori_ori_n692_), .Y(ori_ori_n700_));
  INV        o672(.A(ori_ori_n236_), .Y(ori_ori_n701_));
  NA2        o673(.A(ori_ori_n701_), .B(ori_ori_n700_), .Y(ori_ori_n702_));
  OR2        o674(.A(ori_ori_n702_), .B(ori_ori_n699_), .Y(ori_ori_n703_));
  NO4        o675(.A(ori_ori_n703_), .B(ori_ori_n696_), .C(ori_ori_n694_), .D(ori_ori_n691_), .Y(ori_ori_n704_));
  NA4        o676(.A(ori_ori_n704_), .B(ori_ori_n685_), .C(ori_ori_n665_), .D(ori_ori_n655_), .Y(ori13));
  AN2        o677(.A(d), .B(c), .Y(ori_ori_n706_));
  NA2        o678(.A(ori_ori_n706_), .B(ori_ori_n90_), .Y(ori_ori_n707_));
  NAi32      o679(.An(f), .Bn(e), .C(c), .Y(ori_ori_n708_));
  NO3        o680(.A(m), .B(i), .C(h), .Y(ori_ori_n709_));
  NA3        o681(.A(k), .B(j), .C(i), .Y(ori_ori_n710_));
  NO2        o682(.A(f), .B(c), .Y(ori_ori_n711_));
  NOi21      o683(.An(ori_ori_n711_), .B(ori_ori_n318_), .Y(ori_ori_n712_));
  AN3        o684(.A(g), .B(f), .C(c), .Y(ori_ori_n713_));
  NA3        o685(.A(l), .B(k), .C(j), .Y(ori_ori_n714_));
  NA2        o686(.A(i), .B(h), .Y(ori_ori_n715_));
  NO3        o687(.A(ori_ori_n715_), .B(ori_ori_n714_), .C(ori_ori_n100_), .Y(ori_ori_n716_));
  NO3        o688(.A(ori_ori_n108_), .B(ori_ori_n210_), .C(ori_ori_n165_), .Y(ori_ori_n717_));
  NA4        o689(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(g), .D(ori_ori_n164_), .Y(ori_ori_n718_));
  INV        o690(.A(ori_ori_n718_), .Y(ori_ori_n719_));
  NOi41      o691(.An(ori_ori_n551_), .B(ori_ori_n583_), .C(ori_ori_n573_), .D(ori_ori_n495_), .Y(ori_ori_n720_));
  OAI220     o692(.A0(ori_ori_n720_), .A1(ori_ori_n469_), .B0(ori_ori_n718_), .B1(ori_ori_n413_), .Y(ori_ori_n721_));
  NOi31      o693(.An(m), .B(n), .C(f), .Y(ori_ori_n722_));
  NO2        o694(.A(ori_ori_n605_), .B(ori_ori_n307_), .Y(ori_ori_n723_));
  INV        o695(.A(ori_ori_n210_), .Y(ori_ori_n724_));
  NO3        o696(.A(ori_ori_n723_), .B(ori_ori_n721_), .C(ori_ori_n564_), .Y(ori_ori_n725_));
  NA2        o697(.A(c), .B(b), .Y(ori_ori_n726_));
  NO2        o698(.A(ori_ori_n481_), .B(ori_ori_n726_), .Y(ori_ori_n727_));
  INV        o699(.A(ori_ori_n300_), .Y(ori_ori_n728_));
  OAI210     o700(.A0(ori_ori_n728_), .A1(ori_ori_n589_), .B0(ori_ori_n727_), .Y(ori_ori_n729_));
  NAi21      o701(.An(ori_ori_n305_), .B(ori_ori_n727_), .Y(ori_ori_n730_));
  NA2        o702(.A(ori_ori_n390_), .B(ori_ori_n724_), .Y(ori_ori_n731_));
  NA2        o703(.A(ori_ori_n731_), .B(ori_ori_n730_), .Y(ori_ori_n732_));
  INV        o704(.A(ori_ori_n732_), .Y(ori_ori_n733_));
  NA2        o705(.A(ori_ori_n400_), .B(ori_ori_n297_), .Y(ori_ori_n734_));
  NO2        o706(.A(ori_ori_n267_), .B(ori_ori_n266_), .Y(ori_ori_n735_));
  NA4        o707(.A(ori_ori_n734_), .B(ori_ori_n733_), .C(ori_ori_n729_), .D(ori_ori_n725_), .Y(ori00));
  NA2        o708(.A(ori_ori_n614_), .B(ori_ori_n647_), .Y(ori_ori_n737_));
  INV        o709(.A(ori_ori_n737_), .Y(ori_ori_n738_));
  NA2        o710(.A(ori_ori_n365_), .B(f), .Y(ori_ori_n739_));
  OAI210     o711(.A0(ori_ori_n687_), .A1(ori_ori_n35_), .B0(ori_ori_n439_), .Y(ori_ori_n740_));
  NA3        o712(.A(ori_ori_n740_), .B(ori_ori_n201_), .C(n), .Y(ori_ori_n741_));
  AOI210     o713(.A0(ori_ori_n741_), .A1(ori_ori_n739_), .B0(ori_ori_n707_), .Y(ori_ori_n742_));
  NO2        o714(.A(ori_ori_n742_), .B(ori_ori_n738_), .Y(ori_ori_n743_));
  NA3        o715(.A(ori_ori_n124_), .B(ori_ori_n38_), .C(ori_ori_n37_), .Y(ori_ori_n744_));
  NA3        o716(.A(d), .B(ori_ori_n47_), .C(b), .Y(ori_ori_n745_));
  NO2        o717(.A(ori_ori_n745_), .B(ori_ori_n744_), .Y(ori_ori_n746_));
  INV        o718(.A(ori_ori_n407_), .Y(ori_ori_n747_));
  NO3        o719(.A(ori_ori_n747_), .B(ori_ori_n746_), .C(ori_ori_n735_), .Y(ori_ori_n748_));
  NA3        o720(.A(ori_ori_n276_), .B(ori_ori_n172_), .C(g), .Y(ori_ori_n749_));
  OR2        o721(.A(ori_ori_n749_), .B(ori_ori_n745_), .Y(ori_ori_n750_));
  NO2        o722(.A(h), .B(g), .Y(ori_ori_n751_));
  NA4        o723(.A(ori_ori_n357_), .B(e), .C(ori_ori_n751_), .D(b), .Y(ori_ori_n752_));
  NO2        o724(.A(ori_ori_n72_), .B(ori_ori_n71_), .Y(ori_ori_n753_));
  AOI220     o725(.A0(ori_ori_n753_), .A1(ori_ori_n383_), .B0(ori_ori_n651_), .B1(ori_ori_n406_), .Y(ori_ori_n754_));
  NA2        o726(.A(ori_ori_n223_), .B(ori_ori_n192_), .Y(ori_ori_n755_));
  NA4        o727(.A(ori_ori_n755_), .B(ori_ori_n754_), .C(ori_ori_n752_), .D(ori_ori_n750_), .Y(ori_ori_n756_));
  INV        o728(.A(ori_ori_n756_), .Y(ori_ori_n757_));
  AOI210     o729(.A0(ori_ori_n192_), .A1(ori_ori_n251_), .B0(ori_ori_n409_), .Y(ori_ori_n758_));
  AN3        o730(.A(ori_ori_n758_), .B(ori_ori_n757_), .C(ori_ori_n748_), .Y(ori_ori_n759_));
  NA3        o731(.A(ori_ori_n722_), .B(ori_ori_n419_), .C(ori_ori_n344_), .Y(ori_ori_n760_));
  INV        o732(.A(ori_ori_n760_), .Y(ori_ori_n761_));
  NA2        o733(.A(ori_ori_n719_), .B(ori_ori_n383_), .Y(ori_ori_n762_));
  NA4        o734(.A(ori_ori_n442_), .B(ori_ori_n159_), .C(ori_ori_n172_), .D(ori_ori_n123_), .Y(ori_ori_n763_));
  NA2        o735(.A(ori_ori_n763_), .B(ori_ori_n762_), .Y(ori_ori_n764_));
  NA2        o736(.A(ori_ori_n400_), .B(ori_ori_n297_), .Y(ori_ori_n765_));
  NA2        o737(.A(n), .B(e), .Y(ori_ori_n766_));
  NO2        o738(.A(ori_ori_n766_), .B(ori_ori_n112_), .Y(ori_ori_n767_));
  NA2        o739(.A(ori_ori_n767_), .B(ori_ori_n206_), .Y(ori_ori_n768_));
  NA2        o740(.A(ori_ori_n768_), .B(ori_ori_n765_), .Y(ori_ori_n769_));
  NA2        o741(.A(ori_ori_n767_), .B(ori_ori_n580_), .Y(ori_ori_n770_));
  AOI220     o742(.A0(ori_ori_n657_), .A1(ori_ori_n406_), .B0(ori_ori_n442_), .B1(ori_ori_n189_), .Y(ori_ori_n771_));
  NA3        o743(.A(ori_ori_n771_), .B(ori_ori_n770_), .C(ori_ori_n590_), .Y(ori_ori_n772_));
  NO4        o744(.A(ori_ori_n772_), .B(ori_ori_n769_), .C(ori_ori_n764_), .D(ori_ori_n761_), .Y(ori_ori_n773_));
  NA3        o745(.A(ori_ori_n773_), .B(ori_ori_n759_), .C(ori_ori_n743_), .Y(ori01));
  INV        o746(.A(ori_ori_n209_), .Y(ori_ori_n775_));
  NA2        o747(.A(ori_ori_n287_), .B(i), .Y(ori_ori_n776_));
  NA3        o748(.A(ori_ori_n776_), .B(ori_ori_n775_), .C(ori_ori_n697_), .Y(ori_ori_n777_));
  NA2        o749(.A(ori_ori_n414_), .B(ori_ori_n70_), .Y(ori_ori_n778_));
  NA2        o750(.A(ori_ori_n394_), .B(ori_ori_n205_), .Y(ori_ori_n779_));
  NA2        o751(.A(ori_ori_n661_), .B(ori_ori_n779_), .Y(ori_ori_n780_));
  NA4        o752(.A(ori_ori_n780_), .B(ori_ori_n778_), .C(ori_ori_n627_), .D(ori_ori_n238_), .Y(ori_ori_n781_));
  NA2        o753(.A(ori_ori_n763_), .B(ori_ori_n613_), .Y(ori_ori_n782_));
  NO2        o754(.A(ori_ori_n456_), .B(ori_ori_n368_), .Y(ori_ori_n783_));
  NA2        o755(.A(ori_ori_n783_), .B(ori_ori_n104_), .Y(ori_ori_n784_));
  NO4        o756(.A(ori_ori_n784_), .B(ori_ori_n782_), .C(ori_ori_n781_), .D(ori_ori_n777_), .Y(ori_ori_n785_));
  AOI210     o757(.A0(ori_ori_n158_), .A1(ori_ori_n69_), .B0(ori_ori_n164_), .Y(ori_ori_n786_));
  OAI210     o758(.A0(ori_ori_n554_), .A1(ori_ori_n308_), .B0(ori_ori_n786_), .Y(ori_ori_n787_));
  OAI210     o759(.A0(ori_ori_n260_), .A1(ori_ori_n31_), .B0(m), .Y(ori_ori_n788_));
  OR2        o760(.A(ori_ori_n788_), .B(ori_ori_n237_), .Y(ori_ori_n789_));
  NA2        o761(.A(ori_ori_n789_), .B(ori_ori_n787_), .Y(ori_ori_n790_));
  NA2        o762(.A(ori_ori_n208_), .B(ori_ori_n149_), .Y(ori_ori_n791_));
  NA2        o763(.A(ori_ori_n791_), .B(ori_ori_n452_), .Y(ori_ori_n792_));
  NA2        o764(.A(ori_ori_n231_), .B(ori_ori_n457_), .Y(ori_ori_n793_));
  NA3        o765(.A(ori_ori_n793_), .B(ori_ori_n792_), .C(ori_ori_n535_), .Y(ori_ori_n794_));
  NO2        o766(.A(ori_ori_n794_), .B(ori_ori_n790_), .Y(ori_ori_n795_));
  NO2        o767(.A(ori_ori_n160_), .B(ori_ori_n86_), .Y(ori_ori_n796_));
  NO2        o768(.A(ori_ori_n796_), .B(ori_ori_n746_), .Y(ori_ori_n797_));
  INV        o769(.A(ori_ori_n797_), .Y(ori_ori_n798_));
  NO2        o770(.A(ori_ori_n667_), .B(ori_ori_n181_), .Y(ori_ori_n799_));
  NO2        o771(.A(ori_ori_n668_), .B(ori_ori_n396_), .Y(ori_ori_n800_));
  OAI210     o772(.A0(ori_ori_n800_), .A1(ori_ori_n799_), .B0(ori_ori_n246_), .Y(ori_ori_n801_));
  NO3        o773(.A(ori_ori_n61_), .B(ori_ori_n213_), .C(ori_ori_n37_), .Y(ori_ori_n802_));
  NA2        o774(.A(ori_ori_n802_), .B(ori_ori_n393_), .Y(ori_ori_n803_));
  INV        o775(.A(ori_ori_n803_), .Y(ori_ori_n804_));
  OR2        o776(.A(ori_ori_n749_), .B(ori_ori_n745_), .Y(ori_ori_n805_));
  NA2        o777(.A(ori_ori_n802_), .B(ori_ori_n557_), .Y(ori_ori_n806_));
  NA3        o778(.A(ori_ori_n806_), .B(ori_ori_n805_), .C(ori_ori_n279_), .Y(ori_ori_n807_));
  NOi41      o779(.An(ori_ori_n801_), .B(ori_ori_n807_), .C(ori_ori_n804_), .D(ori_ori_n798_), .Y(ori_ori_n808_));
  NO2        o780(.A(ori_ori_n99_), .B(ori_ori_n37_), .Y(ori_ori_n809_));
  NO2        o781(.A(ori_ori_n37_), .B(ori_ori_n35_), .Y(ori_ori_n810_));
  AO220      o782(.A0(ori_ori_n810_), .A1(ori_ori_n425_), .B0(ori_ori_n809_), .B1(ori_ori_n486_), .Y(ori_ori_n811_));
  NA2        o783(.A(ori_ori_n811_), .B(ori_ori_n246_), .Y(ori_ori_n812_));
  NO3        o784(.A(ori_ori_n715_), .B(ori_ori_n131_), .C(ori_ori_n67_), .Y(ori_ori_n813_));
  NA2        o785(.A(ori_ori_n802_), .B(ori_ori_n671_), .Y(ori_ori_n814_));
  NA2        o786(.A(ori_ori_n814_), .B(ori_ori_n812_), .Y(ori_ori_n815_));
  NO2        o787(.A(ori_ori_n422_), .B(ori_ori_n421_), .Y(ori_ori_n816_));
  NO4        o788(.A(ori_ori_n715_), .B(ori_ori_n816_), .C(ori_ori_n129_), .D(ori_ori_n67_), .Y(ori_ori_n817_));
  NO3        o789(.A(ori_ori_n817_), .B(ori_ori_n815_), .C(ori_ori_n432_), .Y(ori_ori_n818_));
  NA4        o790(.A(ori_ori_n818_), .B(ori_ori_n808_), .C(ori_ori_n795_), .D(ori_ori_n785_), .Y(ori06));
  NO2        o791(.A(ori_ori_n174_), .B(ori_ori_n79_), .Y(ori_ori_n820_));
  OAI210     o792(.A0(ori_ori_n820_), .A1(ori_ori_n813_), .B0(ori_ori_n275_), .Y(ori_ori_n821_));
  NA2        o793(.A(ori_ori_n821_), .B(ori_ori_n801_), .Y(ori_ori_n822_));
  NO3        o794(.A(ori_ori_n822_), .B(ori_ori_n804_), .C(ori_ori_n200_), .Y(ori_ori_n823_));
  NO2        o795(.A(ori_ori_n213_), .B(ori_ori_n37_), .Y(ori_ori_n824_));
  NA2        o796(.A(ori_ori_n824_), .B(ori_ori_n672_), .Y(ori_ori_n825_));
  AOI210     o797(.A0(ori_ori_n824_), .A1(ori_ori_n397_), .B0(ori_ori_n811_), .Y(ori_ori_n826_));
  AOI210     o798(.A0(ori_ori_n826_), .A1(ori_ori_n825_), .B0(ori_ori_n243_), .Y(ori_ori_n827_));
  INV        o799(.A(ori_ori_n69_), .Y(ori_ori_n828_));
  NA2        o800(.A(ori_ori_n828_), .B(ori_ori_n435_), .Y(ori_ori_n829_));
  OAI210     o801(.A0(ori_ori_n338_), .A1(ori_ori_n193_), .B0(ori_ori_n622_), .Y(ori_ori_n830_));
  INV        o802(.A(ori_ori_n830_), .Y(ori_ori_n831_));
  NA2        o803(.A(ori_ori_n831_), .B(ori_ori_n829_), .Y(ori_ori_n832_));
  NO2        o804(.A(ori_ori_n512_), .B(ori_ori_n922_), .Y(ori_ori_n833_));
  INV        o805(.A(ori_ori_n457_), .Y(ori_ori_n834_));
  NOi21      o806(.An(ori_ori_n833_), .B(ori_ori_n834_), .Y(ori_ori_n835_));
  AN2        o807(.A(ori_ori_n657_), .B(ori_ori_n438_), .Y(ori_ori_n836_));
  NO4        o808(.A(ori_ori_n836_), .B(ori_ori_n835_), .C(ori_ori_n832_), .D(ori_ori_n827_), .Y(ori_ori_n837_));
  NO2        o809(.A(ori_ori_n504_), .B(ori_ori_n39_), .Y(ori_ori_n838_));
  NA2        o810(.A(ori_ori_n261_), .B(ori_ori_n838_), .Y(ori_ori_n839_));
  NO3        o811(.A(ori_ori_n188_), .B(ori_ori_n79_), .C(ori_ori_n210_), .Y(ori_ori_n840_));
  OAI220     o812(.A0(ori_ori_n478_), .A1(ori_ori_n193_), .B0(ori_ori_n367_), .B1(ori_ori_n370_), .Y(ori_ori_n841_));
  INV        o813(.A(k), .Y(ori_ori_n842_));
  NO3        o814(.A(ori_ori_n842_), .B(ori_ori_n416_), .C(j), .Y(ori_ori_n843_));
  NO3        o815(.A(ori_ori_n841_), .B(ori_ori_n840_), .C(ori_ori_n723_), .Y(ori_ori_n844_));
  NA3        o816(.A(ori_ori_n844_), .B(ori_ori_n839_), .C(ori_ori_n771_), .Y(ori_ori_n845_));
  NA2        o817(.A(ori_ori_n843_), .B(ori_ori_n537_), .Y(ori_ori_n846_));
  INV        o818(.A(ori_ori_n846_), .Y(ori_ori_n847_));
  AN2        o819(.A(ori_ori_n636_), .B(ori_ori_n635_), .Y(ori_ori_n848_));
  NO2        o820(.A(ori_ori_n848_), .B(ori_ori_n359_), .Y(ori_ori_n849_));
  NA2        o821(.A(ori_ori_n849_), .B(ori_ori_n806_), .Y(ori_ori_n850_));
  NAi21      o822(.An(j), .B(i), .Y(ori_ori_n851_));
  NO4        o823(.A(ori_ori_n816_), .B(ori_ori_n851_), .C(ori_ori_n318_), .D(ori_ori_n183_), .Y(ori_ori_n852_));
  NO4        o824(.A(ori_ori_n852_), .B(ori_ori_n850_), .C(ori_ori_n847_), .D(ori_ori_n845_), .Y(ori_ori_n853_));
  NA4        o825(.A(ori_ori_n853_), .B(ori_ori_n837_), .C(ori_ori_n823_), .D(ori_ori_n818_), .Y(ori07));
  NAi32      o826(.An(m), .Bn(b), .C(n), .Y(ori_ori_n855_));
  NO3        o827(.A(ori_ori_n855_), .B(g), .C(f), .Y(ori_ori_n856_));
  NOi31      o828(.An(n), .B(m), .C(b), .Y(ori_ori_n857_));
  NO3        o829(.A(ori_ori_n100_), .B(ori_ori_n326_), .C(h), .Y(ori_ori_n858_));
  NO2        o830(.A(ori_ori_n708_), .B(ori_ori_n318_), .Y(ori_ori_n859_));
  NO2        o831(.A(ori_ori_n710_), .B(ori_ori_n216_), .Y(ori_ori_n860_));
  NO2        o832(.A(ori_ori_n859_), .B(ori_ori_n856_), .Y(ori_ori_n861_));
  NA3        o833(.A(ori_ori_n475_), .B(ori_ori_n461_), .C(ori_ori_n87_), .Y(ori_ori_n862_));
  NO3        o834(.A(ori_ori_n318_), .B(d), .C(c), .Y(ori_ori_n863_));
  NO2        o835(.A(ori_ori_n329_), .B(a), .Y(ori_ori_n864_));
  NA2        o836(.A(ori_ori_n864_), .B(ori_ori_n88_), .Y(ori_ori_n865_));
  NOi31      o837(.An(m), .B(n), .C(b), .Y(ori_ori_n866_));
  NOi31      o838(.An(f), .B(d), .C(c), .Y(ori_ori_n867_));
  NA2        o839(.A(ori_ori_n867_), .B(ori_ori_n866_), .Y(ori_ori_n868_));
  NA2        o840(.A(ori_ori_n713_), .B(e), .Y(ori_ori_n869_));
  NO2        o841(.A(ori_ori_n869_), .B(ori_ori_n318_), .Y(ori_ori_n870_));
  NO2        o842(.A(i), .B(h), .Y(ori_ori_n871_));
  NO2        o843(.A(ori_ori_n709_), .B(ori_ori_n870_), .Y(ori_ori_n872_));
  AN3        o844(.A(ori_ori_n872_), .B(ori_ori_n868_), .C(ori_ori_n865_), .Y(ori_ori_n873_));
  NA2        o845(.A(ori_ori_n857_), .B(ori_ori_n272_), .Y(ori_ori_n874_));
  INV        o846(.A(ori_ori_n874_), .Y(ori_ori_n875_));
  INV        o847(.A(ori_ori_n716_), .Y(ori_ori_n876_));
  NAi21      o848(.An(ori_ori_n875_), .B(ori_ori_n876_), .Y(ori_ori_n877_));
  NO4        o849(.A(ori_ori_n100_), .B(g), .C(f), .D(e), .Y(ori_ori_n878_));
  NA2        o850(.A(ori_ori_n722_), .B(ori_ori_n295_), .Y(ori_ori_n879_));
  INV        o851(.A(ori_ori_n879_), .Y(ori_ori_n880_));
  NO2        o852(.A(ori_ori_n880_), .B(ori_ori_n877_), .Y(ori_ori_n881_));
  NA4        o853(.A(ori_ori_n881_), .B(ori_ori_n873_), .C(ori_ori_n862_), .D(ori_ori_n861_), .Y(ori_ori_n882_));
  NO2        o854(.A(ori_ori_n726_), .B(ori_ori_n85_), .Y(ori_ori_n883_));
  NO2        o855(.A(ori_ori_n284_), .B(j), .Y(ori_ori_n884_));
  NA2        o856(.A(ori_ori_n871_), .B(ori_ori_n722_), .Y(ori_ori_n885_));
  NA2        o857(.A(ori_ori_n712_), .B(ori_ori_n115_), .Y(ori_ori_n886_));
  NA2        o858(.A(ori_ori_n886_), .B(ori_ori_n885_), .Y(ori_ori_n887_));
  NA2        o859(.A(ori_ori_n884_), .B(ori_ori_n120_), .Y(ori_ori_n888_));
  INV        o860(.A(ori_ori_n888_), .Y(ori_ori_n889_));
  NO2        o861(.A(ori_ori_n889_), .B(ori_ori_n887_), .Y(ori_ori_n890_));
  INV        o862(.A(ori_ori_n40_), .Y(ori_ori_n891_));
  NA2        o863(.A(ori_ori_n891_), .B(ori_ori_n751_), .Y(ori_ori_n892_));
  INV        o864(.A(ori_ori_n892_), .Y(ori_ori_n893_));
  NO2        o865(.A(ori_ori_n174_), .B(ori_ori_n131_), .Y(ori_ori_n894_));
  NO2        o866(.A(ori_ori_n894_), .B(ori_ori_n893_), .Y(ori_ori_n895_));
  NA2        o867(.A(ori_ori_n883_), .B(f), .Y(ori_ori_n896_));
  NO2        o868(.A(ori_ori_n921_), .B(ori_ori_n896_), .Y(ori_ori_n897_));
  NO2        o869(.A(ori_ori_n851_), .B(ori_ori_n129_), .Y(ori_ori_n898_));
  NA2        o870(.A(h), .B(ori_ori_n898_), .Y(ori_ori_n899_));
  INV        o871(.A(ori_ori_n213_), .Y(ori_ori_n900_));
  NA2        o872(.A(ori_ori_n900_), .B(ori_ori_n386_), .Y(ori_ori_n901_));
  NA2        o873(.A(ori_ori_n901_), .B(ori_ori_n899_), .Y(ori_ori_n902_));
  NO2        o874(.A(ori_ori_n902_), .B(ori_ori_n897_), .Y(ori_ori_n903_));
  NA3        o875(.A(ori_ori_n903_), .B(ori_ori_n895_), .C(ori_ori_n890_), .Y(ori_ori_n904_));
  NA2        o876(.A(h), .B(ori_ori_n860_), .Y(ori_ori_n905_));
  OAI210     o877(.A0(ori_ori_n878_), .A1(ori_ori_n857_), .B0(ori_ori_n602_), .Y(ori_ori_n906_));
  NA2        o878(.A(ori_ori_n906_), .B(ori_ori_n905_), .Y(ori_ori_n907_));
  NA2        o879(.A(ori_ori_n85_), .B(ori_ori_n866_), .Y(ori_ori_n908_));
  INV        o880(.A(ori_ori_n908_), .Y(ori_ori_n909_));
  NO2        o881(.A(ori_ori_n909_), .B(ori_ori_n907_), .Y(ori_ori_n910_));
  INV        o882(.A(ori_ori_n428_), .Y(ori_ori_n911_));
  OR2        o883(.A(h), .B(ori_ori_n384_), .Y(ori_ori_n912_));
  NO2        o884(.A(ori_ori_n912_), .B(ori_ori_n129_), .Y(ori_ori_n913_));
  NA2        o885(.A(ori_ori_n717_), .B(ori_ori_n172_), .Y(ori_ori_n914_));
  INV        o886(.A(ori_ori_n914_), .Y(ori_ori_n915_));
  NO3        o887(.A(ori_ori_n915_), .B(ori_ori_n913_), .C(ori_ori_n863_), .Y(ori_ori_n916_));
  NA3        o888(.A(ori_ori_n916_), .B(ori_ori_n911_), .C(ori_ori_n910_), .Y(ori_ori_n917_));
  OR4        o889(.A(ori_ori_n858_), .B(ori_ori_n917_), .C(ori_ori_n904_), .D(ori_ori_n882_), .Y(ori04));
  INV        o890(.A(ori_ori_n88_), .Y(ori_ori_n921_));
  INV        o891(.A(k), .Y(ori_ori_n922_));
  INV        o892(.A(ori_ori_n468_), .Y(ori_ori_n923_));
  INV        o893(.A(ori_ori_n415_), .Y(ori_ori_n924_));
  ZERO       o894(.Y(ori02));
  ZERO       o895(.Y(ori03));
  ZERO       o896(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(g), .Y(mai_mai_n50_));
  INV        m0022(.A(mai_mai_n50_), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0024(.A0(mai_mai_n49_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n53_));
  INV        m0025(.A(c), .Y(mai_mai_n54_));
  NA2        m0026(.A(e), .B(b), .Y(mai_mai_n55_));
  NO2        m0027(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  INV        m0028(.A(d), .Y(mai_mai_n57_));
  NA3        m0029(.A(g), .B(mai_mai_n57_), .C(a), .Y(mai_mai_n58_));
  NAi21      m0030(.An(i), .B(h), .Y(mai_mai_n59_));
  NAi31      m0031(.An(i), .B(l), .C(j), .Y(mai_mai_n60_));
  OAI210     m0032(.A0(mai_mai_n60_), .A1(mai_mai_n49_), .B0(mai_mai_n44_), .Y(mai_mai_n61_));
  NAi31      m0033(.An(mai_mai_n58_), .B(mai_mai_n61_), .C(mai_mai_n56_), .Y(mai_mai_n62_));
  NAi41      m0034(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n63_));
  NA2        m0035(.A(g), .B(f), .Y(mai_mai_n64_));
  NO2        m0036(.A(mai_mai_n64_), .B(mai_mai_n63_), .Y(mai_mai_n65_));
  NAi21      m0037(.An(i), .B(j), .Y(mai_mai_n66_));
  NAi32      m0038(.An(n), .Bn(k), .C(m), .Y(mai_mai_n67_));
  NO2        m0039(.A(mai_mai_n67_), .B(mai_mai_n66_), .Y(mai_mai_n68_));
  NAi31      m0040(.An(l), .B(m), .C(k), .Y(mai_mai_n69_));
  NAi41      m0041(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n68_), .B(mai_mai_n65_), .Y(mai_mai_n71_));
  INV        m0043(.A(m), .Y(mai_mai_n72_));
  NOi21      m0044(.An(k), .B(l), .Y(mai_mai_n73_));
  AN4        m0045(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n74_));
  NOi32      m0046(.An(h), .Bn(g), .C(f), .Y(mai_mai_n75_));
  NA2        m0047(.A(mai_mai_n71_), .B(mai_mai_n62_), .Y(mai_mai_n76_));
  INV        m0048(.A(n), .Y(mai_mai_n77_));
  NOi32      m0049(.An(e), .Bn(b), .C(d), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n77_), .Y(mai_mai_n79_));
  INV        m0051(.A(j), .Y(mai_mai_n80_));
  AN3        m0052(.A(m), .B(k), .C(i), .Y(mai_mai_n81_));
  NA3        m0053(.A(mai_mai_n81_), .B(mai_mai_n80_), .C(g), .Y(mai_mai_n82_));
  NAi32      m0054(.An(g), .Bn(f), .C(h), .Y(mai_mai_n83_));
  NAi31      m0055(.An(j), .B(m), .C(l), .Y(mai_mai_n84_));
  NA2        m0056(.A(m), .B(l), .Y(mai_mai_n85_));
  NAi31      m0057(.An(k), .B(j), .C(g), .Y(mai_mai_n86_));
  NO3        m0058(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(f), .Y(mai_mai_n87_));
  AN2        m0059(.A(j), .B(g), .Y(mai_mai_n88_));
  NOi32      m0060(.An(m), .Bn(l), .C(i), .Y(mai_mai_n89_));
  NOi21      m0061(.An(g), .B(i), .Y(mai_mai_n90_));
  NOi32      m0062(.An(m), .Bn(j), .C(k), .Y(mai_mai_n91_));
  AOI220     m0063(.A0(mai_mai_n91_), .A1(mai_mai_n90_), .B0(mai_mai_n89_), .B1(mai_mai_n88_), .Y(mai_mai_n92_));
  NO2        m0064(.A(mai_mai_n92_), .B(f), .Y(mai_mai_n93_));
  NO2        m0065(.A(mai_mai_n93_), .B(mai_mai_n87_), .Y(mai_mai_n94_));
  NAi41      m0066(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n95_));
  AN2        m0067(.A(e), .B(b), .Y(mai_mai_n96_));
  NOi31      m0068(.An(c), .B(h), .C(f), .Y(mai_mai_n97_));
  NA2        m0069(.A(mai_mai_n97_), .B(mai_mai_n96_), .Y(mai_mai_n98_));
  NOi21      m0070(.An(g), .B(f), .Y(mai_mai_n99_));
  NOi21      m0071(.An(i), .B(h), .Y(mai_mai_n100_));
  NA3        m0072(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(mai_mai_n36_), .Y(mai_mai_n101_));
  INV        m0073(.A(a), .Y(mai_mai_n102_));
  NA2        m0074(.A(mai_mai_n96_), .B(mai_mai_n102_), .Y(mai_mai_n103_));
  INV        m0075(.A(l), .Y(mai_mai_n104_));
  NOi21      m0076(.An(m), .B(n), .Y(mai_mai_n105_));
  AN2        m0077(.A(k), .B(h), .Y(mai_mai_n106_));
  NO2        m0078(.A(mai_mai_n101_), .B(mai_mai_n79_), .Y(mai_mai_n107_));
  INV        m0079(.A(b), .Y(mai_mai_n108_));
  NA2        m0080(.A(l), .B(j), .Y(mai_mai_n109_));
  AN2        m0081(.A(k), .B(i), .Y(mai_mai_n110_));
  NA2        m0082(.A(mai_mai_n110_), .B(mai_mai_n109_), .Y(mai_mai_n111_));
  NA2        m0083(.A(g), .B(e), .Y(mai_mai_n112_));
  NOi32      m0084(.An(c), .Bn(a), .C(d), .Y(mai_mai_n113_));
  NA2        m0085(.A(mai_mai_n113_), .B(mai_mai_n105_), .Y(mai_mai_n114_));
  NO4        m0086(.A(mai_mai_n114_), .B(mai_mai_n112_), .C(mai_mai_n111_), .D(mai_mai_n108_), .Y(mai_mai_n115_));
  NO2        m0087(.A(mai_mai_n115_), .B(mai_mai_n107_), .Y(mai_mai_n116_));
  OAI210     m0088(.A0(mai_mai_n94_), .A1(mai_mai_n79_), .B0(mai_mai_n116_), .Y(mai_mai_n117_));
  NOi31      m0089(.An(k), .B(m), .C(j), .Y(mai_mai_n118_));
  NOi31      m0090(.An(k), .B(m), .C(i), .Y(mai_mai_n119_));
  NA3        m0091(.A(mai_mai_n119_), .B(mai_mai_n75_), .C(mai_mai_n74_), .Y(mai_mai_n120_));
  INV        m0092(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NOi32      m0093(.An(f), .Bn(b), .C(e), .Y(mai_mai_n122_));
  NAi21      m0094(.An(g), .B(h), .Y(mai_mai_n123_));
  NAi21      m0095(.An(m), .B(n), .Y(mai_mai_n124_));
  NAi41      m0096(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n125_));
  NAi31      m0097(.An(j), .B(k), .C(h), .Y(mai_mai_n126_));
  NO3        m0098(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n124_), .Y(mai_mai_n127_));
  INV        m0099(.A(mai_mai_n127_), .Y(mai_mai_n128_));
  NO2        m0100(.A(k), .B(j), .Y(mai_mai_n129_));
  AN2        m0101(.A(k), .B(j), .Y(mai_mai_n130_));
  NAi21      m0102(.An(c), .B(b), .Y(mai_mai_n131_));
  NA2        m0103(.A(f), .B(d), .Y(mai_mai_n132_));
  NA2        m0104(.A(h), .B(c), .Y(mai_mai_n133_));
  NAi31      m0105(.An(f), .B(e), .C(b), .Y(mai_mai_n134_));
  NA2        m0106(.A(d), .B(b), .Y(mai_mai_n135_));
  NAi21      m0107(.An(e), .B(f), .Y(mai_mai_n136_));
  NO2        m0108(.A(mai_mai_n136_), .B(mai_mai_n135_), .Y(mai_mai_n137_));
  NA2        m0109(.A(b), .B(a), .Y(mai_mai_n138_));
  NAi21      m0110(.An(e), .B(g), .Y(mai_mai_n139_));
  NAi21      m0111(.An(c), .B(d), .Y(mai_mai_n140_));
  NAi31      m0112(.An(l), .B(k), .C(h), .Y(mai_mai_n141_));
  NO2        m0113(.A(mai_mai_n124_), .B(mai_mai_n141_), .Y(mai_mai_n142_));
  NA2        m0114(.A(mai_mai_n142_), .B(mai_mai_n137_), .Y(mai_mai_n143_));
  NAi31      m0115(.An(mai_mai_n121_), .B(mai_mai_n143_), .C(mai_mai_n128_), .Y(mai_mai_n144_));
  NAi31      m0116(.An(e), .B(f), .C(b), .Y(mai_mai_n145_));
  INV        m0117(.A(mai_mai_n145_), .Y(mai_mai_n146_));
  NOi21      m0118(.An(h), .B(i), .Y(mai_mai_n147_));
  NOi21      m0119(.An(k), .B(m), .Y(mai_mai_n148_));
  NA3        m0120(.A(mai_mai_n148_), .B(mai_mai_n147_), .C(n), .Y(mai_mai_n149_));
  NOi21      m0121(.An(mai_mai_n146_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  NOi21      m0122(.An(h), .B(g), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n152_));
  NA2        m0124(.A(mai_mai_n152_), .B(mai_mai_n151_), .Y(mai_mai_n153_));
  NAi31      m0125(.An(l), .B(j), .C(h), .Y(mai_mai_n154_));
  NO2        m0126(.A(mai_mai_n154_), .B(mai_mai_n49_), .Y(mai_mai_n155_));
  NA2        m0127(.A(mai_mai_n155_), .B(mai_mai_n65_), .Y(mai_mai_n156_));
  NOi32      m0128(.An(n), .Bn(k), .C(m), .Y(mai_mai_n157_));
  NA2        m0129(.A(l), .B(i), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OAI210     m0131(.A0(mai_mai_n159_), .A1(mai_mai_n153_), .B0(mai_mai_n156_), .Y(mai_mai_n160_));
  NAi31      m0132(.An(d), .B(f), .C(c), .Y(mai_mai_n161_));
  NAi31      m0133(.An(e), .B(f), .C(c), .Y(mai_mai_n162_));
  NA2        m0134(.A(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  NA2        m0135(.A(j), .B(h), .Y(mai_mai_n164_));
  OR3        m0136(.A(n), .B(m), .C(k), .Y(mai_mai_n165_));
  NO2        m0137(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  NAi32      m0138(.An(m), .Bn(k), .C(n), .Y(mai_mai_n167_));
  NO2        m0139(.A(mai_mai_n167_), .B(mai_mai_n164_), .Y(mai_mai_n168_));
  AOI220     m0140(.A0(mai_mai_n168_), .A1(mai_mai_n146_), .B0(mai_mai_n166_), .B1(mai_mai_n163_), .Y(mai_mai_n169_));
  NO2        m0141(.A(n), .B(m), .Y(mai_mai_n170_));
  NAi21      m0142(.An(f), .B(e), .Y(mai_mai_n171_));
  NA2        m0143(.A(d), .B(c), .Y(mai_mai_n172_));
  NAi21      m0144(.An(d), .B(c), .Y(mai_mai_n173_));
  NAi31      m0145(.An(m), .B(n), .C(b), .Y(mai_mai_n174_));
  NA2        m0146(.A(k), .B(i), .Y(mai_mai_n175_));
  NAi21      m0147(.An(h), .B(f), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  NO2        m0149(.A(mai_mai_n174_), .B(mai_mai_n140_), .Y(mai_mai_n178_));
  NA2        m0150(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  NOi32      m0151(.An(f), .Bn(c), .C(d), .Y(mai_mai_n180_));
  NOi32      m0152(.An(f), .Bn(c), .C(e), .Y(mai_mai_n181_));
  NO2        m0153(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NO3        m0154(.A(n), .B(m), .C(j), .Y(mai_mai_n183_));
  NA2        m0155(.A(mai_mai_n183_), .B(mai_mai_n106_), .Y(mai_mai_n184_));
  OR2        m0156(.A(mai_mai_n184_), .B(mai_mai_n182_), .Y(mai_mai_n185_));
  NA3        m0157(.A(mai_mai_n185_), .B(mai_mai_n179_), .C(mai_mai_n169_), .Y(mai_mai_n186_));
  OR4        m0158(.A(mai_mai_n186_), .B(mai_mai_n160_), .C(mai_mai_n150_), .D(mai_mai_n144_), .Y(mai_mai_n187_));
  NO4        m0159(.A(mai_mai_n187_), .B(mai_mai_n117_), .C(mai_mai_n76_), .D(mai_mai_n53_), .Y(mai_mai_n188_));
  NAi31      m0160(.An(n), .B(h), .C(g), .Y(mai_mai_n189_));
  NOi32      m0161(.An(m), .Bn(k), .C(l), .Y(mai_mai_n190_));
  NA3        m0162(.A(mai_mai_n190_), .B(mai_mai_n80_), .C(g), .Y(mai_mai_n191_));
  NO2        m0163(.A(mai_mai_n191_), .B(n), .Y(mai_mai_n192_));
  NA4        m0164(.A(k), .B(mai_mai_n105_), .C(i), .D(g), .Y(mai_mai_n193_));
  AN2        m0165(.A(i), .B(g), .Y(mai_mai_n194_));
  INV        m0166(.A(mai_mai_n193_), .Y(mai_mai_n195_));
  NAi41      m0167(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n196_));
  INV        m0168(.A(mai_mai_n196_), .Y(mai_mai_n197_));
  INV        m0169(.A(f), .Y(mai_mai_n198_));
  INV        m0170(.A(g), .Y(mai_mai_n199_));
  NOi31      m0171(.An(i), .B(j), .C(h), .Y(mai_mai_n200_));
  NOi21      m0172(.An(l), .B(m), .Y(mai_mai_n201_));
  NA2        m0173(.A(mai_mai_n201_), .B(mai_mai_n200_), .Y(mai_mai_n202_));
  NOi21      m0174(.An(n), .B(m), .Y(mai_mai_n203_));
  NOi32      m0175(.An(l), .Bn(i), .C(j), .Y(mai_mai_n204_));
  NA2        m0176(.A(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  OR2        m0177(.A(mai_mai_n205_), .B(mai_mai_n98_), .Y(mai_mai_n206_));
  NAi21      m0178(.An(j), .B(h), .Y(mai_mai_n207_));
  XN2        m0179(.A(i), .B(h), .Y(mai_mai_n208_));
  NA2        m0180(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n209_));
  NOi31      m0181(.An(k), .B(n), .C(m), .Y(mai_mai_n210_));
  NOi31      m0182(.An(mai_mai_n210_), .B(mai_mai_n172_), .C(mai_mai_n171_), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n209_), .Y(mai_mai_n212_));
  NAi31      m0184(.An(f), .B(e), .C(c), .Y(mai_mai_n213_));
  NO4        m0185(.A(mai_mai_n213_), .B(mai_mai_n165_), .C(mai_mai_n164_), .D(mai_mai_n57_), .Y(mai_mai_n214_));
  NA4        m0186(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n215_));
  NAi32      m0187(.An(m), .Bn(i), .C(k), .Y(mai_mai_n216_));
  NO3        m0188(.A(mai_mai_n216_), .B(mai_mai_n83_), .C(mai_mai_n215_), .Y(mai_mai_n217_));
  INV        m0189(.A(k), .Y(mai_mai_n218_));
  NO2        m0190(.A(mai_mai_n217_), .B(mai_mai_n214_), .Y(mai_mai_n219_));
  NAi21      m0191(.An(n), .B(a), .Y(mai_mai_n220_));
  NO2        m0192(.A(mai_mai_n220_), .B(mai_mai_n135_), .Y(mai_mai_n221_));
  NAi41      m0193(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n222_));
  NO2        m0194(.A(mai_mai_n222_), .B(e), .Y(mai_mai_n223_));
  NO3        m0195(.A(mai_mai_n136_), .B(mai_mai_n86_), .C(mai_mai_n85_), .Y(mai_mai_n224_));
  OAI210     m0196(.A0(mai_mai_n224_), .A1(mai_mai_n223_), .B0(mai_mai_n221_), .Y(mai_mai_n225_));
  AN4        m0197(.A(mai_mai_n225_), .B(mai_mai_n219_), .C(mai_mai_n212_), .D(mai_mai_n206_), .Y(mai_mai_n226_));
  NO2        m0198(.A(h), .B(mai_mai_n95_), .Y(mai_mai_n227_));
  NA2        m0199(.A(mai_mai_n227_), .B(mai_mai_n122_), .Y(mai_mai_n228_));
  NAi41      m0200(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n229_), .B(mai_mai_n198_), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n148_), .B(mai_mai_n100_), .Y(mai_mai_n231_));
  NAi21      m0203(.An(mai_mai_n231_), .B(mai_mai_n230_), .Y(mai_mai_n232_));
  NO2        m0204(.A(n), .B(a), .Y(mai_mai_n233_));
  NAi31      m0205(.An(mai_mai_n222_), .B(mai_mai_n233_), .C(mai_mai_n96_), .Y(mai_mai_n234_));
  AN2        m0206(.A(mai_mai_n234_), .B(mai_mai_n232_), .Y(mai_mai_n235_));
  NAi21      m0207(.An(h), .B(i), .Y(mai_mai_n236_));
  NA2        m0208(.A(mai_mai_n170_), .B(k), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  NA2        m0210(.A(mai_mai_n238_), .B(mai_mai_n180_), .Y(mai_mai_n239_));
  NA3        m0211(.A(mai_mai_n239_), .B(mai_mai_n235_), .C(mai_mai_n228_), .Y(mai_mai_n240_));
  NOi21      m0212(.An(g), .B(e), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n242_));
  NA2        m0214(.A(mai_mai_n242_), .B(mai_mai_n241_), .Y(mai_mai_n243_));
  NOi32      m0215(.An(l), .Bn(j), .C(i), .Y(mai_mai_n244_));
  AOI210     m0216(.A0(mai_mai_n73_), .A1(mai_mai_n80_), .B0(mai_mai_n244_), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n236_), .B(mai_mai_n44_), .Y(mai_mai_n246_));
  NAi21      m0218(.An(f), .B(g), .Y(mai_mai_n247_));
  NO2        m0219(.A(mai_mai_n247_), .B(mai_mai_n63_), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n67_), .B(mai_mai_n109_), .Y(mai_mai_n249_));
  AOI220     m0221(.A0(mai_mai_n249_), .A1(mai_mai_n248_), .B0(mai_mai_n246_), .B1(mai_mai_n65_), .Y(mai_mai_n250_));
  OAI210     m0222(.A0(mai_mai_n245_), .A1(mai_mai_n243_), .B0(mai_mai_n250_), .Y(mai_mai_n251_));
  NO2        m0223(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n252_));
  NOi31      m0224(.An(mai_mai_n226_), .B(mai_mai_n251_), .C(mai_mai_n240_), .Y(mai_mai_n253_));
  NO3        m0225(.A(mai_mai_n48_), .B(mai_mai_n43_), .C(mai_mai_n39_), .Y(mai_mai_n254_));
  NO2        m0226(.A(mai_mai_n254_), .B(mai_mai_n103_), .Y(mai_mai_n255_));
  NAi21      m0227(.An(h), .B(g), .Y(mai_mai_n256_));
  OR4        m0228(.A(mai_mai_n256_), .B(mai_mai_n1386_), .C(mai_mai_n205_), .D(e), .Y(mai_mai_n257_));
  NAi31      m0229(.An(g), .B(k), .C(h), .Y(mai_mai_n258_));
  NO3        m0230(.A(mai_mai_n124_), .B(mai_mai_n258_), .C(l), .Y(mai_mai_n259_));
  NAi31      m0231(.An(e), .B(d), .C(a), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n259_), .B(mai_mai_n122_), .Y(mai_mai_n261_));
  NA2        m0233(.A(mai_mai_n261_), .B(mai_mai_n257_), .Y(mai_mai_n262_));
  NA3        m0234(.A(mai_mai_n148_), .B(mai_mai_n147_), .C(mai_mai_n77_), .Y(mai_mai_n263_));
  NO2        m0235(.A(mai_mai_n263_), .B(mai_mai_n182_), .Y(mai_mai_n264_));
  INV        m0236(.A(mai_mai_n264_), .Y(mai_mai_n265_));
  NA3        m0237(.A(e), .B(c), .C(b), .Y(mai_mai_n266_));
  NO2        m0238(.A(mai_mai_n58_), .B(mai_mai_n266_), .Y(mai_mai_n267_));
  NAi32      m0239(.An(k), .Bn(i), .C(j), .Y(mai_mai_n268_));
  NAi31      m0240(.An(h), .B(l), .C(i), .Y(mai_mai_n269_));
  NA3        m0241(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n154_), .Y(mai_mai_n270_));
  NOi21      m0242(.An(mai_mai_n270_), .B(mai_mai_n49_), .Y(mai_mai_n271_));
  OAI210     m0243(.A0(mai_mai_n248_), .A1(mai_mai_n267_), .B0(mai_mai_n271_), .Y(mai_mai_n272_));
  NAi21      m0244(.An(l), .B(k), .Y(mai_mai_n273_));
  NO2        m0245(.A(mai_mai_n273_), .B(mai_mai_n49_), .Y(mai_mai_n274_));
  NOi21      m0246(.An(l), .B(j), .Y(mai_mai_n275_));
  NA2        m0247(.A(mai_mai_n151_), .B(mai_mai_n275_), .Y(mai_mai_n276_));
  NA3        m0248(.A(mai_mai_n110_), .B(mai_mai_n109_), .C(g), .Y(mai_mai_n277_));
  OR3        m0249(.A(mai_mai_n70_), .B(mai_mai_n72_), .C(e), .Y(mai_mai_n278_));
  AOI210     m0250(.A0(mai_mai_n277_), .A1(mai_mai_n276_), .B0(mai_mai_n278_), .Y(mai_mai_n279_));
  INV        m0251(.A(mai_mai_n279_), .Y(mai_mai_n280_));
  NAi32      m0252(.An(j), .Bn(h), .C(i), .Y(mai_mai_n281_));
  NAi21      m0253(.An(m), .B(l), .Y(mai_mai_n282_));
  NO3        m0254(.A(mai_mai_n282_), .B(mai_mai_n281_), .C(mai_mai_n77_), .Y(mai_mai_n283_));
  NA2        m0255(.A(h), .B(g), .Y(mai_mai_n284_));
  NA2        m0256(.A(mai_mai_n157_), .B(mai_mai_n45_), .Y(mai_mai_n285_));
  NO2        m0257(.A(mai_mai_n285_), .B(mai_mai_n284_), .Y(mai_mai_n286_));
  OAI210     m0258(.A0(mai_mai_n286_), .A1(mai_mai_n283_), .B0(mai_mai_n152_), .Y(mai_mai_n287_));
  NA4        m0259(.A(mai_mai_n287_), .B(mai_mai_n280_), .C(mai_mai_n272_), .D(mai_mai_n265_), .Y(mai_mai_n288_));
  NO2        m0260(.A(mai_mai_n134_), .B(d), .Y(mai_mai_n289_));
  NA2        m0261(.A(mai_mai_n289_), .B(mai_mai_n52_), .Y(mai_mai_n290_));
  NAi32      m0262(.An(n), .Bn(m), .C(l), .Y(mai_mai_n291_));
  NO2        m0263(.A(mai_mai_n291_), .B(mai_mai_n281_), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n114_), .B(mai_mai_n108_), .Y(mai_mai_n293_));
  NAi31      m0265(.An(k), .B(l), .C(j), .Y(mai_mai_n294_));
  OAI210     m0266(.A0(mai_mai_n273_), .A1(j), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  NOi21      m0267(.An(mai_mai_n295_), .B(mai_mai_n112_), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n296_), .B(mai_mai_n293_), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n297_), .B(mai_mai_n290_), .Y(mai_mai_n298_));
  NO4        m0270(.A(mai_mai_n298_), .B(mai_mai_n288_), .C(mai_mai_n262_), .D(mai_mai_n255_), .Y(mai_mai_n299_));
  NA2        m0271(.A(mai_mai_n238_), .B(mai_mai_n181_), .Y(mai_mai_n300_));
  NAi21      m0272(.An(m), .B(k), .Y(mai_mai_n301_));
  NO2        m0273(.A(mai_mai_n208_), .B(mai_mai_n301_), .Y(mai_mai_n302_));
  NAi41      m0274(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n303_), .B(mai_mai_n139_), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n304_), .B(mai_mai_n302_), .Y(mai_mai_n305_));
  NAi31      m0277(.An(i), .B(l), .C(h), .Y(mai_mai_n306_));
  NO4        m0278(.A(mai_mai_n306_), .B(mai_mai_n139_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n307_));
  NA2        m0279(.A(e), .B(c), .Y(mai_mai_n308_));
  NO3        m0280(.A(mai_mai_n308_), .B(n), .C(d), .Y(mai_mai_n309_));
  NOi21      m0281(.An(f), .B(h), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n310_), .B(mai_mai_n110_), .Y(mai_mai_n311_));
  NO2        m0283(.A(mai_mai_n311_), .B(mai_mai_n199_), .Y(mai_mai_n312_));
  NAi31      m0284(.An(d), .B(e), .C(b), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n124_), .B(mai_mai_n313_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n314_), .B(mai_mai_n312_), .Y(mai_mai_n315_));
  NAi41      m0287(.An(mai_mai_n307_), .B(mai_mai_n315_), .C(mai_mai_n305_), .D(mai_mai_n300_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n233_), .B(mai_mai_n96_), .Y(mai_mai_n317_));
  OR2        m0289(.A(mai_mai_n317_), .B(mai_mai_n191_), .Y(mai_mai_n318_));
  NOi31      m0290(.An(l), .B(n), .C(m), .Y(mai_mai_n319_));
  INV        m0291(.A(mai_mai_n318_), .Y(mai_mai_n320_));
  NAi32      m0292(.An(m), .Bn(j), .C(k), .Y(mai_mai_n321_));
  NAi41      m0293(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n322_));
  NA2        m0294(.A(mai_mai_n196_), .B(mai_mai_n322_), .Y(mai_mai_n323_));
  NOi31      m0295(.An(j), .B(m), .C(k), .Y(mai_mai_n324_));
  NO2        m0296(.A(mai_mai_n118_), .B(mai_mai_n324_), .Y(mai_mai_n325_));
  AN3        m0297(.A(h), .B(g), .C(f), .Y(mai_mai_n326_));
  NAi31      m0298(.An(mai_mai_n325_), .B(mai_mai_n326_), .C(mai_mai_n323_), .Y(mai_mai_n327_));
  NOi32      m0299(.An(m), .Bn(j), .C(l), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n328_), .B(mai_mai_n89_), .Y(mai_mai_n329_));
  NAi32      m0301(.An(mai_mai_n329_), .Bn(mai_mai_n189_), .C(mai_mai_n289_), .Y(mai_mai_n330_));
  NO2        m0302(.A(mai_mai_n282_), .B(mai_mai_n281_), .Y(mai_mai_n331_));
  NO2        m0303(.A(mai_mai_n202_), .B(g), .Y(mai_mai_n332_));
  INV        m0304(.A(mai_mai_n145_), .Y(mai_mai_n333_));
  INV        m0305(.A(mai_mai_n216_), .Y(mai_mai_n334_));
  NA3        m0306(.A(mai_mai_n334_), .B(mai_mai_n326_), .C(mai_mai_n197_), .Y(mai_mai_n335_));
  NA3        m0307(.A(mai_mai_n335_), .B(mai_mai_n330_), .C(mai_mai_n327_), .Y(mai_mai_n336_));
  NA3        m0308(.A(h), .B(g), .C(f), .Y(mai_mai_n337_));
  NA2        m0309(.A(mai_mai_n151_), .B(e), .Y(mai_mai_n338_));
  NO2        m0310(.A(mai_mai_n338_), .B(mai_mai_n41_), .Y(mai_mai_n339_));
  NA2        m0311(.A(mai_mai_n339_), .B(mai_mai_n293_), .Y(mai_mai_n340_));
  NOi32      m0312(.An(j), .Bn(g), .C(i), .Y(mai_mai_n341_));
  NA3        m0313(.A(mai_mai_n341_), .B(mai_mai_n273_), .C(mai_mai_n105_), .Y(mai_mai_n342_));
  OR2        m0314(.A(mai_mai_n103_), .B(mai_mai_n342_), .Y(mai_mai_n343_));
  NOi32      m0315(.An(e), .Bn(b), .C(a), .Y(mai_mai_n344_));
  AN2        m0316(.A(l), .B(j), .Y(mai_mai_n345_));
  NA2        m0317(.A(mai_mai_n193_), .B(mai_mai_n35_), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n346_), .B(mai_mai_n344_), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n313_), .B(n), .Y(mai_mai_n348_));
  NA2        m0320(.A(mai_mai_n194_), .B(k), .Y(mai_mai_n349_));
  NA3        m0321(.A(m), .B(mai_mai_n104_), .C(mai_mai_n198_), .Y(mai_mai_n350_));
  NA4        m0322(.A(mai_mai_n190_), .B(mai_mai_n80_), .C(g), .D(mai_mai_n198_), .Y(mai_mai_n351_));
  OAI210     m0323(.A0(mai_mai_n350_), .A1(mai_mai_n349_), .B0(mai_mai_n351_), .Y(mai_mai_n352_));
  NAi41      m0324(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n50_), .B(mai_mai_n105_), .Y(mai_mai_n354_));
  NO2        m0326(.A(mai_mai_n354_), .B(mai_mai_n353_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n352_), .B(mai_mai_n348_), .Y(mai_mai_n356_));
  NA4        m0328(.A(mai_mai_n356_), .B(mai_mai_n347_), .C(mai_mai_n343_), .D(mai_mai_n340_), .Y(mai_mai_n357_));
  NO4        m0329(.A(mai_mai_n357_), .B(mai_mai_n336_), .C(mai_mai_n320_), .D(mai_mai_n316_), .Y(mai_mai_n358_));
  NA4        m0330(.A(mai_mai_n358_), .B(mai_mai_n299_), .C(mai_mai_n253_), .D(mai_mai_n188_), .Y(mai10));
  NA3        m0331(.A(m), .B(k), .C(i), .Y(mai_mai_n360_));
  NO3        m0332(.A(mai_mai_n360_), .B(j), .C(mai_mai_n199_), .Y(mai_mai_n361_));
  NOi21      m0333(.An(e), .B(f), .Y(mai_mai_n362_));
  NO4        m0334(.A(mai_mai_n140_), .B(mai_mai_n362_), .C(n), .D(mai_mai_n102_), .Y(mai_mai_n363_));
  NAi31      m0335(.An(b), .B(f), .C(c), .Y(mai_mai_n364_));
  INV        m0336(.A(mai_mai_n364_), .Y(mai_mai_n365_));
  NOi32      m0337(.An(k), .Bn(h), .C(j), .Y(mai_mai_n366_));
  NA2        m0338(.A(mai_mai_n366_), .B(mai_mai_n203_), .Y(mai_mai_n367_));
  OR2        m0339(.A(m), .B(k), .Y(mai_mai_n368_));
  NO2        m0340(.A(mai_mai_n164_), .B(mai_mai_n368_), .Y(mai_mai_n369_));
  NA4        m0341(.A(n), .B(f), .C(c), .D(mai_mai_n108_), .Y(mai_mai_n370_));
  NOi32      m0342(.An(d), .Bn(a), .C(c), .Y(mai_mai_n371_));
  NA2        m0343(.A(mai_mai_n371_), .B(mai_mai_n171_), .Y(mai_mai_n372_));
  NAi21      m0344(.An(i), .B(g), .Y(mai_mai_n373_));
  NAi31      m0345(.An(k), .B(m), .C(j), .Y(mai_mai_n374_));
  NO3        m0346(.A(mai_mai_n374_), .B(mai_mai_n373_), .C(n), .Y(mai_mai_n375_));
  NOi21      m0347(.An(mai_mai_n375_), .B(mai_mai_n372_), .Y(mai_mai_n376_));
  INV        m0348(.A(mai_mai_n376_), .Y(mai_mai_n377_));
  NO2        m0349(.A(mai_mai_n370_), .B(mai_mai_n282_), .Y(mai_mai_n378_));
  NOi32      m0350(.An(f), .Bn(d), .C(c), .Y(mai_mai_n379_));
  AOI220     m0351(.A0(mai_mai_n379_), .A1(mai_mai_n292_), .B0(mai_mai_n378_), .B1(mai_mai_n200_), .Y(mai_mai_n380_));
  NA2        m0352(.A(mai_mai_n380_), .B(mai_mai_n377_), .Y(mai_mai_n381_));
  NO2        m0353(.A(mai_mai_n57_), .B(mai_mai_n108_), .Y(mai_mai_n382_));
  NA2        m0354(.A(mai_mai_n233_), .B(mai_mai_n382_), .Y(mai_mai_n383_));
  INV        m0355(.A(e), .Y(mai_mai_n384_));
  NA2        m0356(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n385_));
  AN2        m0357(.A(g), .B(e), .Y(mai_mai_n386_));
  NA3        m0358(.A(mai_mai_n386_), .B(mai_mai_n190_), .C(i), .Y(mai_mai_n387_));
  INV        m0359(.A(mai_mai_n387_), .Y(mai_mai_n388_));
  NO2        m0360(.A(mai_mai_n92_), .B(mai_mai_n384_), .Y(mai_mai_n389_));
  NO2        m0361(.A(mai_mai_n389_), .B(mai_mai_n388_), .Y(mai_mai_n390_));
  NOi32      m0362(.An(h), .Bn(e), .C(g), .Y(mai_mai_n391_));
  NA3        m0363(.A(mai_mai_n391_), .B(mai_mai_n275_), .C(m), .Y(mai_mai_n392_));
  AN3        m0364(.A(m), .B(l), .C(i), .Y(mai_mai_n393_));
  NA3        m0365(.A(mai_mai_n393_), .B(g), .C(e), .Y(mai_mai_n394_));
  AN3        m0366(.A(h), .B(g), .C(e), .Y(mai_mai_n395_));
  NA2        m0367(.A(mai_mai_n395_), .B(mai_mai_n89_), .Y(mai_mai_n396_));
  AN3        m0368(.A(mai_mai_n396_), .B(mai_mai_n394_), .C(mai_mai_n392_), .Y(mai_mai_n397_));
  AOI210     m0369(.A0(mai_mai_n397_), .A1(mai_mai_n390_), .B0(mai_mai_n383_), .Y(mai_mai_n398_));
  NA3        m0370(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n399_));
  NA3        m0371(.A(mai_mai_n371_), .B(mai_mai_n171_), .C(mai_mai_n77_), .Y(mai_mai_n400_));
  NAi31      m0372(.An(b), .B(c), .C(a), .Y(mai_mai_n401_));
  NO2        m0373(.A(mai_mai_n401_), .B(n), .Y(mai_mai_n402_));
  NA2        m0374(.A(mai_mai_n50_), .B(m), .Y(mai_mai_n403_));
  NO2        m0375(.A(mai_mai_n403_), .B(mai_mai_n136_), .Y(mai_mai_n404_));
  NA2        m0376(.A(mai_mai_n404_), .B(mai_mai_n402_), .Y(mai_mai_n405_));
  INV        m0377(.A(mai_mai_n405_), .Y(mai_mai_n406_));
  NO3        m0378(.A(mai_mai_n406_), .B(mai_mai_n398_), .C(mai_mai_n381_), .Y(mai_mai_n407_));
  NA2        m0379(.A(i), .B(g), .Y(mai_mai_n408_));
  NO3        m0380(.A(mai_mai_n260_), .B(mai_mai_n408_), .C(c), .Y(mai_mai_n409_));
  NOi21      m0381(.An(a), .B(n), .Y(mai_mai_n410_));
  NOi21      m0382(.An(d), .B(c), .Y(mai_mai_n411_));
  NA2        m0383(.A(mai_mai_n411_), .B(mai_mai_n410_), .Y(mai_mai_n412_));
  NA3        m0384(.A(i), .B(g), .C(f), .Y(mai_mai_n413_));
  OR2        m0385(.A(mai_mai_n413_), .B(mai_mai_n69_), .Y(mai_mai_n414_));
  NA3        m0386(.A(mai_mai_n393_), .B(g), .C(mai_mai_n171_), .Y(mai_mai_n415_));
  AOI210     m0387(.A0(mai_mai_n415_), .A1(mai_mai_n414_), .B0(mai_mai_n412_), .Y(mai_mai_n416_));
  AOI210     m0388(.A0(mai_mai_n409_), .A1(mai_mai_n274_), .B0(mai_mai_n416_), .Y(mai_mai_n417_));
  OR2        m0389(.A(n), .B(m), .Y(mai_mai_n418_));
  NO2        m0390(.A(mai_mai_n172_), .B(mai_mai_n136_), .Y(mai_mai_n419_));
  NA2        m0391(.A(mai_mai_n166_), .B(mai_mai_n419_), .Y(mai_mai_n420_));
  INV        m0392(.A(mai_mai_n354_), .Y(mai_mai_n421_));
  NA3        m0393(.A(mai_mai_n421_), .B(mai_mai_n344_), .C(d), .Y(mai_mai_n422_));
  NO2        m0394(.A(mai_mai_n401_), .B(mai_mai_n49_), .Y(mai_mai_n423_));
  NAi21      m0395(.An(k), .B(j), .Y(mai_mai_n424_));
  NAi21      m0396(.An(e), .B(d), .Y(mai_mai_n425_));
  INV        m0397(.A(mai_mai_n425_), .Y(mai_mai_n426_));
  NO2        m0398(.A(mai_mai_n237_), .B(mai_mai_n198_), .Y(mai_mai_n427_));
  NA3        m0399(.A(mai_mai_n427_), .B(mai_mai_n426_), .C(mai_mai_n209_), .Y(mai_mai_n428_));
  NA3        m0400(.A(mai_mai_n428_), .B(mai_mai_n422_), .C(mai_mai_n420_), .Y(mai_mai_n429_));
  NAi31      m0401(.An(g), .B(f), .C(c), .Y(mai_mai_n430_));
  NOi31      m0402(.An(mai_mai_n417_), .B(mai_mai_n429_), .C(mai_mai_n251_), .Y(mai_mai_n431_));
  NOi32      m0403(.An(c), .Bn(a), .C(b), .Y(mai_mai_n432_));
  NA2        m0404(.A(mai_mai_n432_), .B(mai_mai_n105_), .Y(mai_mai_n433_));
  INV        m0405(.A(mai_mai_n258_), .Y(mai_mai_n434_));
  AN2        m0406(.A(e), .B(d), .Y(mai_mai_n435_));
  NA2        m0407(.A(mai_mai_n435_), .B(mai_mai_n434_), .Y(mai_mai_n436_));
  INV        m0408(.A(mai_mai_n136_), .Y(mai_mai_n437_));
  NO2        m0409(.A(mai_mai_n123_), .B(mai_mai_n41_), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n64_), .B(e), .Y(mai_mai_n439_));
  NOi31      m0411(.An(j), .B(k), .C(i), .Y(mai_mai_n440_));
  NOi21      m0412(.An(mai_mai_n154_), .B(mai_mai_n440_), .Y(mai_mai_n441_));
  NA4        m0413(.A(mai_mai_n306_), .B(mai_mai_n441_), .C(mai_mai_n245_), .D(mai_mai_n111_), .Y(mai_mai_n442_));
  AOI220     m0414(.A0(mai_mai_n442_), .A1(mai_mai_n439_), .B0(mai_mai_n438_), .B1(mai_mai_n437_), .Y(mai_mai_n443_));
  AOI210     m0415(.A0(mai_mai_n443_), .A1(mai_mai_n436_), .B0(mai_mai_n433_), .Y(mai_mai_n444_));
  NO2        m0416(.A(mai_mai_n195_), .B(mai_mai_n192_), .Y(mai_mai_n445_));
  NOi21      m0417(.An(a), .B(b), .Y(mai_mai_n446_));
  NA3        m0418(.A(e), .B(d), .C(c), .Y(mai_mai_n447_));
  NAi21      m0419(.An(mai_mai_n447_), .B(mai_mai_n446_), .Y(mai_mai_n448_));
  NO2        m0420(.A(mai_mai_n400_), .B(mai_mai_n191_), .Y(mai_mai_n449_));
  NOi21      m0421(.An(mai_mai_n448_), .B(mai_mai_n449_), .Y(mai_mai_n450_));
  AOI210     m0422(.A0(mai_mai_n254_), .A1(mai_mai_n445_), .B0(mai_mai_n450_), .Y(mai_mai_n451_));
  NO4        m0423(.A(mai_mai_n176_), .B(mai_mai_n95_), .C(mai_mai_n54_), .D(b), .Y(mai_mai_n452_));
  NA2        m0424(.A(mai_mai_n365_), .B(mai_mai_n142_), .Y(mai_mai_n453_));
  OR2        m0425(.A(k), .B(j), .Y(mai_mai_n454_));
  NA2        m0426(.A(l), .B(k), .Y(mai_mai_n455_));
  NA2        m0427(.A(mai_mai_n454_), .B(mai_mai_n203_), .Y(mai_mai_n456_));
  AOI210     m0428(.A0(mai_mai_n216_), .A1(mai_mai_n321_), .B0(mai_mai_n77_), .Y(mai_mai_n457_));
  BUFFER     m0429(.A(mai_mai_n456_), .Y(mai_mai_n458_));
  OR3        m0430(.A(mai_mai_n458_), .B(mai_mai_n133_), .C(mai_mai_n125_), .Y(mai_mai_n459_));
  INV        m0431(.A(mai_mai_n120_), .Y(mai_mai_n460_));
  NA2        m0432(.A(mai_mai_n371_), .B(mai_mai_n105_), .Y(mai_mai_n461_));
  NO4        m0433(.A(mai_mai_n461_), .B(mai_mai_n86_), .C(mai_mai_n104_), .D(e), .Y(mai_mai_n462_));
  NO3        m0434(.A(mai_mai_n400_), .B(mai_mai_n84_), .C(mai_mai_n123_), .Y(mai_mai_n463_));
  NO4        m0435(.A(mai_mai_n463_), .B(mai_mai_n462_), .C(mai_mai_n460_), .D(mai_mai_n307_), .Y(mai_mai_n464_));
  NA3        m0436(.A(mai_mai_n464_), .B(mai_mai_n459_), .C(mai_mai_n453_), .Y(mai_mai_n465_));
  NO3        m0437(.A(mai_mai_n465_), .B(mai_mai_n451_), .C(mai_mai_n444_), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n68_), .B(mai_mai_n65_), .Y(mai_mai_n467_));
  NOi21      m0439(.An(d), .B(e), .Y(mai_mai_n468_));
  NAi31      m0440(.An(j), .B(l), .C(i), .Y(mai_mai_n469_));
  OAI210     m0441(.A0(mai_mai_n469_), .A1(mai_mai_n124_), .B0(mai_mai_n95_), .Y(mai_mai_n470_));
  NO3        m0442(.A(mai_mai_n372_), .B(mai_mai_n329_), .C(mai_mai_n189_), .Y(mai_mai_n471_));
  NO2        m0443(.A(mai_mai_n372_), .B(mai_mai_n354_), .Y(mai_mai_n472_));
  NO2        m0444(.A(mai_mai_n472_), .B(mai_mai_n471_), .Y(mai_mai_n473_));
  NA3        m0445(.A(mai_mai_n473_), .B(mai_mai_n467_), .C(mai_mai_n226_), .Y(mai_mai_n474_));
  OAI210     m0446(.A0(mai_mai_n119_), .A1(mai_mai_n118_), .B0(n), .Y(mai_mai_n475_));
  NO2        m0447(.A(mai_mai_n475_), .B(mai_mai_n123_), .Y(mai_mai_n476_));
  OA210      m0448(.A0(mai_mai_n227_), .A1(mai_mai_n476_), .B0(mai_mai_n181_), .Y(mai_mai_n477_));
  XO2        m0449(.A(i), .B(h), .Y(mai_mai_n478_));
  NAi31      m0450(.An(c), .B(f), .C(d), .Y(mai_mai_n479_));
  AOI210     m0451(.A0(mai_mai_n263_), .A1(mai_mai_n184_), .B0(mai_mai_n479_), .Y(mai_mai_n480_));
  INV        m0452(.A(mai_mai_n480_), .Y(mai_mai_n481_));
  NA3        m0453(.A(mai_mai_n363_), .B(mai_mai_n89_), .C(mai_mai_n88_), .Y(mai_mai_n482_));
  NA2        m0454(.A(mai_mai_n210_), .B(mai_mai_n100_), .Y(mai_mai_n483_));
  NO2        m0455(.A(mai_mai_n483_), .B(mai_mai_n479_), .Y(mai_mai_n484_));
  AOI210     m0456(.A0(mai_mai_n342_), .A1(mai_mai_n35_), .B0(mai_mai_n448_), .Y(mai_mai_n485_));
  NOi31      m0457(.An(mai_mai_n482_), .B(mai_mai_n485_), .C(mai_mai_n484_), .Y(mai_mai_n486_));
  AO220      m0458(.A0(mai_mai_n271_), .A1(mai_mai_n248_), .B0(mai_mai_n155_), .B1(mai_mai_n65_), .Y(mai_mai_n487_));
  NA3        m0459(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n488_));
  NO2        m0460(.A(mai_mai_n488_), .B(mai_mai_n412_), .Y(mai_mai_n489_));
  INV        m0461(.A(mai_mai_n279_), .Y(mai_mai_n490_));
  NAi41      m0462(.An(mai_mai_n487_), .B(mai_mai_n490_), .C(mai_mai_n486_), .D(mai_mai_n481_), .Y(mai_mai_n491_));
  NO3        m0463(.A(mai_mai_n491_), .B(mai_mai_n477_), .C(mai_mai_n474_), .Y(mai_mai_n492_));
  NA4        m0464(.A(mai_mai_n492_), .B(mai_mai_n466_), .C(mai_mai_n431_), .D(mai_mai_n407_), .Y(mai11));
  NO2        m0465(.A(mai_mai_n70_), .B(f), .Y(mai_mai_n494_));
  NA2        m0466(.A(j), .B(g), .Y(mai_mai_n495_));
  NAi31      m0467(.An(i), .B(m), .C(l), .Y(mai_mai_n496_));
  NA3        m0468(.A(m), .B(k), .C(j), .Y(mai_mai_n497_));
  OAI220     m0469(.A0(mai_mai_n497_), .A1(mai_mai_n123_), .B0(mai_mai_n496_), .B1(mai_mai_n495_), .Y(mai_mai_n498_));
  NA2        m0470(.A(mai_mai_n498_), .B(mai_mai_n494_), .Y(mai_mai_n499_));
  NOi32      m0471(.An(e), .Bn(b), .C(f), .Y(mai_mai_n500_));
  NA2        m0472(.A(mai_mai_n244_), .B(mai_mai_n105_), .Y(mai_mai_n501_));
  NA2        m0473(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n502_));
  NO2        m0474(.A(mai_mai_n502_), .B(mai_mai_n285_), .Y(mai_mai_n503_));
  NAi31      m0475(.An(d), .B(e), .C(a), .Y(mai_mai_n504_));
  NO2        m0476(.A(mai_mai_n504_), .B(n), .Y(mai_mai_n505_));
  AOI220     m0477(.A0(mai_mai_n505_), .A1(mai_mai_n93_), .B0(mai_mai_n503_), .B1(mai_mai_n500_), .Y(mai_mai_n506_));
  NAi41      m0478(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n507_));
  AN2        m0479(.A(mai_mai_n507_), .B(mai_mai_n353_), .Y(mai_mai_n508_));
  AOI210     m0480(.A0(mai_mai_n508_), .A1(mai_mai_n372_), .B0(mai_mai_n256_), .Y(mai_mai_n509_));
  NA2        m0481(.A(j), .B(i), .Y(mai_mai_n510_));
  NAi31      m0482(.An(n), .B(m), .C(k), .Y(mai_mai_n511_));
  NO3        m0483(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n104_), .Y(mai_mai_n512_));
  NO4        m0484(.A(n), .B(d), .C(mai_mai_n108_), .D(a), .Y(mai_mai_n513_));
  OR2        m0485(.A(n), .B(c), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n514_), .B(mai_mai_n138_), .Y(mai_mai_n515_));
  NO2        m0487(.A(mai_mai_n515_), .B(mai_mai_n513_), .Y(mai_mai_n516_));
  NOi32      m0488(.An(g), .Bn(f), .C(i), .Y(mai_mai_n517_));
  AOI220     m0489(.A0(mai_mai_n517_), .A1(mai_mai_n91_), .B0(mai_mai_n498_), .B1(f), .Y(mai_mai_n518_));
  NO2        m0490(.A(mai_mai_n518_), .B(mai_mai_n516_), .Y(mai_mai_n519_));
  AOI210     m0491(.A0(mai_mai_n512_), .A1(mai_mai_n509_), .B0(mai_mai_n519_), .Y(mai_mai_n520_));
  NA2        m0492(.A(mai_mai_n130_), .B(mai_mai_n34_), .Y(mai_mai_n521_));
  OAI220     m0493(.A0(mai_mai_n521_), .A1(m), .B0(mai_mai_n502_), .B1(mai_mai_n216_), .Y(mai_mai_n522_));
  NOi41      m0494(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n523_));
  NAi32      m0495(.An(e), .Bn(b), .C(c), .Y(mai_mai_n524_));
  AN2        m0496(.A(mai_mai_n523_), .B(mai_mai_n522_), .Y(mai_mai_n525_));
  OAI220     m0497(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n496_), .B1(mai_mai_n495_), .Y(mai_mai_n526_));
  NAi31      m0498(.An(d), .B(c), .C(a), .Y(mai_mai_n527_));
  NO2        m0499(.A(mai_mai_n527_), .B(n), .Y(mai_mai_n528_));
  NA3        m0500(.A(mai_mai_n528_), .B(mai_mai_n526_), .C(e), .Y(mai_mai_n529_));
  NO3        m0501(.A(mai_mai_n60_), .B(mai_mai_n49_), .C(mai_mai_n199_), .Y(mai_mai_n530_));
  NO2        m0502(.A(mai_mai_n213_), .B(mai_mai_n102_), .Y(mai_mai_n531_));
  OAI210     m0503(.A0(mai_mai_n530_), .A1(mai_mai_n375_), .B0(mai_mai_n531_), .Y(mai_mai_n532_));
  NA2        m0504(.A(mai_mai_n532_), .B(mai_mai_n529_), .Y(mai_mai_n533_));
  NO2        m0505(.A(mai_mai_n260_), .B(n), .Y(mai_mai_n534_));
  NO2        m0506(.A(mai_mai_n402_), .B(mai_mai_n534_), .Y(mai_mai_n535_));
  NA2        m0507(.A(mai_mai_n526_), .B(f), .Y(mai_mai_n536_));
  NAi32      m0508(.An(d), .Bn(a), .C(b), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n537_), .B(mai_mai_n49_), .Y(mai_mai_n538_));
  NA2        m0510(.A(h), .B(f), .Y(mai_mai_n539_));
  NO2        m0511(.A(mai_mai_n539_), .B(mai_mai_n86_), .Y(mai_mai_n540_));
  NA2        m0512(.A(mai_mai_n540_), .B(mai_mai_n538_), .Y(mai_mai_n541_));
  OAI210     m0513(.A0(mai_mai_n536_), .A1(mai_mai_n535_), .B0(mai_mai_n541_), .Y(mai_mai_n542_));
  AN3        m0514(.A(j), .B(h), .C(g), .Y(mai_mai_n543_));
  NO2        m0515(.A(mai_mai_n135_), .B(c), .Y(mai_mai_n544_));
  NA3        m0516(.A(f), .B(d), .C(b), .Y(mai_mai_n545_));
  NO3        m0517(.A(mai_mai_n542_), .B(mai_mai_n533_), .C(mai_mai_n525_), .Y(mai_mai_n546_));
  AN4        m0518(.A(mai_mai_n546_), .B(mai_mai_n520_), .C(mai_mai_n506_), .D(mai_mai_n499_), .Y(mai_mai_n547_));
  INV        m0519(.A(k), .Y(mai_mai_n548_));
  NA3        m0520(.A(l), .B(mai_mai_n548_), .C(i), .Y(mai_mai_n549_));
  INV        m0521(.A(mai_mai_n549_), .Y(mai_mai_n550_));
  NA4        m0522(.A(mai_mai_n371_), .B(g), .C(mai_mai_n171_), .D(mai_mai_n105_), .Y(mai_mai_n551_));
  NAi32      m0523(.An(h), .Bn(f), .C(g), .Y(mai_mai_n552_));
  NAi41      m0524(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n553_));
  OAI210     m0525(.A0(mai_mai_n504_), .A1(n), .B0(mai_mai_n553_), .Y(mai_mai_n554_));
  NA2        m0526(.A(mai_mai_n554_), .B(m), .Y(mai_mai_n555_));
  NAi31      m0527(.An(h), .B(g), .C(f), .Y(mai_mai_n556_));
  OR3        m0528(.A(mai_mai_n556_), .B(mai_mai_n260_), .C(mai_mai_n49_), .Y(mai_mai_n557_));
  NA4        m0529(.A(g), .B(mai_mai_n113_), .C(mai_mai_n105_), .D(e), .Y(mai_mai_n558_));
  AN2        m0530(.A(mai_mai_n558_), .B(mai_mai_n557_), .Y(mai_mai_n559_));
  OA210      m0531(.A0(mai_mai_n555_), .A1(mai_mai_n552_), .B0(mai_mai_n559_), .Y(mai_mai_n560_));
  NO3        m0532(.A(mai_mai_n552_), .B(mai_mai_n70_), .C(mai_mai_n72_), .Y(mai_mai_n561_));
  NO4        m0533(.A(mai_mai_n556_), .B(mai_mai_n514_), .C(mai_mai_n138_), .D(mai_mai_n72_), .Y(mai_mai_n562_));
  OR2        m0534(.A(mai_mai_n562_), .B(mai_mai_n561_), .Y(mai_mai_n563_));
  NAi31      m0535(.An(mai_mai_n563_), .B(mai_mai_n560_), .C(mai_mai_n551_), .Y(mai_mai_n564_));
  NAi31      m0536(.An(f), .B(h), .C(g), .Y(mai_mai_n565_));
  NOi32      m0537(.An(b), .Bn(a), .C(c), .Y(mai_mai_n566_));
  NOi32      m0538(.An(d), .Bn(a), .C(e), .Y(mai_mai_n567_));
  NA2        m0539(.A(mai_mai_n567_), .B(mai_mai_n105_), .Y(mai_mai_n568_));
  NO2        m0540(.A(n), .B(c), .Y(mai_mai_n569_));
  NA3        m0541(.A(mai_mai_n569_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n570_));
  NOi32      m0542(.An(e), .Bn(a), .C(d), .Y(mai_mai_n571_));
  AOI210     m0543(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n571_), .Y(mai_mai_n572_));
  AOI210     m0544(.A0(mai_mai_n572_), .A1(mai_mai_n198_), .B0(mai_mai_n521_), .Y(mai_mai_n573_));
  NA2        m0545(.A(mai_mai_n573_), .B(mai_mai_n105_), .Y(mai_mai_n574_));
  OAI210     m0546(.A0(mai_mai_n232_), .A1(mai_mai_n80_), .B0(mai_mai_n574_), .Y(mai_mai_n575_));
  AOI210     m0547(.A0(mai_mai_n564_), .A1(mai_mai_n550_), .B0(mai_mai_n575_), .Y(mai_mai_n576_));
  NO3        m0548(.A(mai_mai_n301_), .B(mai_mai_n59_), .C(n), .Y(mai_mai_n577_));
  NA3        m0549(.A(mai_mai_n479_), .B(mai_mai_n162_), .C(mai_mai_n161_), .Y(mai_mai_n578_));
  NA2        m0550(.A(mai_mai_n430_), .B(mai_mai_n213_), .Y(mai_mai_n579_));
  OR2        m0551(.A(mai_mai_n579_), .B(mai_mai_n578_), .Y(mai_mai_n580_));
  NA2        m0552(.A(mai_mai_n73_), .B(mai_mai_n105_), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n581_), .B(mai_mai_n45_), .Y(mai_mai_n582_));
  AOI220     m0554(.A0(mai_mai_n582_), .A1(mai_mai_n509_), .B0(mai_mai_n580_), .B1(mai_mai_n577_), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n583_), .B(mai_mai_n80_), .Y(mai_mai_n584_));
  NOi32      m0556(.An(e), .Bn(c), .C(f), .Y(mai_mai_n585_));
  NOi21      m0557(.An(f), .B(g), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n586_), .B(mai_mai_n196_), .Y(mai_mai_n587_));
  AOI220     m0559(.A0(mai_mai_n587_), .A1(mai_mai_n369_), .B0(mai_mai_n585_), .B1(mai_mai_n166_), .Y(mai_mai_n588_));
  NA2        m0560(.A(mai_mai_n588_), .B(mai_mai_n169_), .Y(mai_mai_n589_));
  AOI210     m0561(.A0(mai_mai_n508_), .A1(mai_mai_n372_), .B0(mai_mai_n284_), .Y(mai_mai_n590_));
  NAi21      m0562(.An(k), .B(h), .Y(mai_mai_n591_));
  NO2        m0563(.A(mai_mai_n591_), .B(mai_mai_n247_), .Y(mai_mai_n592_));
  NA2        m0564(.A(mai_mai_n592_), .B(j), .Y(mai_mai_n593_));
  OR2        m0565(.A(mai_mai_n593_), .B(mai_mai_n555_), .Y(mai_mai_n594_));
  NOi31      m0566(.An(m), .B(n), .C(k), .Y(mai_mai_n595_));
  NA2        m0567(.A(j), .B(mai_mai_n595_), .Y(mai_mai_n596_));
  NO2        m0568(.A(mai_mai_n260_), .B(mai_mai_n49_), .Y(mai_mai_n597_));
  NO2        m0569(.A(mai_mai_n504_), .B(mai_mai_n49_), .Y(mai_mai_n598_));
  NA2        m0570(.A(mai_mai_n597_), .B(mai_mai_n540_), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n599_), .B(mai_mai_n594_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n100_), .B(mai_mai_n36_), .Y(mai_mai_n601_));
  NO2        m0573(.A(k), .B(mai_mai_n199_), .Y(mai_mai_n602_));
  NO2        m0574(.A(mai_mai_n500_), .B(mai_mai_n344_), .Y(mai_mai_n603_));
  NO2        m0575(.A(mai_mai_n603_), .B(n), .Y(mai_mai_n604_));
  NAi31      m0576(.An(mai_mai_n601_), .B(mai_mai_n604_), .C(mai_mai_n602_), .Y(mai_mai_n605_));
  AN3        m0577(.A(f), .B(d), .C(b), .Y(mai_mai_n606_));
  NO2        m0578(.A(mai_mai_n606_), .B(mai_mai_n122_), .Y(mai_mai_n607_));
  NA3        m0579(.A(mai_mai_n478_), .B(mai_mai_n148_), .C(mai_mai_n199_), .Y(mai_mai_n608_));
  AOI210     m0580(.A0(mai_mai_n607_), .A1(mai_mai_n215_), .B0(mai_mai_n608_), .Y(mai_mai_n609_));
  NAi31      m0581(.An(m), .B(n), .C(k), .Y(mai_mai_n610_));
  OR2        m0582(.A(mai_mai_n125_), .B(mai_mai_n59_), .Y(mai_mai_n611_));
  OAI210     m0583(.A0(mai_mai_n611_), .A1(mai_mai_n610_), .B0(mai_mai_n234_), .Y(mai_mai_n612_));
  OAI210     m0584(.A0(mai_mai_n612_), .A1(mai_mai_n609_), .B0(j), .Y(mai_mai_n613_));
  NA2        m0585(.A(mai_mai_n613_), .B(mai_mai_n605_), .Y(mai_mai_n614_));
  NO4        m0586(.A(mai_mai_n614_), .B(mai_mai_n600_), .C(mai_mai_n589_), .D(mai_mai_n584_), .Y(mai_mai_n615_));
  NA2        m0587(.A(mai_mai_n363_), .B(mai_mai_n151_), .Y(mai_mai_n616_));
  NAi31      m0588(.An(g), .B(h), .C(f), .Y(mai_mai_n617_));
  OR3        m0589(.A(mai_mai_n617_), .B(mai_mai_n260_), .C(n), .Y(mai_mai_n618_));
  OA210      m0590(.A0(mai_mai_n504_), .A1(n), .B0(mai_mai_n553_), .Y(mai_mai_n619_));
  NA3        m0591(.A(mai_mai_n391_), .B(mai_mai_n113_), .C(mai_mai_n77_), .Y(mai_mai_n620_));
  OAI210     m0592(.A0(mai_mai_n619_), .A1(mai_mai_n83_), .B0(mai_mai_n620_), .Y(mai_mai_n621_));
  NOi21      m0593(.An(mai_mai_n618_), .B(mai_mai_n621_), .Y(mai_mai_n622_));
  AOI210     m0594(.A0(mai_mai_n622_), .A1(mai_mai_n616_), .B0(mai_mai_n497_), .Y(mai_mai_n623_));
  NO3        m0595(.A(g), .B(mai_mai_n198_), .C(mai_mai_n54_), .Y(mai_mai_n624_));
  NO2        m0596(.A(mai_mai_n483_), .B(mai_mai_n80_), .Y(mai_mai_n625_));
  OAI210     m0597(.A0(mai_mai_n625_), .A1(mai_mai_n369_), .B0(mai_mai_n624_), .Y(mai_mai_n626_));
  OR2        m0598(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n627_));
  NA2        m0599(.A(mai_mai_n566_), .B(mai_mai_n326_), .Y(mai_mai_n628_));
  OA220      m0600(.A0(mai_mai_n596_), .A1(mai_mai_n628_), .B0(mai_mai_n593_), .B1(mai_mai_n627_), .Y(mai_mai_n629_));
  NA3        m0601(.A(mai_mai_n494_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n630_));
  AN2        m0602(.A(h), .B(f), .Y(mai_mai_n631_));
  NA2        m0603(.A(mai_mai_n631_), .B(mai_mai_n37_), .Y(mai_mai_n632_));
  NA2        m0604(.A(mai_mai_n91_), .B(mai_mai_n46_), .Y(mai_mai_n633_));
  OAI220     m0605(.A0(mai_mai_n633_), .A1(mai_mai_n317_), .B0(mai_mai_n632_), .B1(mai_mai_n433_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(mai_mai_n537_), .A1(mai_mai_n401_), .B0(mai_mai_n49_), .Y(mai_mai_n635_));
  NO2        m0607(.A(mai_mai_n556_), .B(mai_mai_n549_), .Y(mai_mai_n636_));
  AOI210     m0608(.A0(mai_mai_n636_), .A1(mai_mai_n635_), .B0(mai_mai_n634_), .Y(mai_mai_n637_));
  NA4        m0609(.A(mai_mai_n637_), .B(mai_mai_n630_), .C(mai_mai_n629_), .D(mai_mai_n626_), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n236_), .B(f), .Y(mai_mai_n639_));
  NO2        m0611(.A(mai_mai_n586_), .B(mai_mai_n59_), .Y(mai_mai_n640_));
  NO3        m0612(.A(mai_mai_n640_), .B(mai_mai_n639_), .C(mai_mai_n34_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n314_), .B(mai_mai_n130_), .Y(mai_mai_n642_));
  NA2        m0614(.A(mai_mai_n124_), .B(mai_mai_n49_), .Y(mai_mai_n643_));
  NA2        m0615(.A(mai_mai_n344_), .B(mai_mai_n105_), .Y(mai_mai_n644_));
  OA220      m0616(.A0(mai_mai_n644_), .A1(mai_mai_n521_), .B0(mai_mai_n342_), .B1(mai_mai_n103_), .Y(mai_mai_n645_));
  OAI210     m0617(.A0(mai_mai_n642_), .A1(mai_mai_n641_), .B0(mai_mai_n645_), .Y(mai_mai_n646_));
  NO3        m0618(.A(mai_mai_n379_), .B(mai_mai_n181_), .C(mai_mai_n180_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n647_), .B(mai_mai_n213_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n648_), .B(mai_mai_n238_), .C(j), .Y(mai_mai_n649_));
  NA2        m0621(.A(mai_mai_n432_), .B(mai_mai_n77_), .Y(mai_mai_n650_));
  NA3        m0622(.A(mai_mai_n649_), .B(mai_mai_n482_), .C(mai_mai_n377_), .Y(mai_mai_n651_));
  NO4        m0623(.A(mai_mai_n651_), .B(mai_mai_n646_), .C(mai_mai_n638_), .D(mai_mai_n623_), .Y(mai_mai_n652_));
  NA4        m0624(.A(mai_mai_n652_), .B(mai_mai_n615_), .C(mai_mai_n576_), .D(mai_mai_n547_), .Y(mai08));
  NO2        m0625(.A(k), .B(h), .Y(mai_mai_n654_));
  AO210      m0626(.A0(mai_mai_n236_), .A1(mai_mai_n424_), .B0(mai_mai_n654_), .Y(mai_mai_n655_));
  NO2        m0627(.A(mai_mai_n655_), .B(mai_mai_n282_), .Y(mai_mai_n656_));
  NA2        m0628(.A(mai_mai_n585_), .B(mai_mai_n77_), .Y(mai_mai_n657_));
  NA2        m0629(.A(mai_mai_n657_), .B(mai_mai_n430_), .Y(mai_mai_n658_));
  AOI210     m0630(.A0(mai_mai_n658_), .A1(mai_mai_n656_), .B0(mai_mai_n463_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n77_), .B(mai_mai_n102_), .Y(mai_mai_n660_));
  NO2        m0632(.A(mai_mai_n660_), .B(mai_mai_n55_), .Y(mai_mai_n661_));
  NA2        m0633(.A(mai_mai_n545_), .B(mai_mai_n215_), .Y(mai_mai_n662_));
  NA2        m0634(.A(mai_mai_n662_), .B(mai_mai_n332_), .Y(mai_mai_n663_));
  NA4        m0635(.A(mai_mai_n201_), .B(mai_mai_n130_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n664_));
  AN2        m0636(.A(l), .B(k), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n663_), .B(mai_mai_n659_), .Y(mai_mai_n666_));
  AN2        m0638(.A(mai_mai_n505_), .B(mai_mai_n87_), .Y(mai_mai_n667_));
  NO4        m0639(.A(mai_mai_n164_), .B(mai_mai_n368_), .C(mai_mai_n104_), .D(g), .Y(mai_mai_n668_));
  INV        m0640(.A(mai_mai_n489_), .Y(mai_mai_n669_));
  INV        m0641(.A(mai_mai_n38_), .Y(mai_mai_n670_));
  NA2        m0642(.A(mai_mai_n670_), .B(mai_mai_n534_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n671_), .B(mai_mai_n669_), .Y(mai_mai_n672_));
  NO2        m0644(.A(mai_mai_n508_), .B(mai_mai_n35_), .Y(mai_mai_n673_));
  OAI210     m0645(.A0(mai_mai_n524_), .A1(mai_mai_n47_), .B0(mai_mai_n611_), .Y(mai_mai_n674_));
  NO2        m0646(.A(mai_mai_n455_), .B(mai_mai_n124_), .Y(mai_mai_n675_));
  AOI210     m0647(.A0(mai_mai_n675_), .A1(mai_mai_n674_), .B0(mai_mai_n673_), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n655_), .B(mai_mai_n126_), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n677_), .B(mai_mai_n378_), .Y(mai_mai_n678_));
  NA2        m0650(.A(mai_mai_n676_), .B(mai_mai_n678_), .Y(mai_mai_n679_));
  NA2        m0651(.A(mai_mai_n344_), .B(mai_mai_n43_), .Y(mai_mai_n680_));
  NA3        m0652(.A(mai_mai_n648_), .B(mai_mai_n319_), .C(mai_mai_n366_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n665_), .B(mai_mai_n203_), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n682_), .B(mai_mai_n313_), .Y(mai_mai_n683_));
  AOI210     m0655(.A0(mai_mai_n683_), .A1(mai_mai_n639_), .B0(mai_mai_n462_), .Y(mai_mai_n684_));
  NA3        m0656(.A(m), .B(l), .C(k), .Y(mai_mai_n685_));
  AOI210     m0657(.A0(mai_mai_n620_), .A1(mai_mai_n618_), .B0(mai_mai_n685_), .Y(mai_mai_n686_));
  NO2        m0658(.A(mai_mai_n507_), .B(mai_mai_n256_), .Y(mai_mai_n687_));
  NOi21      m0659(.An(mai_mai_n687_), .B(mai_mai_n501_), .Y(mai_mai_n688_));
  NA4        m0660(.A(mai_mai_n105_), .B(l), .C(k), .D(mai_mai_n80_), .Y(mai_mai_n689_));
  NO2        m0661(.A(mai_mai_n688_), .B(mai_mai_n686_), .Y(mai_mai_n690_));
  NA4        m0662(.A(mai_mai_n690_), .B(mai_mai_n684_), .C(mai_mai_n681_), .D(mai_mai_n680_), .Y(mai_mai_n691_));
  NO4        m0663(.A(mai_mai_n691_), .B(mai_mai_n679_), .C(mai_mai_n672_), .D(mai_mai_n666_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n587_), .B(mai_mai_n369_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n598_), .B(g), .Y(mai_mai_n694_));
  NO2        m0666(.A(mai_mai_n372_), .B(mai_mai_n495_), .Y(mai_mai_n695_));
  AOI210     m0667(.A0(mai_mai_n695_), .A1(mai_mai_n105_), .B0(mai_mai_n472_), .Y(mai_mai_n696_));
  NA4        m0668(.A(mai_mai_n696_), .B(mai_mai_n694_), .C(mai_mai_n693_), .D(mai_mai_n235_), .Y(mai_mai_n697_));
  NA2        m0669(.A(mai_mai_n665_), .B(mai_mai_n72_), .Y(mai_mai_n698_));
  NO3        m0670(.A(mai_mai_n647_), .B(mai_mai_n164_), .C(i), .Y(mai_mai_n699_));
  NOi21      m0671(.An(h), .B(j), .Y(mai_mai_n700_));
  NA2        m0672(.A(mai_mai_n700_), .B(f), .Y(mai_mai_n701_));
  NO2        m0673(.A(mai_mai_n701_), .B(mai_mai_n229_), .Y(mai_mai_n702_));
  NO2        m0674(.A(mai_mai_n702_), .B(mai_mai_n699_), .Y(mai_mai_n703_));
  OAI220     m0675(.A0(mai_mai_n703_), .A1(mai_mai_n698_), .B0(mai_mai_n559_), .B1(mai_mai_n60_), .Y(mai_mai_n704_));
  AOI210     m0676(.A0(mai_mai_n697_), .A1(l), .B0(mai_mai_n704_), .Y(mai_mai_n705_));
  NO2        m0677(.A(j), .B(i), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n75_), .B(l), .Y(mai_mai_n707_));
  NA2        m0679(.A(mai_mai_n706_), .B(mai_mai_n33_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n395_), .B(mai_mai_n113_), .Y(mai_mai_n709_));
  OA220      m0681(.A0(mai_mai_n709_), .A1(mai_mai_n708_), .B0(mai_mai_n707_), .B1(mai_mai_n555_), .Y(mai_mai_n710_));
  NO3        m0682(.A(mai_mai_n140_), .B(mai_mai_n49_), .C(mai_mai_n102_), .Y(mai_mai_n711_));
  NO3        m0683(.A(mai_mai_n514_), .B(mai_mai_n138_), .C(mai_mai_n72_), .Y(mai_mai_n712_));
  NO2        m0684(.A(mai_mai_n455_), .B(mai_mai_n413_), .Y(mai_mai_n713_));
  OAI210     m0685(.A0(mai_mai_n712_), .A1(mai_mai_n711_), .B0(mai_mai_n713_), .Y(mai_mai_n714_));
  OAI210     m0686(.A0(mai_mai_n694_), .A1(mai_mai_n60_), .B0(mai_mai_n714_), .Y(mai_mai_n715_));
  NA2        m0687(.A(k), .B(j), .Y(mai_mai_n716_));
  NO3        m0688(.A(mai_mai_n164_), .B(mai_mai_n368_), .C(mai_mai_n104_), .Y(mai_mai_n717_));
  NA2        m0689(.A(mai_mai_n717_), .B(mai_mai_n230_), .Y(mai_mai_n718_));
  INV        m0690(.A(mai_mai_n718_), .Y(mai_mai_n719_));
  NO2        m0691(.A(mai_mai_n282_), .B(mai_mai_n126_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n720_), .B(mai_mai_n587_), .Y(mai_mai_n721_));
  NO2        m0693(.A(mai_mai_n685_), .B(mai_mai_n83_), .Y(mai_mai_n722_));
  NA2        m0694(.A(mai_mai_n722_), .B(mai_mai_n554_), .Y(mai_mai_n723_));
  NA2        m0695(.A(mai_mai_n713_), .B(mai_mai_n635_), .Y(mai_mai_n724_));
  NA3        m0696(.A(mai_mai_n724_), .B(mai_mai_n723_), .C(mai_mai_n721_), .Y(mai_mai_n725_));
  OR3        m0697(.A(mai_mai_n725_), .B(mai_mai_n719_), .C(mai_mai_n715_), .Y(mai_mai_n726_));
  NO3        m0698(.A(mai_mai_n455_), .B(mai_mai_n408_), .C(f), .Y(mai_mai_n727_));
  OAI220     m0699(.A0(mai_mai_n664_), .A1(mai_mai_n657_), .B0(mai_mai_n317_), .B1(mai_mai_n38_), .Y(mai_mai_n728_));
  AOI210     m0700(.A0(mai_mai_n727_), .A1(mai_mai_n242_), .B0(mai_mai_n728_), .Y(mai_mai_n729_));
  NA3        m0701(.A(mai_mai_n517_), .B(mai_mai_n275_), .C(h), .Y(mai_mai_n730_));
  NOi21      m0702(.An(mai_mai_n635_), .B(mai_mai_n730_), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n84_), .B(mai_mai_n47_), .Y(mai_mai_n732_));
  OAI220     m0704(.A0(mai_mai_n730_), .A1(mai_mai_n570_), .B0(mai_mai_n707_), .B1(mai_mai_n627_), .Y(mai_mai_n733_));
  AOI210     m0705(.A0(mai_mai_n732_), .A1(mai_mai_n604_), .B0(mai_mai_n733_), .Y(mai_mai_n734_));
  NAi31      m0706(.An(mai_mai_n731_), .B(mai_mai_n734_), .C(mai_mai_n729_), .Y(mai_mai_n735_));
  AOI220     m0707(.A0(mai_mai_n722_), .A1(mai_mai_n221_), .B0(mai_mai_n713_), .B1(mai_mai_n597_), .Y(mai_mai_n736_));
  OAI210     m0708(.A0(mai_mai_n685_), .A1(mai_mai_n617_), .B0(mai_mai_n488_), .Y(mai_mai_n737_));
  NA3        m0709(.A(mai_mai_n233_), .B(mai_mai_n57_), .C(b), .Y(mai_mai_n738_));
  AOI220     m0710(.A0(mai_mai_n569_), .A1(mai_mai_n29_), .B0(mai_mai_n432_), .B1(mai_mai_n77_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n739_), .B(mai_mai_n738_), .Y(mai_mai_n740_));
  NO2        m0712(.A(mai_mai_n730_), .B(mai_mai_n461_), .Y(mai_mai_n741_));
  AOI210     m0713(.A0(mai_mai_n740_), .A1(mai_mai_n737_), .B0(mai_mai_n741_), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n742_), .B(mai_mai_n736_), .Y(mai_mai_n743_));
  NOi41      m0715(.An(mai_mai_n710_), .B(mai_mai_n743_), .C(mai_mai_n735_), .D(mai_mai_n726_), .Y(mai_mai_n744_));
  OR3        m0716(.A(mai_mai_n664_), .B(mai_mai_n215_), .C(g), .Y(mai_mai_n745_));
  NO3        m0717(.A(mai_mai_n325_), .B(mai_mai_n284_), .C(mai_mai_n104_), .Y(mai_mai_n746_));
  INV        m0718(.A(mai_mai_n46_), .Y(mai_mai_n747_));
  NO3        m0719(.A(mai_mai_n747_), .B(mai_mai_n708_), .C(mai_mai_n260_), .Y(mai_mai_n748_));
  NO3        m0720(.A(mai_mai_n495_), .B(mai_mai_n85_), .C(h), .Y(mai_mai_n749_));
  AOI210     m0721(.A0(mai_mai_n749_), .A1(mai_mai_n661_), .B0(mai_mai_n748_), .Y(mai_mai_n750_));
  NA3        m0722(.A(mai_mai_n750_), .B(mai_mai_n745_), .C(mai_mai_n380_), .Y(mai_mai_n751_));
  OR2        m0723(.A(mai_mai_n617_), .B(mai_mai_n84_), .Y(mai_mai_n752_));
  NOi31      m0724(.An(b), .B(d), .C(a), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n753_), .B(mai_mai_n567_), .Y(mai_mai_n754_));
  NO2        m0726(.A(mai_mai_n754_), .B(n), .Y(mai_mai_n755_));
  NOi21      m0727(.An(mai_mai_n739_), .B(mai_mai_n755_), .Y(mai_mai_n756_));
  NO2        m0728(.A(mai_mai_n756_), .B(mai_mai_n752_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n524_), .B(mai_mai_n77_), .Y(mai_mai_n758_));
  NO3        m0730(.A(mai_mai_n586_), .B(mai_mai_n313_), .C(mai_mai_n109_), .Y(mai_mai_n759_));
  NOi21      m0731(.An(mai_mai_n759_), .B(mai_mai_n149_), .Y(mai_mai_n760_));
  AOI210     m0732(.A0(mai_mai_n746_), .A1(mai_mai_n758_), .B0(mai_mai_n760_), .Y(mai_mai_n761_));
  OAI210     m0733(.A0(mai_mai_n664_), .A1(mai_mai_n370_), .B0(mai_mai_n761_), .Y(mai_mai_n762_));
  NO2        m0734(.A(mai_mai_n647_), .B(n), .Y(mai_mai_n763_));
  AOI220     m0735(.A0(mai_mai_n720_), .A1(mai_mai_n624_), .B0(mai_mai_n763_), .B1(mai_mai_n656_), .Y(mai_mai_n764_));
  NO2        m0736(.A(mai_mai_n308_), .B(mai_mai_n220_), .Y(mai_mai_n765_));
  NA2        m0737(.A(mai_mai_n87_), .B(mai_mai_n765_), .Y(mai_mai_n766_));
  NA2        m0738(.A(mai_mai_n113_), .B(mai_mai_n77_), .Y(mai_mai_n767_));
  AOI210     m0739(.A0(mai_mai_n399_), .A1(mai_mai_n392_), .B0(mai_mai_n767_), .Y(mai_mai_n768_));
  NAi21      m0740(.An(mai_mai_n768_), .B(mai_mai_n766_), .Y(mai_mai_n769_));
  NA2        m0741(.A(mai_mai_n683_), .B(mai_mai_n34_), .Y(mai_mai_n770_));
  NAi21      m0742(.An(mai_mai_n689_), .B(mai_mai_n409_), .Y(mai_mai_n771_));
  NO2        m0743(.A(mai_mai_n256_), .B(i), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n668_), .B(mai_mai_n333_), .Y(mai_mai_n773_));
  OAI210     m0745(.A0(mai_mai_n562_), .A1(mai_mai_n561_), .B0(mai_mai_n345_), .Y(mai_mai_n774_));
  AN3        m0746(.A(mai_mai_n774_), .B(mai_mai_n773_), .C(mai_mai_n771_), .Y(mai_mai_n775_));
  NAi41      m0747(.An(mai_mai_n769_), .B(mai_mai_n775_), .C(mai_mai_n770_), .D(mai_mai_n764_), .Y(mai_mai_n776_));
  NO4        m0748(.A(mai_mai_n776_), .B(mai_mai_n762_), .C(mai_mai_n757_), .D(mai_mai_n751_), .Y(mai_mai_n777_));
  NA4        m0749(.A(mai_mai_n777_), .B(mai_mai_n744_), .C(mai_mai_n705_), .D(mai_mai_n692_), .Y(mai09));
  INV        m0750(.A(mai_mai_n114_), .Y(mai_mai_n779_));
  NA2        m0751(.A(f), .B(e), .Y(mai_mai_n780_));
  NO2        m0752(.A(mai_mai_n208_), .B(mai_mai_n104_), .Y(mai_mai_n781_));
  NA2        m0753(.A(mai_mai_n781_), .B(g), .Y(mai_mai_n782_));
  NA4        m0754(.A(mai_mai_n294_), .B(mai_mai_n441_), .C(mai_mai_n245_), .D(mai_mai_n111_), .Y(mai_mai_n783_));
  AOI210     m0755(.A0(mai_mai_n783_), .A1(g), .B0(mai_mai_n438_), .Y(mai_mai_n784_));
  AOI210     m0756(.A0(mai_mai_n784_), .A1(mai_mai_n782_), .B0(mai_mai_n780_), .Y(mai_mai_n785_));
  NA2        m0757(.A(mai_mai_n785_), .B(mai_mai_n779_), .Y(mai_mai_n786_));
  NO2        m0758(.A(mai_mai_n191_), .B(mai_mai_n198_), .Y(mai_mai_n787_));
  NA3        m0759(.A(m), .B(l), .C(i), .Y(mai_mai_n788_));
  OAI220     m0760(.A0(mai_mai_n556_), .A1(mai_mai_n788_), .B0(mai_mai_n337_), .B1(mai_mai_n496_), .Y(mai_mai_n789_));
  NA4        m0761(.A(mai_mai_n81_), .B(mai_mai_n80_), .C(g), .D(f), .Y(mai_mai_n790_));
  NAi31      m0762(.An(mai_mai_n789_), .B(mai_mai_n790_), .C(mai_mai_n414_), .Y(mai_mai_n791_));
  OR2        m0763(.A(mai_mai_n791_), .B(mai_mai_n787_), .Y(mai_mai_n792_));
  NA3        m0764(.A(mai_mai_n752_), .B(mai_mai_n536_), .C(mai_mai_n488_), .Y(mai_mai_n793_));
  OA210      m0765(.A0(mai_mai_n793_), .A1(mai_mai_n792_), .B0(mai_mai_n755_), .Y(mai_mai_n794_));
  INV        m0766(.A(mai_mai_n322_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n796_));
  NA2        m0768(.A(mai_mai_n738_), .B(mai_mai_n317_), .Y(mai_mai_n797_));
  NA2        m0769(.A(mai_mai_n326_), .B(mai_mai_n328_), .Y(mai_mai_n798_));
  OAI210     m0770(.A0(mai_mai_n191_), .A1(mai_mai_n198_), .B0(mai_mai_n798_), .Y(mai_mai_n799_));
  NA2        m0771(.A(mai_mai_n799_), .B(mai_mai_n797_), .Y(mai_mai_n800_));
  NA2        m0772(.A(mai_mai_n158_), .B(mai_mai_n106_), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n801_), .B(mai_mai_n655_), .Y(mai_mai_n802_));
  NA3        m0774(.A(mai_mai_n802_), .B(mai_mai_n178_), .C(mai_mai_n31_), .Y(mai_mai_n803_));
  NA3        m0775(.A(mai_mai_n803_), .B(mai_mai_n800_), .C(mai_mai_n588_), .Y(mai_mai_n804_));
  NO2        m0776(.A(mai_mai_n552_), .B(mai_mai_n469_), .Y(mai_mai_n805_));
  NA2        m0777(.A(mai_mai_n805_), .B(mai_mai_n178_), .Y(mai_mai_n806_));
  NOi21      m0778(.An(f), .B(d), .Y(mai_mai_n807_));
  NA2        m0779(.A(mai_mai_n807_), .B(m), .Y(mai_mai_n808_));
  NO2        m0780(.A(mai_mai_n808_), .B(mai_mai_n51_), .Y(mai_mai_n809_));
  NOi32      m0781(.An(g), .Bn(f), .C(d), .Y(mai_mai_n810_));
  NA4        m0782(.A(mai_mai_n810_), .B(mai_mai_n569_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n811_));
  NOi21      m0783(.An(mai_mai_n295_), .B(mai_mai_n811_), .Y(mai_mai_n812_));
  AOI210     m0784(.A0(mai_mai_n809_), .A1(mai_mai_n515_), .B0(mai_mai_n812_), .Y(mai_mai_n813_));
  NA2        m0785(.A(mai_mai_n245_), .B(mai_mai_n111_), .Y(mai_mai_n814_));
  AN2        m0786(.A(f), .B(d), .Y(mai_mai_n815_));
  NA3        m0787(.A(mai_mai_n446_), .B(mai_mai_n815_), .C(mai_mai_n77_), .Y(mai_mai_n816_));
  NO3        m0788(.A(mai_mai_n816_), .B(mai_mai_n72_), .C(mai_mai_n199_), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n268_), .B(mai_mai_n54_), .Y(mai_mai_n818_));
  NA2        m0790(.A(mai_mai_n814_), .B(mai_mai_n817_), .Y(mai_mai_n819_));
  NAi41      m0791(.An(mai_mai_n460_), .B(mai_mai_n819_), .C(mai_mai_n813_), .D(mai_mai_n806_), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n610_), .B(mai_mai_n313_), .Y(mai_mai_n821_));
  AN2        m0793(.A(mai_mai_n821_), .B(mai_mai_n639_), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n822_), .B(mai_mai_n217_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n567_), .B(mai_mai_n77_), .Y(mai_mai_n824_));
  NO2        m0796(.A(mai_mai_n798_), .B(mai_mai_n824_), .Y(mai_mai_n825_));
  NA3        m0797(.A(mai_mai_n148_), .B(mai_mai_n100_), .C(mai_mai_n99_), .Y(mai_mai_n826_));
  OAI220     m0798(.A0(mai_mai_n816_), .A1(mai_mai_n403_), .B0(mai_mai_n322_), .B1(mai_mai_n826_), .Y(mai_mai_n827_));
  NOi31      m0799(.An(mai_mai_n206_), .B(mai_mai_n827_), .C(mai_mai_n825_), .Y(mai_mai_n828_));
  NA2        m0800(.A(c), .B(mai_mai_n108_), .Y(mai_mai_n829_));
  NO2        m0801(.A(mai_mai_n829_), .B(mai_mai_n384_), .Y(mai_mai_n830_));
  NA2        m0802(.A(mai_mai_n830_), .B(mai_mai_n283_), .Y(mai_mai_n831_));
  OR2        m0803(.A(mai_mai_n617_), .B(mai_mai_n511_), .Y(mai_mai_n832_));
  INV        m0804(.A(mai_mai_n832_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n754_), .B(mai_mai_n103_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n834_), .B(mai_mai_n833_), .Y(mai_mai_n835_));
  NA4        m0807(.A(mai_mai_n835_), .B(mai_mai_n831_), .C(mai_mai_n828_), .D(mai_mai_n823_), .Y(mai_mai_n836_));
  NO4        m0808(.A(mai_mai_n836_), .B(mai_mai_n820_), .C(mai_mai_n804_), .D(mai_mai_n794_), .Y(mai_mai_n837_));
  OR2        m0809(.A(mai_mai_n816_), .B(mai_mai_n72_), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n781_), .B(g), .Y(mai_mai_n839_));
  AOI210     m0811(.A0(mai_mai_n839_), .A1(mai_mai_n276_), .B0(mai_mai_n838_), .Y(mai_mai_n840_));
  NO2        m0812(.A(mai_mai_n317_), .B(mai_mai_n790_), .Y(mai_mai_n841_));
  NO2        m0813(.A(mai_mai_n403_), .B(mai_mai_n780_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n842_), .B(mai_mai_n528_), .Y(mai_mai_n843_));
  INV        m0815(.A(mai_mai_n843_), .Y(mai_mai_n844_));
  NA2        m0816(.A(e), .B(d), .Y(mai_mai_n845_));
  OAI220     m0817(.A0(mai_mai_n845_), .A1(c), .B0(mai_mai_n308_), .B1(d), .Y(mai_mai_n846_));
  NA3        m0818(.A(mai_mai_n846_), .B(mai_mai_n427_), .C(mai_mai_n478_), .Y(mai_mai_n847_));
  NO2        m0819(.A(mai_mai_n483_), .B(mai_mai_n213_), .Y(mai_mai_n848_));
  INV        m0820(.A(mai_mai_n848_), .Y(mai_mai_n849_));
  NA2        m0821(.A(mai_mai_n268_), .B(mai_mai_n154_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n817_), .B(mai_mai_n850_), .Y(mai_mai_n851_));
  NA3        m0823(.A(mai_mai_n157_), .B(mai_mai_n78_), .C(mai_mai_n34_), .Y(mai_mai_n852_));
  NA4        m0824(.A(mai_mai_n852_), .B(mai_mai_n851_), .C(mai_mai_n849_), .D(mai_mai_n847_), .Y(mai_mai_n853_));
  NO4        m0825(.A(mai_mai_n853_), .B(mai_mai_n844_), .C(mai_mai_n841_), .D(mai_mai_n840_), .Y(mai_mai_n854_));
  NA2        m0826(.A(mai_mai_n795_), .B(mai_mai_n31_), .Y(mai_mai_n855_));
  OR2        m0827(.A(mai_mai_n855_), .B(mai_mai_n202_), .Y(mai_mai_n856_));
  OAI220     m0828(.A0(mai_mai_n586_), .A1(mai_mai_n59_), .B0(mai_mai_n284_), .B1(j), .Y(mai_mai_n857_));
  AOI220     m0829(.A0(mai_mai_n857_), .A1(mai_mai_n821_), .B0(mai_mai_n577_), .B1(mai_mai_n585_), .Y(mai_mai_n858_));
  INV        m0830(.A(mai_mai_n858_), .Y(mai_mai_n859_));
  OAI210     m0831(.A0(mai_mai_n781_), .A1(mai_mai_n850_), .B0(mai_mai_n810_), .Y(mai_mai_n860_));
  NO2        m0832(.A(mai_mai_n860_), .B(mai_mai_n570_), .Y(mai_mai_n861_));
  AOI210     m0833(.A0(mai_mai_n110_), .A1(mai_mai_n109_), .B0(mai_mai_n244_), .Y(mai_mai_n862_));
  NO2        m0834(.A(mai_mai_n862_), .B(mai_mai_n811_), .Y(mai_mai_n863_));
  AO210      m0835(.A0(mai_mai_n797_), .A1(mai_mai_n789_), .B0(mai_mai_n863_), .Y(mai_mai_n864_));
  NOi31      m0836(.An(mai_mai_n515_), .B(mai_mai_n808_), .C(mai_mai_n276_), .Y(mai_mai_n865_));
  NO4        m0837(.A(mai_mai_n865_), .B(mai_mai_n864_), .C(mai_mai_n861_), .D(mai_mai_n859_), .Y(mai_mai_n866_));
  AO220      m0838(.A0(mai_mai_n427_), .A1(mai_mai_n700_), .B0(mai_mai_n166_), .B1(f), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n867_), .B(mai_mai_n846_), .Y(mai_mai_n868_));
  NO2        m0840(.A(mai_mai_n413_), .B(mai_mai_n69_), .Y(mai_mai_n869_));
  OAI210     m0841(.A0(mai_mai_n793_), .A1(mai_mai_n869_), .B0(mai_mai_n661_), .Y(mai_mai_n870_));
  AN4        m0842(.A(mai_mai_n870_), .B(mai_mai_n868_), .C(mai_mai_n866_), .D(mai_mai_n856_), .Y(mai_mai_n871_));
  NA4        m0843(.A(mai_mai_n871_), .B(mai_mai_n854_), .C(mai_mai_n837_), .D(mai_mai_n786_), .Y(mai12));
  NO2        m0844(.A(mai_mai_n425_), .B(c), .Y(mai_mai_n873_));
  NO4        m0845(.A(mai_mai_n418_), .B(mai_mai_n236_), .C(mai_mai_n548_), .D(mai_mai_n199_), .Y(mai_mai_n874_));
  NA2        m0846(.A(mai_mai_n874_), .B(mai_mai_n873_), .Y(mai_mai_n875_));
  NA2        m0847(.A(mai_mai_n515_), .B(mai_mai_n869_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n425_), .B(mai_mai_n108_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n796_), .B(mai_mai_n337_), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n617_), .B(mai_mai_n360_), .Y(mai_mai_n879_));
  AOI220     m0851(.A0(mai_mai_n879_), .A1(mai_mai_n513_), .B0(mai_mai_n878_), .B1(mai_mai_n877_), .Y(mai_mai_n880_));
  NA4        m0852(.A(mai_mai_n880_), .B(mai_mai_n876_), .C(mai_mai_n875_), .D(mai_mai_n417_), .Y(mai_mai_n881_));
  AOI210     m0853(.A0(mai_mai_n216_), .A1(mai_mai_n321_), .B0(mai_mai_n189_), .Y(mai_mai_n882_));
  OR2        m0854(.A(mai_mai_n882_), .B(mai_mai_n874_), .Y(mai_mai_n883_));
  NA2        m0855(.A(mai_mai_n883_), .B(mai_mai_n379_), .Y(mai_mai_n884_));
  NO2        m0856(.A(mai_mai_n601_), .B(mai_mai_n247_), .Y(mai_mai_n885_));
  NO2        m0857(.A(mai_mai_n556_), .B(mai_mai_n788_), .Y(mai_mai_n886_));
  AOI220     m0858(.A0(mai_mai_n886_), .A1(mai_mai_n534_), .B0(mai_mai_n765_), .B1(mai_mai_n885_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n140_), .B(mai_mai_n220_), .Y(mai_mai_n888_));
  NA3        m0860(.A(mai_mai_n888_), .B(mai_mai_n223_), .C(i), .Y(mai_mai_n889_));
  NA3        m0861(.A(mai_mai_n889_), .B(mai_mai_n887_), .C(mai_mai_n884_), .Y(mai_mai_n890_));
  NO3        m0862(.A(mai_mai_n622_), .B(mai_mai_n84_), .C(mai_mai_n45_), .Y(mai_mai_n891_));
  NO3        m0863(.A(mai_mai_n891_), .B(mai_mai_n890_), .C(mai_mai_n881_), .Y(mai_mai_n892_));
  NO2        m0864(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n553_), .B(mai_mai_n70_), .Y(mai_mai_n894_));
  NOi21      m0866(.An(mai_mai_n34_), .B(mai_mai_n610_), .Y(mai_mai_n895_));
  NA2        m0867(.A(mai_mai_n894_), .B(mai_mai_n893_), .Y(mai_mai_n896_));
  OAI210     m0868(.A0(mai_mai_n234_), .A1(mai_mai_n45_), .B0(mai_mai_n896_), .Y(mai_mai_n897_));
  NA2        m0869(.A(mai_mai_n409_), .B(mai_mai_n249_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n898_), .B(mai_mai_n305_), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n475_), .B(mai_mai_n284_), .Y(mai_mai_n900_));
  INV        m0872(.A(mai_mai_n900_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n901_), .B(mai_mai_n134_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n595_), .B(mai_mai_n345_), .Y(mai_mai_n903_));
  INV        m0875(.A(mai_mai_n347_), .Y(mai_mai_n904_));
  NO4        m0876(.A(mai_mai_n904_), .B(mai_mai_n902_), .C(mai_mai_n899_), .D(mai_mai_n897_), .Y(mai_mai_n905_));
  NA2        m0877(.A(mai_mai_n331_), .B(g), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n151_), .B(i), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n907_), .B(mai_mai_n84_), .Y(mai_mai_n908_));
  AOI210     m0880(.A0(mai_mai_n393_), .A1(mai_mai_n37_), .B0(mai_mai_n908_), .Y(mai_mai_n909_));
  NA2        m0881(.A(mai_mai_n524_), .B(mai_mai_n364_), .Y(mai_mai_n910_));
  AOI210     m0882(.A0(mai_mai_n910_), .A1(n), .B0(mai_mai_n523_), .Y(mai_mai_n911_));
  OAI220     m0883(.A0(mai_mai_n911_), .A1(mai_mai_n906_), .B0(mai_mai_n909_), .B1(mai_mai_n317_), .Y(mai_mai_n912_));
  NO2        m0884(.A(mai_mai_n617_), .B(mai_mai_n469_), .Y(mai_mai_n913_));
  NA3        m0885(.A(mai_mai_n326_), .B(j), .C(i), .Y(mai_mai_n914_));
  INV        m0886(.A(mai_mai_n914_), .Y(mai_mai_n915_));
  OAI220     m0887(.A0(mai_mai_n915_), .A1(mai_mai_n913_), .B0(mai_mai_n635_), .B1(mai_mai_n712_), .Y(mai_mai_n916_));
  NA2        m0888(.A(mai_mai_n571_), .B(mai_mai_n105_), .Y(mai_mai_n917_));
  OR3        m0889(.A(mai_mai_n294_), .B(mai_mai_n408_), .C(f), .Y(mai_mai_n918_));
  NA3        m0890(.A(j), .B(mai_mai_n75_), .C(i), .Y(mai_mai_n919_));
  OA220      m0891(.A0(mai_mai_n919_), .A1(mai_mai_n917_), .B0(mai_mai_n918_), .B1(mai_mai_n555_), .Y(mai_mai_n920_));
  NA3        m0892(.A(mai_mai_n310_), .B(mai_mai_n110_), .C(g), .Y(mai_mai_n921_));
  AOI210     m0893(.A0(mai_mai_n632_), .A1(mai_mai_n921_), .B0(m), .Y(mai_mai_n922_));
  OAI210     m0894(.A0(mai_mai_n922_), .A1(mai_mai_n878_), .B0(mai_mai_n309_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n650_), .B(mai_mai_n824_), .Y(mai_mai_n924_));
  NA2        m0896(.A(mai_mai_n790_), .B(mai_mai_n414_), .Y(mai_mai_n925_));
  NA2        m0897(.A(mai_mai_n204_), .B(h), .Y(mai_mai_n926_));
  NA3        m0898(.A(mai_mai_n926_), .B(mai_mai_n919_), .C(mai_mai_n918_), .Y(mai_mai_n927_));
  AOI220     m0899(.A0(mai_mai_n927_), .A1(mai_mai_n242_), .B0(mai_mai_n925_), .B1(mai_mai_n924_), .Y(mai_mai_n928_));
  NA4        m0900(.A(mai_mai_n928_), .B(mai_mai_n923_), .C(mai_mai_n920_), .D(mai_mai_n916_), .Y(mai_mai_n929_));
  NO2        m0901(.A(mai_mai_n360_), .B(mai_mai_n83_), .Y(mai_mai_n930_));
  OAI210     m0902(.A0(mai_mai_n930_), .A1(mai_mai_n885_), .B0(mai_mai_n221_), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n621_), .B(mai_mai_n81_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n932_), .B(mai_mai_n931_), .Y(mai_mai_n933_));
  OAI210     m0905(.A0(mai_mai_n925_), .A1(mai_mai_n886_), .B0(mai_mai_n513_), .Y(mai_mai_n934_));
  AOI210     m0906(.A0(mai_mai_n394_), .A1(mai_mai_n387_), .B0(mai_mai_n767_), .Y(mai_mai_n935_));
  OAI210     m0907(.A0(mai_mai_n350_), .A1(mai_mai_n349_), .B0(mai_mai_n101_), .Y(mai_mai_n936_));
  AOI210     m0908(.A0(mai_mai_n936_), .A1(mai_mai_n505_), .B0(mai_mai_n935_), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n922_), .B(mai_mai_n877_), .Y(mai_mai_n938_));
  NO3        m0910(.A(l), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n939_));
  NA2        m0911(.A(mai_mai_n939_), .B(mai_mai_n590_), .Y(mai_mai_n940_));
  NA4        m0912(.A(mai_mai_n940_), .B(mai_mai_n938_), .C(mai_mai_n937_), .D(mai_mai_n934_), .Y(mai_mai_n941_));
  NO4        m0913(.A(mai_mai_n941_), .B(mai_mai_n933_), .C(mai_mai_n929_), .D(mai_mai_n912_), .Y(mai_mai_n942_));
  NAi31      m0914(.An(mai_mai_n131_), .B(mai_mai_n395_), .C(n), .Y(mai_mai_n943_));
  NO3        m0915(.A(mai_mai_n256_), .B(mai_mai_n131_), .C(mai_mai_n384_), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n944_), .B(mai_mai_n470_), .Y(mai_mai_n945_));
  NA2        m0917(.A(mai_mai_n463_), .B(i), .Y(mai_mai_n946_));
  NA2        m0918(.A(mai_mai_n946_), .B(mai_mai_n945_), .Y(mai_mai_n947_));
  NA2        m0919(.A(mai_mai_n213_), .B(mai_mai_n162_), .Y(mai_mai_n948_));
  INV        m0920(.A(mai_mai_n166_), .Y(mai_mai_n949_));
  NOi31      m0921(.An(mai_mai_n948_), .B(mai_mai_n949_), .C(mai_mai_n199_), .Y(mai_mai_n950_));
  INV        m0922(.A(mai_mai_n1385_), .Y(mai_mai_n951_));
  OAI220     m0923(.A0(mai_mai_n943_), .A1(mai_mai_n216_), .B0(mai_mai_n914_), .B1(mai_mai_n568_), .Y(mai_mai_n952_));
  NO2        m0924(.A(mai_mai_n618_), .B(mai_mai_n360_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n882_), .B(mai_mai_n873_), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n514_), .B(mai_mai_n138_), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n955_), .B(mai_mai_n361_), .Y(mai_mai_n956_));
  OAI220     m0928(.A0(mai_mai_n879_), .A1(mai_mai_n886_), .B0(mai_mai_n515_), .B1(mai_mai_n402_), .Y(mai_mai_n957_));
  NA3        m0929(.A(mai_mai_n957_), .B(mai_mai_n956_), .C(mai_mai_n954_), .Y(mai_mai_n958_));
  OAI210     m0930(.A0(mai_mai_n882_), .A1(mai_mai_n874_), .B0(mai_mai_n948_), .Y(mai_mai_n959_));
  NA3        m0931(.A(mai_mai_n910_), .B(mai_mai_n457_), .C(mai_mai_n46_), .Y(mai_mai_n960_));
  NA3        m0932(.A(mai_mai_n960_), .B(mai_mai_n959_), .C(mai_mai_n257_), .Y(mai_mai_n961_));
  OR4        m0933(.A(mai_mai_n961_), .B(mai_mai_n958_), .C(mai_mai_n953_), .D(mai_mai_n952_), .Y(mai_mai_n962_));
  NO4        m0934(.A(mai_mai_n962_), .B(mai_mai_n951_), .C(mai_mai_n950_), .D(mai_mai_n947_), .Y(mai_mai_n963_));
  NA4        m0935(.A(mai_mai_n963_), .B(mai_mai_n942_), .C(mai_mai_n905_), .D(mai_mai_n892_), .Y(mai13));
  AN2        m0936(.A(c), .B(b), .Y(mai_mai_n965_));
  NA3        m0937(.A(mai_mai_n233_), .B(mai_mai_n965_), .C(m), .Y(mai_mai_n966_));
  NA2        m0938(.A(mai_mai_n468_), .B(f), .Y(mai_mai_n967_));
  NO3        m0939(.A(mai_mai_n967_), .B(mai_mai_n966_), .C(mai_mai_n549_), .Y(mai_mai_n968_));
  NAi32      m0940(.An(d), .Bn(c), .C(e), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n130_), .B(mai_mai_n45_), .Y(mai_mai_n970_));
  NO4        m0942(.A(mai_mai_n970_), .B(mai_mai_n969_), .C(mai_mai_n556_), .D(mai_mai_n291_), .Y(mai_mai_n971_));
  NA2        m0943(.A(mai_mai_n386_), .B(mai_mai_n198_), .Y(mai_mai_n972_));
  AN2        m0944(.A(d), .B(c), .Y(mai_mai_n973_));
  NA2        m0945(.A(mai_mai_n973_), .B(mai_mai_n108_), .Y(mai_mai_n974_));
  NO4        m0946(.A(mai_mai_n974_), .B(mai_mai_n972_), .C(mai_mai_n167_), .D(mai_mai_n158_), .Y(mai_mai_n975_));
  NA2        m0947(.A(mai_mai_n468_), .B(c), .Y(mai_mai_n976_));
  NO4        m0948(.A(mai_mai_n970_), .B(mai_mai_n552_), .C(mai_mai_n976_), .D(mai_mai_n291_), .Y(mai_mai_n977_));
  OR2        m0949(.A(mai_mai_n975_), .B(mai_mai_n977_), .Y(mai_mai_n978_));
  OR3        m0950(.A(mai_mai_n978_), .B(mai_mai_n971_), .C(mai_mai_n968_), .Y(mai_mai_n979_));
  NAi32      m0951(.An(f), .Bn(e), .C(c), .Y(mai_mai_n980_));
  OR3        m0952(.A(mai_mai_n207_), .B(mai_mai_n167_), .C(mai_mai_n158_), .Y(mai_mai_n981_));
  NO2        m0953(.A(mai_mai_n981_), .B(mai_mai_n980_), .Y(mai_mai_n982_));
  NO2        m0954(.A(mai_mai_n976_), .B(mai_mai_n291_), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n592_), .B(mai_mai_n1383_), .Y(mai_mai_n984_));
  NOi21      m0956(.An(mai_mai_n983_), .B(mai_mai_n984_), .Y(mai_mai_n985_));
  NO2        m0957(.A(mai_mai_n716_), .B(mai_mai_n104_), .Y(mai_mai_n986_));
  NOi41      m0958(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n987_), .B(mai_mai_n986_), .Y(mai_mai_n988_));
  NO2        m0960(.A(mai_mai_n988_), .B(mai_mai_n980_), .Y(mai_mai_n989_));
  NA3        m0961(.A(k), .B(j), .C(i), .Y(mai_mai_n990_));
  NO3        m0962(.A(mai_mai_n990_), .B(mai_mai_n291_), .C(mai_mai_n83_), .Y(mai_mai_n991_));
  BUFFER     m0963(.A(mai_mai_n991_), .Y(mai_mai_n992_));
  OR4        m0964(.A(mai_mai_n992_), .B(mai_mai_n989_), .C(mai_mai_n985_), .D(mai_mai_n982_), .Y(mai_mai_n993_));
  NA3        m0965(.A(mai_mai_n435_), .B(mai_mai_n319_), .C(mai_mai_n54_), .Y(mai_mai_n994_));
  NO2        m0966(.A(mai_mai_n994_), .B(mai_mai_n984_), .Y(mai_mai_n995_));
  NO3        m0967(.A(mai_mai_n994_), .B(mai_mai_n552_), .C(mai_mai_n424_), .Y(mai_mai_n996_));
  NO2        m0968(.A(f), .B(c), .Y(mai_mai_n997_));
  NOi21      m0969(.An(mai_mai_n997_), .B(mai_mai_n418_), .Y(mai_mai_n998_));
  NA2        m0970(.A(mai_mai_n998_), .B(mai_mai_n57_), .Y(mai_mai_n999_));
  OR2        m0971(.A(k), .B(i), .Y(mai_mai_n1000_));
  NO3        m0972(.A(mai_mai_n1000_), .B(h), .C(l), .Y(mai_mai_n1001_));
  NOi31      m0973(.An(mai_mai_n1001_), .B(mai_mai_n999_), .C(j), .Y(mai_mai_n1002_));
  OR3        m0974(.A(mai_mai_n1002_), .B(mai_mai_n996_), .C(mai_mai_n995_), .Y(mai_mai_n1003_));
  OR3        m0975(.A(mai_mai_n1003_), .B(mai_mai_n993_), .C(mai_mai_n979_), .Y(mai02));
  OR2        m0976(.A(l), .B(k), .Y(mai_mai_n1005_));
  OR3        m0977(.A(h), .B(g), .C(f), .Y(mai_mai_n1006_));
  OR3        m0978(.A(n), .B(m), .C(i), .Y(mai_mai_n1007_));
  NO4        m0979(.A(mai_mai_n1007_), .B(mai_mai_n1006_), .C(mai_mai_n1005_), .D(e), .Y(mai_mai_n1008_));
  NO2        m0980(.A(mai_mai_n991_), .B(mai_mai_n971_), .Y(mai_mai_n1009_));
  AN3        m0981(.A(g), .B(f), .C(c), .Y(mai_mai_n1010_));
  NA2        m0982(.A(mai_mai_n1010_), .B(mai_mai_n435_), .Y(mai_mai_n1011_));
  OR2        m0983(.A(mai_mai_n990_), .B(mai_mai_n291_), .Y(mai_mai_n1012_));
  OR2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .Y(mai_mai_n1013_));
  NO3        m0985(.A(mai_mai_n994_), .B(mai_mai_n970_), .C(mai_mai_n552_), .Y(mai_mai_n1014_));
  NO2        m0986(.A(mai_mai_n1014_), .B(mai_mai_n982_), .Y(mai_mai_n1015_));
  NA3        m0987(.A(l), .B(k), .C(j), .Y(mai_mai_n1016_));
  NA2        m0988(.A(i), .B(h), .Y(mai_mai_n1017_));
  NO3        m0989(.A(mai_mai_n1017_), .B(mai_mai_n1016_), .C(mai_mai_n124_), .Y(mai_mai_n1018_));
  NO3        m0990(.A(mai_mai_n132_), .B(mai_mai_n266_), .C(mai_mai_n199_), .Y(mai_mai_n1019_));
  AOI210     m0991(.A0(mai_mai_n1019_), .A1(mai_mai_n1018_), .B0(mai_mai_n985_), .Y(mai_mai_n1020_));
  NA3        m0992(.A(c), .B(b), .C(a), .Y(mai_mai_n1021_));
  NO3        m0993(.A(mai_mai_n1021_), .B(mai_mai_n845_), .C(mai_mai_n198_), .Y(mai_mai_n1022_));
  NO2        m0994(.A(mai_mai_n284_), .B(mai_mai_n49_), .Y(mai_mai_n1023_));
  AOI210     m0995(.A0(mai_mai_n1023_), .A1(mai_mai_n1022_), .B0(mai_mai_n995_), .Y(mai_mai_n1024_));
  AN4        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1020_), .C(mai_mai_n1015_), .D(mai_mai_n1013_), .Y(mai_mai_n1025_));
  NO2        m0997(.A(mai_mai_n974_), .B(mai_mai_n972_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n988_), .B(mai_mai_n981_), .Y(mai_mai_n1027_));
  AOI210     m0999(.A0(mai_mai_n1027_), .A1(mai_mai_n1026_), .B0(mai_mai_n968_), .Y(mai_mai_n1028_));
  NAi41      m1000(.An(mai_mai_n1008_), .B(mai_mai_n1028_), .C(mai_mai_n1025_), .D(mai_mai_n1009_), .Y(mai03));
  NO2        m1001(.A(mai_mai_n496_), .B(mai_mai_n565_), .Y(mai_mai_n1030_));
  NA4        m1002(.A(mai_mai_n543_), .B(m), .C(mai_mai_n104_), .D(mai_mai_n198_), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n1031_), .B(mai_mai_n351_), .Y(mai_mai_n1032_));
  NO3        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1030_), .C(mai_mai_n936_), .Y(mai_mai_n1033_));
  NOi31      m1005(.An(mai_mai_n752_), .B(mai_mai_n799_), .C(mai_mai_n791_), .Y(mai_mai_n1034_));
  OAI220     m1006(.A0(mai_mai_n1034_), .A1(mai_mai_n650_), .B0(mai_mai_n1033_), .B1(mai_mai_n553_), .Y(mai_mai_n1035_));
  NOi31      m1007(.An(i), .B(k), .C(j), .Y(mai_mai_n1036_));
  NA4        m1008(.A(mai_mai_n1036_), .B(e), .C(mai_mai_n326_), .D(mai_mai_n319_), .Y(mai_mai_n1037_));
  OAI210     m1009(.A0(mai_mai_n767_), .A1(mai_mai_n396_), .B0(mai_mai_n1037_), .Y(mai_mai_n1038_));
  NOi31      m1010(.An(m), .B(n), .C(f), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n1039_), .B(mai_mai_n50_), .Y(mai_mai_n1040_));
  NA2        m1012(.A(c), .B(a), .Y(mai_mai_n1041_));
  OAI220     m1013(.A0(mai_mai_n1041_), .A1(mai_mai_n1040_), .B0(mai_mai_n832_), .B1(mai_mai_n401_), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n478_), .B(l), .Y(mai_mai_n1043_));
  NOi31      m1015(.An(mai_mai_n810_), .B(mai_mai_n966_), .C(mai_mai_n1043_), .Y(mai_mai_n1044_));
  NO4        m1016(.A(mai_mai_n1044_), .B(mai_mai_n1042_), .C(mai_mai_n1038_), .D(mai_mai_n935_), .Y(mai_mai_n1045_));
  INV        m1017(.A(mai_mai_n971_), .Y(mai_mai_n1046_));
  NO2        m1018(.A(mai_mai_n1017_), .B(mai_mai_n455_), .Y(mai_mai_n1047_));
  NO2        m1019(.A(mai_mai_n80_), .B(g), .Y(mai_mai_n1048_));
  AOI210     m1020(.A0(mai_mai_n1048_), .A1(mai_mai_n1047_), .B0(mai_mai_n1001_), .Y(mai_mai_n1049_));
  OR2        m1021(.A(mai_mai_n1049_), .B(mai_mai_n999_), .Y(mai_mai_n1050_));
  NA3        m1022(.A(mai_mai_n1050_), .B(mai_mai_n1046_), .C(mai_mai_n1045_), .Y(mai_mai_n1051_));
  NO4        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1035_), .C(mai_mai_n769_), .D(mai_mai_n533_), .Y(mai_mai_n1052_));
  NA2        m1024(.A(c), .B(b), .Y(mai_mai_n1053_));
  NO2        m1025(.A(mai_mai_n660_), .B(mai_mai_n1053_), .Y(mai_mai_n1054_));
  OAI210     m1026(.A0(mai_mai_n808_), .A1(mai_mai_n784_), .B0(mai_mai_n390_), .Y(mai_mai_n1055_));
  OAI210     m1027(.A0(mai_mai_n1055_), .A1(mai_mai_n809_), .B0(mai_mai_n1054_), .Y(mai_mai_n1056_));
  NAi21      m1028(.An(mai_mai_n397_), .B(mai_mai_n1054_), .Y(mai_mai_n1057_));
  NA3        m1029(.A(mai_mai_n402_), .B(mai_mai_n526_), .C(f), .Y(mai_mai_n1058_));
  NA2        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1057_), .Y(mai_mai_n1059_));
  NA2        m1031(.A(mai_mai_n245_), .B(mai_mai_n111_), .Y(mai_mai_n1060_));
  OAI210     m1032(.A0(mai_mai_n1060_), .A1(mai_mai_n270_), .B0(g), .Y(mai_mai_n1061_));
  NAi21      m1033(.An(f), .B(d), .Y(mai_mai_n1062_));
  NO2        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1021_), .Y(mai_mai_n1063_));
  INV        m1035(.A(mai_mai_n1063_), .Y(mai_mai_n1064_));
  AOI210     m1036(.A0(mai_mai_n1061_), .A1(mai_mai_n276_), .B0(mai_mai_n1064_), .Y(mai_mai_n1065_));
  AOI210     m1037(.A0(mai_mai_n1065_), .A1(mai_mai_n105_), .B0(mai_mai_n1059_), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n438_), .B(mai_mai_n437_), .Y(mai_mai_n1067_));
  NO2        m1039(.A(mai_mai_n172_), .B(mai_mai_n220_), .Y(mai_mai_n1068_));
  NA2        m1040(.A(mai_mai_n1068_), .B(m), .Y(mai_mai_n1069_));
  NA3        m1041(.A(mai_mai_n862_), .B(mai_mai_n1043_), .C(mai_mai_n441_), .Y(mai_mai_n1070_));
  OAI210     m1042(.A0(mai_mai_n1070_), .A1(mai_mai_n295_), .B0(mai_mai_n439_), .Y(mai_mai_n1071_));
  AOI210     m1043(.A0(mai_mai_n1071_), .A1(mai_mai_n1067_), .B0(mai_mai_n1069_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n147_), .B(mai_mai_n33_), .Y(mai_mai_n1073_));
  AOI210     m1045(.A0(mai_mai_n903_), .A1(mai_mai_n1073_), .B0(mai_mai_n199_), .Y(mai_mai_n1074_));
  NA2        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1063_), .Y(mai_mai_n1075_));
  NA2        m1047(.A(mai_mai_n1068_), .B(mai_mai_n404_), .Y(mai_mai_n1076_));
  NA2        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1075_), .Y(mai_mai_n1077_));
  NO2        m1049(.A(mai_mai_n1077_), .B(mai_mai_n1072_), .Y(mai_mai_n1078_));
  NA4        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1066_), .C(mai_mai_n1056_), .D(mai_mai_n1052_), .Y(mai00));
  NO2        m1051(.A(mai_mai_n283_), .B(mai_mai_n259_), .Y(mai_mai_n1080_));
  NO2        m1052(.A(mai_mai_n1080_), .B(mai_mai_n545_), .Y(mai_mai_n1081_));
  AOI210     m1053(.A0(mai_mai_n842_), .A1(mai_mai_n888_), .B0(mai_mai_n1038_), .Y(mai_mai_n1082_));
  NO2        m1054(.A(mai_mai_n1014_), .B(mai_mai_n667_), .Y(mai_mai_n1083_));
  NA3        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1082_), .C(mai_mai_n937_), .Y(mai_mai_n1084_));
  NA2        m1056(.A(mai_mai_n283_), .B(f), .Y(mai_mai_n1085_));
  NO2        m1057(.A(mai_mai_n1085_), .B(mai_mai_n974_), .Y(mai_mai_n1086_));
  NO4        m1058(.A(mai_mai_n1086_), .B(mai_mai_n1084_), .C(mai_mai_n1081_), .D(mai_mai_n993_), .Y(mai_mai_n1087_));
  NA3        m1059(.A(mai_mai_n157_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1088_));
  NA3        m1060(.A(d), .B(mai_mai_n54_), .C(b), .Y(mai_mai_n1089_));
  NOi31      m1061(.An(n), .B(m), .C(i), .Y(mai_mai_n1090_));
  NA3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n606_), .C(mai_mai_n50_), .Y(mai_mai_n1091_));
  OAI210     m1063(.A0(mai_mai_n1089_), .A1(mai_mai_n1088_), .B0(mai_mai_n1091_), .Y(mai_mai_n1092_));
  NO2        m1064(.A(mai_mai_n1092_), .B(mai_mai_n865_), .Y(mai_mai_n1093_));
  NO4        m1065(.A(mai_mai_n458_), .B(mai_mai_n338_), .C(mai_mai_n1053_), .D(mai_mai_n57_), .Y(mai_mai_n1094_));
  OR2        m1066(.A(mai_mai_n367_), .B(mai_mai_n125_), .Y(mai_mai_n1095_));
  NO2        m1067(.A(h), .B(g), .Y(mai_mai_n1096_));
  NO2        m1068(.A(mai_mai_n496_), .B(mai_mai_n565_), .Y(mai_mai_n1097_));
  NA2        m1069(.A(mai_mai_n1097_), .B(mai_mai_n505_), .Y(mai_mai_n1098_));
  NA2        m1070(.A(mai_mai_n168_), .B(mai_mai_n137_), .Y(mai_mai_n1099_));
  NA3        m1071(.A(mai_mai_n1099_), .B(mai_mai_n1098_), .C(mai_mai_n1095_), .Y(mai_mai_n1100_));
  NO3        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1094_), .C(mai_mai_n251_), .Y(mai_mai_n1101_));
  INV        m1073(.A(mai_mai_n307_), .Y(mai_mai_n1102_));
  NA2        m1074(.A(mai_mai_n1102_), .B(mai_mai_n143_), .Y(mai_mai_n1103_));
  NO2        m1075(.A(mai_mai_n222_), .B(mai_mai_n171_), .Y(mai_mai_n1104_));
  NA2        m1076(.A(mai_mai_n1104_), .B(mai_mai_n402_), .Y(mai_mai_n1105_));
  NA3        m1077(.A(mai_mai_n170_), .B(mai_mai_n104_), .C(g), .Y(mai_mai_n1106_));
  NA2        m1078(.A(mai_mai_n435_), .B(f), .Y(mai_mai_n1107_));
  NOi31      m1079(.An(mai_mai_n818_), .B(mai_mai_n1107_), .C(mai_mai_n1106_), .Y(mai_mai_n1108_));
  NAi31      m1080(.An(mai_mai_n174_), .B(mai_mai_n805_), .C(mai_mai_n435_), .Y(mai_mai_n1109_));
  NAi31      m1081(.An(mai_mai_n1108_), .B(mai_mai_n1109_), .C(mai_mai_n1105_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n258_), .B(mai_mai_n72_), .Y(mai_mai_n1111_));
  NO3        m1083(.A(mai_mai_n401_), .B(mai_mai_n780_), .C(n), .Y(mai_mai_n1112_));
  AOI210     m1084(.A0(mai_mai_n1112_), .A1(mai_mai_n1111_), .B0(mai_mai_n1008_), .Y(mai_mai_n1113_));
  NAi31      m1085(.An(mai_mai_n977_), .B(mai_mai_n1113_), .C(mai_mai_n71_), .Y(mai_mai_n1114_));
  NO4        m1086(.A(mai_mai_n1114_), .B(mai_mai_n1110_), .C(mai_mai_n1103_), .D(mai_mai_n487_), .Y(mai_mai_n1115_));
  AN3        m1087(.A(mai_mai_n1115_), .B(mai_mai_n1101_), .C(mai_mai_n1093_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(mai_mai_n505_), .B(mai_mai_n93_), .Y(mai_mai_n1117_));
  NA3        m1089(.A(mai_mai_n1039_), .B(mai_mai_n571_), .C(mai_mai_n434_), .Y(mai_mai_n1118_));
  NA4        m1090(.A(mai_mai_n1118_), .B(mai_mai_n529_), .C(mai_mai_n1117_), .D(mai_mai_n225_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n1032_), .B(mai_mai_n505_), .Y(mai_mai_n1120_));
  NA2        m1092(.A(mai_mai_n1120_), .B(mai_mai_n280_), .Y(mai_mai_n1121_));
  OAI210     m1093(.A0(mai_mai_n433_), .A1(mai_mai_n112_), .B0(mai_mai_n811_), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n1122_), .B(mai_mai_n1070_), .Y(mai_mai_n1123_));
  OR3        m1095(.A(mai_mai_n974_), .B(mai_mai_n256_), .C(mai_mai_n205_), .Y(mai_mai_n1124_));
  NO2        m1096(.A(mai_mai_n202_), .B(mai_mai_n199_), .Y(mai_mai_n1125_));
  NA2        m1097(.A(mai_mai_n795_), .B(mai_mai_n1125_), .Y(mai_mai_n1126_));
  OAI210     m1098(.A0(mai_mai_n339_), .A1(mai_mai_n296_), .B0(mai_mai_n423_), .Y(mai_mai_n1127_));
  NA4        m1099(.A(mai_mai_n1127_), .B(mai_mai_n1126_), .C(mai_mai_n1124_), .D(mai_mai_n1123_), .Y(mai_mai_n1128_));
  INV        m1100(.A(mai_mai_n768_), .Y(mai_mai_n1129_));
  AOI220     m1101(.A0(mai_mai_n895_), .A1(mai_mai_n544_), .B0(mai_mai_n606_), .B1(mai_mai_n227_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n66_), .B(h), .Y(mai_mai_n1131_));
  NO3        m1103(.A(mai_mai_n974_), .B(mai_mai_n972_), .C(mai_mai_n682_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n1005_), .B(mai_mai_n124_), .Y(mai_mai_n1133_));
  AN2        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1019_), .Y(mai_mai_n1134_));
  OAI210     m1106(.A0(mai_mai_n1134_), .A1(mai_mai_n1132_), .B0(mai_mai_n1131_), .Y(mai_mai_n1135_));
  NA4        m1107(.A(mai_mai_n1135_), .B(mai_mai_n1130_), .C(mai_mai_n1129_), .D(mai_mai_n813_), .Y(mai_mai_n1136_));
  NO4        m1108(.A(mai_mai_n1136_), .B(mai_mai_n1128_), .C(mai_mai_n1121_), .D(mai_mai_n1119_), .Y(mai_mai_n1137_));
  NA2        m1109(.A(mai_mai_n785_), .B(mai_mai_n711_), .Y(mai_mai_n1138_));
  NA4        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1137_), .C(mai_mai_n1116_), .D(mai_mai_n1087_), .Y(mai01));
  AN2        m1111(.A(mai_mai_n956_), .B(mai_mai_n954_), .Y(mai_mai_n1140_));
  NO4        m1112(.A(mai_mai_n748_), .B(mai_mai_n741_), .C(mai_mai_n449_), .D(mai_mai_n264_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1140_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n858_), .B(mai_mai_n318_), .Y(mai_mai_n1143_));
  NA2        m1115(.A(mai_mai_n665_), .B(mai_mai_n88_), .Y(mai_mai_n1144_));
  INV        m1116(.A(mai_mai_n1144_), .Y(mai_mai_n1145_));
  NA2        m1117(.A(mai_mai_n1145_), .B(mai_mai_n597_), .Y(mai_mai_n1146_));
  INV        m1118(.A(mai_mai_n110_), .Y(mai_mai_n1147_));
  OA220      m1119(.A0(mai_mai_n1147_), .A1(mai_mai_n551_), .B0(mai_mai_n619_), .B1(mai_mai_n351_), .Y(mai_mai_n1148_));
  NAi31      m1120(.An(mai_mai_n150_), .B(mai_mai_n1148_), .C(mai_mai_n1146_), .Y(mai_mai_n1149_));
  NO3        m1121(.A(mai_mai_n731_), .B(mai_mai_n634_), .C(mai_mai_n480_), .Y(mai_mai_n1150_));
  NA4        m1122(.A(mai_mai_n665_), .B(mai_mai_n88_), .C(mai_mai_n45_), .D(mai_mai_n198_), .Y(mai_mai_n1151_));
  OR2        m1123(.A(mai_mai_n184_), .B(mai_mai_n182_), .Y(mai_mai_n1152_));
  NA3        m1124(.A(mai_mai_n1152_), .B(mai_mai_n1150_), .C(mai_mai_n128_), .Y(mai_mai_n1153_));
  NO4        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1149_), .C(mai_mai_n1143_), .D(mai_mai_n1142_), .Y(mai_mai_n1154_));
  NA2        m1126(.A(mai_mai_n286_), .B(mai_mai_n500_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n508_), .B(mai_mai_n372_), .Y(mai_mai_n1156_));
  NA2        m1128(.A(mai_mai_n530_), .B(mai_mai_n1156_), .Y(mai_mai_n1157_));
  AOI210     m1129(.A0(mai_mai_n191_), .A1(mai_mai_n82_), .B0(mai_mai_n198_), .Y(mai_mai_n1158_));
  OAI210     m1130(.A0(mai_mai_n755_), .A1(mai_mai_n402_), .B0(mai_mai_n1158_), .Y(mai_mai_n1159_));
  AN3        m1131(.A(m), .B(l), .C(k), .Y(mai_mai_n1160_));
  OAI210     m1132(.A0(mai_mai_n341_), .A1(mai_mai_n34_), .B0(mai_mai_n1160_), .Y(mai_mai_n1161_));
  NA2        m1133(.A(mai_mai_n190_), .B(mai_mai_n34_), .Y(mai_mai_n1162_));
  AO210      m1134(.A0(mai_mai_n1162_), .A1(mai_mai_n1161_), .B0(mai_mai_n317_), .Y(mai_mai_n1163_));
  NA4        m1135(.A(mai_mai_n1163_), .B(mai_mai_n1159_), .C(mai_mai_n1157_), .D(mai_mai_n1155_), .Y(mai_mai_n1164_));
  NA2        m1136(.A(mai_mai_n563_), .B(mai_mai_n110_), .Y(mai_mai_n1165_));
  OAI210     m1137(.A0(mai_mai_n1147_), .A1(mai_mai_n560_), .B0(mai_mai_n1165_), .Y(mai_mai_n1166_));
  NO3        m1138(.A(mai_mai_n767_), .B(mai_mai_n191_), .C(mai_mai_n384_), .Y(mai_mai_n1167_));
  INV        m1139(.A(mai_mai_n1167_), .Y(mai_mai_n1168_));
  OAI210     m1140(.A0(mai_mai_n1145_), .A1(mai_mai_n312_), .B0(mai_mai_n635_), .Y(mai_mai_n1169_));
  NA3        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1168_), .C(mai_mai_n734_), .Y(mai_mai_n1170_));
  NO3        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1166_), .C(mai_mai_n1164_), .Y(mai_mai_n1171_));
  NA3        m1143(.A(mai_mai_n569_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1172_));
  NO2        m1144(.A(mai_mai_n1172_), .B(mai_mai_n191_), .Y(mai_mai_n1173_));
  AOI210     m1145(.A0(mai_mai_n476_), .A1(mai_mai_n56_), .B0(mai_mai_n1173_), .Y(mai_mai_n1174_));
  OR2        m1146(.A(mai_mai_n1144_), .B(mai_mai_n570_), .Y(mai_mai_n1175_));
  NO2        m1147(.A(mai_mai_n1151_), .B(mai_mai_n917_), .Y(mai_mai_n1176_));
  NO2        m1148(.A(mai_mai_n1176_), .B(mai_mai_n1092_), .Y(mai_mai_n1177_));
  NA4        m1149(.A(mai_mai_n1177_), .B(mai_mai_n1175_), .C(mai_mai_n1174_), .D(mai_mai_n710_), .Y(mai_mai_n1178_));
  NO2        m1150(.A(mai_mai_n907_), .B(mai_mai_n215_), .Y(mai_mai_n1179_));
  NA2        m1151(.A(mai_mai_n540_), .B(mai_mai_n538_), .Y(mai_mai_n1180_));
  NA2        m1152(.A(mai_mai_n1180_), .B(mai_mai_n629_), .Y(mai_mai_n1181_));
  NO2        m1153(.A(mai_mai_n351_), .B(mai_mai_n70_), .Y(mai_mai_n1182_));
  NO3        m1154(.A(mai_mai_n1182_), .B(mai_mai_n1181_), .C(mai_mai_n1178_), .Y(mai_mai_n1183_));
  NO2        m1155(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1184_));
  AN2        m1156(.A(mai_mai_n1184_), .B(mai_mai_n587_), .Y(mai_mai_n1185_));
  NA2        m1157(.A(mai_mai_n1185_), .B(mai_mai_n324_), .Y(mai_mai_n1186_));
  INV        m1158(.A(mai_mai_n125_), .Y(mai_mai_n1187_));
  NO3        m1159(.A(mai_mai_n1017_), .B(mai_mai_n167_), .C(mai_mai_n80_), .Y(mai_mai_n1188_));
  NA2        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1187_), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n1189_), .B(mai_mai_n1186_), .Y(mai_mai_n1190_));
  NO2        m1162(.A(mai_mai_n579_), .B(mai_mai_n578_), .Y(mai_mai_n1191_));
  NO4        m1163(.A(mai_mai_n1017_), .B(mai_mai_n1191_), .C(mai_mai_n165_), .D(mai_mai_n80_), .Y(mai_mai_n1192_));
  NO3        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1190_), .C(mai_mai_n600_), .Y(mai_mai_n1193_));
  NA4        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1183_), .C(mai_mai_n1171_), .D(mai_mai_n1154_), .Y(mai06));
  NO2        m1166(.A(mai_mai_n385_), .B(mai_mai_n527_), .Y(mai_mai_n1195_));
  NA2        m1167(.A(mai_mai_n252_), .B(mai_mai_n1195_), .Y(mai_mai_n1196_));
  NO3        m1168(.A(mai_mai_n566_), .B(mai_mai_n753_), .C(mai_mai_n567_), .Y(mai_mai_n1197_));
  OR2        m1169(.A(mai_mai_n1197_), .B(mai_mai_n832_), .Y(mai_mai_n1198_));
  NA2        m1170(.A(mai_mai_n1198_), .B(mai_mai_n1196_), .Y(mai_mai_n1199_));
  NO3        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1181_), .C(mai_mai_n240_), .Y(mai_mai_n1200_));
  NO2        m1172(.A(mai_mai_n284_), .B(mai_mai_n45_), .Y(mai_mai_n1201_));
  AOI210     m1173(.A0(mai_mai_n1201_), .A1(mai_mai_n523_), .B0(mai_mai_n1179_), .Y(mai_mai_n1202_));
  INV        m1174(.A(mai_mai_n1185_), .Y(mai_mai_n1203_));
  AOI210     m1175(.A0(mai_mai_n1203_), .A1(mai_mai_n1202_), .B0(mai_mai_n321_), .Y(mai_mai_n1204_));
  INV        m1176(.A(mai_mai_n633_), .Y(mai_mai_n1205_));
  NA2        m1177(.A(mai_mai_n1205_), .B(mai_mai_n604_), .Y(mai_mai_n1206_));
  NO2        m1178(.A(mai_mai_n483_), .B(mai_mai_n162_), .Y(mai_mai_n1207_));
  NOi21      m1179(.An(mai_mai_n127_), .B(mai_mai_n45_), .Y(mai_mai_n1208_));
  NO2        m1180(.A(mai_mai_n572_), .B(mai_mai_n1040_), .Y(mai_mai_n1209_));
  OAI210     m1181(.A0(mai_mai_n430_), .A1(mai_mai_n231_), .B0(mai_mai_n852_), .Y(mai_mai_n1210_));
  NO4        m1182(.A(mai_mai_n1210_), .B(mai_mai_n1209_), .C(mai_mai_n1208_), .D(mai_mai_n1207_), .Y(mai_mai_n1211_));
  NA2        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1206_), .Y(mai_mai_n1212_));
  NO2        m1184(.A(mai_mai_n701_), .B(mai_mai_n349_), .Y(mai_mai_n1213_));
  NO3        m1185(.A(mai_mai_n635_), .B(mai_mai_n712_), .C(mai_mai_n597_), .Y(mai_mai_n1214_));
  NOi21      m1186(.An(mai_mai_n1213_), .B(mai_mai_n1214_), .Y(mai_mai_n1215_));
  NO3        m1187(.A(mai_mai_n1215_), .B(mai_mai_n1212_), .C(mai_mai_n1204_), .Y(mai_mai_n1216_));
  NO2        m1188(.A(mai_mai_n747_), .B(mai_mai_n260_), .Y(mai_mai_n1217_));
  OAI220     m1189(.A0(mai_mai_n689_), .A1(mai_mai_n47_), .B0(mai_mai_n207_), .B1(mai_mai_n581_), .Y(mai_mai_n1218_));
  OAI210     m1190(.A0(mai_mai_n260_), .A1(c), .B0(mai_mai_n603_), .Y(mai_mai_n1219_));
  AOI220     m1191(.A0(mai_mai_n1219_), .A1(mai_mai_n1218_), .B0(mai_mai_n1217_), .B1(mai_mai_n252_), .Y(mai_mai_n1220_));
  OAI220     m1192(.A0(mai_mai_n657_), .A1(mai_mai_n231_), .B0(mai_mai_n479_), .B1(mai_mai_n483_), .Y(mai_mai_n1221_));
  NO2        m1193(.A(mai_mai_n565_), .B(j), .Y(mai_mai_n1222_));
  NOi21      m1194(.An(mai_mai_n1222_), .B(mai_mai_n627_), .Y(mai_mai_n1223_));
  NO3        m1195(.A(mai_mai_n1223_), .B(mai_mai_n1221_), .C(mai_mai_n1042_), .Y(mai_mai_n1224_));
  NA4        m1196(.A(mai_mai_n739_), .B(mai_mai_n738_), .C(mai_mai_n412_), .D(mai_mai_n824_), .Y(mai_mai_n1225_));
  NAi31      m1197(.An(mai_mai_n701_), .B(mai_mai_n1225_), .C(mai_mai_n190_), .Y(mai_mai_n1226_));
  NA4        m1198(.A(mai_mai_n1226_), .B(mai_mai_n1224_), .C(mai_mai_n1220_), .D(mai_mai_n1130_), .Y(mai_mai_n1227_));
  OR2        m1199(.A(mai_mai_n730_), .B(mai_mai_n511_), .Y(mai_mai_n1228_));
  OR3        m1200(.A(mai_mai_n353_), .B(mai_mai_n207_), .C(mai_mai_n581_), .Y(mai_mai_n1229_));
  AOI210     m1201(.A0(mai_mai_n540_), .A1(mai_mai_n423_), .B0(mai_mai_n355_), .Y(mai_mai_n1230_));
  NA3        m1202(.A(mai_mai_n1230_), .B(mai_mai_n1229_), .C(mai_mai_n1228_), .Y(mai_mai_n1231_));
  NA2        m1203(.A(mai_mai_n1213_), .B(mai_mai_n711_), .Y(mai_mai_n1232_));
  AN2        m1204(.A(mai_mai_n874_), .B(mai_mai_n873_), .Y(mai_mai_n1233_));
  NO4        m1205(.A(mai_mai_n1233_), .B(mai_mai_n822_), .C(mai_mai_n472_), .D(mai_mai_n452_), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n1234_), .B(mai_mai_n1232_), .Y(mai_mai_n1235_));
  NAi21      m1207(.An(j), .B(i), .Y(mai_mai_n1236_));
  NO4        m1208(.A(mai_mai_n1191_), .B(mai_mai_n1236_), .C(mai_mai_n418_), .D(mai_mai_n218_), .Y(mai_mai_n1237_));
  NO4        m1209(.A(mai_mai_n1237_), .B(mai_mai_n1235_), .C(mai_mai_n1231_), .D(mai_mai_n1227_), .Y(mai_mai_n1238_));
  NA4        m1210(.A(mai_mai_n1238_), .B(mai_mai_n1216_), .C(mai_mai_n1200_), .D(mai_mai_n1193_), .Y(mai07));
  NOi21      m1211(.An(j), .B(k), .Y(mai_mai_n1240_));
  NA4        m1212(.A(mai_mai_n170_), .B(mai_mai_n100_), .C(mai_mai_n1240_), .D(f), .Y(mai_mai_n1241_));
  NAi21      m1213(.An(f), .B(c), .Y(mai_mai_n1242_));
  OR2        m1214(.A(e), .B(d), .Y(mai_mai_n1243_));
  NO2        m1215(.A(mai_mai_n591_), .B(mai_mai_n308_), .Y(mai_mai_n1244_));
  NA3        m1216(.A(mai_mai_n1244_), .B(mai_mai_n1383_), .C(mai_mai_n170_), .Y(mai_mai_n1245_));
  NOi31      m1217(.An(n), .B(m), .C(b), .Y(mai_mai_n1246_));
  NO3        m1218(.A(mai_mai_n124_), .B(mai_mai_n424_), .C(h), .Y(mai_mai_n1247_));
  NA2        m1219(.A(mai_mai_n1245_), .B(mai_mai_n1241_), .Y(mai_mai_n1248_));
  NOi41      m1220(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1249_));
  NO2        m1221(.A(k), .B(i), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n80_), .B(mai_mai_n45_), .Y(mai_mai_n1251_));
  NO2        m1223(.A(mai_mai_n980_), .B(mai_mai_n418_), .Y(mai_mai_n1252_));
  NA3        m1224(.A(mai_mai_n1252_), .B(mai_mai_n1251_), .C(mai_mai_n199_), .Y(mai_mai_n1253_));
  NO2        m1225(.A(mai_mai_n990_), .B(mai_mai_n291_), .Y(mai_mai_n1254_));
  NA2        m1226(.A(mai_mai_n512_), .B(mai_mai_n75_), .Y(mai_mai_n1255_));
  NA2        m1227(.A(mai_mai_n1131_), .B(mai_mai_n274_), .Y(mai_mai_n1256_));
  NA3        m1228(.A(mai_mai_n1256_), .B(mai_mai_n1255_), .C(mai_mai_n1253_), .Y(mai_mai_n1257_));
  NO2        m1229(.A(mai_mai_n1257_), .B(mai_mai_n1248_), .Y(mai_mai_n1258_));
  NO3        m1230(.A(e), .B(d), .C(c), .Y(mai_mai_n1259_));
  NA2        m1231(.A(mai_mai_n1381_), .B(mai_mai_n1259_), .Y(mai_mai_n1260_));
  NO2        m1232(.A(mai_mai_n1260_), .B(mai_mai_n199_), .Y(mai_mai_n1261_));
  NA3        m1233(.A(mai_mai_n654_), .B(mai_mai_n643_), .C(mai_mai_n104_), .Y(mai_mai_n1262_));
  NO2        m1234(.A(mai_mai_n1262_), .B(mai_mai_n45_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(l), .B(k), .Y(mai_mai_n1264_));
  NOi41      m1236(.An(mai_mai_n517_), .B(mai_mai_n1264_), .C(mai_mai_n447_), .D(mai_mai_n418_), .Y(mai_mai_n1265_));
  NO3        m1237(.A(mai_mai_n1265_), .B(mai_mai_n1263_), .C(mai_mai_n1261_), .Y(mai_mai_n1266_));
  NO2        m1238(.A(mai_mai_n1000_), .B(l), .Y(mai_mai_n1267_));
  NO2        m1239(.A(g), .B(c), .Y(mai_mai_n1268_));
  NA3        m1240(.A(mai_mai_n1268_), .B(mai_mai_n132_), .C(mai_mai_n175_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n1269_), .B(mai_mai_n1267_), .Y(mai_mai_n1270_));
  NA2        m1242(.A(mai_mai_n1270_), .B(mai_mai_n170_), .Y(mai_mai_n1271_));
  NO2        m1243(.A(mai_mai_n425_), .B(a), .Y(mai_mai_n1272_));
  NA3        m1244(.A(mai_mai_n1272_), .B(k), .C(mai_mai_n105_), .Y(mai_mai_n1273_));
  NO2        m1245(.A(i), .B(h), .Y(mai_mai_n1274_));
  NA2        m1246(.A(mai_mai_n1062_), .B(h), .Y(mai_mai_n1275_));
  NA2        m1247(.A(mai_mai_n129_), .B(mai_mai_n203_), .Y(mai_mai_n1276_));
  NO2        m1248(.A(mai_mai_n1276_), .B(mai_mai_n1275_), .Y(mai_mai_n1277_));
  NO2        m1249(.A(mai_mai_n708_), .B(mai_mai_n176_), .Y(mai_mai_n1278_));
  NOi31      m1250(.An(m), .B(n), .C(b), .Y(mai_mai_n1279_));
  NO2        m1251(.A(mai_mai_n1278_), .B(mai_mai_n1277_), .Y(mai_mai_n1280_));
  NA2        m1252(.A(mai_mai_n1010_), .B(mai_mai_n435_), .Y(mai_mai_n1281_));
  NO4        m1253(.A(mai_mai_n1281_), .B(mai_mai_n986_), .C(mai_mai_n418_), .D(mai_mai_n45_), .Y(mai_mai_n1282_));
  OAI210     m1254(.A0(mai_mai_n172_), .A1(mai_mai_n495_), .B0(mai_mai_n987_), .Y(mai_mai_n1283_));
  INV        m1255(.A(mai_mai_n1283_), .Y(mai_mai_n1284_));
  NO2        m1256(.A(mai_mai_n1284_), .B(mai_mai_n1282_), .Y(mai_mai_n1285_));
  AN4        m1257(.A(mai_mai_n1285_), .B(mai_mai_n1280_), .C(mai_mai_n1273_), .D(mai_mai_n1271_), .Y(mai_mai_n1286_));
  NA2        m1258(.A(mai_mai_n1246_), .B(mai_mai_n362_), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n176_), .B(b), .Y(mai_mai_n1288_));
  AOI220     m1260(.A0(mai_mai_n1090_), .A1(mai_mai_n1288_), .B0(mai_mai_n1018_), .B1(mai_mai_n1281_), .Y(mai_mai_n1289_));
  INV        m1261(.A(mai_mai_n1289_), .Y(mai_mai_n1290_));
  NO4        m1262(.A(mai_mai_n124_), .B(g), .C(f), .D(e), .Y(mai_mai_n1291_));
  NA2        m1263(.A(mai_mai_n275_), .B(h), .Y(mai_mai_n1292_));
  OR2        m1264(.A(e), .B(a), .Y(mai_mai_n1293_));
  NO2        m1265(.A(mai_mai_n1243_), .B(mai_mai_n1242_), .Y(mai_mai_n1294_));
  AOI210     m1266(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1294_), .Y(mai_mai_n1295_));
  NO2        m1267(.A(mai_mai_n1295_), .B(mai_mai_n1007_), .Y(mai_mai_n1296_));
  NA2        m1268(.A(mai_mai_n1249_), .B(mai_mai_n1264_), .Y(mai_mai_n1297_));
  INV        m1269(.A(mai_mai_n1297_), .Y(mai_mai_n1298_));
  NA2        m1270(.A(mai_mai_n1039_), .B(mai_mai_n384_), .Y(mai_mai_n1299_));
  NO3        m1271(.A(mai_mai_n1298_), .B(mai_mai_n1296_), .C(mai_mai_n1290_), .Y(mai_mai_n1300_));
  NA4        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1286_), .C(mai_mai_n1266_), .D(mai_mai_n1258_), .Y(mai_mai_n1301_));
  NO3        m1273(.A(mai_mai_n701_), .B(mai_mai_n165_), .C(mai_mai_n386_), .Y(mai_mai_n1302_));
  OR2        m1274(.A(n), .B(i), .Y(mai_mai_n1303_));
  OAI210     m1275(.A0(mai_mai_n1303_), .A1(mai_mai_n997_), .B0(mai_mai_n49_), .Y(mai_mai_n1304_));
  AOI220     m1276(.A0(mai_mai_n1304_), .A1(mai_mai_n1096_), .B0(mai_mai_n772_), .B1(mai_mai_n183_), .Y(mai_mai_n1305_));
  INV        m1277(.A(mai_mai_n1305_), .Y(mai_mai_n1306_));
  NO2        m1278(.A(mai_mai_n124_), .B(l), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n207_), .B(k), .Y(mai_mai_n1308_));
  OAI210     m1280(.A0(mai_mai_n1308_), .A1(mai_mai_n1274_), .B0(mai_mai_n1307_), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n1309_), .B(mai_mai_n31_), .Y(mai_mai_n1310_));
  NO2        m1282(.A(mai_mai_n1310_), .B(mai_mai_n1306_), .Y(mai_mai_n1311_));
  NO2        m1283(.A(mai_mai_n1007_), .B(h), .Y(mai_mai_n1312_));
  NA3        m1284(.A(mai_mai_n1312_), .B(d), .C(mai_mai_n972_), .Y(mai_mai_n1313_));
  NO2        m1285(.A(mai_mai_n1313_), .B(c), .Y(mai_mai_n1314_));
  NOi21      m1286(.An(d), .B(f), .Y(mai_mai_n1315_));
  NO2        m1287(.A(mai_mai_n1243_), .B(f), .Y(mai_mai_n1316_));
  INV        m1288(.A(mai_mai_n1314_), .Y(mai_mai_n1317_));
  NA3        m1289(.A(mai_mai_n1317_), .B(mai_mai_n1311_), .C(mai_mai_n1384_), .Y(mai_mai_n1318_));
  NO3        m1290(.A(mai_mai_n1010_), .B(mai_mai_n997_), .C(mai_mai_n40_), .Y(mai_mai_n1319_));
  NO2        m1291(.A(mai_mai_n435_), .B(mai_mai_n284_), .Y(mai_mai_n1320_));
  OAI210     m1292(.A0(mai_mai_n1320_), .A1(mai_mai_n1319_), .B0(mai_mai_n1254_), .Y(mai_mai_n1321_));
  OAI210     m1293(.A0(mai_mai_n1291_), .A1(mai_mai_n1246_), .B0(mai_mai_n829_), .Y(mai_mai_n1322_));
  NO2        m1294(.A(mai_mai_n969_), .B(mai_mai_n124_), .Y(mai_mai_n1323_));
  NA2        m1295(.A(mai_mai_n1323_), .B(mai_mai_n586_), .Y(mai_mai_n1324_));
  NA3        m1296(.A(mai_mai_n1324_), .B(mai_mai_n1322_), .C(mai_mai_n1321_), .Y(mai_mai_n1325_));
  NA2        m1297(.A(mai_mai_n1268_), .B(mai_mai_n1315_), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n1326_), .B(m), .Y(mai_mai_n1327_));
  NO2        m1299(.A(mai_mai_n140_), .B(mai_mai_n171_), .Y(mai_mai_n1328_));
  OAI210     m1300(.A0(mai_mai_n1328_), .A1(mai_mai_n102_), .B0(mai_mai_n1279_), .Y(mai_mai_n1329_));
  INV        m1301(.A(mai_mai_n1329_), .Y(mai_mai_n1330_));
  NO3        m1302(.A(mai_mai_n1330_), .B(mai_mai_n1327_), .C(mai_mai_n1325_), .Y(mai_mai_n1331_));
  NO2        m1303(.A(mai_mai_n1242_), .B(e), .Y(mai_mai_n1332_));
  INV        m1304(.A(mai_mai_n1332_), .Y(mai_mai_n1333_));
  NA2        m1305(.A(mai_mai_n1048_), .B(mai_mai_n595_), .Y(mai_mai_n1334_));
  OR3        m1306(.A(mai_mai_n1308_), .B(mai_mai_n1131_), .C(mai_mai_n124_), .Y(mai_mai_n1335_));
  OAI220     m1307(.A0(mai_mai_n1335_), .A1(mai_mai_n1333_), .B0(mai_mai_n1334_), .B1(mai_mai_n419_), .Y(mai_mai_n1336_));
  INV        m1308(.A(mai_mai_n1336_), .Y(mai_mai_n1337_));
  NO2        m1309(.A(mai_mai_n171_), .B(c), .Y(mai_mai_n1338_));
  OAI210     m1310(.A0(mai_mai_n1338_), .A1(mai_mai_n1332_), .B0(mai_mai_n170_), .Y(mai_mai_n1339_));
  AOI220     m1311(.A0(mai_mai_n1339_), .A1(mai_mai_n999_), .B0(mai_mai_n502_), .B1(mai_mai_n349_), .Y(mai_mai_n1340_));
  NO2        m1312(.A(mai_mai_n1293_), .B(f), .Y(mai_mai_n1341_));
  AOI210     m1313(.A0(mai_mai_n1048_), .A1(a), .B0(mai_mai_n1341_), .Y(mai_mai_n1342_));
  NO2        m1314(.A(mai_mai_n1342_), .B(mai_mai_n67_), .Y(mai_mai_n1343_));
  NA2        m1315(.A(mai_mai_n1341_), .B(mai_mai_n1251_), .Y(mai_mai_n1344_));
  OAI220     m1316(.A0(mai_mai_n1344_), .A1(mai_mai_n49_), .B0(mai_mai_n1382_), .B1(mai_mai_n165_), .Y(mai_mai_n1345_));
  NA4        m1317(.A(mai_mai_n1019_), .B(mai_mai_n1016_), .C(mai_mai_n203_), .D(mai_mai_n66_), .Y(mai_mai_n1346_));
  NA2        m1318(.A(mai_mai_n1247_), .B(mai_mai_n172_), .Y(mai_mai_n1347_));
  NO2        m1319(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1348_));
  OAI210     m1320(.A0(mai_mai_n1293_), .A1(mai_mai_n807_), .B0(mai_mai_n454_), .Y(mai_mai_n1349_));
  OAI210     m1321(.A0(mai_mai_n1349_), .A1(mai_mai_n1022_), .B0(mai_mai_n1348_), .Y(mai_mai_n1350_));
  NO2        m1322(.A(mai_mai_n236_), .B(g), .Y(mai_mai_n1351_));
  NO2        m1323(.A(m), .B(i), .Y(mai_mai_n1352_));
  NA2        m1324(.A(mai_mai_n998_), .B(mai_mai_n1351_), .Y(mai_mai_n1353_));
  NA4        m1325(.A(mai_mai_n1353_), .B(mai_mai_n1350_), .C(mai_mai_n1347_), .D(mai_mai_n1346_), .Y(mai_mai_n1354_));
  NO4        m1326(.A(mai_mai_n1354_), .B(mai_mai_n1345_), .C(mai_mai_n1343_), .D(mai_mai_n1340_), .Y(mai_mai_n1355_));
  NA3        m1327(.A(mai_mai_n1355_), .B(mai_mai_n1337_), .C(mai_mai_n1331_), .Y(mai_mai_n1356_));
  INV        m1328(.A(mai_mai_n173_), .Y(mai_mai_n1357_));
  NA2        m1329(.A(mai_mai_n1357_), .B(mai_mai_n1312_), .Y(mai_mai_n1358_));
  NOi21      m1330(.An(mai_mai_n1247_), .B(e), .Y(mai_mai_n1359_));
  AN2        m1331(.A(mai_mai_n1019_), .B(mai_mai_n1005_), .Y(mai_mai_n1360_));
  AOI220     m1332(.A0(mai_mai_n1352_), .A1(mai_mai_n602_), .B0(mai_mai_n1383_), .B1(mai_mai_n148_), .Y(mai_mai_n1361_));
  NOi31      m1333(.An(mai_mai_n30_), .B(mai_mai_n1361_), .C(n), .Y(mai_mai_n1362_));
  AOI210     m1334(.A0(mai_mai_n1360_), .A1(mai_mai_n1090_), .B0(mai_mai_n1362_), .Y(mai_mai_n1363_));
  NA2        m1335(.A(mai_mai_n57_), .B(a), .Y(mai_mai_n1364_));
  NO2        m1336(.A(mai_mai_n1250_), .B(mai_mai_n110_), .Y(mai_mai_n1365_));
  OAI220     m1337(.A0(mai_mai_n1365_), .A1(mai_mai_n1287_), .B0(mai_mai_n1299_), .B1(mai_mai_n1364_), .Y(mai_mai_n1366_));
  INV        m1338(.A(mai_mai_n1366_), .Y(mai_mai_n1367_));
  NA4        m1339(.A(mai_mai_n1367_), .B(mai_mai_n1363_), .C(mai_mai_n1387_), .D(mai_mai_n1358_), .Y(mai_mai_n1368_));
  OR4        m1340(.A(mai_mai_n1368_), .B(mai_mai_n1356_), .C(mai_mai_n1318_), .D(mai_mai_n1301_), .Y(mai04));
  NOi31      m1341(.An(mai_mai_n1291_), .B(mai_mai_n1292_), .C(mai_mai_n974_), .Y(mai_mai_n1370_));
  NA2        m1342(.A(mai_mai_n1316_), .B(mai_mai_n772_), .Y(mai_mai_n1371_));
  NO2        m1343(.A(mai_mai_n1371_), .B(mai_mai_n966_), .Y(mai_mai_n1372_));
  OR3        m1344(.A(mai_mai_n1372_), .B(mai_mai_n1370_), .C(mai_mai_n989_), .Y(mai_mai_n1373_));
  NO2        m1345(.A(mai_mai_n1251_), .B(mai_mai_n83_), .Y(mai_mai_n1374_));
  AOI210     m1346(.A0(mai_mai_n1374_), .A1(mai_mai_n983_), .B0(mai_mai_n1108_), .Y(mai_mai_n1375_));
  NA2        m1347(.A(mai_mai_n1375_), .B(mai_mai_n1135_), .Y(mai_mai_n1376_));
  NO4        m1348(.A(mai_mai_n1376_), .B(mai_mai_n1373_), .C(mai_mai_n996_), .D(mai_mai_n979_), .Y(mai_mai_n1377_));
  NA4        m1349(.A(mai_mai_n1377_), .B(mai_mai_n1050_), .C(mai_mai_n1037_), .D(mai_mai_n1025_), .Y(mai05));
  INV        m1350(.A(m), .Y(mai_mai_n1381_));
  INV        m1351(.A(mai_mai_n97_), .Y(mai_mai_n1382_));
  INV        m1352(.A(j), .Y(mai_mai_n1383_));
  INV        m1353(.A(mai_mai_n1302_), .Y(mai_mai_n1384_));
  INV        m1354(.A(mai_mai_n452_), .Y(mai_mai_n1385_));
  INV        m1355(.A(b), .Y(mai_mai_n1386_));
  INV        m1356(.A(mai_mai_n1359_), .Y(mai_mai_n1387_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO3        u0023(.A(men_men_n48_), .B(men_men_n43_), .C(men_men_n39_), .Y(men_men_n52_));
  AOI210     u0024(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n53_));
  INV        u0025(.A(c), .Y(men_men_n54_));
  NA2        u0026(.A(e), .B(b), .Y(men_men_n55_));
  NO2        u0027(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  INV        u0028(.A(d), .Y(men_men_n57_));
  NA2        u0029(.A(g), .B(men_men_n57_), .Y(men_men_n58_));
  NAi21      u0030(.An(i), .B(h), .Y(men_men_n59_));
  NAi31      u0031(.An(i), .B(l), .C(j), .Y(men_men_n60_));
  OAI220     u0032(.A0(men_men_n60_), .A1(men_men_n49_), .B0(men_men_n59_), .B1(men_men_n44_), .Y(men_men_n61_));
  NAi31      u0033(.An(men_men_n58_), .B(men_men_n61_), .C(men_men_n56_), .Y(men_men_n62_));
  NAi41      u0034(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n63_));
  NA2        u0035(.A(g), .B(f), .Y(men_men_n64_));
  NO2        u0036(.A(men_men_n64_), .B(men_men_n63_), .Y(men_men_n65_));
  NAi21      u0037(.An(i), .B(j), .Y(men_men_n66_));
  NAi32      u0038(.An(n), .Bn(k), .C(m), .Y(men_men_n67_));
  NAi31      u0039(.An(l), .B(m), .C(k), .Y(men_men_n68_));
  NAi21      u0040(.An(e), .B(h), .Y(men_men_n69_));
  NAi41      u0041(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n70_));
  INV        u0042(.A(m), .Y(men_men_n71_));
  NOi21      u0043(.An(k), .B(l), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  AN4        u0045(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n74_));
  NOi31      u0046(.An(h), .B(g), .C(f), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NAi32      u0048(.An(m), .Bn(k), .C(j), .Y(men_men_n77_));
  NOi32      u0049(.An(h), .Bn(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n74_), .Y(men_men_n79_));
  OA220      u0051(.A0(men_men_n79_), .A1(men_men_n77_), .B0(men_men_n76_), .B1(men_men_n73_), .Y(men_men_n80_));
  NA2        u0052(.A(men_men_n80_), .B(men_men_n62_), .Y(men_men_n81_));
  INV        u0053(.A(n), .Y(men_men_n82_));
  NOi32      u0054(.An(e), .Bn(b), .C(d), .Y(men_men_n83_));
  NA2        u0055(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n84_));
  INV        u0056(.A(j), .Y(men_men_n85_));
  AN3        u0057(.A(m), .B(k), .C(i), .Y(men_men_n86_));
  NA3        u0058(.A(men_men_n86_), .B(men_men_n85_), .C(g), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(f), .Y(men_men_n88_));
  NAi32      u0060(.An(g), .Bn(f), .C(h), .Y(men_men_n89_));
  NAi31      u0061(.An(j), .B(m), .C(l), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n91_));
  NA2        u0063(.A(m), .B(l), .Y(men_men_n92_));
  NAi31      u0064(.An(k), .B(j), .C(g), .Y(men_men_n93_));
  NO3        u0065(.A(men_men_n93_), .B(men_men_n92_), .C(f), .Y(men_men_n94_));
  AN2        u0066(.A(j), .B(g), .Y(men_men_n95_));
  NOi32      u0067(.An(m), .Bn(l), .C(i), .Y(men_men_n96_));
  NOi21      u0068(.An(g), .B(i), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(j), .C(k), .Y(men_men_n98_));
  AOI220     u0070(.A0(men_men_n98_), .A1(men_men_n97_), .B0(men_men_n96_), .B1(men_men_n95_), .Y(men_men_n99_));
  NO2        u0071(.A(men_men_n99_), .B(f), .Y(men_men_n100_));
  NO4        u0072(.A(men_men_n100_), .B(men_men_n94_), .C(men_men_n91_), .D(men_men_n88_), .Y(men_men_n101_));
  NAi41      u0073(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n102_));
  AN2        u0074(.A(e), .B(b), .Y(men_men_n103_));
  NOi31      u0075(.An(c), .B(h), .C(f), .Y(men_men_n104_));
  NA2        u0076(.A(men_men_n104_), .B(men_men_n103_), .Y(men_men_n105_));
  NOi21      u0077(.An(i), .B(h), .Y(men_men_n106_));
  NA3        u0078(.A(men_men_n106_), .B(g), .C(men_men_n36_), .Y(men_men_n107_));
  INV        u0079(.A(a), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n103_), .B(men_men_n108_), .Y(men_men_n109_));
  INV        u0081(.A(l), .Y(men_men_n110_));
  NOi21      u0082(.An(m), .B(n), .Y(men_men_n111_));
  AN2        u0083(.A(k), .B(h), .Y(men_men_n112_));
  NO2        u0084(.A(men_men_n107_), .B(men_men_n84_), .Y(men_men_n113_));
  INV        u0085(.A(b), .Y(men_men_n114_));
  NA2        u0086(.A(l), .B(j), .Y(men_men_n115_));
  AN2        u0087(.A(k), .B(i), .Y(men_men_n116_));
  NA2        u0088(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NA2        u0089(.A(g), .B(e), .Y(men_men_n118_));
  NOi32      u0090(.An(c), .Bn(a), .C(d), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n111_), .Y(men_men_n120_));
  NO4        u0092(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n117_), .D(men_men_n114_), .Y(men_men_n121_));
  NO2        u0093(.A(men_men_n121_), .B(men_men_n113_), .Y(men_men_n122_));
  OAI210     u0094(.A0(men_men_n101_), .A1(men_men_n84_), .B0(men_men_n122_), .Y(men_men_n123_));
  NOi31      u0095(.An(k), .B(m), .C(j), .Y(men_men_n124_));
  NA3        u0096(.A(men_men_n124_), .B(men_men_n75_), .C(men_men_n74_), .Y(men_men_n125_));
  NOi31      u0097(.An(k), .B(m), .C(i), .Y(men_men_n126_));
  NA3        u0098(.A(men_men_n126_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n127_));
  NA2        u0099(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n128_));
  NOi32      u0100(.An(f), .Bn(b), .C(e), .Y(men_men_n129_));
  NAi21      u0101(.An(g), .B(h), .Y(men_men_n130_));
  NAi21      u0102(.An(m), .B(n), .Y(men_men_n131_));
  NAi21      u0103(.An(j), .B(k), .Y(men_men_n132_));
  NO3        u0104(.A(men_men_n132_), .B(men_men_n131_), .C(men_men_n130_), .Y(men_men_n133_));
  NAi41      u0105(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n134_));
  NAi31      u0106(.An(j), .B(k), .C(h), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n131_), .Y(men_men_n136_));
  AOI210     u0108(.A0(men_men_n133_), .A1(men_men_n129_), .B0(men_men_n136_), .Y(men_men_n137_));
  NO2        u0109(.A(k), .B(j), .Y(men_men_n138_));
  NO2        u0110(.A(men_men_n138_), .B(men_men_n131_), .Y(men_men_n139_));
  AN2        u0111(.A(k), .B(j), .Y(men_men_n140_));
  NAi21      u0112(.An(c), .B(b), .Y(men_men_n141_));
  NA2        u0113(.A(f), .B(d), .Y(men_men_n142_));
  NO3        u0114(.A(men_men_n142_), .B(men_men_n141_), .C(men_men_n130_), .Y(men_men_n143_));
  NA2        u0115(.A(h), .B(c), .Y(men_men_n144_));
  NAi31      u0116(.An(f), .B(e), .C(b), .Y(men_men_n145_));
  NA2        u0117(.A(men_men_n143_), .B(men_men_n139_), .Y(men_men_n146_));
  NA2        u0118(.A(d), .B(b), .Y(men_men_n147_));
  NAi21      u0119(.An(e), .B(f), .Y(men_men_n148_));
  NO2        u0120(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n149_));
  NA2        u0121(.A(b), .B(a), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(g), .Y(men_men_n151_));
  NAi21      u0123(.An(c), .B(d), .Y(men_men_n152_));
  NAi31      u0124(.An(l), .B(k), .C(h), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n131_), .B(men_men_n153_), .Y(men_men_n154_));
  NA2        u0126(.A(men_men_n154_), .B(men_men_n149_), .Y(men_men_n155_));
  NAi41      u0127(.An(men_men_n128_), .B(men_men_n155_), .C(men_men_n146_), .D(men_men_n137_), .Y(men_men_n156_));
  NAi31      u0128(.An(e), .B(f), .C(b), .Y(men_men_n157_));
  NOi21      u0129(.An(g), .B(d), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NOi21      u0131(.An(h), .B(i), .Y(men_men_n160_));
  NOi21      u0132(.An(k), .B(m), .Y(men_men_n161_));
  NA3        u0133(.A(men_men_n161_), .B(men_men_n160_), .C(n), .Y(men_men_n162_));
  NOi21      u0134(.An(men_men_n159_), .B(men_men_n162_), .Y(men_men_n163_));
  NOi21      u0135(.An(h), .B(g), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n142_), .B(men_men_n141_), .Y(men_men_n165_));
  NAi31      u0137(.An(l), .B(j), .C(h), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n166_), .B(men_men_n49_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n65_), .Y(men_men_n168_));
  NOi32      u0140(.An(n), .Bn(k), .C(m), .Y(men_men_n169_));
  NA2        u0141(.A(l), .B(i), .Y(men_men_n170_));
  INV        u0142(.A(men_men_n168_), .Y(men_men_n171_));
  NAi31      u0143(.An(d), .B(f), .C(c), .Y(men_men_n172_));
  NAi31      u0144(.An(e), .B(f), .C(c), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NA2        u0146(.A(j), .B(h), .Y(men_men_n175_));
  OR3        u0147(.A(n), .B(m), .C(k), .Y(men_men_n176_));
  NO2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  NAi32      u0149(.An(m), .Bn(k), .C(n), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n175_), .Y(men_men_n179_));
  AOI220     u0151(.A0(men_men_n179_), .A1(men_men_n159_), .B0(men_men_n177_), .B1(men_men_n174_), .Y(men_men_n180_));
  NO2        u0152(.A(n), .B(m), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n50_), .Y(men_men_n182_));
  NAi21      u0154(.An(f), .B(e), .Y(men_men_n183_));
  NA2        u0155(.A(d), .B(c), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NOi21      u0157(.An(men_men_n185_), .B(men_men_n182_), .Y(men_men_n186_));
  NAi31      u0158(.An(m), .B(n), .C(b), .Y(men_men_n187_));
  NAi21      u0159(.An(h), .B(f), .Y(men_men_n188_));
  NO2        u0160(.A(men_men_n187_), .B(men_men_n152_), .Y(men_men_n189_));
  NOi32      u0161(.An(f), .Bn(c), .C(d), .Y(men_men_n190_));
  NOi32      u0162(.An(f), .Bn(c), .C(e), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NO3        u0164(.A(n), .B(m), .C(j), .Y(men_men_n193_));
  NA2        u0165(.A(men_men_n193_), .B(men_men_n112_), .Y(men_men_n194_));
  AO210      u0166(.A0(men_men_n194_), .A1(men_men_n182_), .B0(men_men_n192_), .Y(men_men_n195_));
  NAi31      u0167(.An(men_men_n186_), .B(men_men_n195_), .C(men_men_n180_), .Y(men_men_n196_));
  OR4        u0168(.A(men_men_n196_), .B(men_men_n171_), .C(men_men_n163_), .D(men_men_n156_), .Y(men_men_n197_));
  NO4        u0169(.A(men_men_n197_), .B(men_men_n123_), .C(men_men_n81_), .D(men_men_n53_), .Y(men_men_n198_));
  NA3        u0170(.A(m), .B(men_men_n110_), .C(j), .Y(men_men_n199_));
  NAi31      u0171(.An(n), .B(h), .C(g), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n200_), .B(men_men_n199_), .Y(men_men_n201_));
  NOi32      u0173(.An(m), .Bn(k), .C(l), .Y(men_men_n202_));
  NA3        u0174(.A(men_men_n202_), .B(men_men_n85_), .C(g), .Y(men_men_n203_));
  NO2        u0175(.A(men_men_n203_), .B(n), .Y(men_men_n204_));
  NOi21      u0176(.An(k), .B(j), .Y(men_men_n205_));
  NA4        u0177(.A(men_men_n205_), .B(men_men_n111_), .C(i), .D(g), .Y(men_men_n206_));
  AN2        u0178(.A(i), .B(g), .Y(men_men_n207_));
  NA3        u0179(.A(men_men_n72_), .B(men_men_n207_), .C(men_men_n111_), .Y(men_men_n208_));
  NA2        u0180(.A(men_men_n208_), .B(men_men_n206_), .Y(men_men_n209_));
  NO3        u0181(.A(men_men_n209_), .B(men_men_n204_), .C(men_men_n201_), .Y(men_men_n210_));
  NAi41      u0182(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n211_));
  INV        u0183(.A(men_men_n211_), .Y(men_men_n212_));
  INV        u0184(.A(f), .Y(men_men_n213_));
  INV        u0185(.A(g), .Y(men_men_n214_));
  NOi31      u0186(.An(i), .B(j), .C(h), .Y(men_men_n215_));
  NOi21      u0187(.An(l), .B(m), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NO3        u0189(.A(men_men_n217_), .B(men_men_n214_), .C(men_men_n213_), .Y(men_men_n218_));
  NA2        u0190(.A(men_men_n218_), .B(men_men_n212_), .Y(men_men_n219_));
  OAI210     u0191(.A0(men_men_n210_), .A1(men_men_n32_), .B0(men_men_n219_), .Y(men_men_n220_));
  NOi21      u0192(.An(n), .B(m), .Y(men_men_n221_));
  NA2        u0193(.A(i), .B(men_men_n221_), .Y(men_men_n222_));
  OA220      u0194(.A0(men_men_n222_), .A1(men_men_n105_), .B0(men_men_n77_), .B1(men_men_n76_), .Y(men_men_n223_));
  NAi21      u0195(.An(j), .B(h), .Y(men_men_n224_));
  XN2        u0196(.A(i), .B(h), .Y(men_men_n225_));
  NOi31      u0197(.An(k), .B(n), .C(m), .Y(men_men_n226_));
  NAi31      u0198(.An(f), .B(e), .C(c), .Y(men_men_n227_));
  NO4        u0199(.A(men_men_n227_), .B(men_men_n176_), .C(men_men_n175_), .D(men_men_n57_), .Y(men_men_n228_));
  NA4        u0200(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n229_));
  NAi32      u0201(.An(m), .Bn(i), .C(k), .Y(men_men_n230_));
  NO3        u0202(.A(men_men_n230_), .B(men_men_n89_), .C(men_men_n229_), .Y(men_men_n231_));
  INV        u0203(.A(k), .Y(men_men_n232_));
  NO2        u0204(.A(men_men_n231_), .B(men_men_n228_), .Y(men_men_n233_));
  NAi21      u0205(.An(n), .B(a), .Y(men_men_n234_));
  NO2        u0206(.A(men_men_n234_), .B(men_men_n147_), .Y(men_men_n235_));
  NAi41      u0207(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n236_));
  NO2        u0208(.A(men_men_n236_), .B(e), .Y(men_men_n237_));
  NO3        u0209(.A(men_men_n148_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n238_));
  OAI210     u0210(.A0(men_men_n238_), .A1(men_men_n237_), .B0(men_men_n235_), .Y(men_men_n239_));
  AN3        u0211(.A(men_men_n239_), .B(men_men_n233_), .C(men_men_n223_), .Y(men_men_n240_));
  OR2        u0212(.A(h), .B(g), .Y(men_men_n241_));
  NAi41      u0213(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n242_), .B(men_men_n213_), .Y(men_men_n243_));
  NA2        u0215(.A(men_men_n161_), .B(men_men_n106_), .Y(men_men_n244_));
  NAi21      u0216(.An(men_men_n244_), .B(men_men_n243_), .Y(men_men_n245_));
  NO2        u0217(.A(n), .B(a), .Y(men_men_n246_));
  NAi21      u0218(.An(h), .B(i), .Y(men_men_n247_));
  NA2        u0219(.A(men_men_n181_), .B(k), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n248_), .B(men_men_n247_), .Y(men_men_n249_));
  INV        u0221(.A(men_men_n245_), .Y(men_men_n250_));
  NOi21      u0222(.An(g), .B(e), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n70_), .B(men_men_n71_), .Y(men_men_n252_));
  NOi32      u0224(.An(l), .Bn(j), .C(i), .Y(men_men_n253_));
  AOI210     u0225(.A0(men_men_n72_), .A1(men_men_n85_), .B0(men_men_n253_), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n247_), .B(men_men_n44_), .Y(men_men_n255_));
  NAi21      u0227(.An(f), .B(g), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n63_), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n67_), .B(men_men_n115_), .Y(men_men_n258_));
  AOI220     u0230(.A0(men_men_n258_), .A1(men_men_n257_), .B0(men_men_n255_), .B1(men_men_n65_), .Y(men_men_n259_));
  INV        u0231(.A(men_men_n259_), .Y(men_men_n260_));
  NO3        u0232(.A(men_men_n132_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n261_));
  NOi41      u0233(.An(men_men_n240_), .B(men_men_n260_), .C(men_men_n250_), .D(men_men_n220_), .Y(men_men_n262_));
  NO4        u0234(.A(men_men_n201_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n263_), .B(men_men_n109_), .Y(men_men_n264_));
  NA3        u0236(.A(men_men_n57_), .B(c), .C(b), .Y(men_men_n265_));
  NAi21      u0237(.An(h), .B(g), .Y(men_men_n266_));
  OR4        u0238(.A(men_men_n266_), .B(men_men_n265_), .C(men_men_n222_), .D(e), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n244_), .B(men_men_n256_), .Y(men_men_n268_));
  NAi31      u0240(.An(g), .B(k), .C(h), .Y(men_men_n269_));
  NO3        u0241(.A(men_men_n131_), .B(men_men_n269_), .C(l), .Y(men_men_n270_));
  NAi31      u0242(.An(e), .B(d), .C(a), .Y(men_men_n271_));
  NA2        u0243(.A(men_men_n270_), .B(men_men_n129_), .Y(men_men_n272_));
  NA2        u0244(.A(men_men_n272_), .B(men_men_n267_), .Y(men_men_n273_));
  NA4        u0245(.A(men_men_n161_), .B(men_men_n78_), .C(men_men_n74_), .D(men_men_n115_), .Y(men_men_n274_));
  NA3        u0246(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n82_), .Y(men_men_n275_));
  NA3        u0247(.A(e), .B(c), .C(b), .Y(men_men_n276_));
  NO2        u0248(.A(men_men_n58_), .B(men_men_n276_), .Y(men_men_n277_));
  NAi32      u0249(.An(k), .Bn(i), .C(j), .Y(men_men_n278_));
  NAi31      u0250(.An(h), .B(l), .C(i), .Y(men_men_n279_));
  NA3        u0251(.A(men_men_n279_), .B(men_men_n278_), .C(men_men_n166_), .Y(men_men_n280_));
  NOi21      u0252(.An(men_men_n280_), .B(men_men_n49_), .Y(men_men_n281_));
  OAI210     u0253(.A0(men_men_n257_), .A1(men_men_n277_), .B0(men_men_n281_), .Y(men_men_n282_));
  NAi21      u0254(.An(l), .B(k), .Y(men_men_n283_));
  NO2        u0255(.A(men_men_n283_), .B(men_men_n49_), .Y(men_men_n284_));
  NOi21      u0256(.An(l), .B(j), .Y(men_men_n285_));
  NA2        u0257(.A(men_men_n164_), .B(men_men_n285_), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n116_), .B(men_men_n115_), .C(g), .Y(men_men_n287_));
  OR3        u0259(.A(men_men_n70_), .B(men_men_n71_), .C(e), .Y(men_men_n288_));
  AOI210     u0260(.A0(men_men_n287_), .A1(men_men_n286_), .B0(men_men_n288_), .Y(men_men_n289_));
  INV        u0261(.A(men_men_n289_), .Y(men_men_n290_));
  NAi32      u0262(.An(j), .Bn(h), .C(i), .Y(men_men_n291_));
  NAi21      u0263(.An(m), .B(l), .Y(men_men_n292_));
  NO3        u0264(.A(men_men_n292_), .B(men_men_n291_), .C(men_men_n82_), .Y(men_men_n293_));
  NA2        u0265(.A(h), .B(g), .Y(men_men_n294_));
  NA2        u0266(.A(men_men_n169_), .B(men_men_n45_), .Y(men_men_n295_));
  NO2        u0267(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n296_));
  OAI210     u0268(.A0(men_men_n296_), .A1(men_men_n293_), .B0(men_men_n165_), .Y(men_men_n297_));
  NA4        u0269(.A(men_men_n297_), .B(men_men_n290_), .C(men_men_n282_), .D(men_men_n274_), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n145_), .B(d), .Y(men_men_n299_));
  NAi32      u0271(.An(n), .Bn(m), .C(l), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n300_), .B(men_men_n291_), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n301_), .B(men_men_n185_), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n120_), .B(men_men_n114_), .Y(men_men_n303_));
  NAi31      u0275(.An(k), .B(l), .C(j), .Y(men_men_n304_));
  OAI210     u0276(.A0(men_men_n283_), .A1(j), .B0(men_men_n304_), .Y(men_men_n305_));
  NOi21      u0277(.An(men_men_n305_), .B(men_men_n118_), .Y(men_men_n306_));
  NA2        u0278(.A(men_men_n306_), .B(men_men_n303_), .Y(men_men_n307_));
  NA2        u0279(.A(men_men_n307_), .B(men_men_n302_), .Y(men_men_n308_));
  NO4        u0280(.A(men_men_n308_), .B(men_men_n298_), .C(men_men_n273_), .D(men_men_n264_), .Y(men_men_n309_));
  NAi21      u0281(.An(m), .B(k), .Y(men_men_n310_));
  NO2        u0282(.A(men_men_n225_), .B(men_men_n310_), .Y(men_men_n311_));
  NAi41      u0283(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n312_));
  NO4        u0284(.A(i), .B(men_men_n151_), .C(men_men_n70_), .D(men_men_n71_), .Y(men_men_n313_));
  NA2        u0285(.A(e), .B(c), .Y(men_men_n314_));
  NO3        u0286(.A(men_men_n314_), .B(n), .C(d), .Y(men_men_n315_));
  NAi31      u0287(.An(d), .B(e), .C(b), .Y(men_men_n316_));
  NO2        u0288(.A(men_men_n131_), .B(men_men_n316_), .Y(men_men_n317_));
  NO4        u0289(.A(men_men_n312_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n214_), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n246_), .B(men_men_n103_), .Y(men_men_n319_));
  NOi31      u0291(.An(l), .B(n), .C(m), .Y(men_men_n320_));
  NA2        u0292(.A(men_men_n320_), .B(men_men_n215_), .Y(men_men_n321_));
  NO2        u0293(.A(men_men_n321_), .B(men_men_n192_), .Y(men_men_n322_));
  OR2        u0294(.A(men_men_n322_), .B(men_men_n318_), .Y(men_men_n323_));
  NAi32      u0295(.An(m), .Bn(j), .C(k), .Y(men_men_n324_));
  NAi41      u0296(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n325_));
  NOi31      u0297(.An(j), .B(m), .C(k), .Y(men_men_n326_));
  NO2        u0298(.A(men_men_n124_), .B(men_men_n326_), .Y(men_men_n327_));
  AN3        u0299(.A(h), .B(g), .C(f), .Y(men_men_n328_));
  NOi32      u0300(.An(m), .Bn(j), .C(l), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n329_), .B(men_men_n96_), .Y(men_men_n330_));
  NAi32      u0302(.An(men_men_n330_), .Bn(men_men_n200_), .C(men_men_n299_), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n292_), .B(men_men_n291_), .Y(men_men_n332_));
  NO2        u0304(.A(men_men_n217_), .B(g), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n157_), .B(men_men_n82_), .Y(men_men_n334_));
  AOI220     u0306(.A0(men_men_n334_), .A1(men_men_n333_), .B0(men_men_n243_), .B1(men_men_n332_), .Y(men_men_n335_));
  INV        u0307(.A(men_men_n230_), .Y(men_men_n336_));
  NA3        u0308(.A(men_men_n336_), .B(men_men_n328_), .C(men_men_n212_), .Y(men_men_n337_));
  NA3        u0309(.A(men_men_n337_), .B(men_men_n335_), .C(men_men_n331_), .Y(men_men_n338_));
  NA3        u0310(.A(h), .B(g), .C(f), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n339_), .B(men_men_n73_), .Y(men_men_n340_));
  NA2        u0312(.A(men_men_n325_), .B(men_men_n211_), .Y(men_men_n341_));
  NA2        u0313(.A(men_men_n164_), .B(e), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n342_), .B(men_men_n41_), .Y(men_men_n343_));
  AOI220     u0315(.A0(men_men_n343_), .A1(men_men_n303_), .B0(men_men_n341_), .B1(men_men_n340_), .Y(men_men_n344_));
  NOi32      u0316(.An(j), .Bn(g), .C(i), .Y(men_men_n345_));
  NA3        u0317(.A(men_men_n345_), .B(men_men_n283_), .C(men_men_n111_), .Y(men_men_n346_));
  AO210      u0318(.A0(men_men_n109_), .A1(men_men_n32_), .B0(men_men_n346_), .Y(men_men_n347_));
  NOi32      u0319(.An(e), .Bn(b), .C(a), .Y(men_men_n348_));
  INV        u0320(.A(men_men_n310_), .Y(men_men_n349_));
  NO3        u0321(.A(men_men_n312_), .B(men_men_n69_), .C(men_men_n214_), .Y(men_men_n350_));
  NA3        u0322(.A(men_men_n208_), .B(men_men_n206_), .C(men_men_n35_), .Y(men_men_n351_));
  AOI220     u0323(.A0(men_men_n351_), .A1(men_men_n348_), .B0(men_men_n350_), .B1(men_men_n349_), .Y(men_men_n352_));
  NO2        u0324(.A(men_men_n316_), .B(n), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n207_), .B(k), .Y(men_men_n354_));
  NA3        u0326(.A(m), .B(men_men_n110_), .C(men_men_n213_), .Y(men_men_n355_));
  NA4        u0327(.A(men_men_n202_), .B(men_men_n85_), .C(g), .D(men_men_n213_), .Y(men_men_n356_));
  OAI210     u0328(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n356_), .Y(men_men_n357_));
  NAi41      u0329(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n358_));
  NA2        u0330(.A(men_men_n51_), .B(men_men_n111_), .Y(men_men_n359_));
  NO2        u0331(.A(men_men_n359_), .B(men_men_n358_), .Y(men_men_n360_));
  AOI220     u0332(.A0(men_men_n360_), .A1(b), .B0(men_men_n357_), .B1(men_men_n353_), .Y(men_men_n361_));
  NA4        u0333(.A(men_men_n361_), .B(men_men_n352_), .C(men_men_n347_), .D(men_men_n344_), .Y(men_men_n362_));
  NO4        u0334(.A(men_men_n362_), .B(men_men_n338_), .C(men_men_n323_), .D(men_men_n313_), .Y(men_men_n363_));
  NA4        u0335(.A(men_men_n363_), .B(men_men_n309_), .C(men_men_n262_), .D(men_men_n198_), .Y(men10));
  NA3        u0336(.A(m), .B(k), .C(i), .Y(men_men_n365_));
  NO3        u0337(.A(men_men_n365_), .B(j), .C(men_men_n214_), .Y(men_men_n366_));
  NOi21      u0338(.An(e), .B(f), .Y(men_men_n367_));
  NO4        u0339(.A(men_men_n152_), .B(men_men_n367_), .C(n), .D(men_men_n108_), .Y(men_men_n368_));
  NAi31      u0340(.An(b), .B(f), .C(c), .Y(men_men_n369_));
  INV        u0341(.A(men_men_n369_), .Y(men_men_n370_));
  NOi32      u0342(.An(k), .Bn(h), .C(j), .Y(men_men_n371_));
  NA2        u0343(.A(men_men_n371_), .B(men_men_n221_), .Y(men_men_n372_));
  NA2        u0344(.A(men_men_n162_), .B(men_men_n372_), .Y(men_men_n373_));
  AOI220     u0345(.A0(men_men_n373_), .A1(men_men_n370_), .B0(men_men_n368_), .B1(men_men_n366_), .Y(men_men_n374_));
  AN2        u0346(.A(j), .B(h), .Y(men_men_n375_));
  NO3        u0347(.A(n), .B(m), .C(k), .Y(men_men_n376_));
  NA2        u0348(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n377_));
  NO3        u0349(.A(men_men_n377_), .B(men_men_n152_), .C(men_men_n213_), .Y(men_men_n378_));
  OR2        u0350(.A(m), .B(k), .Y(men_men_n379_));
  NO2        u0351(.A(men_men_n175_), .B(men_men_n379_), .Y(men_men_n380_));
  NA4        u0352(.A(n), .B(f), .C(c), .D(men_men_n114_), .Y(men_men_n381_));
  NOi21      u0353(.An(men_men_n380_), .B(men_men_n381_), .Y(men_men_n382_));
  NOi32      u0354(.An(d), .Bn(a), .C(c), .Y(men_men_n383_));
  NA2        u0355(.A(men_men_n383_), .B(men_men_n183_), .Y(men_men_n384_));
  NAi21      u0356(.An(i), .B(g), .Y(men_men_n385_));
  NAi31      u0357(.An(k), .B(m), .C(j), .Y(men_men_n386_));
  NO3        u0358(.A(men_men_n386_), .B(men_men_n385_), .C(n), .Y(men_men_n387_));
  NOi21      u0359(.An(men_men_n387_), .B(men_men_n384_), .Y(men_men_n388_));
  NO3        u0360(.A(men_men_n388_), .B(men_men_n382_), .C(men_men_n378_), .Y(men_men_n389_));
  NO2        u0361(.A(men_men_n381_), .B(men_men_n292_), .Y(men_men_n390_));
  NOi32      u0362(.An(f), .Bn(d), .C(c), .Y(men_men_n391_));
  AOI220     u0363(.A0(men_men_n391_), .A1(men_men_n301_), .B0(men_men_n390_), .B1(men_men_n215_), .Y(men_men_n392_));
  NA3        u0364(.A(men_men_n392_), .B(men_men_n389_), .C(men_men_n374_), .Y(men_men_n393_));
  NO2        u0365(.A(men_men_n57_), .B(men_men_n114_), .Y(men_men_n394_));
  NA2        u0366(.A(men_men_n246_), .B(men_men_n394_), .Y(men_men_n395_));
  INV        u0367(.A(e), .Y(men_men_n396_));
  NA2        u0368(.A(men_men_n46_), .B(e), .Y(men_men_n397_));
  OAI220     u0369(.A0(men_men_n397_), .A1(men_men_n199_), .B0(men_men_n203_), .B1(men_men_n396_), .Y(men_men_n398_));
  AN2        u0370(.A(g), .B(e), .Y(men_men_n399_));
  NA3        u0371(.A(men_men_n399_), .B(men_men_n202_), .C(i), .Y(men_men_n400_));
  NA2        u0372(.A(men_men_n87_), .B(men_men_n400_), .Y(men_men_n401_));
  NO2        u0373(.A(men_men_n401_), .B(men_men_n398_), .Y(men_men_n402_));
  NOi32      u0374(.An(h), .Bn(e), .C(g), .Y(men_men_n403_));
  NA3        u0375(.A(men_men_n403_), .B(men_men_n285_), .C(m), .Y(men_men_n404_));
  NOi21      u0376(.An(g), .B(h), .Y(men_men_n405_));
  AN3        u0377(.A(m), .B(l), .C(i), .Y(men_men_n406_));
  AN3        u0378(.A(h), .B(g), .C(e), .Y(men_men_n407_));
  NA2        u0379(.A(men_men_n407_), .B(men_men_n96_), .Y(men_men_n408_));
  AOI210     u0380(.A0(men_men_n404_), .A1(men_men_n402_), .B0(men_men_n395_), .Y(men_men_n409_));
  NA3        u0381(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n410_));
  NO2        u0382(.A(men_men_n410_), .B(men_men_n395_), .Y(men_men_n411_));
  NA3        u0383(.A(men_men_n383_), .B(men_men_n183_), .C(men_men_n82_), .Y(men_men_n412_));
  NAi31      u0384(.An(b), .B(c), .C(a), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n413_), .B(n), .Y(men_men_n414_));
  OAI210     u0386(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n415_));
  NO2        u0387(.A(men_men_n415_), .B(men_men_n148_), .Y(men_men_n416_));
  NO3        u0388(.A(men_men_n411_), .B(men_men_n409_), .C(men_men_n393_), .Y(men_men_n417_));
  NA2        u0389(.A(i), .B(g), .Y(men_men_n418_));
  NO3        u0390(.A(men_men_n271_), .B(men_men_n418_), .C(c), .Y(men_men_n419_));
  NOi21      u0391(.An(a), .B(n), .Y(men_men_n420_));
  NOi21      u0392(.An(d), .B(c), .Y(men_men_n421_));
  NA2        u0393(.A(men_men_n421_), .B(men_men_n420_), .Y(men_men_n422_));
  NA3        u0394(.A(i), .B(g), .C(f), .Y(men_men_n423_));
  OR2        u0395(.A(men_men_n423_), .B(men_men_n68_), .Y(men_men_n424_));
  NA3        u0396(.A(men_men_n406_), .B(men_men_n405_), .C(men_men_n183_), .Y(men_men_n425_));
  AOI210     u0397(.A0(men_men_n425_), .A1(men_men_n424_), .B0(men_men_n422_), .Y(men_men_n426_));
  AOI210     u0398(.A0(men_men_n419_), .A1(men_men_n284_), .B0(men_men_n426_), .Y(men_men_n427_));
  OR2        u0399(.A(n), .B(m), .Y(men_men_n428_));
  NO2        u0400(.A(men_men_n428_), .B(men_men_n153_), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n184_), .B(men_men_n148_), .Y(men_men_n430_));
  OAI210     u0402(.A0(men_men_n429_), .A1(men_men_n177_), .B0(men_men_n430_), .Y(men_men_n431_));
  NO2        u0403(.A(men_men_n413_), .B(men_men_n49_), .Y(men_men_n432_));
  NO3        u0404(.A(men_men_n64_), .B(men_men_n110_), .C(e), .Y(men_men_n433_));
  NAi21      u0405(.An(k), .B(j), .Y(men_men_n434_));
  NA2        u0406(.A(men_men_n433_), .B(men_men_n432_), .Y(men_men_n435_));
  NAi21      u0407(.An(e), .B(d), .Y(men_men_n436_));
  INV        u0408(.A(men_men_n436_), .Y(men_men_n437_));
  NO2        u0409(.A(men_men_n248_), .B(men_men_n213_), .Y(men_men_n438_));
  NA2        u0410(.A(men_men_n435_), .B(men_men_n431_), .Y(men_men_n439_));
  NO2        u0411(.A(men_men_n321_), .B(men_men_n213_), .Y(men_men_n440_));
  NA2        u0412(.A(men_men_n440_), .B(men_men_n437_), .Y(men_men_n441_));
  NOi31      u0413(.An(n), .B(m), .C(k), .Y(men_men_n442_));
  AOI220     u0414(.A0(men_men_n442_), .A1(men_men_n375_), .B0(men_men_n221_), .B1(men_men_n50_), .Y(men_men_n443_));
  NAi31      u0415(.An(g), .B(f), .C(c), .Y(men_men_n444_));
  OR3        u0416(.A(men_men_n444_), .B(men_men_n443_), .C(e), .Y(men_men_n445_));
  NA3        u0417(.A(men_men_n445_), .B(men_men_n441_), .C(men_men_n302_), .Y(men_men_n446_));
  NOi41      u0418(.An(men_men_n427_), .B(men_men_n446_), .C(men_men_n439_), .D(men_men_n260_), .Y(men_men_n447_));
  NOi32      u0419(.An(c), .Bn(a), .C(b), .Y(men_men_n448_));
  NA2        u0420(.A(men_men_n448_), .B(men_men_n111_), .Y(men_men_n449_));
  INV        u0421(.A(men_men_n269_), .Y(men_men_n450_));
  AN2        u0422(.A(e), .B(d), .Y(men_men_n451_));
  NA2        u0423(.A(men_men_n451_), .B(men_men_n450_), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n148_), .Y(men_men_n453_));
  NO2        u0425(.A(men_men_n130_), .B(men_men_n41_), .Y(men_men_n454_));
  NO2        u0426(.A(men_men_n64_), .B(e), .Y(men_men_n455_));
  NOi31      u0427(.An(j), .B(k), .C(i), .Y(men_men_n456_));
  NOi21      u0428(.An(men_men_n166_), .B(men_men_n456_), .Y(men_men_n457_));
  INV        u0429(.A(men_men_n457_), .Y(men_men_n458_));
  NA2        u0430(.A(men_men_n458_), .B(men_men_n455_), .Y(men_men_n459_));
  AOI210     u0431(.A0(men_men_n459_), .A1(men_men_n452_), .B0(men_men_n449_), .Y(men_men_n460_));
  NO2        u0432(.A(men_men_n209_), .B(men_men_n204_), .Y(men_men_n461_));
  NOi21      u0433(.An(a), .B(b), .Y(men_men_n462_));
  NA3        u0434(.A(e), .B(d), .C(c), .Y(men_men_n463_));
  NAi21      u0435(.An(men_men_n463_), .B(men_men_n462_), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n412_), .B(men_men_n203_), .Y(men_men_n465_));
  NOi21      u0437(.An(men_men_n464_), .B(men_men_n465_), .Y(men_men_n466_));
  AOI210     u0438(.A0(men_men_n263_), .A1(men_men_n461_), .B0(men_men_n466_), .Y(men_men_n467_));
  NO4        u0439(.A(men_men_n188_), .B(men_men_n102_), .C(men_men_n54_), .D(b), .Y(men_men_n468_));
  NA2        u0440(.A(men_men_n370_), .B(men_men_n154_), .Y(men_men_n469_));
  OR2        u0441(.A(k), .B(j), .Y(men_men_n470_));
  NA2        u0442(.A(l), .B(k), .Y(men_men_n471_));
  NA3        u0443(.A(men_men_n471_), .B(men_men_n470_), .C(men_men_n221_), .Y(men_men_n472_));
  AOI210     u0444(.A0(men_men_n230_), .A1(men_men_n324_), .B0(men_men_n82_), .Y(men_men_n473_));
  NOi21      u0445(.An(men_men_n472_), .B(men_men_n473_), .Y(men_men_n474_));
  OR3        u0446(.A(men_men_n474_), .B(men_men_n144_), .C(men_men_n134_), .Y(men_men_n475_));
  NA3        u0447(.A(men_men_n274_), .B(men_men_n127_), .C(men_men_n125_), .Y(men_men_n476_));
  NA2        u0448(.A(men_men_n383_), .B(men_men_n111_), .Y(men_men_n477_));
  NO4        u0449(.A(men_men_n477_), .B(men_men_n93_), .C(men_men_n110_), .D(e), .Y(men_men_n478_));
  NO3        u0450(.A(men_men_n412_), .B(men_men_n90_), .C(men_men_n130_), .Y(men_men_n479_));
  NO4        u0451(.A(men_men_n479_), .B(men_men_n478_), .C(men_men_n476_), .D(men_men_n313_), .Y(men_men_n480_));
  NA3        u0452(.A(men_men_n480_), .B(men_men_n475_), .C(men_men_n469_), .Y(men_men_n481_));
  NO4        u0453(.A(men_men_n481_), .B(men_men_n468_), .C(men_men_n467_), .D(men_men_n460_), .Y(men_men_n482_));
  NOi21      u0454(.An(d), .B(e), .Y(men_men_n483_));
  NO2        u0455(.A(men_men_n188_), .B(men_men_n54_), .Y(men_men_n484_));
  NAi31      u0456(.An(j), .B(l), .C(i), .Y(men_men_n485_));
  OAI210     u0457(.A0(men_men_n485_), .A1(men_men_n131_), .B0(men_men_n102_), .Y(men_men_n486_));
  NA3        u0458(.A(men_men_n486_), .B(men_men_n484_), .C(men_men_n483_), .Y(men_men_n487_));
  NO3        u0459(.A(men_men_n384_), .B(men_men_n330_), .C(men_men_n200_), .Y(men_men_n488_));
  NO2        u0460(.A(men_men_n488_), .B(men_men_n186_), .Y(men_men_n489_));
  NA3        u0461(.A(men_men_n489_), .B(men_men_n487_), .C(men_men_n240_), .Y(men_men_n490_));
  OAI210     u0462(.A0(men_men_n126_), .A1(men_men_n124_), .B0(n), .Y(men_men_n491_));
  NO2        u0463(.A(men_men_n491_), .B(men_men_n130_), .Y(men_men_n492_));
  OA210      u0464(.A0(men_men_n293_), .A1(men_men_n492_), .B0(men_men_n191_), .Y(men_men_n493_));
  XO2        u0465(.A(i), .B(h), .Y(men_men_n494_));
  NA3        u0466(.A(men_men_n494_), .B(men_men_n161_), .C(n), .Y(men_men_n495_));
  NAi41      u0467(.An(men_men_n293_), .B(men_men_n495_), .C(men_men_n443_), .D(men_men_n372_), .Y(men_men_n496_));
  NOi32      u0468(.An(men_men_n496_), .Bn(men_men_n455_), .C(men_men_n265_), .Y(men_men_n497_));
  NAi31      u0469(.An(c), .B(f), .C(d), .Y(men_men_n498_));
  AOI210     u0470(.A0(men_men_n275_), .A1(men_men_n194_), .B0(men_men_n498_), .Y(men_men_n499_));
  NOi21      u0471(.An(men_men_n80_), .B(men_men_n499_), .Y(men_men_n500_));
  NA3        u0472(.A(men_men_n368_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n501_));
  NA2        u0473(.A(men_men_n226_), .B(men_men_n106_), .Y(men_men_n502_));
  NO2        u0474(.A(men_men_n182_), .B(men_men_n498_), .Y(men_men_n503_));
  AOI210     u0475(.A0(men_men_n346_), .A1(men_men_n35_), .B0(men_men_n464_), .Y(men_men_n504_));
  NOi31      u0476(.An(men_men_n501_), .B(men_men_n504_), .C(men_men_n503_), .Y(men_men_n505_));
  AO220      u0477(.A0(men_men_n281_), .A1(men_men_n257_), .B0(men_men_n167_), .B1(men_men_n65_), .Y(men_men_n506_));
  NA3        u0478(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n507_));
  NO2        u0479(.A(men_men_n507_), .B(men_men_n422_), .Y(men_men_n508_));
  NO2        u0480(.A(men_men_n508_), .B(men_men_n289_), .Y(men_men_n509_));
  NAi41      u0481(.An(men_men_n506_), .B(men_men_n509_), .C(men_men_n505_), .D(men_men_n500_), .Y(men_men_n510_));
  NO4        u0482(.A(men_men_n510_), .B(men_men_n497_), .C(men_men_n493_), .D(men_men_n490_), .Y(men_men_n511_));
  NA4        u0483(.A(men_men_n511_), .B(men_men_n482_), .C(men_men_n447_), .D(men_men_n417_), .Y(men11));
  NO2        u0484(.A(men_men_n70_), .B(f), .Y(men_men_n513_));
  NA2        u0485(.A(j), .B(g), .Y(men_men_n514_));
  NAi31      u0486(.An(i), .B(m), .C(l), .Y(men_men_n515_));
  NA3        u0487(.A(m), .B(k), .C(j), .Y(men_men_n516_));
  OAI220     u0488(.A0(men_men_n516_), .A1(men_men_n130_), .B0(men_men_n515_), .B1(men_men_n514_), .Y(men_men_n517_));
  NA2        u0489(.A(men_men_n517_), .B(men_men_n513_), .Y(men_men_n518_));
  NOi32      u0490(.An(e), .Bn(b), .C(f), .Y(men_men_n519_));
  NA2        u0491(.A(men_men_n253_), .B(men_men_n111_), .Y(men_men_n520_));
  NA2        u0492(.A(men_men_n46_), .B(j), .Y(men_men_n521_));
  NO2        u0493(.A(men_men_n521_), .B(men_men_n295_), .Y(men_men_n522_));
  NAi31      u0494(.An(d), .B(e), .C(a), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n523_), .B(n), .Y(men_men_n524_));
  AOI220     u0496(.A0(men_men_n524_), .A1(men_men_n100_), .B0(men_men_n522_), .B1(men_men_n519_), .Y(men_men_n525_));
  NAi41      u0497(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n526_));
  AN2        u0498(.A(men_men_n526_), .B(men_men_n358_), .Y(men_men_n527_));
  AOI210     u0499(.A0(men_men_n527_), .A1(men_men_n384_), .B0(men_men_n266_), .Y(men_men_n528_));
  NA2        u0500(.A(j), .B(i), .Y(men_men_n529_));
  NAi31      u0501(.An(n), .B(m), .C(k), .Y(men_men_n530_));
  NO3        u0502(.A(men_men_n530_), .B(men_men_n529_), .C(men_men_n110_), .Y(men_men_n531_));
  NO4        u0503(.A(n), .B(d), .C(men_men_n114_), .D(a), .Y(men_men_n532_));
  OR2        u0504(.A(n), .B(c), .Y(men_men_n533_));
  NO2        u0505(.A(men_men_n533_), .B(men_men_n150_), .Y(men_men_n534_));
  NO2        u0506(.A(men_men_n534_), .B(men_men_n532_), .Y(men_men_n535_));
  NOi32      u0507(.An(g), .Bn(f), .C(i), .Y(men_men_n536_));
  AOI220     u0508(.A0(men_men_n536_), .A1(men_men_n98_), .B0(men_men_n517_), .B1(f), .Y(men_men_n537_));
  NO2        u0509(.A(men_men_n269_), .B(men_men_n49_), .Y(men_men_n538_));
  NO2        u0510(.A(men_men_n537_), .B(men_men_n535_), .Y(men_men_n539_));
  AOI210     u0511(.A0(men_men_n531_), .A1(men_men_n528_), .B0(men_men_n539_), .Y(men_men_n540_));
  NA2        u0512(.A(men_men_n140_), .B(men_men_n34_), .Y(men_men_n541_));
  OAI220     u0513(.A0(men_men_n541_), .A1(m), .B0(men_men_n521_), .B1(men_men_n230_), .Y(men_men_n542_));
  NOi41      u0514(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n543_));
  NAi32      u0515(.An(e), .Bn(b), .C(c), .Y(men_men_n544_));
  OR2        u0516(.A(men_men_n544_), .B(men_men_n82_), .Y(men_men_n545_));
  AN2        u0517(.A(men_men_n325_), .B(men_men_n312_), .Y(men_men_n546_));
  NA2        u0518(.A(men_men_n546_), .B(men_men_n545_), .Y(men_men_n547_));
  AN2        u0519(.A(men_men_n547_), .B(men_men_n542_), .Y(men_men_n548_));
  OAI220     u0520(.A0(men_men_n386_), .A1(men_men_n385_), .B0(men_men_n515_), .B1(men_men_n514_), .Y(men_men_n549_));
  NAi31      u0521(.An(d), .B(c), .C(a), .Y(men_men_n550_));
  NO2        u0522(.A(men_men_n550_), .B(n), .Y(men_men_n551_));
  NA3        u0523(.A(men_men_n551_), .B(men_men_n549_), .C(e), .Y(men_men_n552_));
  NO3        u0524(.A(men_men_n60_), .B(men_men_n49_), .C(men_men_n214_), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n227_), .B(men_men_n108_), .Y(men_men_n554_));
  OAI210     u0526(.A0(men_men_n553_), .A1(men_men_n387_), .B0(men_men_n554_), .Y(men_men_n555_));
  NA2        u0527(.A(men_men_n555_), .B(men_men_n552_), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n271_), .B(n), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n414_), .B(men_men_n557_), .Y(men_men_n558_));
  NA2        u0530(.A(men_men_n549_), .B(f), .Y(men_men_n559_));
  NAi32      u0531(.An(d), .Bn(a), .C(b), .Y(men_men_n560_));
  NO2        u0532(.A(men_men_n560_), .B(men_men_n49_), .Y(men_men_n561_));
  NA2        u0533(.A(h), .B(f), .Y(men_men_n562_));
  NO2        u0534(.A(men_men_n562_), .B(men_men_n93_), .Y(men_men_n563_));
  NO3        u0535(.A(men_men_n178_), .B(men_men_n175_), .C(g), .Y(men_men_n564_));
  AOI220     u0536(.A0(men_men_n564_), .A1(men_men_n56_), .B0(men_men_n563_), .B1(men_men_n561_), .Y(men_men_n565_));
  OAI210     u0537(.A0(men_men_n559_), .A1(men_men_n558_), .B0(men_men_n565_), .Y(men_men_n566_));
  AN3        u0538(.A(j), .B(h), .C(g), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n147_), .B(c), .Y(men_men_n568_));
  NA3        u0540(.A(men_men_n568_), .B(men_men_n567_), .C(men_men_n442_), .Y(men_men_n569_));
  NA3        u0541(.A(f), .B(d), .C(b), .Y(men_men_n570_));
  NO4        u0542(.A(men_men_n570_), .B(men_men_n178_), .C(men_men_n175_), .D(g), .Y(men_men_n571_));
  NAi21      u0543(.An(men_men_n571_), .B(men_men_n569_), .Y(men_men_n572_));
  NO4        u0544(.A(men_men_n572_), .B(men_men_n566_), .C(men_men_n556_), .D(men_men_n548_), .Y(men_men_n573_));
  AN4        u0545(.A(men_men_n573_), .B(men_men_n540_), .C(men_men_n525_), .D(men_men_n518_), .Y(men_men_n574_));
  INV        u0546(.A(k), .Y(men_men_n575_));
  NA3        u0547(.A(l), .B(men_men_n575_), .C(i), .Y(men_men_n576_));
  INV        u0548(.A(men_men_n576_), .Y(men_men_n577_));
  NA4        u0549(.A(men_men_n383_), .B(men_men_n405_), .C(men_men_n183_), .D(men_men_n111_), .Y(men_men_n578_));
  NAi32      u0550(.An(h), .Bn(f), .C(g), .Y(men_men_n579_));
  NAi41      u0551(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n580_));
  OAI210     u0552(.A0(men_men_n523_), .A1(n), .B0(men_men_n580_), .Y(men_men_n581_));
  NA2        u0553(.A(men_men_n581_), .B(m), .Y(men_men_n582_));
  NAi31      u0554(.An(h), .B(g), .C(f), .Y(men_men_n583_));
  OR3        u0555(.A(men_men_n583_), .B(men_men_n271_), .C(men_men_n49_), .Y(men_men_n584_));
  NA4        u0556(.A(men_men_n405_), .B(men_men_n119_), .C(men_men_n111_), .D(e), .Y(men_men_n585_));
  AN2        u0557(.A(men_men_n585_), .B(men_men_n584_), .Y(men_men_n586_));
  OA210      u0558(.A0(men_men_n582_), .A1(men_men_n579_), .B0(men_men_n586_), .Y(men_men_n587_));
  NO3        u0559(.A(men_men_n579_), .B(men_men_n70_), .C(men_men_n71_), .Y(men_men_n588_));
  NO4        u0560(.A(men_men_n583_), .B(men_men_n533_), .C(men_men_n150_), .D(men_men_n71_), .Y(men_men_n589_));
  OR2        u0561(.A(men_men_n589_), .B(men_men_n588_), .Y(men_men_n590_));
  NAi31      u0562(.An(men_men_n590_), .B(men_men_n587_), .C(men_men_n578_), .Y(men_men_n591_));
  NAi31      u0563(.An(f), .B(h), .C(g), .Y(men_men_n592_));
  NO4        u0564(.A(men_men_n304_), .B(men_men_n592_), .C(men_men_n70_), .D(men_men_n71_), .Y(men_men_n593_));
  NOi32      u0565(.An(b), .Bn(a), .C(c), .Y(men_men_n594_));
  NOi41      u0566(.An(men_men_n594_), .B(men_men_n339_), .C(men_men_n67_), .D(men_men_n115_), .Y(men_men_n595_));
  OR2        u0567(.A(men_men_n595_), .B(men_men_n593_), .Y(men_men_n596_));
  NOi32      u0568(.An(d), .Bn(a), .C(e), .Y(men_men_n597_));
  NA2        u0569(.A(men_men_n597_), .B(men_men_n111_), .Y(men_men_n598_));
  NO2        u0570(.A(n), .B(c), .Y(men_men_n599_));
  NA3        u0571(.A(men_men_n599_), .B(men_men_n29_), .C(m), .Y(men_men_n600_));
  NAi32      u0572(.An(n), .Bn(f), .C(m), .Y(men_men_n601_));
  NA3        u0573(.A(men_men_n601_), .B(men_men_n600_), .C(men_men_n598_), .Y(men_men_n602_));
  NOi32      u0574(.An(e), .Bn(a), .C(d), .Y(men_men_n603_));
  AOI210     u0575(.A0(men_men_n29_), .A1(d), .B0(men_men_n603_), .Y(men_men_n604_));
  AOI210     u0576(.A0(men_men_n604_), .A1(men_men_n213_), .B0(men_men_n541_), .Y(men_men_n605_));
  AOI210     u0577(.A0(men_men_n605_), .A1(men_men_n602_), .B0(men_men_n596_), .Y(men_men_n606_));
  INV        u0578(.A(men_men_n606_), .Y(men_men_n607_));
  AOI210     u0579(.A0(men_men_n591_), .A1(men_men_n577_), .B0(men_men_n607_), .Y(men_men_n608_));
  NO3        u0580(.A(men_men_n310_), .B(men_men_n59_), .C(n), .Y(men_men_n609_));
  NA3        u0581(.A(men_men_n498_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n610_));
  NA2        u0582(.A(men_men_n444_), .B(men_men_n227_), .Y(men_men_n611_));
  OR2        u0583(.A(men_men_n611_), .B(men_men_n610_), .Y(men_men_n612_));
  NA2        u0584(.A(men_men_n72_), .B(men_men_n111_), .Y(men_men_n613_));
  NO2        u0585(.A(men_men_n613_), .B(men_men_n45_), .Y(men_men_n614_));
  AOI220     u0586(.A0(men_men_n614_), .A1(men_men_n528_), .B0(men_men_n612_), .B1(men_men_n609_), .Y(men_men_n615_));
  NO2        u0587(.A(men_men_n615_), .B(men_men_n85_), .Y(men_men_n616_));
  NA3        u0588(.A(men_men_n543_), .B(men_men_n326_), .C(men_men_n46_), .Y(men_men_n617_));
  NOi32      u0589(.An(e), .Bn(c), .C(f), .Y(men_men_n618_));
  NOi21      u0590(.An(f), .B(g), .Y(men_men_n619_));
  NO2        u0591(.A(men_men_n619_), .B(men_men_n211_), .Y(men_men_n620_));
  NA2        u0592(.A(men_men_n617_), .B(men_men_n180_), .Y(men_men_n621_));
  AOI210     u0593(.A0(men_men_n527_), .A1(men_men_n384_), .B0(men_men_n294_), .Y(men_men_n622_));
  NA2        u0594(.A(men_men_n622_), .B(men_men_n258_), .Y(men_men_n623_));
  NOi21      u0595(.An(j), .B(l), .Y(men_men_n624_));
  NO2        u0596(.A(k), .B(men_men_n256_), .Y(men_men_n625_));
  NA2        u0597(.A(men_men_n625_), .B(men_men_n624_), .Y(men_men_n626_));
  OR2        u0598(.A(men_men_n626_), .B(men_men_n582_), .Y(men_men_n627_));
  NOi31      u0599(.An(m), .B(n), .C(k), .Y(men_men_n628_));
  NA2        u0600(.A(men_men_n624_), .B(men_men_n628_), .Y(men_men_n629_));
  AOI210     u0601(.A0(men_men_n384_), .A1(men_men_n358_), .B0(men_men_n294_), .Y(men_men_n630_));
  NAi21      u0602(.An(men_men_n629_), .B(men_men_n630_), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n271_), .B(men_men_n49_), .Y(men_men_n632_));
  NO2        u0604(.A(men_men_n304_), .B(men_men_n592_), .Y(men_men_n633_));
  NO2        u0605(.A(men_men_n523_), .B(men_men_n49_), .Y(men_men_n634_));
  AOI220     u0606(.A0(men_men_n634_), .A1(men_men_n633_), .B0(men_men_n632_), .B1(men_men_n563_), .Y(men_men_n635_));
  NA4        u0607(.A(men_men_n635_), .B(men_men_n631_), .C(men_men_n627_), .D(men_men_n623_), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n106_), .B(men_men_n36_), .Y(men_men_n637_));
  NO2        u0609(.A(k), .B(men_men_n214_), .Y(men_men_n638_));
  NO2        u0610(.A(men_men_n519_), .B(men_men_n348_), .Y(men_men_n639_));
  NO2        u0611(.A(men_men_n639_), .B(n), .Y(men_men_n640_));
  NO2        u0612(.A(men_men_n521_), .B(men_men_n178_), .Y(men_men_n641_));
  NA3        u0613(.A(men_men_n544_), .B(men_men_n265_), .C(men_men_n145_), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n494_), .B(men_men_n161_), .Y(men_men_n643_));
  NO3        u0615(.A(men_men_n381_), .B(men_men_n643_), .C(men_men_n85_), .Y(men_men_n644_));
  AOI210     u0616(.A0(men_men_n642_), .A1(men_men_n641_), .B0(men_men_n644_), .Y(men_men_n645_));
  AN3        u0617(.A(f), .B(d), .C(b), .Y(men_men_n646_));
  OAI210     u0618(.A0(men_men_n646_), .A1(men_men_n129_), .B0(n), .Y(men_men_n647_));
  NA3        u0619(.A(men_men_n494_), .B(men_men_n161_), .C(men_men_n214_), .Y(men_men_n648_));
  AOI210     u0620(.A0(men_men_n647_), .A1(men_men_n229_), .B0(men_men_n648_), .Y(men_men_n649_));
  NAi31      u0621(.An(m), .B(n), .C(k), .Y(men_men_n650_));
  NO2        u0622(.A(men_men_n134_), .B(men_men_n650_), .Y(men_men_n651_));
  OAI210     u0623(.A0(men_men_n651_), .A1(men_men_n649_), .B0(j), .Y(men_men_n652_));
  NA2        u0624(.A(men_men_n652_), .B(men_men_n645_), .Y(men_men_n653_));
  NO4        u0625(.A(men_men_n653_), .B(men_men_n636_), .C(men_men_n621_), .D(men_men_n616_), .Y(men_men_n654_));
  NAi31      u0626(.An(g), .B(h), .C(f), .Y(men_men_n655_));
  OR3        u0627(.A(men_men_n655_), .B(men_men_n271_), .C(n), .Y(men_men_n656_));
  OA210      u0628(.A0(men_men_n523_), .A1(n), .B0(men_men_n580_), .Y(men_men_n657_));
  NA3        u0629(.A(men_men_n403_), .B(men_men_n119_), .C(men_men_n82_), .Y(men_men_n658_));
  OAI210     u0630(.A0(men_men_n657_), .A1(men_men_n89_), .B0(men_men_n658_), .Y(men_men_n659_));
  NOi21      u0631(.An(men_men_n656_), .B(men_men_n659_), .Y(men_men_n660_));
  NO2        u0632(.A(men_men_n660_), .B(men_men_n516_), .Y(men_men_n661_));
  NO3        u0633(.A(g), .B(men_men_n213_), .C(men_men_n54_), .Y(men_men_n662_));
  NAi21      u0634(.An(h), .B(j), .Y(men_men_n663_));
  NA2        u0635(.A(men_men_n594_), .B(men_men_n328_), .Y(men_men_n664_));
  OA220      u0636(.A0(men_men_n629_), .A1(men_men_n664_), .B0(men_men_n626_), .B1(men_men_n70_), .Y(men_men_n665_));
  NA3        u0637(.A(men_men_n513_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n666_));
  NA2        u0638(.A(h), .B(men_men_n37_), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n98_), .B(men_men_n46_), .Y(men_men_n668_));
  NO2        u0640(.A(men_men_n668_), .B(men_men_n319_), .Y(men_men_n669_));
  AOI210     u0641(.A0(men_men_n560_), .A1(men_men_n413_), .B0(men_men_n49_), .Y(men_men_n670_));
  INV        u0642(.A(men_men_n669_), .Y(men_men_n671_));
  NA3        u0643(.A(men_men_n671_), .B(men_men_n666_), .C(men_men_n665_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n247_), .B(f), .Y(men_men_n673_));
  NA2        u0645(.A(men_men_n317_), .B(men_men_n140_), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n131_), .B(men_men_n49_), .Y(men_men_n675_));
  AOI220     u0647(.A0(men_men_n675_), .A1(men_men_n519_), .B0(men_men_n348_), .B1(men_men_n111_), .Y(men_men_n676_));
  OA220      u0648(.A0(men_men_n676_), .A1(men_men_n541_), .B0(men_men_n346_), .B1(men_men_n109_), .Y(men_men_n677_));
  OAI210     u0649(.A0(men_men_n674_), .A1(men_men_n247_), .B0(men_men_n677_), .Y(men_men_n678_));
  NO3        u0650(.A(men_men_n391_), .B(men_men_n191_), .C(men_men_n190_), .Y(men_men_n679_));
  NA2        u0651(.A(men_men_n679_), .B(men_men_n227_), .Y(men_men_n680_));
  NA3        u0652(.A(men_men_n680_), .B(men_men_n249_), .C(j), .Y(men_men_n681_));
  NO3        u0653(.A(men_men_n444_), .B(men_men_n175_), .C(i), .Y(men_men_n682_));
  NA2        u0654(.A(men_men_n448_), .B(men_men_n82_), .Y(men_men_n683_));
  NO4        u0655(.A(men_men_n516_), .B(men_men_n683_), .C(men_men_n130_), .D(men_men_n213_), .Y(men_men_n684_));
  INV        u0656(.A(men_men_n684_), .Y(men_men_n685_));
  NA4        u0657(.A(men_men_n685_), .B(men_men_n681_), .C(men_men_n501_), .D(men_men_n389_), .Y(men_men_n686_));
  NO4        u0658(.A(men_men_n686_), .B(men_men_n678_), .C(men_men_n672_), .D(men_men_n661_), .Y(men_men_n687_));
  NA4        u0659(.A(men_men_n687_), .B(men_men_n654_), .C(men_men_n608_), .D(men_men_n574_), .Y(men08));
  NO2        u0660(.A(k), .B(h), .Y(men_men_n689_));
  AO210      u0661(.A0(men_men_n247_), .A1(men_men_n434_), .B0(men_men_n689_), .Y(men_men_n690_));
  NO2        u0662(.A(men_men_n690_), .B(men_men_n292_), .Y(men_men_n691_));
  NA2        u0663(.A(men_men_n618_), .B(men_men_n82_), .Y(men_men_n692_));
  INV        u0664(.A(men_men_n479_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n82_), .B(men_men_n108_), .Y(men_men_n694_));
  NO2        u0666(.A(men_men_n694_), .B(men_men_n55_), .Y(men_men_n695_));
  NO4        u0667(.A(men_men_n365_), .B(men_men_n110_), .C(j), .D(men_men_n214_), .Y(men_men_n696_));
  NA2        u0668(.A(men_men_n570_), .B(men_men_n229_), .Y(men_men_n697_));
  AOI220     u0669(.A0(men_men_n697_), .A1(men_men_n333_), .B0(men_men_n696_), .B1(men_men_n695_), .Y(men_men_n698_));
  AOI210     u0670(.A0(men_men_n570_), .A1(men_men_n157_), .B0(men_men_n82_), .Y(men_men_n699_));
  NA4        u0671(.A(men_men_n216_), .B(men_men_n140_), .C(men_men_n45_), .D(h), .Y(men_men_n700_));
  AN2        u0672(.A(l), .B(k), .Y(men_men_n701_));
  NA4        u0673(.A(men_men_n701_), .B(men_men_n106_), .C(men_men_n71_), .D(men_men_n214_), .Y(men_men_n702_));
  OAI210     u0674(.A0(men_men_n700_), .A1(g), .B0(men_men_n702_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n703_), .B(men_men_n699_), .Y(men_men_n704_));
  NA4        u0676(.A(men_men_n704_), .B(men_men_n698_), .C(men_men_n693_), .D(men_men_n335_), .Y(men_men_n705_));
  AN2        u0677(.A(men_men_n524_), .B(men_men_n94_), .Y(men_men_n706_));
  NO4        u0678(.A(men_men_n175_), .B(men_men_n379_), .C(men_men_n110_), .D(g), .Y(men_men_n707_));
  AOI210     u0679(.A0(men_men_n707_), .A1(men_men_n697_), .B0(men_men_n508_), .Y(men_men_n708_));
  NO2        u0680(.A(men_men_n38_), .B(men_men_n213_), .Y(men_men_n709_));
  AOI220     u0681(.A0(men_men_n620_), .A1(men_men_n332_), .B0(men_men_n709_), .B1(men_men_n557_), .Y(men_men_n710_));
  NAi31      u0682(.An(men_men_n706_), .B(men_men_n710_), .C(men_men_n708_), .Y(men_men_n711_));
  NO2        u0683(.A(men_men_n527_), .B(men_men_n35_), .Y(men_men_n712_));
  OAI210     u0684(.A0(men_men_n544_), .A1(men_men_n47_), .B0(men_men_n134_), .Y(men_men_n713_));
  NO2        u0685(.A(men_men_n471_), .B(men_men_n131_), .Y(men_men_n714_));
  AOI210     u0686(.A0(men_men_n714_), .A1(men_men_n713_), .B0(men_men_n712_), .Y(men_men_n715_));
  NO3        u0687(.A(men_men_n310_), .B(men_men_n130_), .C(men_men_n41_), .Y(men_men_n716_));
  NAi21      u0688(.An(men_men_n716_), .B(men_men_n702_), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n690_), .B(men_men_n135_), .Y(men_men_n718_));
  AOI220     u0690(.A0(men_men_n718_), .A1(men_men_n390_), .B0(men_men_n717_), .B1(men_men_n74_), .Y(men_men_n719_));
  OAI210     u0691(.A0(men_men_n715_), .A1(men_men_n85_), .B0(men_men_n719_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n348_), .B(men_men_n43_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n680_), .B(men_men_n320_), .C(men_men_n371_), .Y(men_men_n722_));
  NA2        u0694(.A(men_men_n701_), .B(men_men_n221_), .Y(men_men_n723_));
  NO2        u0695(.A(men_men_n723_), .B(men_men_n316_), .Y(men_men_n724_));
  AOI210     u0696(.A0(men_men_n724_), .A1(men_men_n673_), .B0(men_men_n478_), .Y(men_men_n725_));
  NA3        u0697(.A(m), .B(l), .C(k), .Y(men_men_n726_));
  AOI210     u0698(.A0(men_men_n658_), .A1(men_men_n656_), .B0(men_men_n726_), .Y(men_men_n727_));
  NO2        u0699(.A(men_men_n526_), .B(men_men_n266_), .Y(men_men_n728_));
  NOi21      u0700(.An(men_men_n728_), .B(men_men_n520_), .Y(men_men_n729_));
  NA4        u0701(.A(men_men_n111_), .B(l), .C(k), .D(men_men_n85_), .Y(men_men_n730_));
  NA3        u0702(.A(men_men_n119_), .B(men_men_n399_), .C(i), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n731_), .B(men_men_n730_), .Y(men_men_n732_));
  NO3        u0704(.A(men_men_n732_), .B(men_men_n729_), .C(men_men_n727_), .Y(men_men_n733_));
  NA4        u0705(.A(men_men_n733_), .B(men_men_n725_), .C(men_men_n722_), .D(men_men_n721_), .Y(men_men_n734_));
  NO4        u0706(.A(men_men_n734_), .B(men_men_n720_), .C(men_men_n711_), .D(men_men_n705_), .Y(men_men_n735_));
  NOi31      u0707(.An(g), .B(h), .C(f), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n634_), .B(men_men_n736_), .Y(men_men_n737_));
  AO210      u0709(.A0(men_men_n737_), .A1(men_men_n584_), .B0(men_men_n529_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n384_), .B(men_men_n514_), .C(h), .Y(men_men_n739_));
  NA2        u0711(.A(men_men_n739_), .B(men_men_n111_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n740_), .B(men_men_n738_), .Y(men_men_n741_));
  NA2        u0713(.A(men_men_n701_), .B(men_men_n71_), .Y(men_men_n742_));
  NO4        u0714(.A(men_men_n679_), .B(men_men_n175_), .C(n), .D(i), .Y(men_men_n743_));
  NOi21      u0715(.An(h), .B(j), .Y(men_men_n744_));
  NA2        u0716(.A(men_men_n744_), .B(f), .Y(men_men_n745_));
  NO2        u0717(.A(men_men_n745_), .B(men_men_n242_), .Y(men_men_n746_));
  NO3        u0718(.A(men_men_n746_), .B(men_men_n743_), .C(men_men_n682_), .Y(men_men_n747_));
  OAI220     u0719(.A0(men_men_n747_), .A1(men_men_n742_), .B0(men_men_n586_), .B1(men_men_n60_), .Y(men_men_n748_));
  AOI210     u0720(.A0(men_men_n741_), .A1(l), .B0(men_men_n748_), .Y(men_men_n749_));
  NO2        u0721(.A(j), .B(i), .Y(men_men_n750_));
  NA3        u0722(.A(men_men_n750_), .B(men_men_n78_), .C(l), .Y(men_men_n751_));
  NA2        u0723(.A(men_men_n750_), .B(men_men_n33_), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n407_), .B(men_men_n119_), .Y(men_men_n753_));
  OA220      u0725(.A0(men_men_n753_), .A1(men_men_n752_), .B0(men_men_n751_), .B1(men_men_n582_), .Y(men_men_n754_));
  NO3        u0726(.A(men_men_n152_), .B(men_men_n49_), .C(men_men_n108_), .Y(men_men_n755_));
  NO3        u0727(.A(men_men_n533_), .B(men_men_n150_), .C(men_men_n71_), .Y(men_men_n756_));
  NO3        u0728(.A(men_men_n471_), .B(men_men_n423_), .C(j), .Y(men_men_n757_));
  OAI210     u0729(.A0(men_men_n756_), .A1(men_men_n755_), .B0(men_men_n757_), .Y(men_men_n758_));
  OAI210     u0730(.A0(men_men_n737_), .A1(men_men_n60_), .B0(men_men_n758_), .Y(men_men_n759_));
  NA2        u0731(.A(k), .B(j), .Y(men_men_n760_));
  NO3        u0732(.A(men_men_n292_), .B(men_men_n760_), .C(men_men_n40_), .Y(men_men_n761_));
  AOI210     u0733(.A0(men_men_n519_), .A1(n), .B0(men_men_n543_), .Y(men_men_n762_));
  NA2        u0734(.A(men_men_n762_), .B(men_men_n546_), .Y(men_men_n763_));
  AN3        u0735(.A(men_men_n763_), .B(men_men_n761_), .C(men_men_n97_), .Y(men_men_n764_));
  NO3        u0736(.A(men_men_n175_), .B(men_men_n379_), .C(men_men_n110_), .Y(men_men_n765_));
  AOI220     u0737(.A0(men_men_n765_), .A1(men_men_n243_), .B0(men_men_n611_), .B1(men_men_n301_), .Y(men_men_n766_));
  NAi31      u0738(.An(men_men_n604_), .B(men_men_n91_), .C(men_men_n82_), .Y(men_men_n767_));
  NA2        u0739(.A(men_men_n767_), .B(men_men_n766_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n716_), .B(men_men_n699_), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n726_), .B(men_men_n89_), .Y(men_men_n770_));
  NO2        u0742(.A(men_men_n583_), .B(men_men_n115_), .Y(men_men_n771_));
  OAI210     u0743(.A0(men_men_n771_), .A1(men_men_n757_), .B0(men_men_n670_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n772_), .B(men_men_n769_), .Y(men_men_n773_));
  OR4        u0745(.A(men_men_n773_), .B(men_men_n768_), .C(men_men_n764_), .D(men_men_n759_), .Y(men_men_n774_));
  NA3        u0746(.A(men_men_n762_), .B(men_men_n546_), .C(men_men_n545_), .Y(men_men_n775_));
  NA4        u0747(.A(men_men_n775_), .B(men_men_n216_), .C(men_men_n434_), .D(men_men_n34_), .Y(men_men_n776_));
  NO4        u0748(.A(men_men_n471_), .B(men_men_n418_), .C(j), .D(f), .Y(men_men_n777_));
  OAI220     u0749(.A0(men_men_n700_), .A1(men_men_n692_), .B0(men_men_n319_), .B1(men_men_n38_), .Y(men_men_n778_));
  AOI210     u0750(.A0(men_men_n777_), .A1(men_men_n252_), .B0(men_men_n778_), .Y(men_men_n779_));
  NA3        u0751(.A(men_men_n536_), .B(men_men_n285_), .C(h), .Y(men_men_n780_));
  NOi21      u0752(.An(men_men_n670_), .B(men_men_n780_), .Y(men_men_n781_));
  OAI220     u0753(.A0(men_men_n780_), .A1(men_men_n600_), .B0(men_men_n751_), .B1(men_men_n70_), .Y(men_men_n782_));
  INV        u0754(.A(men_men_n782_), .Y(men_men_n783_));
  NAi41      u0755(.An(men_men_n781_), .B(men_men_n783_), .C(men_men_n779_), .D(men_men_n776_), .Y(men_men_n784_));
  OR2        u0756(.A(men_men_n770_), .B(men_men_n94_), .Y(men_men_n785_));
  AOI220     u0757(.A0(men_men_n785_), .A1(men_men_n235_), .B0(men_men_n757_), .B1(men_men_n632_), .Y(men_men_n786_));
  NO2        u0758(.A(men_men_n657_), .B(men_men_n71_), .Y(men_men_n787_));
  AOI210     u0759(.A0(men_men_n777_), .A1(men_men_n787_), .B0(men_men_n322_), .Y(men_men_n788_));
  NO2        u0760(.A(men_men_n780_), .B(men_men_n477_), .Y(men_men_n789_));
  INV        u0761(.A(men_men_n789_), .Y(men_men_n790_));
  NA3        u0762(.A(men_men_n790_), .B(men_men_n788_), .C(men_men_n786_), .Y(men_men_n791_));
  NOi41      u0763(.An(men_men_n754_), .B(men_men_n791_), .C(men_men_n784_), .D(men_men_n774_), .Y(men_men_n792_));
  OR2        u0764(.A(men_men_n700_), .B(men_men_n229_), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n327_), .B(men_men_n294_), .C(men_men_n110_), .Y(men_men_n794_));
  NA2        u0766(.A(men_men_n794_), .B(men_men_n763_), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n46_), .B(men_men_n54_), .Y(men_men_n796_));
  NO3        u0768(.A(men_men_n796_), .B(men_men_n752_), .C(men_men_n271_), .Y(men_men_n797_));
  INV        u0769(.A(men_men_n797_), .Y(men_men_n798_));
  NA4        u0770(.A(men_men_n798_), .B(men_men_n795_), .C(men_men_n793_), .D(men_men_n392_), .Y(men_men_n799_));
  OR2        u0771(.A(men_men_n655_), .B(men_men_n90_), .Y(men_men_n800_));
  NOi31      u0772(.An(b), .B(d), .C(a), .Y(men_men_n801_));
  NO2        u0773(.A(men_men_n801_), .B(men_men_n597_), .Y(men_men_n802_));
  NO2        u0774(.A(men_men_n802_), .B(n), .Y(men_men_n803_));
  INV        u0775(.A(men_men_n803_), .Y(men_men_n804_));
  OAI220     u0776(.A0(men_men_n804_), .A1(men_men_n800_), .B0(men_men_n780_), .B1(men_men_n598_), .Y(men_men_n805_));
  NO2        u0777(.A(men_men_n544_), .B(men_men_n82_), .Y(men_men_n806_));
  NO2        u0778(.A(men_men_n316_), .B(men_men_n115_), .Y(men_men_n807_));
  NOi21      u0779(.An(men_men_n807_), .B(men_men_n162_), .Y(men_men_n808_));
  AOI210     u0780(.A0(men_men_n794_), .A1(men_men_n806_), .B0(men_men_n808_), .Y(men_men_n809_));
  INV        u0781(.A(men_men_n809_), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n679_), .B(n), .Y(men_men_n811_));
  NA2        u0783(.A(men_men_n811_), .B(men_men_n691_), .Y(men_men_n812_));
  NO2        u0784(.A(men_men_n314_), .B(men_men_n234_), .Y(men_men_n813_));
  OAI210     u0785(.A0(men_men_n94_), .A1(men_men_n91_), .B0(men_men_n813_), .Y(men_men_n814_));
  NA2        u0786(.A(men_men_n119_), .B(men_men_n82_), .Y(men_men_n815_));
  AOI210     u0787(.A0(men_men_n410_), .A1(men_men_n404_), .B0(men_men_n815_), .Y(men_men_n816_));
  NAi21      u0788(.An(men_men_n816_), .B(men_men_n814_), .Y(men_men_n817_));
  NA2        u0789(.A(men_men_n724_), .B(men_men_n34_), .Y(men_men_n818_));
  NAi21      u0790(.An(men_men_n730_), .B(men_men_n419_), .Y(men_men_n819_));
  NO2        u0791(.A(men_men_n266_), .B(i), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n707_), .B(men_men_n334_), .Y(men_men_n821_));
  OAI210     u0793(.A0(men_men_n589_), .A1(men_men_n588_), .B0(j), .Y(men_men_n822_));
  AN3        u0794(.A(men_men_n822_), .B(men_men_n821_), .C(men_men_n819_), .Y(men_men_n823_));
  NAi41      u0795(.An(men_men_n817_), .B(men_men_n823_), .C(men_men_n818_), .D(men_men_n812_), .Y(men_men_n824_));
  NO4        u0796(.A(men_men_n824_), .B(men_men_n810_), .C(men_men_n805_), .D(men_men_n799_), .Y(men_men_n825_));
  NA4        u0797(.A(men_men_n825_), .B(men_men_n792_), .C(men_men_n749_), .D(men_men_n735_), .Y(men09));
  INV        u0798(.A(men_men_n120_), .Y(men_men_n827_));
  NA2        u0799(.A(f), .B(e), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n225_), .B(men_men_n110_), .Y(men_men_n829_));
  NA2        u0801(.A(men_men_n829_), .B(g), .Y(men_men_n830_));
  NA4        u0802(.A(men_men_n304_), .B(men_men_n457_), .C(men_men_n254_), .D(men_men_n117_), .Y(men_men_n831_));
  AOI210     u0803(.A0(men_men_n831_), .A1(g), .B0(men_men_n454_), .Y(men_men_n832_));
  AOI210     u0804(.A0(men_men_n832_), .A1(men_men_n830_), .B0(men_men_n828_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n429_), .B(e), .Y(men_men_n834_));
  NO2        u0806(.A(men_men_n834_), .B(men_men_n498_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n833_), .A1(men_men_n827_), .B0(men_men_n835_), .Y(men_men_n836_));
  NO2        u0808(.A(men_men_n203_), .B(men_men_n213_), .Y(men_men_n837_));
  NA3        u0809(.A(m), .B(l), .C(i), .Y(men_men_n838_));
  NA4        u0810(.A(men_men_n86_), .B(men_men_n85_), .C(g), .D(f), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n839_), .B(men_men_n424_), .Y(men_men_n840_));
  OR2        u0812(.A(men_men_n840_), .B(men_men_n837_), .Y(men_men_n841_));
  NA3        u0813(.A(men_men_n800_), .B(men_men_n559_), .C(men_men_n507_), .Y(men_men_n842_));
  OA210      u0814(.A0(men_men_n842_), .A1(men_men_n841_), .B0(men_men_n803_), .Y(men_men_n843_));
  INV        u0815(.A(men_men_n325_), .Y(men_men_n844_));
  NO2        u0816(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n845_));
  NOi31      u0817(.An(k), .B(m), .C(l), .Y(men_men_n846_));
  NO2        u0818(.A(men_men_n326_), .B(men_men_n846_), .Y(men_men_n847_));
  AOI210     u0819(.A0(men_men_n847_), .A1(men_men_n845_), .B0(men_men_n592_), .Y(men_men_n848_));
  NA2        u0820(.A(men_men_n328_), .B(men_men_n329_), .Y(men_men_n849_));
  NA2        u0821(.A(men_men_n848_), .B(men_men_n844_), .Y(men_men_n850_));
  NA3        u0822(.A(men_men_n112_), .B(men_men_n189_), .C(men_men_n31_), .Y(men_men_n851_));
  NA3        u0823(.A(men_men_n851_), .B(men_men_n850_), .C(men_men_n80_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n579_), .B(men_men_n485_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n853_), .B(men_men_n189_), .Y(men_men_n854_));
  NOi21      u0826(.An(f), .B(d), .Y(men_men_n855_));
  NA2        u0827(.A(men_men_n855_), .B(m), .Y(men_men_n856_));
  NOi32      u0828(.An(g), .Bn(f), .C(d), .Y(men_men_n857_));
  NA4        u0829(.A(men_men_n857_), .B(men_men_n599_), .C(men_men_n29_), .D(m), .Y(men_men_n858_));
  NA3        u0830(.A(men_men_n304_), .B(men_men_n254_), .C(men_men_n117_), .Y(men_men_n859_));
  AN2        u0831(.A(f), .B(d), .Y(men_men_n860_));
  NA3        u0832(.A(men_men_n462_), .B(men_men_n860_), .C(men_men_n82_), .Y(men_men_n861_));
  NO3        u0833(.A(men_men_n861_), .B(men_men_n71_), .C(men_men_n214_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n859_), .B(men_men_n862_), .Y(men_men_n863_));
  NAi41      u0835(.An(men_men_n476_), .B(men_men_n863_), .C(men_men_n858_), .D(men_men_n854_), .Y(men_men_n864_));
  NO4        u0836(.A(men_men_n619_), .B(men_men_n131_), .C(men_men_n316_), .D(men_men_n153_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n650_), .B(men_men_n316_), .Y(men_men_n866_));
  AN2        u0838(.A(men_men_n866_), .B(men_men_n673_), .Y(men_men_n867_));
  NO3        u0839(.A(men_men_n867_), .B(men_men_n865_), .C(men_men_n231_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n597_), .B(men_men_n82_), .Y(men_men_n869_));
  NO2        u0841(.A(men_men_n849_), .B(men_men_n869_), .Y(men_men_n870_));
  NOi21      u0842(.An(men_men_n223_), .B(men_men_n870_), .Y(men_men_n871_));
  NA2        u0843(.A(c), .B(men_men_n114_), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n872_), .B(men_men_n396_), .Y(men_men_n873_));
  NA3        u0845(.A(men_men_n873_), .B(men_men_n496_), .C(f), .Y(men_men_n874_));
  OR2        u0846(.A(men_men_n655_), .B(men_men_n530_), .Y(men_men_n875_));
  NA3        u0847(.A(men_men_n874_), .B(men_men_n871_), .C(men_men_n868_), .Y(men_men_n876_));
  NO4        u0848(.A(men_men_n876_), .B(men_men_n864_), .C(men_men_n852_), .D(men_men_n843_), .Y(men_men_n877_));
  OR2        u0849(.A(men_men_n861_), .B(men_men_n71_), .Y(men_men_n878_));
  NA2        u0850(.A(men_men_n110_), .B(j), .Y(men_men_n879_));
  NA2        u0851(.A(men_men_n829_), .B(g), .Y(men_men_n880_));
  AOI210     u0852(.A0(men_men_n880_), .A1(men_men_n286_), .B0(men_men_n878_), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n319_), .B(men_men_n839_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n135_), .B(men_men_n131_), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n227_), .B(men_men_n224_), .Y(men_men_n884_));
  AOI220     u0856(.A0(men_men_n884_), .A1(men_men_n226_), .B0(men_men_n299_), .B1(men_men_n883_), .Y(men_men_n885_));
  NA2        u0857(.A(e), .B(d), .Y(men_men_n886_));
  OAI220     u0858(.A0(men_men_n886_), .A1(c), .B0(men_men_n314_), .B1(d), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n182_), .B(men_men_n227_), .Y(men_men_n888_));
  AOI210     u0860(.A0(men_men_n620_), .A1(men_men_n332_), .B0(men_men_n888_), .Y(men_men_n889_));
  INV        u0861(.A(men_men_n278_), .Y(men_men_n890_));
  NA2        u0862(.A(men_men_n862_), .B(men_men_n890_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n891_), .B(men_men_n889_), .Y(men_men_n892_));
  NO4        u0864(.A(men_men_n892_), .B(men_men_n1483_), .C(men_men_n882_), .D(men_men_n881_), .Y(men_men_n893_));
  NA2        u0865(.A(men_men_n844_), .B(men_men_n31_), .Y(men_men_n894_));
  AO210      u0866(.A0(men_men_n894_), .A1(men_men_n692_), .B0(men_men_n217_), .Y(men_men_n895_));
  NA2        u0867(.A(men_men_n609_), .B(men_men_n618_), .Y(men_men_n896_));
  OAI210     u0868(.A0(men_men_n834_), .A1(men_men_n172_), .B0(men_men_n896_), .Y(men_men_n897_));
  AOI210     u0869(.A0(men_men_n116_), .A1(men_men_n115_), .B0(men_men_n253_), .Y(men_men_n898_));
  NOi31      u0870(.An(men_men_n534_), .B(men_men_n856_), .C(men_men_n286_), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n899_), .B(men_men_n897_), .Y(men_men_n900_));
  AO220      u0872(.A0(men_men_n438_), .A1(men_men_n744_), .B0(men_men_n177_), .B1(f), .Y(men_men_n901_));
  OAI210     u0873(.A0(men_men_n901_), .A1(men_men_n440_), .B0(men_men_n887_), .Y(men_men_n902_));
  NO2        u0874(.A(men_men_n423_), .B(men_men_n68_), .Y(men_men_n903_));
  OAI210     u0875(.A0(men_men_n842_), .A1(men_men_n903_), .B0(men_men_n695_), .Y(men_men_n904_));
  AN4        u0876(.A(men_men_n904_), .B(men_men_n902_), .C(men_men_n900_), .D(men_men_n895_), .Y(men_men_n905_));
  NA4        u0877(.A(men_men_n905_), .B(men_men_n893_), .C(men_men_n877_), .D(men_men_n836_), .Y(men12));
  NA2        u0878(.A(men_men_n534_), .B(men_men_n903_), .Y(men_men_n907_));
  NO2        u0879(.A(men_men_n436_), .B(men_men_n114_), .Y(men_men_n908_));
  NO2        u0880(.A(men_men_n845_), .B(men_men_n339_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n655_), .B(men_men_n365_), .Y(men_men_n910_));
  NA2        u0882(.A(men_men_n909_), .B(men_men_n908_), .Y(men_men_n911_));
  NA3        u0883(.A(men_men_n911_), .B(men_men_n907_), .C(men_men_n427_), .Y(men_men_n912_));
  AOI210     u0884(.A0(men_men_n321_), .A1(men_men_n377_), .B0(men_men_n214_), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n913_), .B(men_men_n391_), .Y(men_men_n914_));
  NO2        u0886(.A(men_men_n637_), .B(men_men_n256_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n583_), .B(men_men_n838_), .Y(men_men_n916_));
  AOI220     u0888(.A0(men_men_n916_), .A1(men_men_n557_), .B0(men_men_n813_), .B1(men_men_n915_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n152_), .B(men_men_n234_), .Y(men_men_n918_));
  NA2        u0890(.A(men_men_n918_), .B(men_men_n237_), .Y(men_men_n919_));
  NA3        u0891(.A(men_men_n919_), .B(men_men_n917_), .C(men_men_n914_), .Y(men_men_n920_));
  OR2        u0892(.A(men_men_n315_), .B(men_men_n908_), .Y(men_men_n921_));
  NO3        u0893(.A(men_men_n131_), .B(men_men_n153_), .C(men_men_n214_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n922_), .B(men_men_n519_), .Y(men_men_n923_));
  NA4        u0895(.A(men_men_n429_), .B(men_men_n421_), .C(men_men_n183_), .D(g), .Y(men_men_n924_));
  NA2        u0896(.A(men_men_n924_), .B(men_men_n923_), .Y(men_men_n925_));
  NO3        u0897(.A(men_men_n660_), .B(men_men_n90_), .C(men_men_n45_), .Y(men_men_n926_));
  NO4        u0898(.A(men_men_n926_), .B(men_men_n925_), .C(men_men_n920_), .D(men_men_n912_), .Y(men_men_n927_));
  NO2        u0899(.A(men_men_n355_), .B(men_men_n354_), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n580_), .B(men_men_n70_), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n544_), .B(men_men_n145_), .Y(men_men_n930_));
  NOi21      u0902(.An(men_men_n34_), .B(men_men_n650_), .Y(men_men_n931_));
  AOI220     u0903(.A0(men_men_n931_), .A1(men_men_n930_), .B0(men_men_n929_), .B1(men_men_n928_), .Y(men_men_n932_));
  INV        u0904(.A(men_men_n932_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n419_), .B(men_men_n258_), .Y(men_men_n934_));
  NO3        u0906(.A(men_men_n815_), .B(men_men_n87_), .C(men_men_n396_), .Y(men_men_n935_));
  NAi21      u0907(.An(men_men_n935_), .B(men_men_n934_), .Y(men_men_n936_));
  NO2        u0908(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n491_), .B(men_men_n294_), .Y(men_men_n938_));
  INV        u0910(.A(men_men_n352_), .Y(men_men_n939_));
  NO3        u0911(.A(men_men_n939_), .B(men_men_n936_), .C(men_men_n933_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n332_), .B(g), .Y(men_men_n941_));
  NA2        u0913(.A(men_men_n164_), .B(i), .Y(men_men_n942_));
  NA2        u0914(.A(men_men_n46_), .B(i), .Y(men_men_n943_));
  OAI220     u0915(.A0(men_men_n943_), .A1(men_men_n199_), .B0(men_men_n942_), .B1(men_men_n90_), .Y(men_men_n944_));
  AOI210     u0916(.A0(men_men_n406_), .A1(men_men_n37_), .B0(men_men_n944_), .Y(men_men_n945_));
  NO2        u0917(.A(men_men_n145_), .B(men_men_n82_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n544_), .B(men_men_n369_), .Y(men_men_n947_));
  AOI210     u0919(.A0(men_men_n947_), .A1(n), .B0(men_men_n946_), .Y(men_men_n948_));
  OAI220     u0920(.A0(men_men_n948_), .A1(men_men_n941_), .B0(men_men_n945_), .B1(men_men_n319_), .Y(men_men_n949_));
  NO2        u0921(.A(men_men_n655_), .B(men_men_n485_), .Y(men_men_n950_));
  NA3        u0922(.A(men_men_n328_), .B(men_men_n624_), .C(i), .Y(men_men_n951_));
  OAI210     u0923(.A0(men_men_n423_), .A1(men_men_n304_), .B0(men_men_n951_), .Y(men_men_n952_));
  OAI220     u0924(.A0(men_men_n952_), .A1(men_men_n950_), .B0(men_men_n670_), .B1(men_men_n756_), .Y(men_men_n953_));
  NA2        u0925(.A(men_men_n603_), .B(men_men_n111_), .Y(men_men_n954_));
  OR3        u0926(.A(men_men_n304_), .B(men_men_n418_), .C(f), .Y(men_men_n955_));
  NA3        u0927(.A(men_men_n624_), .B(men_men_n78_), .C(i), .Y(men_men_n956_));
  OA220      u0928(.A0(men_men_n956_), .A1(men_men_n954_), .B0(men_men_n955_), .B1(men_men_n582_), .Y(men_men_n957_));
  NA3        u0929(.A(f), .B(men_men_n116_), .C(g), .Y(men_men_n958_));
  AOI210     u0930(.A0(men_men_n667_), .A1(men_men_n958_), .B0(m), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n959_), .A1(men_men_n909_), .B0(men_men_n315_), .Y(men_men_n960_));
  NA2        u0932(.A(men_men_n683_), .B(men_men_n869_), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n839_), .B(men_men_n424_), .Y(men_men_n962_));
  NA2        u0934(.A(i), .B(men_men_n75_), .Y(men_men_n963_));
  NA3        u0935(.A(men_men_n963_), .B(men_men_n956_), .C(men_men_n955_), .Y(men_men_n964_));
  AOI220     u0936(.A0(men_men_n964_), .A1(men_men_n252_), .B0(men_men_n962_), .B1(men_men_n961_), .Y(men_men_n965_));
  NA4        u0937(.A(men_men_n965_), .B(men_men_n960_), .C(men_men_n957_), .D(men_men_n953_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n915_), .B(men_men_n235_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n659_), .B(men_men_n86_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n443_), .B(men_men_n214_), .Y(men_men_n969_));
  AOI220     u0941(.A0(men_men_n969_), .A1(men_men_n370_), .B0(men_men_n921_), .B1(men_men_n218_), .Y(men_men_n970_));
  AOI220     u0942(.A0(men_men_n910_), .A1(men_men_n918_), .B0(men_men_n581_), .B1(men_men_n88_), .Y(men_men_n971_));
  NA4        u0943(.A(men_men_n971_), .B(men_men_n970_), .C(men_men_n968_), .D(men_men_n967_), .Y(men_men_n972_));
  NO2        u0944(.A(men_men_n400_), .B(men_men_n815_), .Y(men_men_n973_));
  OAI210     u0945(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n107_), .Y(men_men_n974_));
  AOI210     u0946(.A0(men_men_n974_), .A1(men_men_n524_), .B0(men_men_n973_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n959_), .B(men_men_n908_), .Y(men_men_n976_));
  NO3        u0948(.A(men_men_n879_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n977_));
  AOI220     u0949(.A0(men_men_n977_), .A1(men_men_n622_), .B0(men_men_n641_), .B1(men_men_n519_), .Y(men_men_n978_));
  NA3        u0950(.A(men_men_n978_), .B(men_men_n976_), .C(men_men_n975_), .Y(men_men_n979_));
  NO4        u0951(.A(men_men_n979_), .B(men_men_n972_), .C(men_men_n966_), .D(men_men_n949_), .Y(men_men_n980_));
  NAi31      u0952(.An(men_men_n141_), .B(men_men_n407_), .C(n), .Y(men_men_n981_));
  NO3        u0953(.A(men_men_n124_), .B(men_men_n326_), .C(men_men_n846_), .Y(men_men_n982_));
  NO2        u0954(.A(men_men_n982_), .B(men_men_n981_), .Y(men_men_n983_));
  INV        u0955(.A(men_men_n983_), .Y(men_men_n984_));
  INV        u0956(.A(men_men_n479_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n985_), .B(men_men_n984_), .Y(men_men_n986_));
  NA2        u0958(.A(men_men_n227_), .B(men_men_n173_), .Y(men_men_n987_));
  NO3        u0959(.A(men_men_n301_), .B(men_men_n429_), .C(men_men_n177_), .Y(men_men_n988_));
  NOi31      u0960(.An(men_men_n987_), .B(men_men_n988_), .C(men_men_n214_), .Y(men_men_n989_));
  NAi21      u0961(.An(men_men_n544_), .B(men_men_n969_), .Y(men_men_n990_));
  NO3        u0962(.A(men_men_n423_), .B(men_men_n304_), .C(men_men_n71_), .Y(men_men_n991_));
  AOI220     u0963(.A0(men_men_n991_), .A1(men_men_n420_), .B0(men_men_n468_), .B1(g), .Y(men_men_n992_));
  NA2        u0964(.A(men_men_n992_), .B(men_men_n990_), .Y(men_men_n993_));
  OAI220     u0965(.A0(men_men_n981_), .A1(men_men_n230_), .B0(men_men_n951_), .B1(men_men_n598_), .Y(men_men_n994_));
  NO2        u0966(.A(men_men_n656_), .B(men_men_n365_), .Y(men_men_n995_));
  NO3        u0967(.A(men_men_n533_), .B(men_men_n150_), .C(men_men_n213_), .Y(men_men_n996_));
  OAI210     u0968(.A0(men_men_n996_), .A1(men_men_n513_), .B0(men_men_n366_), .Y(men_men_n997_));
  NA2        u0969(.A(men_men_n997_), .B(men_men_n617_), .Y(men_men_n998_));
  NA3        u0970(.A(men_men_n947_), .B(men_men_n473_), .C(men_men_n46_), .Y(men_men_n999_));
  AOI210     u0971(.A0(men_men_n368_), .A1(men_men_n366_), .B0(men_men_n318_), .Y(men_men_n1000_));
  NA3        u0972(.A(men_men_n1000_), .B(men_men_n999_), .C(men_men_n267_), .Y(men_men_n1001_));
  OR4        u0973(.A(men_men_n1001_), .B(men_men_n998_), .C(men_men_n995_), .D(men_men_n994_), .Y(men_men_n1002_));
  NO4        u0974(.A(men_men_n1002_), .B(men_men_n993_), .C(men_men_n989_), .D(men_men_n986_), .Y(men_men_n1003_));
  NA4        u0975(.A(men_men_n1003_), .B(men_men_n980_), .C(men_men_n940_), .D(men_men_n927_), .Y(men13));
  NA2        u0976(.A(men_men_n46_), .B(men_men_n85_), .Y(men_men_n1005_));
  AN2        u0977(.A(c), .B(b), .Y(men_men_n1006_));
  NA3        u0978(.A(men_men_n246_), .B(men_men_n1006_), .C(m), .Y(men_men_n1007_));
  NO4        u0979(.A(e), .B(men_men_n1007_), .C(men_men_n1005_), .D(men_men_n576_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n258_), .B(men_men_n1006_), .Y(men_men_n1009_));
  NO4        u0981(.A(men_men_n1009_), .B(e), .C(men_men_n942_), .D(a), .Y(men_men_n1010_));
  NAi32      u0982(.An(d), .Bn(c), .C(e), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n140_), .B(men_men_n45_), .Y(men_men_n1012_));
  NO4        u0984(.A(men_men_n1012_), .B(men_men_n1011_), .C(men_men_n583_), .D(men_men_n300_), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n663_), .B(men_men_n224_), .Y(men_men_n1014_));
  NA2        u0986(.A(men_men_n399_), .B(men_men_n213_), .Y(men_men_n1015_));
  AN2        u0987(.A(d), .B(c), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n1016_), .B(men_men_n114_), .Y(men_men_n1017_));
  NO4        u0989(.A(men_men_n1017_), .B(men_men_n1015_), .C(men_men_n178_), .D(men_men_n170_), .Y(men_men_n1018_));
  NA2        u0990(.A(men_men_n483_), .B(c), .Y(men_men_n1019_));
  NO4        u0991(.A(men_men_n1012_), .B(men_men_n579_), .C(men_men_n1019_), .D(men_men_n300_), .Y(men_men_n1020_));
  AO210      u0992(.A0(men_men_n1018_), .A1(men_men_n1014_), .B0(men_men_n1020_), .Y(men_men_n1021_));
  OR4        u0993(.A(men_men_n1021_), .B(men_men_n1013_), .C(men_men_n1010_), .D(men_men_n1008_), .Y(men_men_n1022_));
  NAi32      u0994(.An(f), .Bn(e), .C(c), .Y(men_men_n1023_));
  NO2        u0995(.A(men_men_n1023_), .B(men_men_n147_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n1024_), .B(g), .Y(men_men_n1025_));
  OR3        u0997(.A(men_men_n224_), .B(men_men_n178_), .C(men_men_n170_), .Y(men_men_n1026_));
  NO2        u0998(.A(men_men_n1026_), .B(men_men_n1025_), .Y(men_men_n1027_));
  NO2        u0999(.A(men_men_n1019_), .B(men_men_n300_), .Y(men_men_n1028_));
  NA2        u1000(.A(men_men_n625_), .B(i), .Y(men_men_n1029_));
  NOi21      u1001(.An(men_men_n1028_), .B(men_men_n1029_), .Y(men_men_n1030_));
  NO2        u1002(.A(men_men_n760_), .B(men_men_n110_), .Y(men_men_n1031_));
  NOi41      u1003(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1032_));
  NA2        u1004(.A(men_men_n1032_), .B(men_men_n1031_), .Y(men_men_n1033_));
  NO2        u1005(.A(men_men_n1033_), .B(men_men_n1025_), .Y(men_men_n1034_));
  OR3        u1006(.A(e), .B(d), .C(c), .Y(men_men_n1035_));
  NA3        u1007(.A(k), .B(j), .C(i), .Y(men_men_n1036_));
  NO3        u1008(.A(men_men_n1036_), .B(men_men_n300_), .C(men_men_n89_), .Y(men_men_n1037_));
  NOi21      u1009(.An(men_men_n1037_), .B(men_men_n1035_), .Y(men_men_n1038_));
  OR4        u1010(.A(men_men_n1038_), .B(men_men_n1034_), .C(men_men_n1030_), .D(men_men_n1027_), .Y(men_men_n1039_));
  NA3        u1011(.A(men_men_n451_), .B(men_men_n320_), .C(men_men_n54_), .Y(men_men_n1040_));
  NO2        u1012(.A(men_men_n1040_), .B(men_men_n1029_), .Y(men_men_n1041_));
  NO2        u1013(.A(f), .B(c), .Y(men_men_n1042_));
  NOi21      u1014(.An(men_men_n1042_), .B(men_men_n428_), .Y(men_men_n1043_));
  NA2        u1015(.A(men_men_n1043_), .B(men_men_n57_), .Y(men_men_n1044_));
  NO3        u1016(.A(i), .B(men_men_n241_), .C(l), .Y(men_men_n1045_));
  NOi21      u1017(.An(men_men_n1045_), .B(men_men_n1044_), .Y(men_men_n1046_));
  OR2        u1018(.A(men_men_n1046_), .B(men_men_n1041_), .Y(men_men_n1047_));
  OR3        u1019(.A(men_men_n1047_), .B(men_men_n1039_), .C(men_men_n1022_), .Y(men02));
  OR3        u1020(.A(h), .B(g), .C(f), .Y(men_men_n1049_));
  OR3        u1021(.A(n), .B(m), .C(i), .Y(men_men_n1050_));
  NO4        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .C(l), .D(men_men_n1035_), .Y(men_men_n1051_));
  NOi31      u1023(.An(e), .B(d), .C(c), .Y(men_men_n1052_));
  AOI210     u1024(.A0(men_men_n1037_), .A1(men_men_n1052_), .B0(men_men_n1013_), .Y(men_men_n1053_));
  NA3        u1025(.A(g), .B(men_men_n451_), .C(h), .Y(men_men_n1054_));
  OR2        u1026(.A(men_men_n1036_), .B(men_men_n300_), .Y(men_men_n1055_));
  OR2        u1027(.A(men_men_n1055_), .B(men_men_n1054_), .Y(men_men_n1056_));
  NO3        u1028(.A(men_men_n1040_), .B(men_men_n1012_), .C(men_men_n579_), .Y(men_men_n1057_));
  NO2        u1029(.A(men_men_n1057_), .B(men_men_n1027_), .Y(men_men_n1058_));
  NA2        u1030(.A(i), .B(h), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n1059_), .B(men_men_n131_), .Y(men_men_n1060_));
  NO3        u1032(.A(men_men_n142_), .B(men_men_n276_), .C(men_men_n214_), .Y(men_men_n1061_));
  AOI210     u1033(.A0(men_men_n1061_), .A1(men_men_n1060_), .B0(men_men_n1030_), .Y(men_men_n1062_));
  NA3        u1034(.A(c), .B(b), .C(a), .Y(men_men_n1063_));
  NO3        u1035(.A(men_men_n1063_), .B(men_men_n886_), .C(men_men_n213_), .Y(men_men_n1064_));
  NO3        u1036(.A(men_men_n1036_), .B(men_men_n49_), .C(men_men_n110_), .Y(men_men_n1065_));
  AOI210     u1037(.A0(men_men_n1065_), .A1(men_men_n1064_), .B0(men_men_n1041_), .Y(men_men_n1066_));
  AN4        u1038(.A(men_men_n1066_), .B(men_men_n1062_), .C(men_men_n1058_), .D(men_men_n1056_), .Y(men_men_n1067_));
  NO2        u1039(.A(men_men_n1017_), .B(men_men_n1015_), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n1033_), .B(men_men_n1026_), .Y(men_men_n1069_));
  AOI210     u1041(.A0(men_men_n1069_), .A1(men_men_n1068_), .B0(men_men_n1008_), .Y(men_men_n1070_));
  NAi41      u1042(.An(men_men_n1051_), .B(men_men_n1070_), .C(men_men_n1067_), .D(men_men_n1053_), .Y(men03));
  NO2        u1043(.A(men_men_n515_), .B(men_men_n592_), .Y(men_men_n1072_));
  NA4        u1044(.A(men_men_n86_), .B(men_men_n85_), .C(g), .D(men_men_n213_), .Y(men_men_n1073_));
  NA4        u1045(.A(men_men_n567_), .B(m), .C(men_men_n110_), .D(men_men_n213_), .Y(men_men_n1074_));
  NA3        u1046(.A(men_men_n1074_), .B(men_men_n356_), .C(men_men_n1073_), .Y(men_men_n1075_));
  NO3        u1047(.A(men_men_n1075_), .B(men_men_n1072_), .C(men_men_n974_), .Y(men_men_n1076_));
  NO2        u1048(.A(men_men_n840_), .B(men_men_n709_), .Y(men_men_n1077_));
  OAI220     u1049(.A0(men_men_n1077_), .A1(men_men_n683_), .B0(men_men_n1076_), .B1(men_men_n580_), .Y(men_men_n1078_));
  NA4        u1050(.A(i), .B(men_men_n1052_), .C(men_men_n328_), .D(men_men_n320_), .Y(men_men_n1079_));
  OAI210     u1051(.A0(men_men_n815_), .A1(men_men_n408_), .B0(men_men_n1079_), .Y(men_men_n1080_));
  NOi31      u1052(.An(m), .B(n), .C(f), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n1081_), .B(men_men_n51_), .Y(men_men_n1082_));
  AN2        u1054(.A(e), .B(c), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n1083_), .B(a), .Y(men_men_n1084_));
  NO2        u1056(.A(men_men_n1084_), .B(men_men_n1082_), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n494_), .B(l), .Y(men_men_n1086_));
  NOi31      u1058(.An(men_men_n857_), .B(men_men_n1007_), .C(men_men_n1086_), .Y(men_men_n1087_));
  NO4        u1059(.A(men_men_n1087_), .B(men_men_n1085_), .C(men_men_n1080_), .D(men_men_n973_), .Y(men_men_n1088_));
  NO2        u1060(.A(men_men_n276_), .B(a), .Y(men_men_n1089_));
  INV        u1061(.A(men_men_n1013_), .Y(men_men_n1090_));
  NO2        u1062(.A(men_men_n85_), .B(g), .Y(men_men_n1091_));
  AOI210     u1063(.A0(men_men_n1091_), .A1(l), .B0(men_men_n1045_), .Y(men_men_n1092_));
  OR2        u1064(.A(men_men_n1092_), .B(men_men_n1044_), .Y(men_men_n1093_));
  NA3        u1065(.A(men_men_n1093_), .B(men_men_n1090_), .C(men_men_n1088_), .Y(men_men_n1094_));
  NO4        u1066(.A(men_men_n1094_), .B(men_men_n1078_), .C(men_men_n817_), .D(men_men_n556_), .Y(men_men_n1095_));
  NA2        u1067(.A(c), .B(b), .Y(men_men_n1096_));
  NO2        u1068(.A(men_men_n694_), .B(men_men_n1096_), .Y(men_men_n1097_));
  OAI210     u1069(.A0(men_men_n856_), .A1(men_men_n832_), .B0(men_men_n402_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n1098_), .B(men_men_n1097_), .Y(men_men_n1099_));
  NAi21      u1071(.An(men_men_n404_), .B(men_men_n1097_), .Y(men_men_n1100_));
  NA3        u1072(.A(men_men_n414_), .B(men_men_n549_), .C(f), .Y(men_men_n1101_));
  OAI210     u1073(.A0(men_men_n538_), .A1(men_men_n39_), .B0(men_men_n1089_), .Y(men_men_n1102_));
  NA3        u1074(.A(men_men_n1102_), .B(men_men_n1101_), .C(men_men_n1100_), .Y(men_men_n1103_));
  NAi21      u1075(.An(f), .B(d), .Y(men_men_n1104_));
  NO2        u1076(.A(men_men_n1104_), .B(men_men_n1063_), .Y(men_men_n1105_));
  AOI210     u1077(.A0(men_men_n1105_), .A1(men_men_n111_), .B0(men_men_n1103_), .Y(men_men_n1106_));
  NA2        u1078(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n184_), .B(men_men_n234_), .Y(men_men_n1108_));
  NA2        u1080(.A(men_men_n1108_), .B(m), .Y(men_men_n1109_));
  NA3        u1081(.A(men_men_n898_), .B(men_men_n1086_), .C(men_men_n457_), .Y(men_men_n1110_));
  INV        u1082(.A(men_men_n455_), .Y(men_men_n1111_));
  AOI210     u1083(.A0(men_men_n1111_), .A1(men_men_n1107_), .B0(men_men_n1109_), .Y(men_men_n1112_));
  NA2        u1084(.A(men_men_n551_), .B(men_men_n398_), .Y(men_men_n1113_));
  NO2        u1085(.A(men_men_n359_), .B(men_men_n358_), .Y(men_men_n1114_));
  AOI210     u1086(.A0(men_men_n1108_), .A1(men_men_n416_), .B0(men_men_n935_), .Y(men_men_n1115_));
  NAi31      u1087(.An(men_men_n1114_), .B(men_men_n1115_), .C(men_men_n1113_), .Y(men_men_n1116_));
  NO2        u1088(.A(men_men_n1116_), .B(men_men_n1112_), .Y(men_men_n1117_));
  NA4        u1089(.A(men_men_n1117_), .B(men_men_n1106_), .C(men_men_n1099_), .D(men_men_n1095_), .Y(men00));
  AOI210     u1090(.A0(men_men_n293_), .A1(men_men_n214_), .B0(men_men_n270_), .Y(men_men_n1119_));
  NO2        u1091(.A(men_men_n1119_), .B(men_men_n570_), .Y(men_men_n1120_));
  INV        u1092(.A(men_men_n1080_), .Y(men_men_n1121_));
  NO3        u1093(.A(men_men_n1057_), .B(men_men_n935_), .C(men_men_n706_), .Y(men_men_n1122_));
  NA3        u1094(.A(men_men_n1122_), .B(men_men_n1121_), .C(men_men_n975_), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n496_), .B(f), .Y(men_men_n1124_));
  OAI210     u1096(.A0(men_men_n982_), .A1(men_men_n40_), .B0(men_men_n643_), .Y(men_men_n1125_));
  NA3        u1097(.A(men_men_n1125_), .B(men_men_n251_), .C(n), .Y(men_men_n1126_));
  AOI210     u1098(.A0(men_men_n1126_), .A1(men_men_n1124_), .B0(men_men_n1017_), .Y(men_men_n1127_));
  NO4        u1099(.A(men_men_n1127_), .B(men_men_n1123_), .C(men_men_n1120_), .D(men_men_n1039_), .Y(men_men_n1128_));
  NA3        u1100(.A(d), .B(men_men_n54_), .C(b), .Y(men_men_n1129_));
  NOi31      u1101(.An(n), .B(m), .C(i), .Y(men_men_n1130_));
  NA3        u1102(.A(men_men_n1130_), .B(men_men_n646_), .C(men_men_n51_), .Y(men_men_n1131_));
  INV        u1103(.A(men_men_n1131_), .Y(men_men_n1132_));
  INV        u1104(.A(men_men_n569_), .Y(men_men_n1133_));
  NO4        u1105(.A(men_men_n1133_), .B(men_men_n1132_), .C(men_men_n1114_), .D(men_men_n899_), .Y(men_men_n1134_));
  NO4        u1106(.A(men_men_n474_), .B(men_men_n342_), .C(men_men_n1096_), .D(men_men_n57_), .Y(men_men_n1135_));
  NA3        u1107(.A(men_men_n371_), .B(men_men_n221_), .C(g), .Y(men_men_n1136_));
  OA220      u1108(.A0(men_men_n1136_), .A1(men_men_n1129_), .B0(men_men_n372_), .B1(men_men_n134_), .Y(men_men_n1137_));
  NO2        u1109(.A(h), .B(g), .Y(men_men_n1138_));
  NA4        u1110(.A(men_men_n486_), .B(men_men_n451_), .C(men_men_n1138_), .D(men_men_n1006_), .Y(men_men_n1139_));
  OAI220     u1111(.A0(men_men_n515_), .A1(men_men_n592_), .B0(men_men_n90_), .B1(men_men_n89_), .Y(men_men_n1140_));
  AOI220     u1112(.A0(men_men_n1140_), .A1(men_men_n524_), .B0(men_men_n922_), .B1(men_men_n568_), .Y(men_men_n1141_));
  AOI220     u1113(.A0(men_men_n311_), .A1(men_men_n243_), .B0(men_men_n179_), .B1(men_men_n149_), .Y(men_men_n1142_));
  NA4        u1114(.A(men_men_n1142_), .B(men_men_n1141_), .C(men_men_n1139_), .D(men_men_n1137_), .Y(men_men_n1143_));
  NO3        u1115(.A(men_men_n1143_), .B(men_men_n1135_), .C(men_men_n260_), .Y(men_men_n1144_));
  INV        u1116(.A(men_men_n313_), .Y(men_men_n1145_));
  AOI210     u1117(.A0(men_men_n243_), .A1(men_men_n332_), .B0(men_men_n571_), .Y(men_men_n1146_));
  NA3        u1118(.A(men_men_n1146_), .B(men_men_n1145_), .C(men_men_n155_), .Y(men_men_n1147_));
  NO2        u1119(.A(men_men_n236_), .B(men_men_n183_), .Y(men_men_n1148_));
  NA2        u1120(.A(men_men_n1148_), .B(men_men_n414_), .Y(men_men_n1149_));
  NA3        u1121(.A(men_men_n181_), .B(men_men_n110_), .C(g), .Y(men_men_n1150_));
  NA3        u1122(.A(men_men_n451_), .B(men_men_n40_), .C(f), .Y(men_men_n1151_));
  NOi31      u1123(.An(j), .B(men_men_n1151_), .C(men_men_n1150_), .Y(men_men_n1152_));
  NAi31      u1124(.An(men_men_n187_), .B(men_men_n853_), .C(men_men_n451_), .Y(men_men_n1153_));
  NAi31      u1125(.An(men_men_n1152_), .B(men_men_n1153_), .C(men_men_n1149_), .Y(men_men_n1154_));
  NO2        u1126(.A(men_men_n269_), .B(men_men_n71_), .Y(men_men_n1155_));
  NO3        u1127(.A(men_men_n413_), .B(men_men_n828_), .C(n), .Y(men_men_n1156_));
  AOI210     u1128(.A0(men_men_n1156_), .A1(men_men_n1155_), .B0(men_men_n1051_), .Y(men_men_n1157_));
  NAi21      u1129(.An(men_men_n1020_), .B(men_men_n1157_), .Y(men_men_n1158_));
  NO4        u1130(.A(men_men_n1158_), .B(men_men_n1154_), .C(men_men_n1147_), .D(men_men_n506_), .Y(men_men_n1159_));
  AN3        u1131(.A(men_men_n1159_), .B(men_men_n1144_), .C(men_men_n1134_), .Y(men_men_n1160_));
  NA2        u1132(.A(men_men_n524_), .B(men_men_n100_), .Y(men_men_n1161_));
  NA3        u1133(.A(men_men_n552_), .B(men_men_n1161_), .C(men_men_n239_), .Y(men_men_n1162_));
  NA2        u1134(.A(men_men_n1075_), .B(men_men_n524_), .Y(men_men_n1163_));
  NA4        u1135(.A(men_men_n646_), .B(men_men_n205_), .C(men_men_n221_), .D(men_men_n164_), .Y(men_men_n1164_));
  NA3        u1136(.A(men_men_n1164_), .B(men_men_n1163_), .C(men_men_n290_), .Y(men_men_n1165_));
  OAI210     u1137(.A0(men_men_n449_), .A1(men_men_n118_), .B0(men_men_n858_), .Y(men_men_n1166_));
  AOI220     u1138(.A0(men_men_n1166_), .A1(men_men_n1110_), .B0(men_men_n551_), .B1(men_men_n398_), .Y(men_men_n1167_));
  OR4        u1139(.A(men_men_n1017_), .B(men_men_n266_), .C(men_men_n222_), .D(e), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n217_), .B(men_men_n214_), .Y(men_men_n1169_));
  NA2        u1141(.A(n), .B(e), .Y(men_men_n1170_));
  NO2        u1142(.A(men_men_n1170_), .B(men_men_n147_), .Y(men_men_n1171_));
  AOI220     u1143(.A0(men_men_n1171_), .A1(men_men_n268_), .B0(men_men_n844_), .B1(men_men_n1169_), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n343_), .A1(men_men_n306_), .B0(men_men_n432_), .Y(men_men_n1173_));
  NA4        u1145(.A(men_men_n1173_), .B(men_men_n1172_), .C(men_men_n1168_), .D(men_men_n1167_), .Y(men_men_n1174_));
  AOI210     u1146(.A0(men_men_n1171_), .A1(men_men_n848_), .B0(men_men_n816_), .Y(men_men_n1175_));
  NO2        u1147(.A(men_men_n66_), .B(h), .Y(men_men_n1176_));
  NO3        u1148(.A(men_men_n1017_), .B(men_men_n1015_), .C(men_men_n723_), .Y(men_men_n1177_));
  OAI210     u1149(.A0(men_men_n1061_), .A1(men_men_n1177_), .B0(men_men_n1176_), .Y(men_men_n1178_));
  NA3        u1150(.A(men_men_n1178_), .B(men_men_n1175_), .C(men_men_n858_), .Y(men_men_n1179_));
  NO4        u1151(.A(men_men_n1179_), .B(men_men_n1174_), .C(men_men_n1165_), .D(men_men_n1162_), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n833_), .B(men_men_n755_), .Y(men_men_n1181_));
  NA4        u1153(.A(men_men_n1181_), .B(men_men_n1180_), .C(men_men_n1160_), .D(men_men_n1128_), .Y(men01));
  NO3        u1154(.A(men_men_n797_), .B(men_men_n789_), .C(men_men_n465_), .Y(men_men_n1183_));
  NA2        u1155(.A(men_men_n382_), .B(i), .Y(men_men_n1184_));
  NA3        u1156(.A(men_men_n1184_), .B(men_men_n1183_), .C(men_men_n997_), .Y(men_men_n1185_));
  NA2        u1157(.A(men_men_n581_), .B(men_men_n88_), .Y(men_men_n1186_));
  NA2        u1158(.A(men_men_n544_), .B(men_men_n265_), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n938_), .B(men_men_n1187_), .Y(men_men_n1188_));
  NA3        u1160(.A(men_men_n1188_), .B(men_men_n1186_), .C(men_men_n896_), .Y(men_men_n1189_));
  NA2        u1161(.A(men_men_n45_), .B(f), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n701_), .B(men_men_n95_), .Y(men_men_n1191_));
  NO2        u1163(.A(men_men_n1191_), .B(men_men_n1190_), .Y(men_men_n1192_));
  OAI210     u1164(.A0(men_men_n780_), .A1(men_men_n598_), .B0(men_men_n1164_), .Y(men_men_n1193_));
  AOI210     u1165(.A0(men_men_n1192_), .A1(men_men_n632_), .B0(men_men_n1193_), .Y(men_men_n1194_));
  INV        u1166(.A(men_men_n116_), .Y(men_men_n1195_));
  OA220      u1167(.A0(men_men_n1195_), .A1(men_men_n578_), .B0(men_men_n657_), .B1(men_men_n356_), .Y(men_men_n1196_));
  NAi41      u1168(.An(men_men_n163_), .B(men_men_n1196_), .C(men_men_n1194_), .D(men_men_n885_), .Y(men_men_n1197_));
  NO3        u1169(.A(men_men_n781_), .B(men_men_n669_), .C(men_men_n499_), .Y(men_men_n1198_));
  NA4        u1170(.A(men_men_n701_), .B(men_men_n95_), .C(men_men_n45_), .D(men_men_n213_), .Y(men_men_n1199_));
  OA220      u1171(.A0(men_men_n1199_), .A1(men_men_n70_), .B0(men_men_n194_), .B1(men_men_n192_), .Y(men_men_n1200_));
  NA3        u1172(.A(men_men_n1200_), .B(men_men_n1198_), .C(men_men_n137_), .Y(men_men_n1201_));
  NO4        u1173(.A(men_men_n1201_), .B(men_men_n1197_), .C(men_men_n1189_), .D(men_men_n1185_), .Y(men_men_n1202_));
  NA2        u1174(.A(men_men_n1136_), .B(men_men_n206_), .Y(men_men_n1203_));
  OAI210     u1175(.A0(men_men_n1203_), .A1(men_men_n296_), .B0(men_men_n519_), .Y(men_men_n1204_));
  NA2        u1176(.A(men_men_n527_), .B(men_men_n384_), .Y(men_men_n1205_));
  NOi21      u1177(.An(men_men_n553_), .B(men_men_n575_), .Y(men_men_n1206_));
  NA2        u1178(.A(men_men_n1206_), .B(men_men_n1205_), .Y(men_men_n1207_));
  NA2        u1179(.A(men_men_n202_), .B(men_men_n34_), .Y(men_men_n1208_));
  OR2        u1180(.A(men_men_n1208_), .B(men_men_n319_), .Y(men_men_n1209_));
  NA3        u1181(.A(men_men_n1209_), .B(men_men_n1207_), .C(men_men_n1204_), .Y(men_men_n1210_));
  AOI210     u1182(.A0(men_men_n590_), .A1(men_men_n116_), .B0(men_men_n596_), .Y(men_men_n1211_));
  OAI210     u1183(.A0(men_men_n1195_), .A1(men_men_n587_), .B0(men_men_n1211_), .Y(men_men_n1212_));
  NA2        u1184(.A(men_men_n275_), .B(men_men_n194_), .Y(men_men_n1213_));
  NA2        u1185(.A(men_men_n1213_), .B(men_men_n662_), .Y(men_men_n1214_));
  NO3        u1186(.A(men_men_n815_), .B(men_men_n203_), .C(men_men_n396_), .Y(men_men_n1215_));
  NO2        u1187(.A(men_men_n1215_), .B(men_men_n935_), .Y(men_men_n1216_));
  NA2        u1188(.A(men_men_n1192_), .B(men_men_n670_), .Y(men_men_n1217_));
  NA4        u1189(.A(men_men_n1217_), .B(men_men_n1216_), .C(men_men_n1214_), .D(men_men_n783_), .Y(men_men_n1218_));
  NO3        u1190(.A(men_men_n1218_), .B(men_men_n1212_), .C(men_men_n1210_), .Y(men_men_n1219_));
  NA3        u1191(.A(men_men_n599_), .B(men_men_n29_), .C(f), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n1220_), .B(men_men_n203_), .Y(men_men_n1221_));
  AOI210     u1193(.A0(men_men_n492_), .A1(men_men_n56_), .B0(men_men_n1221_), .Y(men_men_n1222_));
  OR3        u1194(.A(men_men_n1191_), .B(men_men_n600_), .C(men_men_n1190_), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n1199_), .B(men_men_n954_), .Y(men_men_n1224_));
  NO2        u1196(.A(men_men_n206_), .B(men_men_n109_), .Y(men_men_n1225_));
  NO3        u1197(.A(men_men_n1225_), .B(men_men_n1224_), .C(men_men_n1132_), .Y(men_men_n1226_));
  NA4        u1198(.A(men_men_n1226_), .B(men_men_n1223_), .C(men_men_n1222_), .D(men_men_n754_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n942_), .B(men_men_n229_), .Y(men_men_n1228_));
  NO2        u1200(.A(men_men_n943_), .B(men_men_n546_), .Y(men_men_n1229_));
  OAI210     u1201(.A0(men_men_n1229_), .A1(men_men_n1228_), .B0(men_men_n326_), .Y(men_men_n1230_));
  NA2        u1202(.A(men_men_n563_), .B(men_men_n561_), .Y(men_men_n1231_));
  NO3        u1203(.A(men_men_n77_), .B(men_men_n294_), .C(men_men_n45_), .Y(men_men_n1232_));
  NA2        u1204(.A(men_men_n1232_), .B(men_men_n543_), .Y(men_men_n1233_));
  NA3        u1205(.A(men_men_n1233_), .B(men_men_n1231_), .C(men_men_n665_), .Y(men_men_n1234_));
  OR2        u1206(.A(men_men_n1136_), .B(men_men_n1129_), .Y(men_men_n1235_));
  NO2        u1207(.A(men_men_n356_), .B(men_men_n70_), .Y(men_men_n1236_));
  INV        u1208(.A(men_men_n1236_), .Y(men_men_n1237_));
  NA2        u1209(.A(men_men_n1232_), .B(men_men_n806_), .Y(men_men_n1238_));
  NA4        u1210(.A(men_men_n1238_), .B(men_men_n1237_), .C(men_men_n1235_), .D(men_men_n374_), .Y(men_men_n1239_));
  NOi41      u1211(.An(men_men_n1230_), .B(men_men_n1239_), .C(men_men_n1234_), .D(men_men_n1227_), .Y(men_men_n1240_));
  NO2        u1212(.A(men_men_n130_), .B(men_men_n45_), .Y(men_men_n1241_));
  AN2        u1213(.A(men_men_n1241_), .B(men_men_n699_), .Y(men_men_n1242_));
  NA2        u1214(.A(men_men_n1242_), .B(men_men_n326_), .Y(men_men_n1243_));
  INV        u1215(.A(men_men_n134_), .Y(men_men_n1244_));
  NO3        u1216(.A(men_men_n1059_), .B(men_men_n178_), .C(men_men_n85_), .Y(men_men_n1245_));
  AOI220     u1217(.A0(men_men_n1245_), .A1(men_men_n1244_), .B0(men_men_n1232_), .B1(men_men_n946_), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n1246_), .B(men_men_n1243_), .Y(men_men_n1247_));
  NO2        u1219(.A(men_men_n611_), .B(men_men_n610_), .Y(men_men_n1248_));
  NO4        u1220(.A(men_men_n1059_), .B(men_men_n1248_), .C(men_men_n176_), .D(men_men_n85_), .Y(men_men_n1249_));
  NO3        u1221(.A(men_men_n1249_), .B(men_men_n1247_), .C(men_men_n636_), .Y(men_men_n1250_));
  NA4        u1222(.A(men_men_n1250_), .B(men_men_n1240_), .C(men_men_n1219_), .D(men_men_n1202_), .Y(men06));
  NO2        u1223(.A(men_men_n397_), .B(men_men_n550_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n730_), .B(i), .Y(men_men_n1253_));
  OAI210     u1225(.A0(men_men_n1253_), .A1(men_men_n261_), .B0(men_men_n1252_), .Y(men_men_n1254_));
  NO2        u1226(.A(men_men_n224_), .B(men_men_n102_), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n1255_), .A1(men_men_n1245_), .B0(men_men_n370_), .Y(men_men_n1256_));
  NO3        u1228(.A(men_men_n594_), .B(men_men_n801_), .C(men_men_n597_), .Y(men_men_n1257_));
  OR2        u1229(.A(men_men_n1257_), .B(men_men_n875_), .Y(men_men_n1258_));
  NA4        u1230(.A(men_men_n1258_), .B(men_men_n1256_), .C(men_men_n1254_), .D(men_men_n1230_), .Y(men_men_n1259_));
  NO3        u1231(.A(men_men_n1259_), .B(men_men_n1234_), .C(men_men_n250_), .Y(men_men_n1260_));
  NO2        u1232(.A(men_men_n294_), .B(men_men_n45_), .Y(men_men_n1261_));
  AOI210     u1233(.A0(men_men_n1261_), .A1(men_men_n946_), .B0(men_men_n1228_), .Y(men_men_n1262_));
  AOI210     u1234(.A0(men_men_n1261_), .A1(men_men_n547_), .B0(men_men_n1242_), .Y(men_men_n1263_));
  AOI210     u1235(.A0(men_men_n1263_), .A1(men_men_n1262_), .B0(men_men_n324_), .Y(men_men_n1264_));
  OAI210     u1236(.A0(men_men_n87_), .A1(men_men_n40_), .B0(men_men_n668_), .Y(men_men_n1265_));
  NA2        u1237(.A(men_men_n1265_), .B(men_men_n640_), .Y(men_men_n1266_));
  NO2        u1238(.A(men_men_n502_), .B(men_men_n173_), .Y(men_men_n1267_));
  NO2        u1239(.A(men_men_n604_), .B(men_men_n1082_), .Y(men_men_n1268_));
  NO3        u1240(.A(men_men_n1268_), .B(men_men_n136_), .C(men_men_n1267_), .Y(men_men_n1269_));
  OR2        u1241(.A(men_men_n595_), .B(men_men_n593_), .Y(men_men_n1270_));
  NO2        u1242(.A(men_men_n355_), .B(men_men_n135_), .Y(men_men_n1271_));
  AOI210     u1243(.A0(men_men_n1271_), .A1(men_men_n581_), .B0(men_men_n1270_), .Y(men_men_n1272_));
  NA3        u1244(.A(men_men_n1272_), .B(men_men_n1269_), .C(men_men_n1266_), .Y(men_men_n1273_));
  NO2        u1245(.A(men_men_n745_), .B(men_men_n354_), .Y(men_men_n1274_));
  NOi21      u1246(.An(men_men_n1274_), .B(men_men_n49_), .Y(men_men_n1275_));
  AN2        u1247(.A(men_men_n931_), .B(men_men_n642_), .Y(men_men_n1276_));
  NO4        u1248(.A(men_men_n1276_), .B(men_men_n1275_), .C(men_men_n1273_), .D(men_men_n1264_), .Y(men_men_n1277_));
  NO2        u1249(.A(men_men_n796_), .B(men_men_n271_), .Y(men_men_n1278_));
  OAI220     u1250(.A0(men_men_n730_), .A1(men_men_n47_), .B0(men_men_n224_), .B1(men_men_n613_), .Y(men_men_n1279_));
  NO2        u1251(.A(men_men_n271_), .B(c), .Y(men_men_n1280_));
  AOI220     u1252(.A0(men_men_n1280_), .A1(men_men_n1279_), .B0(men_men_n1278_), .B1(men_men_n261_), .Y(men_men_n1281_));
  NO3        u1253(.A(men_men_n241_), .B(men_men_n102_), .C(men_men_n276_), .Y(men_men_n1282_));
  OAI210     u1254(.A0(l), .A1(i), .B0(k), .Y(men_men_n1283_));
  NO3        u1255(.A(men_men_n1283_), .B(men_men_n592_), .C(j), .Y(men_men_n1284_));
  NOi21      u1256(.An(men_men_n1284_), .B(men_men_n70_), .Y(men_men_n1285_));
  NO3        u1257(.A(men_men_n1285_), .B(men_men_n1282_), .C(men_men_n1085_), .Y(men_men_n1286_));
  NAi31      u1258(.An(men_men_n745_), .B(men_men_n420_), .C(men_men_n202_), .Y(men_men_n1287_));
  NA3        u1259(.A(men_men_n1287_), .B(men_men_n1286_), .C(men_men_n1281_), .Y(men_men_n1288_));
  NOi31      u1260(.An(men_men_n1257_), .B(men_men_n448_), .C(men_men_n383_), .Y(men_men_n1289_));
  OR3        u1261(.A(men_men_n1289_), .B(men_men_n780_), .C(men_men_n530_), .Y(men_men_n1290_));
  AOI210     u1262(.A0(men_men_n563_), .A1(men_men_n432_), .B0(men_men_n360_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n1284_), .B(men_men_n787_), .Y(men_men_n1292_));
  NA3        u1264(.A(men_men_n1292_), .B(men_men_n1291_), .C(men_men_n1290_), .Y(men_men_n1293_));
  NA2        u1265(.A(men_men_n1271_), .B(men_men_n235_), .Y(men_men_n1294_));
  NO2        u1266(.A(men_men_n867_), .B(men_men_n468_), .Y(men_men_n1295_));
  NA3        u1267(.A(men_men_n1295_), .B(men_men_n1294_), .C(men_men_n1238_), .Y(men_men_n1296_));
  NAi21      u1268(.An(j), .B(i), .Y(men_men_n1297_));
  NO4        u1269(.A(men_men_n1248_), .B(men_men_n1297_), .C(men_men_n428_), .D(men_men_n232_), .Y(men_men_n1298_));
  NO4        u1270(.A(men_men_n1298_), .B(men_men_n1296_), .C(men_men_n1293_), .D(men_men_n1288_), .Y(men_men_n1299_));
  NA4        u1271(.A(men_men_n1299_), .B(men_men_n1277_), .C(men_men_n1260_), .D(men_men_n1250_), .Y(men07));
  NOi21      u1272(.An(j), .B(k), .Y(men_men_n1301_));
  NAi32      u1273(.An(m), .Bn(b), .C(n), .Y(men_men_n1302_));
  NO3        u1274(.A(men_men_n1302_), .B(g), .C(f), .Y(men_men_n1303_));
  OAI210     u1275(.A0(i), .A1(men_men_n470_), .B0(men_men_n1303_), .Y(men_men_n1304_));
  NAi21      u1276(.An(f), .B(c), .Y(men_men_n1305_));
  OR2        u1277(.A(e), .B(d), .Y(men_men_n1306_));
  NOi31      u1278(.An(n), .B(m), .C(b), .Y(men_men_n1307_));
  INV        u1279(.A(men_men_n1304_), .Y(men_men_n1308_));
  NOi41      u1280(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1309_));
  NA3        u1281(.A(men_men_n1309_), .B(men_men_n860_), .C(men_men_n399_), .Y(men_men_n1310_));
  INV        u1282(.A(men_men_n1310_), .Y(men_men_n1311_));
  NA2        u1283(.A(men_men_n1061_), .B(men_men_n221_), .Y(men_men_n1312_));
  NO2        u1284(.A(men_men_n1312_), .B(men_men_n59_), .Y(men_men_n1313_));
  NO2        u1285(.A(k), .B(i), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n1176_), .B(men_men_n284_), .Y(men_men_n1315_));
  INV        u1287(.A(men_men_n1315_), .Y(men_men_n1316_));
  NO4        u1288(.A(men_men_n1316_), .B(men_men_n1313_), .C(men_men_n1311_), .D(men_men_n1308_), .Y(men_men_n1317_));
  NO3        u1289(.A(e), .B(d), .C(c), .Y(men_men_n1318_));
  OAI210     u1290(.A0(men_men_n131_), .A1(men_men_n214_), .B0(men_men_n601_), .Y(men_men_n1319_));
  NA2        u1291(.A(men_men_n1319_), .B(men_men_n1318_), .Y(men_men_n1320_));
  INV        u1292(.A(men_men_n1320_), .Y(men_men_n1321_));
  OR2        u1293(.A(h), .B(f), .Y(men_men_n1322_));
  NO3        u1294(.A(n), .B(m), .C(i), .Y(men_men_n1323_));
  OAI210     u1295(.A0(men_men_n1083_), .A1(men_men_n158_), .B0(men_men_n1323_), .Y(men_men_n1324_));
  NO2        u1296(.A(i), .B(g), .Y(men_men_n1325_));
  OR3        u1297(.A(men_men_n1325_), .B(men_men_n1302_), .C(men_men_n69_), .Y(men_men_n1326_));
  OAI220     u1298(.A0(men_men_n1326_), .A1(men_men_n470_), .B0(men_men_n1324_), .B1(men_men_n1322_), .Y(men_men_n1327_));
  NA3        u1299(.A(men_men_n689_), .B(men_men_n675_), .C(men_men_n110_), .Y(men_men_n1328_));
  NA3        u1300(.A(men_men_n1307_), .B(men_men_n1031_), .C(h), .Y(men_men_n1329_));
  AOI210     u1301(.A0(men_men_n1329_), .A1(men_men_n1328_), .B0(men_men_n45_), .Y(men_men_n1330_));
  NA2        u1302(.A(men_men_n1323_), .B(men_men_n638_), .Y(men_men_n1331_));
  NO2        u1303(.A(l), .B(k), .Y(men_men_n1332_));
  NO3        u1304(.A(men_men_n428_), .B(d), .C(c), .Y(men_men_n1333_));
  NO3        u1305(.A(men_men_n1330_), .B(men_men_n1327_), .C(men_men_n1321_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n148_), .B(h), .Y(men_men_n1335_));
  NO2        u1307(.A(g), .B(c), .Y(men_men_n1336_));
  NO2        u1308(.A(men_men_n436_), .B(a), .Y(men_men_n1337_));
  NA3        u1309(.A(men_men_n1337_), .B(men_men_n1482_), .C(men_men_n111_), .Y(men_men_n1338_));
  NO2        u1310(.A(i), .B(h), .Y(men_men_n1339_));
  NA2        u1311(.A(men_men_n1339_), .B(men_men_n221_), .Y(men_men_n1340_));
  AOI210     u1312(.A0(men_men_n251_), .A1(men_men_n114_), .B0(men_men_n519_), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n1341_), .B(men_men_n1340_), .Y(men_men_n1342_));
  NO2        u1314(.A(men_men_n752_), .B(men_men_n188_), .Y(men_men_n1343_));
  NOi31      u1315(.An(m), .B(n), .C(b), .Y(men_men_n1344_));
  NOi31      u1316(.An(f), .B(d), .C(c), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n1345_), .B(men_men_n1344_), .Y(men_men_n1346_));
  INV        u1318(.A(men_men_n1346_), .Y(men_men_n1347_));
  NO3        u1319(.A(men_men_n1347_), .B(men_men_n1343_), .C(men_men_n1342_), .Y(men_men_n1348_));
  OAI210     u1320(.A0(men_men_n184_), .A1(men_men_n514_), .B0(men_men_n1032_), .Y(men_men_n1349_));
  NO3        u1321(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1350_));
  AN3        u1322(.A(men_men_n1349_), .B(men_men_n1348_), .C(men_men_n1338_), .Y(men_men_n1351_));
  NA2        u1323(.A(men_men_n1307_), .B(men_men_n367_), .Y(men_men_n1352_));
  NO2        u1324(.A(men_men_n1352_), .B(men_men_n1014_), .Y(men_men_n1353_));
  NA2        u1325(.A(men_men_n1333_), .B(men_men_n215_), .Y(men_men_n1354_));
  NO2        u1326(.A(men_men_n188_), .B(b), .Y(men_men_n1355_));
  NO2        u1327(.A(i), .B(men_men_n213_), .Y(men_men_n1356_));
  NA4        u1328(.A(men_men_n1108_), .B(men_men_n1356_), .C(men_men_n103_), .D(m), .Y(men_men_n1357_));
  NAi31      u1329(.An(men_men_n1353_), .B(men_men_n1357_), .C(men_men_n1354_), .Y(men_men_n1358_));
  NO4        u1330(.A(men_men_n131_), .B(g), .C(f), .D(e), .Y(men_men_n1359_));
  NA2        u1331(.A(men_men_n1314_), .B(h), .Y(men_men_n1360_));
  NA2        u1332(.A(men_men_n193_), .B(men_men_n97_), .Y(men_men_n1361_));
  NOi41      u1333(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1362_));
  NA2        u1334(.A(men_men_n1362_), .B(men_men_n111_), .Y(men_men_n1363_));
  NA2        u1335(.A(men_men_n1309_), .B(men_men_n1332_), .Y(men_men_n1364_));
  NA2        u1336(.A(men_men_n1364_), .B(men_men_n1363_), .Y(men_men_n1365_));
  OR3        u1337(.A(men_men_n530_), .B(men_men_n529_), .C(men_men_n110_), .Y(men_men_n1366_));
  NA2        u1338(.A(men_men_n1081_), .B(men_men_n396_), .Y(men_men_n1367_));
  OAI220     u1339(.A0(men_men_n1367_), .A1(men_men_n421_), .B0(men_men_n1366_), .B1(men_men_n294_), .Y(men_men_n1368_));
  AO210      u1340(.A0(men_men_n1368_), .A1(men_men_n114_), .B0(men_men_n1365_), .Y(men_men_n1369_));
  NO2        u1341(.A(men_men_n1369_), .B(men_men_n1358_), .Y(men_men_n1370_));
  NA4        u1342(.A(men_men_n1370_), .B(men_men_n1351_), .C(men_men_n1334_), .D(men_men_n1317_), .Y(men_men_n1371_));
  NO2        u1343(.A(men_men_n1096_), .B(men_men_n108_), .Y(men_men_n1372_));
  NA2        u1344(.A(men_men_n367_), .B(men_men_n54_), .Y(men_men_n1373_));
  NO2        u1345(.A(men_men_n1373_), .B(men_men_n1331_), .Y(men_men_n1374_));
  NA2        u1346(.A(men_men_n215_), .B(men_men_n181_), .Y(men_men_n1375_));
  AOI210     u1347(.A0(men_men_n1375_), .A1(men_men_n1150_), .B0(men_men_n1373_), .Y(men_men_n1376_));
  NO2        u1348(.A(men_men_n1054_), .B(men_men_n1050_), .Y(men_men_n1377_));
  NO3        u1349(.A(men_men_n1377_), .B(men_men_n1376_), .C(men_men_n1374_), .Y(men_men_n1378_));
  NO2        u1350(.A(men_men_n379_), .B(j), .Y(men_men_n1379_));
  NA3        u1351(.A(men_men_n1350_), .B(men_men_n1306_), .C(men_men_n1081_), .Y(men_men_n1380_));
  NAi41      u1352(.An(men_men_n1339_), .B(men_men_n1043_), .C(men_men_n170_), .D(men_men_n151_), .Y(men_men_n1381_));
  NA2        u1353(.A(men_men_n1381_), .B(men_men_n1380_), .Y(men_men_n1382_));
  NA3        u1354(.A(g), .B(men_men_n1379_), .C(men_men_n160_), .Y(men_men_n1383_));
  INV        u1355(.A(men_men_n1383_), .Y(men_men_n1384_));
  NO3        u1356(.A(men_men_n745_), .B(men_men_n176_), .C(men_men_n399_), .Y(men_men_n1385_));
  NO3        u1357(.A(men_men_n1385_), .B(men_men_n1384_), .C(men_men_n1382_), .Y(men_men_n1386_));
  NO3        u1358(.A(men_men_n1050_), .B(men_men_n575_), .C(g), .Y(men_men_n1387_));
  NOi21      u1359(.An(men_men_n1375_), .B(men_men_n1387_), .Y(men_men_n1388_));
  AOI210     u1360(.A0(men_men_n1388_), .A1(men_men_n1361_), .B0(men_men_n1023_), .Y(men_men_n1389_));
  OR2        u1361(.A(n), .B(i), .Y(men_men_n1390_));
  OAI210     u1362(.A0(men_men_n1390_), .A1(men_men_n1042_), .B0(men_men_n49_), .Y(men_men_n1391_));
  AOI220     u1363(.A0(men_men_n1391_), .A1(men_men_n1138_), .B0(men_men_n820_), .B1(men_men_n193_), .Y(men_men_n1392_));
  INV        u1364(.A(men_men_n1392_), .Y(men_men_n1393_));
  OAI220     u1365(.A0(men_men_n663_), .A1(g), .B0(men_men_n224_), .B1(c), .Y(men_men_n1394_));
  AOI210     u1366(.A0(men_men_n1355_), .A1(men_men_n41_), .B0(men_men_n1394_), .Y(men_men_n1395_));
  NO2        u1367(.A(men_men_n224_), .B(k), .Y(men_men_n1396_));
  NO2        u1368(.A(men_men_n1395_), .B(men_men_n178_), .Y(men_men_n1397_));
  NO3        u1369(.A(men_men_n1366_), .B(men_men_n451_), .C(men_men_n339_), .Y(men_men_n1398_));
  NO4        u1370(.A(men_men_n1398_), .B(men_men_n1397_), .C(men_men_n1393_), .D(men_men_n1389_), .Y(men_men_n1399_));
  INV        u1371(.A(men_men_n49_), .Y(men_men_n1400_));
  NO3        u1372(.A(men_men_n1063_), .B(men_men_n1306_), .C(men_men_n49_), .Y(men_men_n1401_));
  NA2        u1373(.A(men_men_n1064_), .B(men_men_n1400_), .Y(men_men_n1402_));
  NO2        u1374(.A(men_men_n1402_), .B(j), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1372_), .B(men_men_n451_), .C(f), .Y(men_men_n1404_));
  NA2        u1376(.A(men_men_n181_), .B(men_men_n110_), .Y(men_men_n1405_));
  NO2        u1377(.A(men_men_n1301_), .B(men_men_n42_), .Y(men_men_n1406_));
  AOI210     u1378(.A0(men_men_n111_), .A1(men_men_n40_), .B0(men_men_n1406_), .Y(men_men_n1407_));
  NO2        u1379(.A(men_men_n1407_), .B(men_men_n1404_), .Y(men_men_n1408_));
  AOI210     u1380(.A0(men_men_n514_), .A1(h), .B0(men_men_n67_), .Y(men_men_n1409_));
  NA2        u1381(.A(men_men_n1409_), .B(men_men_n1337_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1297_), .B(men_men_n176_), .Y(men_men_n1411_));
  NOi21      u1383(.An(d), .B(f), .Y(men_men_n1412_));
  NO3        u1384(.A(men_men_n1345_), .B(men_men_n1412_), .C(men_men_n40_), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n1413_), .B(men_men_n1411_), .Y(men_men_n1414_));
  NA2        u1386(.A(men_men_n1337_), .B(men_men_n1406_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n294_), .B(c), .Y(men_men_n1416_));
  NA2        u1388(.A(men_men_n1416_), .B(men_men_n531_), .Y(men_men_n1417_));
  NA4        u1389(.A(men_men_n1417_), .B(men_men_n1415_), .C(men_men_n1414_), .D(men_men_n1410_), .Y(men_men_n1418_));
  NO3        u1390(.A(men_men_n1418_), .B(men_men_n1408_), .C(men_men_n1403_), .Y(men_men_n1419_));
  NA4        u1391(.A(men_men_n1419_), .B(men_men_n1399_), .C(men_men_n1386_), .D(men_men_n1378_), .Y(men_men_n1420_));
  OAI210     u1392(.A0(men_men_n1359_), .A1(men_men_n1307_), .B0(men_men_n872_), .Y(men_men_n1421_));
  OAI220     u1393(.A0(men_men_n1011_), .A1(men_men_n131_), .B0(men_men_n663_), .B1(men_men_n176_), .Y(men_men_n1422_));
  NA2        u1394(.A(men_men_n1422_), .B(men_men_n619_), .Y(men_men_n1423_));
  NA2        u1395(.A(men_men_n1423_), .B(men_men_n1421_), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n1336_), .B(men_men_n1412_), .Y(men_men_n1425_));
  NO2        u1397(.A(men_men_n1425_), .B(m), .Y(men_men_n1426_));
  NA3        u1398(.A(men_men_n1061_), .B(men_men_n106_), .C(men_men_n221_), .Y(men_men_n1427_));
  NO2        u1399(.A(men_men_n152_), .B(men_men_n183_), .Y(men_men_n1428_));
  OAI210     u1400(.A0(men_men_n1428_), .A1(men_men_n108_), .B0(men_men_n1344_), .Y(men_men_n1429_));
  NA2        u1401(.A(men_men_n1429_), .B(men_men_n1427_), .Y(men_men_n1430_));
  NO3        u1402(.A(men_men_n1430_), .B(men_men_n1426_), .C(men_men_n1424_), .Y(men_men_n1431_));
  NO2        u1403(.A(men_men_n1305_), .B(e), .Y(men_men_n1432_));
  NA2        u1404(.A(men_men_n1432_), .B(men_men_n394_), .Y(men_men_n1433_));
  NA2        u1405(.A(men_men_n1091_), .B(men_men_n628_), .Y(men_men_n1434_));
  OR3        u1406(.A(men_men_n1396_), .B(men_men_n1176_), .C(men_men_n131_), .Y(men_men_n1435_));
  OAI220     u1407(.A0(men_men_n1435_), .A1(men_men_n1433_), .B0(men_men_n1434_), .B1(men_men_n430_), .Y(men_men_n1436_));
  NO2        u1408(.A(men_men_n1366_), .B(a), .Y(men_men_n1437_));
  NO2        u1409(.A(men_men_n1437_), .B(men_men_n1436_), .Y(men_men_n1438_));
  NA2        u1410(.A(men_men_n1432_), .B(men_men_n181_), .Y(men_men_n1439_));
  AOI220     u1411(.A0(men_men_n1439_), .A1(men_men_n1044_), .B0(men_men_n521_), .B1(men_men_n354_), .Y(men_men_n1440_));
  NA2        u1412(.A(men_men_n529_), .B(g), .Y(men_men_n1441_));
  AOI210     u1413(.A0(men_men_n1441_), .A1(men_men_n1333_), .B0(men_men_n1401_), .Y(men_men_n1442_));
  NO2        u1414(.A(men_men_n1442_), .B(men_men_n213_), .Y(men_men_n1443_));
  AOI210     u1415(.A0(men_men_n886_), .A1(men_men_n405_), .B0(men_men_n104_), .Y(men_men_n1444_));
  OR2        u1416(.A(men_men_n1444_), .B(men_men_n529_), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n1445_), .B(men_men_n176_), .Y(men_men_n1446_));
  NO2        u1418(.A(men_men_n49_), .B(l), .Y(men_men_n1447_));
  INV        u1419(.A(men_men_n470_), .Y(men_men_n1448_));
  OAI210     u1420(.A0(men_men_n1448_), .A1(men_men_n1064_), .B0(men_men_n1447_), .Y(men_men_n1449_));
  NO2        u1421(.A(m), .B(i), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1450_), .B(men_men_n1335_), .Y(men_men_n1451_));
  NA2        u1423(.A(men_men_n1451_), .B(men_men_n1449_), .Y(men_men_n1452_));
  NO4        u1424(.A(men_men_n1452_), .B(men_men_n1446_), .C(men_men_n1443_), .D(men_men_n1440_), .Y(men_men_n1453_));
  NA3        u1425(.A(men_men_n1453_), .B(men_men_n1438_), .C(men_men_n1431_), .Y(men_men_n1454_));
  NA3        u1426(.A(men_men_n937_), .B(men_men_n138_), .C(men_men_n46_), .Y(men_men_n1455_));
  AOI210     u1427(.A0(men_men_n149_), .A1(c), .B0(men_men_n1455_), .Y(men_men_n1456_));
  AO210      u1428(.A0(men_men_n132_), .A1(l), .B0(men_men_n1352_), .Y(men_men_n1457_));
  NO2        u1429(.A(men_men_n69_), .B(c), .Y(men_men_n1458_));
  NO4        u1430(.A(men_men_n1322_), .B(men_men_n187_), .C(men_men_n434_), .D(men_men_n45_), .Y(men_men_n1459_));
  AOI210     u1431(.A0(men_men_n1411_), .A1(men_men_n1458_), .B0(men_men_n1459_), .Y(men_men_n1460_));
  NA2        u1432(.A(men_men_n1460_), .B(men_men_n1457_), .Y(men_men_n1461_));
  NO2        u1433(.A(men_men_n1461_), .B(men_men_n1456_), .Y(men_men_n1462_));
  NO4        u1434(.A(men_men_n224_), .B(men_men_n187_), .C(men_men_n251_), .D(k), .Y(men_men_n1463_));
  AOI210     u1435(.A0(men_men_n158_), .A1(men_men_n54_), .B0(men_men_n1432_), .Y(men_men_n1464_));
  NO2        u1436(.A(men_men_n1464_), .B(men_men_n1405_), .Y(men_men_n1465_));
  NO2        u1437(.A(men_men_n1455_), .B(men_men_n108_), .Y(men_men_n1466_));
  NO3        u1438(.A(men_men_n1466_), .B(men_men_n1465_), .C(men_men_n1463_), .Y(men_men_n1467_));
  NO2        u1439(.A(men_men_n1404_), .B(men_men_n67_), .Y(men_men_n1468_));
  INV        u1440(.A(men_men_n1468_), .Y(men_men_n1469_));
  NA3        u1441(.A(men_men_n1469_), .B(men_men_n1467_), .C(men_men_n1462_), .Y(men_men_n1470_));
  OR4        u1442(.A(men_men_n1470_), .B(men_men_n1454_), .C(men_men_n1420_), .D(men_men_n1371_), .Y(men04));
  NOi31      u1443(.An(men_men_n1359_), .B(men_men_n1360_), .C(men_men_n1017_), .Y(men_men_n1472_));
  NO4        u1444(.A(men_men_n266_), .B(men_men_n1007_), .C(men_men_n471_), .D(j), .Y(men_men_n1473_));
  OR3        u1445(.A(men_men_n1473_), .B(men_men_n1472_), .C(men_men_n1034_), .Y(men_men_n1474_));
  NO2        u1446(.A(men_men_n89_), .B(k), .Y(men_men_n1475_));
  AOI210     u1447(.A0(men_men_n1475_), .A1(men_men_n1028_), .B0(men_men_n1152_), .Y(men_men_n1476_));
  NA2        u1448(.A(men_men_n1476_), .B(men_men_n1178_), .Y(men_men_n1477_));
  NO3        u1449(.A(men_men_n1477_), .B(men_men_n1474_), .C(men_men_n1022_), .Y(men_men_n1478_));
  NA4        u1450(.A(men_men_n1478_), .B(men_men_n1093_), .C(men_men_n1079_), .D(men_men_n1067_), .Y(men05));
  INV        u1451(.A(i), .Y(men_men_n1482_));
  INV        u1452(.A(men_men_n885_), .Y(men_men_n1483_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule