//Benchmark atmr_alu4_1266_0.25

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n107_, ori_ori_n108_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n325_, ori_ori_n326_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NAi31      o017(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n35_), .Y(ori1));
  INV        o019(.A(i_11_), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n43_));
  INV        o021(.A(i_2_), .Y(ori_ori_n44_));
  INV        o022(.A(i_5_), .Y(ori_ori_n45_));
  NO2        o023(.A(i_7_), .B(i_10_), .Y(ori_ori_n46_));
  AOI210     o024(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n46_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_5_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NA2        o026(.A(i_7_), .B(i_9_), .Y(ori_ori_n49_));
  NA2        o027(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n50_));
  NO2        o028(.A(i_1_), .B(i_6_), .Y(ori_ori_n51_));
  NAi21      o029(.An(i_2_), .B(i_7_), .Y(ori_ori_n52_));
  INV        o030(.A(i_1_), .Y(ori_ori_n53_));
  NA2        o031(.A(ori_ori_n53_), .B(i_6_), .Y(ori_ori_n54_));
  NA3        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .C(ori_ori_n31_), .Y(ori_ori_n55_));
  NA2        o033(.A(i_1_), .B(i_10_), .Y(ori_ori_n56_));
  NO2        o034(.A(ori_ori_n56_), .B(i_6_), .Y(ori_ori_n57_));
  NAi21      o035(.An(ori_ori_n57_), .B(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n47_), .B(i_2_), .Y(ori_ori_n59_));
  AOI210     o037(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n60_));
  NA2        o038(.A(i_1_), .B(i_6_), .Y(ori_ori_n61_));
  NO2        o039(.A(ori_ori_n61_), .B(ori_ori_n25_), .Y(ori_ori_n62_));
  INV        o040(.A(i_0_), .Y(ori_ori_n63_));
  NAi21      o041(.An(i_5_), .B(i_10_), .Y(ori_ori_n64_));
  NA2        o042(.A(i_5_), .B(i_9_), .Y(ori_ori_n65_));
  AOI210     o043(.A0(ori_ori_n65_), .A1(ori_ori_n64_), .B0(ori_ori_n63_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(ori_ori_n62_), .Y(ori_ori_n67_));
  OAI210     o045(.A0(ori_ori_n60_), .A1(ori_ori_n59_), .B0(ori_ori_n67_), .Y(ori_ori_n68_));
  OAI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n58_), .B0(i_0_), .Y(ori_ori_n69_));
  NA2        o047(.A(i_12_), .B(i_5_), .Y(ori_ori_n70_));
  INV        o048(.A(i_6_), .Y(ori_ori_n71_));
  NO2        o049(.A(i_2_), .B(i_7_), .Y(ori_ori_n72_));
  INV        o050(.A(ori_ori_n72_), .Y(ori_ori_n73_));
  NA2        o051(.A(i_1_), .B(ori_ori_n73_), .Y(ori_ori_n74_));
  NAi21      o052(.An(i_6_), .B(i_10_), .Y(ori_ori_n75_));
  NA2        o053(.A(i_6_), .B(i_9_), .Y(ori_ori_n76_));
  AOI210     o054(.A0(ori_ori_n76_), .A1(ori_ori_n75_), .B0(ori_ori_n53_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_2_), .B(i_6_), .Y(ori_ori_n78_));
  INV        o056(.A(ori_ori_n77_), .Y(ori_ori_n79_));
  AOI210     o057(.A0(ori_ori_n79_), .A1(ori_ori_n74_), .B0(ori_ori_n70_), .Y(ori_ori_n80_));
  AN3        o058(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n81_));
  NAi21      o059(.An(i_6_), .B(i_11_), .Y(ori_ori_n82_));
  NA2        o060(.A(ori_ori_n81_), .B(ori_ori_n32_), .Y(ori_ori_n83_));
  INV        o061(.A(i_7_), .Y(ori_ori_n84_));
  NA2        o062(.A(ori_ori_n44_), .B(ori_ori_n84_), .Y(ori_ori_n85_));
  NO2        o063(.A(i_0_), .B(i_5_), .Y(ori_ori_n86_));
  NO2        o064(.A(ori_ori_n86_), .B(ori_ori_n71_), .Y(ori_ori_n87_));
  NA3        o065(.A(i_12_), .B(ori_ori_n87_), .C(ori_ori_n85_), .Y(ori_ori_n88_));
  INV        o066(.A(i_7_), .Y(ori_ori_n89_));
  OR2        o067(.A(ori_ori_n70_), .B(ori_ori_n51_), .Y(ori_ori_n90_));
  NA2        o068(.A(i_12_), .B(i_7_), .Y(ori_ori_n91_));
  NA2        o069(.A(i_11_), .B(i_12_), .Y(ori_ori_n92_));
  NA3        o070(.A(ori_ori_n92_), .B(ori_ori_n88_), .C(ori_ori_n83_), .Y(ori_ori_n93_));
  NOi21      o071(.An(i_1_), .B(i_5_), .Y(ori_ori_n94_));
  NA2        o072(.A(ori_ori_n94_), .B(i_11_), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n84_), .B(ori_ori_n37_), .Y(ori_ori_n96_));
  NA2        o074(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n97_), .B(ori_ori_n96_), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n98_), .B(ori_ori_n44_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n100_));
  INV        o078(.A(ori_ori_n52_), .Y(ori_ori_n101_));
  NOi21      o079(.An(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NO2        o080(.A(i_1_), .B(ori_ori_n71_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n102_), .B(ori_ori_n95_), .Y(ori_ori_n104_));
  NO3        o082(.A(ori_ori_n104_), .B(ori_ori_n93_), .C(ori_ori_n80_), .Y(ori_ori_n105_));
  NA3        o083(.A(ori_ori_n105_), .B(ori_ori_n69_), .C(ori_ori_n50_), .Y(ori2));
  NO2        o084(.A(ori_ori_n53_), .B(ori_ori_n37_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n325_), .B(ori_ori_n107_), .Y(ori_ori_n108_));
  NA4        o086(.A(ori_ori_n108_), .B(ori_ori_n67_), .C(ori_ori_n59_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o087(.A(i_0_), .B(i_1_), .Y(ori_ori_n110_));
  NA2        o088(.A(i_2_), .B(i_3_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(i_4_), .Y(ori_ori_n112_));
  NA2        o090(.A(i_1_), .B(i_5_), .Y(ori_ori_n113_));
  NOi21      o091(.An(i_4_), .B(i_10_), .Y(ori_ori_n114_));
  NOi21      o092(.An(i_4_), .B(i_9_), .Y(ori_ori_n115_));
  NOi21      o093(.An(i_11_), .B(i_13_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n63_), .B(ori_ori_n53_), .Y(ori_ori_n117_));
  NAi21      o095(.An(i_4_), .B(i_12_), .Y(ori_ori_n118_));
  INV        o096(.A(i_8_), .Y(ori_ori_n119_));
  NO3        o097(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n120_));
  NO2        o098(.A(i_13_), .B(i_9_), .Y(ori_ori_n121_));
  NAi21      o099(.An(i_12_), .B(i_3_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n42_), .B(i_5_), .Y(ori_ori_n123_));
  INV        o101(.A(i_13_), .Y(ori_ori_n124_));
  NO2        o102(.A(i_12_), .B(ori_ori_n124_), .Y(ori_ori_n125_));
  NO2        o103(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n126_));
  INV        o104(.A(i_12_), .Y(ori_ori_n127_));
  NO3        o105(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n128_));
  NAi21      o106(.An(i_4_), .B(i_3_), .Y(ori_ori_n129_));
  INV        o107(.A(i_0_), .Y(ori_ori_n130_));
  NO2        o108(.A(i_11_), .B(ori_ori_n124_), .Y(ori_ori_n131_));
  NA2        o109(.A(i_12_), .B(i_6_), .Y(ori_ori_n132_));
  OR2        o110(.A(i_13_), .B(i_9_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n129_), .B(i_2_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_2_), .B(ori_ori_n84_), .Y(ori_ori_n135_));
  AN2        o113(.A(i_3_), .B(i_10_), .Y(ori_ori_n136_));
  NO2        o114(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n44_), .B(ori_ori_n26_), .Y(ori_ori_n138_));
  NO2        o116(.A(i_2_), .B(i_3_), .Y(ori_ori_n139_));
  NO2        o117(.A(i_12_), .B(i_10_), .Y(ori_ori_n140_));
  NOi21      o118(.An(i_5_), .B(i_0_), .Y(ori_ori_n141_));
  NAi21      o119(.An(i_3_), .B(i_4_), .Y(ori_ori_n142_));
  AN2        o120(.A(i_12_), .B(i_5_), .Y(ori_ori_n143_));
  NO2        o121(.A(i_5_), .B(i_10_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n145_));
  NO3        o123(.A(ori_ori_n71_), .B(ori_ori_n45_), .C(i_9_), .Y(ori_ori_n146_));
  NO2        o124(.A(i_0_), .B(i_11_), .Y(ori_ori_n147_));
  NOi21      o125(.An(i_2_), .B(i_12_), .Y(ori_ori_n148_));
  NAi21      o126(.An(i_9_), .B(i_4_), .Y(ori_ori_n149_));
  OR2        o127(.A(i_13_), .B(i_10_), .Y(ori_ori_n150_));
  NO3        o128(.A(ori_ori_n150_), .B(ori_ori_n92_), .C(ori_ori_n149_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n84_), .B(ori_ori_n25_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n63_), .B(i_13_), .Y(ori_ori_n153_));
  NO2        o131(.A(i_10_), .B(i_9_), .Y(ori_ori_n154_));
  NO3        o132(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n132_), .B(ori_ori_n82_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n156_), .B(ori_ori_n155_), .Y(ori_ori_n157_));
  NA2        o135(.A(ori_ori_n131_), .B(ori_ori_n137_), .Y(ori_ori_n158_));
  NO3        o136(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n159_));
  INV        o137(.A(ori_ori_n159_), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n160_), .B(ori_ori_n158_), .Y(ori_ori_n161_));
  INV        o139(.A(ori_ori_n161_), .Y(ori_ori_n162_));
  NO2        o140(.A(i_11_), .B(i_1_), .Y(ori_ori_n163_));
  NA3        o141(.A(ori_ori_n145_), .B(ori_ori_n117_), .C(ori_ori_n112_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n155_), .B(ori_ori_n143_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n159_), .B(ori_ori_n144_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n164_), .B(ori_ori_n162_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n168_));
  AOI210     o146(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n151_), .Y(ori_ori_n169_));
  INV        o147(.A(ori_ori_n169_), .Y(ori_ori_n170_));
  NO3        o148(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n150_), .B(i_1_), .Y(ori_ori_n172_));
  NOi31      o150(.An(ori_ori_n172_), .B(ori_ori_n156_), .C(ori_ori_n63_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n91_), .B(ori_ori_n23_), .Y(ori_ori_n174_));
  NO2        o152(.A(i_12_), .B(ori_ori_n71_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n170_), .B(ori_ori_n167_), .Y(ori_ori_n176_));
  INV        o154(.A(ori_ori_n176_), .Y(ori7));
  NO2        o155(.A(ori_ori_n78_), .B(ori_ori_n49_), .Y(ori_ori_n178_));
  NA2        o156(.A(i_11_), .B(ori_ori_n119_), .Y(ori_ori_n179_));
  NA2        o157(.A(i_2_), .B(ori_ori_n71_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n72_), .B(ori_ori_n120_), .Y(ori_ori_n181_));
  INV        o159(.A(i_10_), .Y(ori_ori_n182_));
  OAI220     o160(.A0(ori_ori_n182_), .A1(ori_ori_n180_), .B0(ori_ori_n181_), .B1(i_13_), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n183_), .B(ori_ori_n178_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n52_), .B(i_10_), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n185_), .A1(ori_ori_n127_), .B0(ori_ori_n114_), .Y(ori_ori_n186_));
  OR2        o164(.A(ori_ori_n186_), .B(ori_ori_n133_), .Y(ori_ori_n187_));
  AOI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n184_), .B0(ori_ori_n53_), .Y(ori_ori_n188_));
  NOi21      o166(.An(i_11_), .B(i_7_), .Y(ori_ori_n189_));
  AO210      o167(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n190_), .B(ori_ori_n189_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n125_), .B(ori_ori_n53_), .Y(ori_ori_n192_));
  NO2        o170(.A(i_1_), .B(i_12_), .Y(ori_ori_n193_));
  INV        o171(.A(ori_ori_n192_), .Y(ori_ori_n194_));
  NA2        o172(.A(ori_ori_n194_), .B(i_6_), .Y(ori_ori_n195_));
  NO2        o173(.A(i_6_), .B(i_11_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n157_), .Y(ori_ori_n197_));
  INV        o175(.A(i_2_), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n107_), .B(i_9_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .Y(ori_ori_n200_));
  AOI210     o178(.A0(ori_ori_n163_), .A1(ori_ori_n152_), .B0(ori_ori_n128_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n180_), .Y(ori_ori_n202_));
  NO2        o180(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n203_));
  OR2        o181(.A(ori_ori_n202_), .B(ori_ori_n200_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(ori_ori_n197_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n127_), .B(ori_ori_n84_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(ori_ori_n189_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_7_), .B(ori_ori_n42_), .Y(ori_ori_n208_));
  NO3        o186(.A(ori_ori_n208_), .B(ori_ori_n138_), .C(i_12_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n92_), .B(ori_ori_n37_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n210_), .B(i_6_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n71_), .B(i_9_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n212_), .B(ori_ori_n53_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n213_), .B(ori_ori_n193_), .Y(ori_ori_n214_));
  NO4        o192(.A(ori_ori_n214_), .B(ori_ori_n211_), .C(ori_ori_n209_), .D(i_4_), .Y(ori_ori_n215_));
  INV        o193(.A(ori_ori_n215_), .Y(ori_ori_n216_));
  NA3        o194(.A(ori_ori_n216_), .B(ori_ori_n205_), .C(ori_ori_n195_), .Y(ori_ori_n217_));
  AOI210     o195(.A0(ori_ori_n132_), .A1(ori_ori_n82_), .B0(i_1_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n142_), .B(i_2_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n219_), .B(ori_ori_n218_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(i_13_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n49_), .B(i_12_), .Y(ori_ori_n222_));
  INV        o200(.A(ori_ori_n222_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(ori_ori_n78_), .Y(ori_ori_n224_));
  INV        o202(.A(ori_ori_n224_), .Y(ori_ori_n225_));
  NA2        o203(.A(ori_ori_n100_), .B(i_13_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(ori_ori_n218_), .Y(ori_ori_n227_));
  INV        o205(.A(ori_ori_n227_), .Y(ori_ori_n228_));
  OR2        o206(.A(i_11_), .B(i_6_), .Y(ori_ori_n229_));
  NA3        o207(.A(ori_ori_n148_), .B(i_10_), .C(ori_ori_n82_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n196_), .B(i_13_), .Y(ori_ori_n231_));
  NA2        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n232_), .B(ori_ori_n53_), .Y(ori_ori_n233_));
  NA3        o211(.A(ori_ori_n233_), .B(ori_ori_n228_), .C(ori_ori_n225_), .Y(ori_ori_n234_));
  OR4        o212(.A(ori_ori_n234_), .B(ori_ori_n221_), .C(ori_ori_n217_), .D(ori_ori_n188_), .Y(ori5));
  NA2        o213(.A(ori_ori_n207_), .B(ori_ori_n134_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n97_), .B(ori_ori_n23_), .Y(ori_ori_n238_));
  INV        o216(.A(ori_ori_n154_), .Y(ori_ori_n239_));
  AOI220     o217(.A0(ori_ori_n139_), .A1(ori_ori_n174_), .B0(i_12_), .B1(ori_ori_n238_), .Y(ori_ori_n240_));
  INV        o218(.A(ori_ori_n240_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n241_), .B(ori_ori_n237_), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n116_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n219_), .B(ori_ori_n89_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(ori_ori_n243_), .Y(ori_ori_n245_));
  INV        o223(.A(ori_ori_n152_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(i_2_), .Y(ori_ori_n247_));
  INV        o225(.A(ori_ori_n247_), .Y(ori_ori_n248_));
  AOI210     o226(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n150_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n249_), .A1(ori_ori_n248_), .B0(ori_ori_n245_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n118_), .B(ori_ori_n98_), .Y(ori_ori_n251_));
  OAI210     o229(.A0(ori_ori_n251_), .A1(ori_ori_n238_), .B0(i_2_), .Y(ori_ori_n252_));
  NO2        o230(.A(ori_ori_n252_), .B(ori_ori_n119_), .Y(ori_ori_n253_));
  OA210      o231(.A0(ori_ori_n191_), .A1(ori_ori_n99_), .B0(i_13_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n122_), .A1(ori_ori_n111_), .B0(ori_ori_n168_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n255_), .B(ori_ori_n152_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n85_), .B(ori_ori_n42_), .Y(ori_ori_n257_));
  INV        o235(.A(ori_ori_n135_), .Y(ori_ori_n258_));
  NA4        o236(.A(ori_ori_n258_), .B(ori_ori_n136_), .C(ori_ori_n97_), .D(ori_ori_n40_), .Y(ori_ori_n259_));
  OAI210     o237(.A0(ori_ori_n259_), .A1(ori_ori_n257_), .B0(ori_ori_n256_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n260_), .B(ori_ori_n254_), .C(ori_ori_n253_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n99_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n263_), .B(ori_ori_n179_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n36_), .Y(ori_ori_n265_));
  NA4        o243(.A(ori_ori_n265_), .B(ori_ori_n261_), .C(ori_ori_n250_), .D(ori_ori_n242_), .Y(ori6));
  INV        o244(.A(ori_ori_n141_), .Y(ori_ori_n267_));
  OR2        o245(.A(ori_ori_n267_), .B(i_12_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n175_), .B(ori_ori_n53_), .Y(ori_ori_n269_));
  INV        o247(.A(ori_ori_n269_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(ori_ori_n63_), .Y(ori_ori_n271_));
  INV        o249(.A(ori_ori_n140_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n65_), .B(ori_ori_n103_), .Y(ori_ori_n273_));
  INV        o251(.A(ori_ori_n97_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n274_), .B(ori_ori_n44_), .Y(ori_ori_n275_));
  AOI210     o253(.A0(ori_ori_n275_), .A1(ori_ori_n273_), .B0(ori_ori_n272_), .Y(ori_ori_n276_));
  NAi32      o254(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n229_), .B(ori_ori_n277_), .Y(ori_ori_n278_));
  OR2        o256(.A(ori_ori_n278_), .B(ori_ori_n276_), .Y(ori_ori_n279_));
  BUFFER     o257(.A(ori_ori_n191_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n110_), .Y(ori_ori_n281_));
  AO210      o259(.A0(ori_ori_n166_), .A1(ori_ori_n239_), .B0(ori_ori_n36_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n281_), .Y(ori_ori_n283_));
  NO2        o261(.A(i_6_), .B(i_11_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n284_), .B(ori_ori_n171_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n146_), .B(ori_ori_n60_), .Y(ori_ori_n286_));
  NA3        o264(.A(ori_ori_n286_), .B(ori_ori_n285_), .C(ori_ori_n181_), .Y(ori_ori_n287_));
  NA2        o265(.A(ori_ori_n90_), .B(ori_ori_n147_), .Y(ori_ori_n288_));
  INV        o266(.A(ori_ori_n288_), .Y(ori_ori_n289_));
  NO4        o267(.A(ori_ori_n289_), .B(ori_ori_n287_), .C(ori_ori_n283_), .D(ori_ori_n279_), .Y(ori_ori_n290_));
  NA3        o268(.A(ori_ori_n290_), .B(ori_ori_n271_), .C(ori_ori_n268_), .Y(ori3));
  NO3        o269(.A(ori_ori_n143_), .B(ori_ori_n38_), .C(i_0_), .Y(ori_ori_n292_));
  NO2        o270(.A(ori_ori_n326_), .B(ori_ori_n53_), .Y(ori_ori_n293_));
  NOi21      o271(.An(i_5_), .B(i_9_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n294_), .B(ori_ori_n153_), .Y(ori_ori_n295_));
  BUFFER     o273(.A(ori_ori_n132_), .Y(ori_ori_n296_));
  NA2        o274(.A(ori_ori_n296_), .B(ori_ori_n163_), .Y(ori_ori_n297_));
  NO2        o275(.A(ori_ori_n297_), .B(ori_ori_n295_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(ori_ori_n293_), .Y(ori_ori_n299_));
  NA2        o277(.A(i_9_), .B(i_0_), .Y(ori_ori_n300_));
  NA2        o278(.A(i_0_), .B(i_10_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n203_), .B(ori_ori_n94_), .Y(ori_ori_n302_));
  NA2        o280(.A(ori_ori_n116_), .B(ori_ori_n86_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n269_), .B(ori_ori_n303_), .Y(ori_ori_n304_));
  INV        o282(.A(ori_ori_n304_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n130_), .B(ori_ori_n126_), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n306_), .A1(ori_ori_n300_), .B0(ori_ori_n113_), .Y(ori_ori_n307_));
  INV        o285(.A(ori_ori_n307_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n308_), .B(ori_ori_n305_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n301_), .B(ori_ori_n294_), .Y(ori_ori_n310_));
  AOI220     o288(.A0(ori_ori_n310_), .A1(i_11_), .B0(ori_ori_n173_), .B1(ori_ori_n65_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n123_), .B(ori_ori_n143_), .C(i_0_), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n66_), .B0(i_13_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n313_), .B(ori_ori_n311_), .Y(ori_ori_n314_));
  NA3        o292(.A(ori_ori_n144_), .B(ori_ori_n116_), .C(ori_ori_n115_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n315_), .B(ori_ori_n165_), .Y(ori_ori_n316_));
  NO3        o294(.A(ori_ori_n316_), .B(ori_ori_n314_), .C(ori_ori_n309_), .Y(ori_ori_n317_));
  INV        o295(.A(ori_ori_n186_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n318_), .B(ori_ori_n121_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n319_), .B(ori_ori_n63_), .Y(ori_ori_n320_));
  INV        o298(.A(ori_ori_n320_), .Y(ori_ori_n321_));
  NA4        o299(.A(ori_ori_n321_), .B(ori_ori_n317_), .C(ori_ori_n302_), .D(ori_ori_n299_), .Y(ori4));
  INV        o300(.A(i_6_), .Y(ori_ori_n325_));
  INV        o301(.A(ori_ori_n292_), .Y(ori_ori_n326_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NOi21      m016(.An(i_12_), .B(i_13_), .Y(mai_mai_n39_));
  INV        m017(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m018(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NO2        m028(.A(mai_mai_n47_), .B(mai_mai_n46_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_0_), .B(i_2_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_7_), .B(i_9_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n51_), .B0(mai_mai_n45_), .Y(mai_mai_n55_));
  NA3        m033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n56_));
  NO2        m034(.A(i_1_), .B(i_6_), .Y(mai_mai_n57_));
  NA2        m035(.A(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  OAI210     m036(.A0(mai_mai_n58_), .A1(mai_mai_n57_), .B0(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n60_));
  NAi21      m038(.An(i_2_), .B(i_7_), .Y(mai_mai_n61_));
  INV        m039(.A(i_1_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n62_), .B(i_6_), .Y(mai_mai_n63_));
  INV        m041(.A(mai_mai_n60_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n65_));
  NA2        m043(.A(i_1_), .B(i_6_), .Y(mai_mai_n66_));
  NO2        m044(.A(mai_mai_n66_), .B(mai_mai_n25_), .Y(mai_mai_n67_));
  INV        m045(.A(i_0_), .Y(mai_mai_n68_));
  NAi21      m046(.An(i_5_), .B(i_10_), .Y(mai_mai_n69_));
  NA2        m047(.A(i_5_), .B(i_9_), .Y(mai_mai_n70_));
  AOI210     m048(.A0(mai_mai_n70_), .A1(mai_mai_n69_), .B0(mai_mai_n68_), .Y(mai_mai_n71_));
  NO2        m049(.A(mai_mai_n71_), .B(mai_mai_n67_), .Y(mai_mai_n72_));
  INV        m050(.A(mai_mai_n72_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(mai_mai_n64_), .B0(i_0_), .Y(mai_mai_n74_));
  NA2        m052(.A(i_12_), .B(i_5_), .Y(mai_mai_n75_));
  NO2        m053(.A(i_3_), .B(i_9_), .Y(mai_mai_n76_));
  NO2        m054(.A(i_3_), .B(i_7_), .Y(mai_mai_n77_));
  INV        m055(.A(i_6_), .Y(mai_mai_n78_));
  OR4        m056(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n79_));
  INV        m057(.A(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m058(.A(i_2_), .B(i_7_), .Y(mai_mai_n81_));
  NAi21      m059(.An(i_6_), .B(i_10_), .Y(mai_mai_n82_));
  NA2        m060(.A(i_6_), .B(i_9_), .Y(mai_mai_n83_));
  AOI210     m061(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n62_), .Y(mai_mai_n84_));
  NA2        m062(.A(i_2_), .B(i_6_), .Y(mai_mai_n85_));
  INV        m063(.A(mai_mai_n84_), .Y(mai_mai_n86_));
  NO2        m064(.A(mai_mai_n86_), .B(mai_mai_n75_), .Y(mai_mai_n87_));
  AN3        m065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n88_));
  NAi21      m066(.An(i_6_), .B(i_11_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_5_), .B(i_8_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  AOI220     m069(.A0(mai_mai_n91_), .A1(mai_mai_n61_), .B0(mai_mai_n88_), .B1(mai_mai_n32_), .Y(mai_mai_n92_));
  INV        m070(.A(i_7_), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n46_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_0_), .B(i_5_), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n95_), .B(mai_mai_n78_), .Y(mai_mai_n96_));
  NA2        m074(.A(i_12_), .B(i_3_), .Y(mai_mai_n97_));
  INV        m075(.A(mai_mai_n97_), .Y(mai_mai_n98_));
  NA3        m076(.A(mai_mai_n98_), .B(mai_mai_n96_), .C(mai_mai_n94_), .Y(mai_mai_n99_));
  NAi21      m077(.An(i_7_), .B(i_11_), .Y(mai_mai_n100_));
  NO3        m078(.A(mai_mai_n100_), .B(mai_mai_n82_), .C(mai_mai_n52_), .Y(mai_mai_n101_));
  AN2        m079(.A(i_2_), .B(i_10_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(i_7_), .Y(mai_mai_n103_));
  OR2        m081(.A(mai_mai_n75_), .B(mai_mai_n57_), .Y(mai_mai_n104_));
  NO2        m082(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n105_));
  NO3        m083(.A(mai_mai_n105_), .B(mai_mai_n104_), .C(mai_mai_n103_), .Y(mai_mai_n106_));
  NA2        m084(.A(i_12_), .B(i_7_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n62_), .B(mai_mai_n26_), .Y(mai_mai_n108_));
  NA2        m086(.A(mai_mai_n108_), .B(i_0_), .Y(mai_mai_n109_));
  NA2        m087(.A(i_11_), .B(i_12_), .Y(mai_mai_n110_));
  OAI210     m088(.A0(mai_mai_n109_), .A1(mai_mai_n107_), .B0(mai_mai_n110_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n111_), .B(mai_mai_n106_), .Y(mai_mai_n112_));
  NAi41      m090(.An(mai_mai_n101_), .B(mai_mai_n112_), .C(mai_mai_n99_), .D(mai_mai_n92_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n93_), .B(mai_mai_n37_), .Y(mai_mai_n114_));
  NA2        m092(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n116_), .B(mai_mai_n46_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n118_));
  NAi21      m096(.An(i_3_), .B(i_8_), .Y(mai_mai_n119_));
  NO2        m097(.A(i_1_), .B(mai_mai_n78_), .Y(mai_mai_n120_));
  NO2        m098(.A(i_6_), .B(i_5_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(i_3_), .Y(mai_mai_n122_));
  AO210      m100(.A0(mai_mai_n122_), .A1(mai_mai_n47_), .B0(mai_mai_n120_), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n123_), .B(mai_mai_n100_), .Y(mai_mai_n124_));
  NO3        m102(.A(mai_mai_n124_), .B(mai_mai_n113_), .C(mai_mai_n87_), .Y(mai_mai_n125_));
  NA3        m103(.A(mai_mai_n125_), .B(mai_mai_n74_), .C(mai_mai_n55_), .Y(mai2));
  NO2        m104(.A(mai_mai_n62_), .B(mai_mai_n37_), .Y(mai_mai_n127_));
  NA2        m105(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n129_));
  NA4        m107(.A(mai_mai_n129_), .B(mai_mai_n72_), .C(mai_mai_n65_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m108(.A(i_8_), .B(i_7_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(i_6_), .Y(mai_mai_n132_));
  NO2        m110(.A(i_12_), .B(i_13_), .Y(mai_mai_n133_));
  NAi21      m111(.An(i_5_), .B(i_11_), .Y(mai_mai_n134_));
  NOi21      m112(.An(mai_mai_n133_), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_0_), .B(i_1_), .Y(mai_mai_n136_));
  NA2        m114(.A(i_2_), .B(i_3_), .Y(mai_mai_n137_));
  NO2        m115(.A(mai_mai_n137_), .B(i_4_), .Y(mai_mai_n138_));
  NA3        m116(.A(mai_mai_n138_), .B(mai_mai_n136_), .C(mai_mai_n135_), .Y(mai_mai_n139_));
  AN2        m117(.A(mai_mai_n133_), .B(mai_mai_n76_), .Y(mai_mai_n140_));
  NA2        m118(.A(i_1_), .B(i_5_), .Y(mai_mai_n141_));
  NO2        m119(.A(mai_mai_n68_), .B(mai_mai_n46_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n142_), .B(mai_mai_n36_), .Y(mai_mai_n143_));
  NO3        m121(.A(mai_mai_n143_), .B(mai_mai_n141_), .C(i_13_), .Y(mai_mai_n144_));
  OR2        m122(.A(i_0_), .B(i_1_), .Y(mai_mai_n145_));
  NO3        m123(.A(mai_mai_n145_), .B(mai_mai_n75_), .C(i_13_), .Y(mai_mai_n146_));
  NAi32      m124(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n147_));
  NAi21      m125(.An(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NOi21      m126(.An(i_4_), .B(i_10_), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n149_), .B(mai_mai_n39_), .Y(mai_mai_n150_));
  NO2        m128(.A(i_3_), .B(i_5_), .Y(mai_mai_n151_));
  NA2        m129(.A(i_0_), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  OAI210     m130(.A0(mai_mai_n152_), .A1(mai_mai_n150_), .B0(mai_mai_n148_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n153_), .B(mai_mai_n144_), .Y(mai_mai_n154_));
  AOI210     m132(.A0(mai_mai_n154_), .A1(mai_mai_n139_), .B0(mai_mai_n132_), .Y(mai_mai_n155_));
  NOi21      m133(.An(i_4_), .B(i_9_), .Y(mai_mai_n156_));
  NOi21      m134(.An(i_11_), .B(i_13_), .Y(mai_mai_n157_));
  NA2        m135(.A(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  BUFFER     m136(.A(mai_mai_n158_), .Y(mai_mai_n159_));
  NO2        m137(.A(i_4_), .B(i_5_), .Y(mai_mai_n160_));
  NAi21      m138(.An(i_12_), .B(i_11_), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n161_), .B(i_13_), .Y(mai_mai_n162_));
  NA3        m140(.A(mai_mai_n162_), .B(mai_mai_n160_), .C(mai_mai_n76_), .Y(mai_mai_n163_));
  AOI210     m141(.A0(mai_mai_n163_), .A1(mai_mai_n159_), .B0(mai_mai_n950_), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n68_), .B(mai_mai_n62_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n166_));
  NAi31      m144(.An(mai_mai_n166_), .B(mai_mai_n140_), .C(i_11_), .Y(mai_mai_n167_));
  NA2        m145(.A(i_3_), .B(i_5_), .Y(mai_mai_n168_));
  AOI210     m146(.A0(mai_mai_n158_), .A1(mai_mai_n167_), .B0(mai_mai_n62_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n68_), .B(i_5_), .Y(mai_mai_n170_));
  NO2        m148(.A(i_13_), .B(i_10_), .Y(mai_mai_n171_));
  NA3        m149(.A(mai_mai_n171_), .B(mai_mai_n170_), .C(mai_mai_n44_), .Y(mai_mai_n172_));
  NO2        m150(.A(i_2_), .B(i_1_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(i_3_), .Y(mai_mai_n174_));
  NAi21      m152(.An(i_4_), .B(i_12_), .Y(mai_mai_n175_));
  NO4        m153(.A(mai_mai_n175_), .B(mai_mai_n174_), .C(mai_mai_n172_), .D(mai_mai_n25_), .Y(mai_mai_n176_));
  NO3        m154(.A(mai_mai_n176_), .B(mai_mai_n169_), .C(mai_mai_n164_), .Y(mai_mai_n177_));
  INV        m155(.A(i_8_), .Y(mai_mai_n178_));
  NA2        m156(.A(i_8_), .B(i_6_), .Y(mai_mai_n179_));
  NO3        m157(.A(i_3_), .B(mai_mai_n78_), .C(mai_mai_n48_), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n180_), .B(mai_mai_n105_), .Y(mai_mai_n181_));
  NO3        m159(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n182_));
  NA3        m160(.A(mai_mai_n182_), .B(mai_mai_n39_), .C(mai_mai_n44_), .Y(mai_mai_n183_));
  NO3        m161(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n184_));
  OAI210     m162(.A0(mai_mai_n88_), .A1(i_12_), .B0(mai_mai_n184_), .Y(mai_mai_n185_));
  AOI210     m163(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(mai_mai_n181_), .Y(mai_mai_n186_));
  NO2        m164(.A(i_3_), .B(i_8_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n188_));
  NA3        m166(.A(mai_mai_n188_), .B(mai_mai_n187_), .C(mai_mai_n39_), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n95_), .B(mai_mai_n57_), .Y(mai_mai_n190_));
  NO2        m168(.A(i_13_), .B(i_9_), .Y(mai_mai_n191_));
  NA3        m169(.A(mai_mai_n191_), .B(i_6_), .C(mai_mai_n178_), .Y(mai_mai_n192_));
  NAi21      m170(.An(i_12_), .B(i_3_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n194_));
  NO3        m172(.A(i_0_), .B(i_2_), .C(mai_mai_n62_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n195_), .B(i_10_), .Y(mai_mai_n196_));
  OAI220     m174(.A0(mai_mai_n196_), .A1(mai_mai_n192_), .B0(mai_mai_n57_), .B1(mai_mai_n189_), .Y(mai_mai_n197_));
  AOI210     m175(.A0(mai_mai_n197_), .A1(i_7_), .B0(mai_mai_n186_), .Y(mai_mai_n198_));
  OAI220     m176(.A0(mai_mai_n198_), .A1(i_4_), .B0(mai_mai_n179_), .B1(mai_mai_n177_), .Y(mai_mai_n199_));
  NA3        m177(.A(i_13_), .B(mai_mai_n178_), .C(i_10_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n200_), .B(i_12_), .Y(mai_mai_n201_));
  NA2        m179(.A(i_0_), .B(i_5_), .Y(mai_mai_n202_));
  OAI220     m180(.A0(mai_mai_n78_), .A1(mai_mai_n174_), .B0(mai_mai_n62_), .B1(mai_mai_n122_), .Y(mai_mai_n203_));
  NAi31      m181(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n46_), .B(mai_mai_n62_), .Y(mai_mai_n206_));
  NA3        m184(.A(mai_mai_n206_), .B(i_0_), .C(mai_mai_n205_), .Y(mai_mai_n207_));
  INV        m185(.A(i_13_), .Y(mai_mai_n208_));
  NO2        m186(.A(i_12_), .B(mai_mai_n208_), .Y(mai_mai_n209_));
  NA3        m187(.A(mai_mai_n209_), .B(mai_mai_n182_), .C(mai_mai_n180_), .Y(mai_mai_n210_));
  OAI210     m188(.A0(mai_mai_n207_), .A1(mai_mai_n204_), .B0(mai_mai_n210_), .Y(mai_mai_n211_));
  AOI220     m189(.A0(mai_mai_n211_), .A1(mai_mai_n131_), .B0(mai_mai_n203_), .B1(mai_mai_n201_), .Y(mai_mai_n212_));
  NO2        m190(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n168_), .B(i_4_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n214_), .B(mai_mai_n213_), .Y(mai_mai_n215_));
  OR2        m193(.A(i_8_), .B(i_7_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n216_), .B(mai_mai_n78_), .Y(mai_mai_n217_));
  INV        m195(.A(i_12_), .Y(mai_mai_n218_));
  NO3        m196(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n219_));
  NA2        m197(.A(i_2_), .B(i_1_), .Y(mai_mai_n220_));
  NO2        m198(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n221_));
  NAi21      m199(.An(i_4_), .B(i_3_), .Y(mai_mai_n222_));
  NO2        m200(.A(i_0_), .B(i_6_), .Y(mai_mai_n223_));
  NOi41      m201(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n225_));
  BUFFER     m203(.A(mai_mai_n225_), .Y(mai_mai_n226_));
  INV        m204(.A(mai_mai_n226_), .Y(mai_mai_n227_));
  AOI220     m205(.A0(mai_mai_n227_), .A1(mai_mai_n39_), .B0(mai_mai_n221_), .B1(mai_mai_n191_), .Y(mai_mai_n228_));
  NO2        m206(.A(i_11_), .B(mai_mai_n208_), .Y(mai_mai_n229_));
  NOi21      m207(.An(i_1_), .B(i_6_), .Y(mai_mai_n230_));
  NAi21      m208(.An(i_3_), .B(i_7_), .Y(mai_mai_n231_));
  NA2        m209(.A(mai_mai_n218_), .B(i_9_), .Y(mai_mai_n232_));
  OR4        m210(.A(mai_mai_n232_), .B(mai_mai_n231_), .C(mai_mai_n230_), .D(mai_mai_n170_), .Y(mai_mai_n233_));
  NO2        m211(.A(i_12_), .B(i_3_), .Y(mai_mai_n234_));
  NA2        m212(.A(i_3_), .B(i_9_), .Y(mai_mai_n235_));
  NAi21      m213(.An(i_7_), .B(i_10_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n237_), .B(mai_mai_n63_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n238_), .B(mai_mai_n233_), .Y(mai_mai_n239_));
  NA3        m217(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n240_));
  INV        m218(.A(mai_mai_n132_), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n218_), .B(i_13_), .Y(mai_mai_n242_));
  NO2        m220(.A(mai_mai_n242_), .B(mai_mai_n70_), .Y(mai_mai_n243_));
  AOI220     m221(.A0(mai_mai_n243_), .A1(mai_mai_n241_), .B0(mai_mai_n239_), .B1(mai_mai_n229_), .Y(mai_mai_n244_));
  NO2        m222(.A(mai_mai_n216_), .B(mai_mai_n37_), .Y(mai_mai_n245_));
  NA2        m223(.A(i_12_), .B(i_6_), .Y(mai_mai_n246_));
  OR2        m224(.A(i_13_), .B(i_9_), .Y(mai_mai_n247_));
  NO3        m225(.A(mai_mai_n247_), .B(mai_mai_n246_), .C(mai_mai_n48_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n222_), .B(i_2_), .Y(mai_mai_n249_));
  NA3        m227(.A(mai_mai_n249_), .B(mai_mai_n248_), .C(mai_mai_n44_), .Y(mai_mai_n250_));
  NA2        m228(.A(mai_mai_n229_), .B(i_9_), .Y(mai_mai_n251_));
  OAI210     m229(.A0(mai_mai_n62_), .A1(mai_mai_n251_), .B0(mai_mai_n250_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n142_), .B(mai_mai_n62_), .Y(mai_mai_n253_));
  NO3        m231(.A(i_11_), .B(mai_mai_n208_), .C(mai_mai_n25_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n231_), .B(i_8_), .Y(mai_mai_n255_));
  NO2        m233(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n255_), .B(mai_mai_n254_), .Y(mai_mai_n257_));
  NA3        m235(.A(i_3_), .B(mai_mai_n245_), .C(mai_mai_n209_), .Y(mai_mai_n258_));
  AOI210     m236(.A0(mai_mai_n258_), .A1(mai_mai_n257_), .B0(mai_mai_n253_), .Y(mai_mai_n259_));
  AOI210     m237(.A0(mai_mai_n252_), .A1(mai_mai_n245_), .B0(mai_mai_n259_), .Y(mai_mai_n260_));
  NA4        m238(.A(mai_mai_n260_), .B(mai_mai_n244_), .C(mai_mai_n228_), .D(mai_mai_n212_), .Y(mai_mai_n261_));
  NO3        m239(.A(i_12_), .B(mai_mai_n208_), .C(mai_mai_n37_), .Y(mai_mai_n262_));
  INV        m240(.A(mai_mai_n262_), .Y(mai_mai_n263_));
  NA2        m241(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n264_));
  NO2        m242(.A(i_3_), .B(mai_mai_n264_), .Y(mai_mai_n265_));
  NO2        m243(.A(mai_mai_n220_), .B(i_0_), .Y(mai_mai_n266_));
  NA2        m244(.A(mai_mai_n256_), .B(mai_mai_n26_), .Y(mai_mai_n267_));
  NO2        m245(.A(mai_mai_n267_), .B(mai_mai_n958_), .Y(mai_mai_n268_));
  NO2        m246(.A(mai_mai_n58_), .B(i_6_), .Y(mai_mai_n269_));
  NA3        m247(.A(mai_mai_n269_), .B(i_1_), .C(mai_mai_n151_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n152_), .A1(mai_mai_n132_), .B0(mai_mai_n270_), .Y(mai_mai_n271_));
  NO3        m249(.A(mai_mai_n271_), .B(mai_mai_n268_), .C(mai_mai_n265_), .Y(mai_mai_n272_));
  NO2        m250(.A(i_3_), .B(i_10_), .Y(mai_mai_n273_));
  NA3        m251(.A(mai_mai_n273_), .B(mai_mai_n39_), .C(mai_mai_n44_), .Y(mai_mai_n274_));
  NA2        m252(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n275_));
  AN2        m253(.A(i_3_), .B(i_10_), .Y(mai_mai_n276_));
  NA4        m254(.A(mai_mai_n276_), .B(mai_mai_n182_), .C(mai_mai_n162_), .D(mai_mai_n160_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n278_));
  OR2        m256(.A(mai_mai_n275_), .B(mai_mai_n274_), .Y(mai_mai_n279_));
  OAI220     m257(.A0(mai_mai_n279_), .A1(i_6_), .B0(mai_mai_n272_), .B1(mai_mai_n263_), .Y(mai_mai_n280_));
  NO4        m258(.A(mai_mai_n280_), .B(mai_mai_n261_), .C(mai_mai_n199_), .D(mai_mai_n155_), .Y(mai_mai_n281_));
  NO3        m259(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n282_));
  NO3        m260(.A(i_6_), .B(mai_mai_n178_), .C(i_7_), .Y(mai_mai_n283_));
  NA2        m261(.A(mai_mai_n283_), .B(mai_mai_n182_), .Y(mai_mai_n284_));
  AOI210     m262(.A0(mai_mai_n284_), .A1(mai_mai_n220_), .B0(i_5_), .Y(mai_mai_n285_));
  NO2        m263(.A(i_2_), .B(i_3_), .Y(mai_mai_n286_));
  OR2        m264(.A(i_0_), .B(i_5_), .Y(mai_mai_n287_));
  NA2        m265(.A(mai_mai_n202_), .B(mai_mai_n287_), .Y(mai_mai_n288_));
  NA4        m266(.A(mai_mai_n288_), .B(mai_mai_n217_), .C(mai_mai_n286_), .D(i_1_), .Y(mai_mai_n289_));
  NA3        m267(.A(mai_mai_n266_), .B(mai_mai_n151_), .C(mai_mai_n105_), .Y(mai_mai_n290_));
  NAi21      m268(.An(i_8_), .B(i_7_), .Y(mai_mai_n291_));
  NA3        m269(.A(i_2_), .B(i_7_), .C(mai_mai_n151_), .Y(mai_mai_n292_));
  NA3        m270(.A(mai_mai_n292_), .B(mai_mai_n290_), .C(mai_mai_n289_), .Y(mai_mai_n293_));
  OAI210     m271(.A0(mai_mai_n293_), .A1(mai_mai_n285_), .B0(i_4_), .Y(mai_mai_n294_));
  NO2        m272(.A(i_12_), .B(i_10_), .Y(mai_mai_n295_));
  NOi21      m273(.An(i_5_), .B(i_0_), .Y(mai_mai_n296_));
  NO3        m274(.A(mai_mai_n275_), .B(mai_mai_n296_), .C(mai_mai_n119_), .Y(mai_mai_n297_));
  NA4        m275(.A(mai_mai_n77_), .B(mai_mai_n36_), .C(mai_mai_n78_), .D(i_8_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n297_), .B(mai_mai_n295_), .Y(mai_mai_n299_));
  NO2        m277(.A(i_6_), .B(i_8_), .Y(mai_mai_n300_));
  AN2        m278(.A(i_0_), .B(mai_mai_n300_), .Y(mai_mai_n301_));
  NO2        m279(.A(i_1_), .B(i_7_), .Y(mai_mai_n302_));
  NA3        m280(.A(mai_mai_n300_), .B(mai_mai_n41_), .C(i_5_), .Y(mai_mai_n303_));
  NA3        m281(.A(mai_mai_n303_), .B(mai_mai_n299_), .C(mai_mai_n294_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n95_), .B(mai_mai_n115_), .Y(mai_mai_n305_));
  NA2        m283(.A(mai_mai_n305_), .B(i_3_), .Y(mai_mai_n306_));
  NO2        m284(.A(mai_mai_n85_), .B(mai_mai_n178_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n178_), .B(i_9_), .Y(mai_mai_n308_));
  AOI210     m286(.A0(mai_mai_n956_), .A1(mai_mai_n306_), .B0(mai_mai_n150_), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n304_), .A1(mai_mai_n282_), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  NOi32      m288(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n311_), .Y(mai_mai_n312_));
  NAi21      m290(.An(i_1_), .B(i_5_), .Y(mai_mai_n313_));
  NA2        m291(.A(mai_mai_n313_), .B(i_0_), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n314_), .B(mai_mai_n25_), .Y(mai_mai_n315_));
  OAI210     m293(.A0(mai_mai_n315_), .A1(mai_mai_n147_), .B0(mai_mai_n225_), .Y(mai_mai_n316_));
  NAi41      m294(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n317_));
  OAI220     m295(.A0(mai_mai_n317_), .A1(mai_mai_n313_), .B0(mai_mai_n204_), .B1(mai_mai_n147_), .Y(mai_mai_n318_));
  AOI210     m296(.A0(mai_mai_n317_), .A1(mai_mai_n147_), .B0(mai_mai_n145_), .Y(mai_mai_n319_));
  NOi32      m297(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n320_));
  NA2        m298(.A(mai_mai_n320_), .B(mai_mai_n46_), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n321_), .B(i_0_), .Y(mai_mai_n322_));
  OR3        m300(.A(mai_mai_n322_), .B(mai_mai_n319_), .C(mai_mai_n318_), .Y(mai_mai_n323_));
  NO2        m301(.A(i_1_), .B(mai_mai_n93_), .Y(mai_mai_n324_));
  NAi21      m302(.An(i_3_), .B(i_4_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n325_), .B(i_9_), .Y(mai_mai_n326_));
  AN2        m304(.A(i_6_), .B(i_7_), .Y(mai_mai_n327_));
  OAI210     m305(.A0(mai_mai_n327_), .A1(mai_mai_n324_), .B0(mai_mai_n326_), .Y(mai_mai_n328_));
  NA2        m306(.A(i_2_), .B(i_7_), .Y(mai_mai_n329_));
  NO2        m307(.A(mai_mai_n325_), .B(i_10_), .Y(mai_mai_n330_));
  NA3        m308(.A(mai_mai_n330_), .B(mai_mai_n329_), .C(mai_mai_n223_), .Y(mai_mai_n331_));
  AOI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n328_), .B0(mai_mai_n170_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n333_));
  OAI210     m311(.A0(mai_mai_n333_), .A1(mai_mai_n173_), .B0(mai_mai_n330_), .Y(mai_mai_n334_));
  AOI220     m312(.A0(mai_mai_n330_), .A1(mai_mai_n302_), .B0(mai_mai_n219_), .B1(mai_mai_n173_), .Y(mai_mai_n335_));
  AOI210     m313(.A0(mai_mai_n335_), .A1(mai_mai_n334_), .B0(i_5_), .Y(mai_mai_n336_));
  NO4        m314(.A(mai_mai_n336_), .B(mai_mai_n332_), .C(mai_mai_n323_), .D(mai_mai_n316_), .Y(mai_mai_n337_));
  NO2        m315(.A(mai_mai_n337_), .B(mai_mai_n312_), .Y(mai_mai_n338_));
  NO2        m316(.A(mai_mai_n58_), .B(mai_mai_n25_), .Y(mai_mai_n339_));
  AN2        m317(.A(i_12_), .B(i_5_), .Y(mai_mai_n340_));
  NO2        m318(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n342_));
  NO2        m320(.A(i_11_), .B(i_6_), .Y(mai_mai_n343_));
  NA3        m321(.A(mai_mai_n343_), .B(i_2_), .C(mai_mai_n208_), .Y(mai_mai_n344_));
  NO2        m322(.A(mai_mai_n344_), .B(mai_mai_n342_), .Y(mai_mai_n345_));
  NO2        m323(.A(mai_mai_n222_), .B(i_5_), .Y(mai_mai_n346_));
  NO2        m324(.A(i_5_), .B(i_10_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n133_), .B(mai_mai_n45_), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(mai_mai_n222_), .Y(mai_mai_n349_));
  OAI210     m327(.A0(mai_mai_n349_), .A1(mai_mai_n345_), .B0(mai_mai_n339_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n139_), .B(mai_mai_n78_), .Y(mai_mai_n352_));
  OAI210     m330(.A0(mai_mai_n352_), .A1(mai_mai_n345_), .B0(mai_mai_n351_), .Y(mai_mai_n353_));
  NO2        m331(.A(i_11_), .B(i_12_), .Y(mai_mai_n354_));
  NA2        m332(.A(mai_mai_n347_), .B(mai_mai_n218_), .Y(mai_mai_n355_));
  OAI220     m333(.A0(mai_mai_n36_), .A1(mai_mai_n204_), .B0(mai_mai_n355_), .B1(mai_mai_n298_), .Y(mai_mai_n356_));
  NAi21      m334(.An(i_13_), .B(i_0_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n357_), .B(mai_mai_n220_), .Y(mai_mai_n358_));
  NA2        m336(.A(mai_mai_n356_), .B(mai_mai_n358_), .Y(mai_mai_n359_));
  NA3        m337(.A(mai_mai_n359_), .B(mai_mai_n353_), .C(mai_mai_n350_), .Y(mai_mai_n360_));
  NO2        m338(.A(i_0_), .B(i_11_), .Y(mai_mai_n361_));
  AN2        m339(.A(i_1_), .B(i_6_), .Y(mai_mai_n362_));
  NOi21      m340(.An(i_2_), .B(i_12_), .Y(mai_mai_n363_));
  NA2        m341(.A(mai_mai_n131_), .B(i_9_), .Y(mai_mai_n364_));
  NO2        m342(.A(mai_mai_n364_), .B(i_4_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n363_), .B(mai_mai_n365_), .Y(mai_mai_n366_));
  NAi21      m344(.An(i_9_), .B(i_4_), .Y(mai_mai_n367_));
  OR2        m345(.A(i_13_), .B(i_10_), .Y(mai_mai_n368_));
  NO2        m346(.A(mai_mai_n158_), .B(mai_mai_n114_), .Y(mai_mai_n369_));
  BUFFER     m347(.A(mai_mai_n200_), .Y(mai_mai_n370_));
  NO2        m348(.A(mai_mai_n93_), .B(mai_mai_n25_), .Y(mai_mai_n371_));
  NA2        m349(.A(mai_mai_n262_), .B(mai_mai_n371_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n256_), .B(mai_mai_n195_), .Y(mai_mai_n373_));
  OAI220     m351(.A0(mai_mai_n373_), .A1(mai_mai_n370_), .B0(mai_mai_n372_), .B1(mai_mai_n95_), .Y(mai_mai_n374_));
  INV        m352(.A(mai_mai_n374_), .Y(mai_mai_n375_));
  AOI210     m353(.A0(mai_mai_n375_), .A1(mai_mai_n366_), .B0(mai_mai_n26_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n290_), .B(mai_mai_n289_), .Y(mai_mai_n377_));
  AOI220     m355(.A0(mai_mai_n269_), .A1(i_2_), .B0(mai_mai_n266_), .B1(i_7_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(i_5_), .Y(mai_mai_n379_));
  AOI220     m357(.A0(i_3_), .A1(i_1_), .B0(i_3_), .B1(mai_mai_n195_), .Y(mai_mai_n380_));
  NO2        m358(.A(mai_mai_n380_), .B(mai_mai_n264_), .Y(mai_mai_n381_));
  NO3        m359(.A(mai_mai_n381_), .B(mai_mai_n379_), .C(mai_mai_n377_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n180_), .B(mai_mai_n88_), .Y(mai_mai_n383_));
  NA3        m361(.A(i_2_), .B(mai_mai_n151_), .C(mai_mai_n78_), .Y(mai_mai_n384_));
  AOI210     m362(.A0(mai_mai_n384_), .A1(mai_mai_n383_), .B0(mai_mai_n291_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n178_), .B(i_10_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n63_), .B(i_2_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n269_), .B(i_2_), .Y(mai_mai_n388_));
  OAI220     m366(.A0(mai_mai_n388_), .A1(mai_mai_n168_), .B0(mai_mai_n387_), .B1(mai_mai_n386_), .Y(mai_mai_n389_));
  NA3        m367(.A(mai_mai_n302_), .B(mai_mai_n301_), .C(i_5_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n283_), .B(mai_mai_n288_), .Y(mai_mai_n391_));
  OAI210     m369(.A0(mai_mai_n391_), .A1(mai_mai_n174_), .B0(mai_mai_n390_), .Y(mai_mai_n392_));
  NO3        m370(.A(mai_mai_n392_), .B(mai_mai_n389_), .C(mai_mai_n385_), .Y(mai_mai_n393_));
  AOI210     m371(.A0(mai_mai_n393_), .A1(mai_mai_n382_), .B0(mai_mai_n251_), .Y(mai_mai_n394_));
  NO4        m372(.A(mai_mai_n394_), .B(mai_mai_n376_), .C(mai_mai_n360_), .D(mai_mai_n338_), .Y(mai_mai_n395_));
  NO2        m373(.A(mai_mai_n68_), .B(i_13_), .Y(mai_mai_n396_));
  NA3        m374(.A(mai_mai_n396_), .B(i_1_), .C(i_2_), .Y(mai_mai_n397_));
  NO2        m375(.A(i_10_), .B(i_9_), .Y(mai_mai_n398_));
  NAi21      m376(.An(i_12_), .B(i_8_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n399_), .B(i_3_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n400_), .B(mai_mai_n398_), .Y(mai_mai_n401_));
  OAI220     m379(.A0(i_4_), .A1(mai_mai_n189_), .B0(mai_mai_n401_), .B1(mai_mai_n397_), .Y(mai_mai_n402_));
  NA2        m380(.A(mai_mai_n278_), .B(i_0_), .Y(mai_mai_n403_));
  NO3        m381(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n404_));
  NA2        m382(.A(mai_mai_n246_), .B(mai_mai_n89_), .Y(mai_mai_n405_));
  NA2        m383(.A(mai_mai_n405_), .B(mai_mai_n404_), .Y(mai_mai_n406_));
  NA2        m384(.A(i_8_), .B(i_9_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n262_), .B(mai_mai_n190_), .Y(mai_mai_n408_));
  OAI220     m386(.A0(mai_mai_n408_), .A1(mai_mai_n407_), .B0(mai_mai_n406_), .B1(mai_mai_n403_), .Y(mai_mai_n409_));
  NO3        m387(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n410_));
  NA3        m388(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n411_));
  NA4        m389(.A(mai_mai_n134_), .B(mai_mai_n108_), .C(mai_mai_n75_), .D(mai_mai_n23_), .Y(mai_mai_n412_));
  NO2        m390(.A(mai_mai_n412_), .B(mai_mai_n411_), .Y(mai_mai_n413_));
  NO3        m391(.A(mai_mai_n413_), .B(mai_mai_n409_), .C(mai_mai_n402_), .Y(mai_mai_n414_));
  OR2        m392(.A(mai_mai_n192_), .B(mai_mai_n215_), .Y(mai_mai_n415_));
  NA2        m393(.A(mai_mai_n88_), .B(i_13_), .Y(mai_mai_n416_));
  NA2        m394(.A(i_3_), .B(mai_mai_n339_), .Y(mai_mai_n417_));
  NO2        m395(.A(i_2_), .B(i_13_), .Y(mai_mai_n418_));
  NA3        m396(.A(mai_mai_n418_), .B(mai_mai_n149_), .C(mai_mai_n91_), .Y(mai_mai_n419_));
  OAI220     m397(.A0(mai_mai_n419_), .A1(mai_mai_n218_), .B0(mai_mai_n417_), .B1(mai_mai_n416_), .Y(mai_mai_n420_));
  NO3        m398(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n421_));
  NO2        m399(.A(i_6_), .B(i_7_), .Y(mai_mai_n422_));
  NA2        m400(.A(mai_mai_n422_), .B(mai_mai_n421_), .Y(mai_mai_n423_));
  OR2        m401(.A(i_11_), .B(i_8_), .Y(mai_mai_n424_));
  NOi21      m402(.An(i_2_), .B(i_7_), .Y(mai_mai_n425_));
  NAi31      m403(.An(mai_mai_n424_), .B(mai_mai_n425_), .C(i_0_), .Y(mai_mai_n426_));
  NO2        m404(.A(mai_mai_n368_), .B(mai_mai_n426_), .Y(mai_mai_n427_));
  NO2        m405(.A(i_6_), .B(i_10_), .Y(mai_mai_n428_));
  NA4        m406(.A(mai_mai_n428_), .B(mai_mai_n282_), .C(i_8_), .D(mai_mai_n218_), .Y(mai_mai_n429_));
  NO2        m407(.A(mai_mai_n429_), .B(mai_mai_n143_), .Y(mai_mai_n430_));
  NA3        m408(.A(mai_mai_n224_), .B(mai_mai_n157_), .C(mai_mai_n121_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n432_));
  NO2        m410(.A(mai_mai_n145_), .B(i_3_), .Y(mai_mai_n433_));
  NAi31      m411(.An(mai_mai_n432_), .B(mai_mai_n433_), .C(mai_mai_n209_), .Y(mai_mai_n434_));
  NA2        m412(.A(mai_mai_n434_), .B(mai_mai_n431_), .Y(mai_mai_n435_));
  NO4        m413(.A(mai_mai_n435_), .B(mai_mai_n430_), .C(mai_mai_n427_), .D(mai_mai_n420_), .Y(mai_mai_n436_));
  NA2        m414(.A(mai_mai_n410_), .B(mai_mai_n347_), .Y(mai_mai_n437_));
  NO2        m415(.A(mai_mai_n437_), .B(mai_mai_n207_), .Y(mai_mai_n438_));
  NAi21      m416(.An(mai_mai_n200_), .B(mai_mai_n354_), .Y(mai_mai_n439_));
  NO2        m417(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n440_));
  NA3        m418(.A(i_6_), .B(mai_mai_n440_), .C(mai_mai_n131_), .Y(mai_mai_n441_));
  OR3        m419(.A(mai_mai_n275_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n442_));
  OAI220     m420(.A0(mai_mai_n442_), .A1(mai_mai_n441_), .B0(i_1_), .B1(mai_mai_n439_), .Y(mai_mai_n443_));
  NA2        m421(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n444_));
  NA2        m422(.A(mai_mai_n282_), .B(mai_mai_n219_), .Y(mai_mai_n445_));
  OAI220     m423(.A0(mai_mai_n445_), .A1(mai_mai_n387_), .B0(mai_mai_n444_), .B1(mai_mai_n416_), .Y(mai_mai_n446_));
  NA4        m424(.A(mai_mai_n276_), .B(mai_mai_n206_), .C(mai_mai_n68_), .D(mai_mai_n218_), .Y(mai_mai_n447_));
  NO2        m425(.A(mai_mai_n447_), .B(mai_mai_n423_), .Y(mai_mai_n448_));
  NO4        m426(.A(mai_mai_n448_), .B(mai_mai_n446_), .C(mai_mai_n443_), .D(mai_mai_n438_), .Y(mai_mai_n449_));
  NA4        m427(.A(mai_mai_n449_), .B(mai_mai_n436_), .C(mai_mai_n415_), .D(mai_mai_n414_), .Y(mai_mai_n450_));
  NA3        m428(.A(mai_mai_n276_), .B(mai_mai_n162_), .C(mai_mai_n160_), .Y(mai_mai_n451_));
  OAI210     m429(.A0(mai_mai_n274_), .A1(mai_mai_n166_), .B0(mai_mai_n451_), .Y(mai_mai_n452_));
  NA2        m430(.A(mai_mai_n217_), .B(mai_mai_n452_), .Y(mai_mai_n453_));
  AN2        m431(.A(mai_mai_n57_), .B(mai_mai_n404_), .Y(mai_mai_n454_));
  NA2        m432(.A(mai_mai_n282_), .B(i_0_), .Y(mai_mai_n455_));
  OAI210     m433(.A0(mai_mai_n455_), .A1(mai_mai_n215_), .B0(mai_mai_n277_), .Y(mai_mai_n456_));
  AOI220     m434(.A0(mai_mai_n456_), .A1(i_7_), .B0(mai_mai_n454_), .B1(mai_mai_n278_), .Y(mai_mai_n457_));
  NA4        m435(.A(mai_mai_n396_), .B(i_1_), .C(mai_mai_n187_), .D(i_2_), .Y(mai_mai_n458_));
  INV        m436(.A(mai_mai_n458_), .Y(mai_mai_n459_));
  NA2        m437(.A(mai_mai_n340_), .B(mai_mai_n208_), .Y(mai_mai_n460_));
  NA2        m438(.A(mai_mai_n311_), .B(mai_mai_n68_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n327_), .B(mai_mai_n320_), .Y(mai_mai_n462_));
  AO210      m440(.A0(mai_mai_n461_), .A1(mai_mai_n460_), .B0(mai_mai_n462_), .Y(mai_mai_n463_));
  INV        m441(.A(mai_mai_n463_), .Y(mai_mai_n464_));
  AOI210     m442(.A0(mai_mai_n459_), .A1(mai_mai_n188_), .B0(mai_mai_n464_), .Y(mai_mai_n465_));
  NO2        m443(.A(i_7_), .B(mai_mai_n183_), .Y(mai_mai_n466_));
  NO2        m444(.A(mai_mai_n168_), .B(mai_mai_n78_), .Y(mai_mai_n467_));
  AOI220     m445(.A0(mai_mai_n467_), .A1(mai_mai_n466_), .B0(mai_mai_n949_), .B1(mai_mai_n369_), .Y(mai_mai_n468_));
  NA4        m446(.A(mai_mai_n468_), .B(mai_mai_n465_), .C(mai_mai_n457_), .D(mai_mai_n453_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n346_), .B(i_1_), .Y(mai_mai_n470_));
  NA2        m448(.A(mai_mai_n342_), .B(mai_mai_n470_), .Y(mai_mai_n471_));
  NO2        m449(.A(i_12_), .B(mai_mai_n178_), .Y(mai_mai_n472_));
  NA2        m450(.A(mai_mai_n472_), .B(mai_mai_n208_), .Y(mai_mai_n473_));
  NO2        m451(.A(i_10_), .B(mai_mai_n473_), .Y(mai_mai_n474_));
  NOi31      m452(.An(mai_mai_n283_), .B(mai_mai_n368_), .C(mai_mai_n38_), .Y(mai_mai_n475_));
  OAI210     m453(.A0(mai_mai_n475_), .A1(mai_mai_n474_), .B0(mai_mai_n471_), .Y(mai_mai_n476_));
  NO2        m454(.A(i_8_), .B(i_7_), .Y(mai_mai_n477_));
  NA2        m455(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n478_));
  NO2        m456(.A(mai_mai_n478_), .B(i_6_), .Y(mai_mai_n479_));
  NA3        m457(.A(mai_mai_n479_), .B(i_2_), .C(mai_mai_n477_), .Y(mai_mai_n480_));
  OAI220     m458(.A0(mai_mai_n168_), .A1(mai_mai_n242_), .B0(mai_mai_n416_), .B1(mai_mai_n122_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n481_), .B(mai_mai_n245_), .Y(mai_mai_n482_));
  NOi31      m460(.An(mai_mai_n266_), .B(mai_mai_n274_), .C(mai_mai_n166_), .Y(mai_mai_n483_));
  NA3        m461(.A(mai_mai_n276_), .B(mai_mai_n160_), .C(mai_mai_n88_), .Y(mai_mai_n484_));
  NO2        m462(.A(mai_mai_n145_), .B(i_5_), .Y(mai_mai_n485_));
  NA2        m463(.A(mai_mai_n485_), .B(mai_mai_n286_), .Y(mai_mai_n486_));
  NA2        m464(.A(mai_mai_n486_), .B(mai_mai_n484_), .Y(mai_mai_n487_));
  OAI210     m465(.A0(mai_mai_n487_), .A1(mai_mai_n483_), .B0(mai_mai_n410_), .Y(mai_mai_n488_));
  NA4        m466(.A(mai_mai_n488_), .B(mai_mai_n482_), .C(mai_mai_n480_), .D(mai_mai_n476_), .Y(mai_mai_n489_));
  NA2        m467(.A(mai_mai_n262_), .B(mai_mai_n77_), .Y(mai_mai_n490_));
  NO2        m468(.A(i_11_), .B(mai_mai_n490_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n269_), .B(i_2_), .Y(mai_mai_n492_));
  NO2        m470(.A(mai_mai_n492_), .B(mai_mai_n159_), .Y(mai_mai_n493_));
  NA2        m471(.A(mai_mai_n206_), .B(i_0_), .Y(mai_mai_n494_));
  NA2        m472(.A(mai_mai_n398_), .B(mai_mai_n205_), .Y(mai_mai_n495_));
  NO2        m473(.A(mai_mai_n494_), .B(mai_mai_n495_), .Y(mai_mai_n496_));
  NA2        m474(.A(i_0_), .B(mai_mai_n48_), .Y(mai_mai_n497_));
  NA3        m475(.A(mai_mai_n472_), .B(mai_mai_n254_), .C(mai_mai_n497_), .Y(mai_mai_n498_));
  INV        m476(.A(mai_mai_n498_), .Y(mai_mai_n499_));
  NO4        m477(.A(mai_mai_n499_), .B(mai_mai_n496_), .C(mai_mai_n493_), .D(mai_mai_n491_), .Y(mai_mai_n500_));
  NO4        m478(.A(mai_mai_n230_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n501_));
  NO3        m479(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n502_));
  NO2        m480(.A(mai_mai_n216_), .B(mai_mai_n36_), .Y(mai_mai_n503_));
  AN2        m481(.A(mai_mai_n503_), .B(mai_mai_n502_), .Y(mai_mai_n504_));
  OA210      m482(.A0(mai_mai_n504_), .A1(mai_mai_n501_), .B0(mai_mai_n311_), .Y(mai_mai_n505_));
  NO2        m483(.A(mai_mai_n368_), .B(i_1_), .Y(mai_mai_n506_));
  AN3        m484(.A(mai_mai_n506_), .B(mai_mai_n365_), .C(i_2_), .Y(mai_mai_n507_));
  NO2        m485(.A(mai_mai_n378_), .B(mai_mai_n163_), .Y(mai_mai_n508_));
  NO3        m486(.A(mai_mai_n508_), .B(mai_mai_n507_), .C(mai_mai_n505_), .Y(mai_mai_n509_));
  NOi21      m487(.An(i_10_), .B(i_6_), .Y(mai_mai_n510_));
  NO2        m488(.A(mai_mai_n78_), .B(mai_mai_n25_), .Y(mai_mai_n511_));
  AOI220     m489(.A0(mai_mai_n262_), .A1(mai_mai_n511_), .B0(mai_mai_n254_), .B1(mai_mai_n510_), .Y(mai_mai_n512_));
  NO2        m490(.A(mai_mai_n512_), .B(mai_mai_n403_), .Y(mai_mai_n513_));
  NO2        m491(.A(mai_mai_n107_), .B(mai_mai_n23_), .Y(mai_mai_n514_));
  NA2        m492(.A(mai_mai_n283_), .B(i_0_), .Y(mai_mai_n515_));
  AOI220     m493(.A0(mai_mai_n515_), .A1(mai_mai_n388_), .B0(mai_mai_n158_), .B1(mai_mai_n167_), .Y(mai_mai_n516_));
  NOi21      m494(.An(mai_mai_n135_), .B(mai_mai_n298_), .Y(mai_mai_n517_));
  NO3        m495(.A(mai_mai_n517_), .B(mai_mai_n516_), .C(mai_mai_n513_), .Y(mai_mai_n518_));
  NO2        m496(.A(mai_mai_n461_), .B(mai_mai_n335_), .Y(mai_mai_n519_));
  INV        m497(.A(mai_mai_n286_), .Y(mai_mai_n520_));
  NO2        m498(.A(i_12_), .B(mai_mai_n78_), .Y(mai_mai_n521_));
  NA3        m499(.A(mai_mai_n521_), .B(mai_mai_n254_), .C(mai_mai_n497_), .Y(mai_mai_n522_));
  NA3        m500(.A(mai_mai_n343_), .B(mai_mai_n262_), .C(mai_mai_n202_), .Y(mai_mai_n523_));
  AOI210     m501(.A0(mai_mai_n523_), .A1(mai_mai_n522_), .B0(mai_mai_n520_), .Y(mai_mai_n524_));
  NO3        m502(.A(i_4_), .B(i_8_), .C(mai_mai_n274_), .Y(mai_mai_n525_));
  OR2        m503(.A(i_5_), .B(mai_mai_n362_), .Y(mai_mai_n526_));
  AOI210     m504(.A0(i_6_), .A1(mai_mai_n526_), .B0(mai_mai_n439_), .Y(mai_mai_n527_));
  NO4        m505(.A(mai_mai_n527_), .B(mai_mai_n525_), .C(mai_mai_n524_), .D(mai_mai_n519_), .Y(mai_mai_n528_));
  NA4        m506(.A(mai_mai_n528_), .B(mai_mai_n518_), .C(mai_mai_n509_), .D(mai_mai_n500_), .Y(mai_mai_n529_));
  NO4        m507(.A(mai_mai_n529_), .B(mai_mai_n489_), .C(mai_mai_n469_), .D(mai_mai_n450_), .Y(mai_mai_n530_));
  NA4        m508(.A(mai_mai_n530_), .B(mai_mai_n395_), .C(mai_mai_n310_), .D(mai_mai_n281_), .Y(mai7));
  NO2        m509(.A(mai_mai_n100_), .B(mai_mai_n82_), .Y(mai_mai_n532_));
  NA2        m510(.A(mai_mai_n341_), .B(mai_mai_n532_), .Y(mai_mai_n533_));
  NA2        m511(.A(mai_mai_n428_), .B(mai_mai_n77_), .Y(mai_mai_n534_));
  NA2        m512(.A(i_11_), .B(mai_mai_n178_), .Y(mai_mai_n535_));
  OAI210     m513(.A0(mai_mai_n951_), .A1(mai_mai_n534_), .B0(mai_mai_n533_), .Y(mai_mai_n536_));
  NA3        m514(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n537_));
  NO2        m515(.A(mai_mai_n218_), .B(i_4_), .Y(mai_mai_n538_));
  NA2        m516(.A(mai_mai_n538_), .B(i_8_), .Y(mai_mai_n539_));
  AOI210     m517(.A0(mai_mai_n539_), .A1(mai_mai_n97_), .B0(mai_mai_n537_), .Y(mai_mai_n540_));
  OAI210     m518(.A0(mai_mai_n81_), .A1(mai_mai_n187_), .B0(mai_mai_n188_), .Y(mai_mai_n541_));
  NO2        m519(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n542_));
  NA2        m520(.A(i_4_), .B(i_8_), .Y(mai_mai_n543_));
  NO2        m521(.A(mai_mai_n541_), .B(i_13_), .Y(mai_mai_n544_));
  NO3        m522(.A(mai_mai_n544_), .B(mai_mai_n540_), .C(mai_mai_n536_), .Y(mai_mai_n545_));
  AOI210     m523(.A0(mai_mai_n119_), .A1(mai_mai_n61_), .B0(i_10_), .Y(mai_mai_n546_));
  AOI210     m524(.A0(mai_mai_n546_), .A1(mai_mai_n218_), .B0(mai_mai_n149_), .Y(mai_mai_n547_));
  OR2        m525(.A(i_6_), .B(i_10_), .Y(mai_mai_n548_));
  NO2        m526(.A(mai_mai_n548_), .B(mai_mai_n23_), .Y(mai_mai_n549_));
  OR3        m527(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n550_));
  NO3        m528(.A(mai_mai_n550_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n551_));
  INV        m529(.A(mai_mai_n184_), .Y(mai_mai_n552_));
  NO2        m530(.A(mai_mai_n551_), .B(mai_mai_n549_), .Y(mai_mai_n553_));
  OA220      m531(.A0(mai_mai_n553_), .A1(mai_mai_n520_), .B0(mai_mai_n547_), .B1(mai_mai_n247_), .Y(mai_mai_n554_));
  AOI210     m532(.A0(mai_mai_n554_), .A1(mai_mai_n545_), .B0(mai_mai_n62_), .Y(mai_mai_n555_));
  NOi21      m533(.An(i_11_), .B(i_7_), .Y(mai_mai_n556_));
  AO210      m534(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n557_));
  NO2        m535(.A(mai_mai_n557_), .B(mai_mai_n556_), .Y(mai_mai_n558_));
  NA2        m536(.A(mai_mai_n558_), .B(mai_mai_n191_), .Y(mai_mai_n559_));
  NA3        m537(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n560_));
  NAi31      m538(.An(mai_mai_n560_), .B(i_12_), .C(i_11_), .Y(mai_mai_n561_));
  AOI210     m539(.A0(mai_mai_n561_), .A1(mai_mai_n559_), .B0(mai_mai_n62_), .Y(mai_mai_n562_));
  NA2        m540(.A(mai_mai_n80_), .B(mai_mai_n62_), .Y(mai_mai_n563_));
  AO210      m541(.A0(mai_mai_n563_), .A1(mai_mai_n335_), .B0(mai_mai_n40_), .Y(mai_mai_n564_));
  NO3        m542(.A(mai_mai_n236_), .B(mai_mai_n193_), .C(mai_mai_n535_), .Y(mai_mai_n565_));
  OAI210     m543(.A0(mai_mai_n565_), .A1(mai_mai_n209_), .B0(mai_mai_n62_), .Y(mai_mai_n566_));
  NA2        m544(.A(mai_mai_n363_), .B(mai_mai_n31_), .Y(mai_mai_n567_));
  OR2        m545(.A(mai_mai_n193_), .B(mai_mai_n100_), .Y(mai_mai_n568_));
  NA2        m546(.A(mai_mai_n568_), .B(mai_mai_n567_), .Y(mai_mai_n569_));
  NO2        m547(.A(mai_mai_n62_), .B(i_9_), .Y(mai_mai_n570_));
  NO2        m548(.A(mai_mai_n570_), .B(i_4_), .Y(mai_mai_n571_));
  NA2        m549(.A(mai_mai_n571_), .B(mai_mai_n569_), .Y(mai_mai_n572_));
  NO2        m550(.A(i_1_), .B(i_12_), .Y(mai_mai_n573_));
  NA3        m551(.A(mai_mai_n572_), .B(mai_mai_n566_), .C(mai_mai_n564_), .Y(mai_mai_n574_));
  OAI210     m552(.A0(mai_mai_n574_), .A1(mai_mai_n562_), .B0(i_6_), .Y(mai_mai_n575_));
  OAI210     m553(.A0(mai_mai_n560_), .A1(mai_mai_n100_), .B0(mai_mai_n411_), .Y(mai_mai_n576_));
  NA2        m554(.A(mai_mai_n576_), .B(mai_mai_n521_), .Y(mai_mai_n577_));
  NO2        m555(.A(mai_mai_n218_), .B(mai_mai_n78_), .Y(mai_mai_n578_));
  NO2        m556(.A(mai_mai_n578_), .B(i_11_), .Y(mai_mai_n579_));
  NA2        m557(.A(mai_mai_n577_), .B(mai_mai_n406_), .Y(mai_mai_n580_));
  NO4        m558(.A(i_12_), .B(mai_mai_n119_), .C(i_13_), .D(mai_mai_n78_), .Y(mai_mai_n581_));
  NA2        m559(.A(mai_mai_n581_), .B(mai_mai_n570_), .Y(mai_mai_n582_));
  NO3        m560(.A(mai_mai_n548_), .B(mai_mai_n216_), .C(mai_mai_n23_), .Y(mai_mai_n583_));
  AOI210     m561(.A0(i_1_), .A1(mai_mai_n237_), .B0(mai_mai_n583_), .Y(mai_mai_n584_));
  OAI210     m562(.A0(mai_mai_n584_), .A1(mai_mai_n44_), .B0(mai_mai_n582_), .Y(mai_mai_n585_));
  NA3        m563(.A(mai_mai_n477_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n586_));
  INV        m564(.A(i_2_), .Y(mai_mai_n587_));
  NA2        m565(.A(mai_mai_n127_), .B(i_9_), .Y(mai_mai_n588_));
  NA3        m566(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n589_));
  NO2        m567(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n590_));
  NA3        m568(.A(mai_mai_n590_), .B(mai_mai_n246_), .C(mai_mai_n44_), .Y(mai_mai_n591_));
  OAI220     m569(.A0(mai_mai_n591_), .A1(mai_mai_n589_), .B0(mai_mai_n588_), .B1(mai_mai_n587_), .Y(mai_mai_n592_));
  NA3        m570(.A(mai_mai_n570_), .B(mai_mai_n286_), .C(i_6_), .Y(mai_mai_n593_));
  NO2        m571(.A(mai_mai_n593_), .B(mai_mai_n23_), .Y(mai_mai_n594_));
  NAi21      m572(.An(mai_mai_n586_), .B(mai_mai_n84_), .Y(mai_mai_n595_));
  INV        m573(.A(mai_mai_n595_), .Y(mai_mai_n596_));
  OR3        m574(.A(mai_mai_n596_), .B(mai_mai_n594_), .C(mai_mai_n592_), .Y(mai_mai_n597_));
  NO3        m575(.A(mai_mai_n597_), .B(mai_mai_n585_), .C(mai_mai_n580_), .Y(mai_mai_n598_));
  NO2        m576(.A(mai_mai_n218_), .B(mai_mai_n93_), .Y(mai_mai_n599_));
  NO2        m577(.A(mai_mai_n599_), .B(mai_mai_n556_), .Y(mai_mai_n600_));
  NA2        m578(.A(mai_mai_n600_), .B(i_1_), .Y(mai_mai_n601_));
  NO2        m579(.A(mai_mai_n601_), .B(mai_mai_n550_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n367_), .B(mai_mai_n78_), .Y(mai_mai_n603_));
  NA2        m581(.A(mai_mai_n602_), .B(mai_mai_n46_), .Y(mai_mai_n604_));
  NA2        m582(.A(i_3_), .B(mai_mai_n178_), .Y(mai_mai_n605_));
  NO2        m583(.A(mai_mai_n605_), .B(mai_mai_n107_), .Y(mai_mai_n606_));
  AN2        m584(.A(mai_mai_n606_), .B(mai_mai_n479_), .Y(mai_mai_n607_));
  NO2        m585(.A(mai_mai_n216_), .B(mai_mai_n44_), .Y(mai_mai_n608_));
  NO2        m586(.A(mai_mai_n78_), .B(i_9_), .Y(mai_mai_n609_));
  NA2        m587(.A(i_1_), .B(i_3_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n407_), .B(mai_mai_n85_), .Y(mai_mai_n611_));
  AOI210     m589(.A0(mai_mai_n608_), .A1(mai_mai_n510_), .B0(mai_mai_n611_), .Y(mai_mai_n612_));
  NO2        m590(.A(mai_mai_n612_), .B(mai_mai_n610_), .Y(mai_mai_n613_));
  NO2        m591(.A(mai_mai_n613_), .B(mai_mai_n607_), .Y(mai_mai_n614_));
  NA4        m592(.A(mai_mai_n614_), .B(mai_mai_n604_), .C(mai_mai_n598_), .D(mai_mai_n575_), .Y(mai_mai_n615_));
  NO3        m593(.A(mai_mai_n424_), .B(i_3_), .C(i_7_), .Y(mai_mai_n616_));
  OA210      m594(.A0(mai_mai_n616_), .A1(mai_mai_n224_), .B0(mai_mai_n78_), .Y(mai_mai_n617_));
  NA2        m595(.A(mai_mai_n327_), .B(mai_mai_n326_), .Y(mai_mai_n618_));
  NA3        m596(.A(mai_mai_n428_), .B(i_4_), .C(mai_mai_n46_), .Y(mai_mai_n619_));
  NO3        m597(.A(mai_mai_n425_), .B(mai_mai_n543_), .C(mai_mai_n78_), .Y(mai_mai_n620_));
  NA2        m598(.A(mai_mai_n620_), .B(mai_mai_n25_), .Y(mai_mai_n621_));
  NA3        m599(.A(mai_mai_n149_), .B(mai_mai_n77_), .C(mai_mai_n78_), .Y(mai_mai_n622_));
  NA4        m600(.A(mai_mai_n622_), .B(mai_mai_n621_), .C(mai_mai_n619_), .D(mai_mai_n618_), .Y(mai_mai_n623_));
  OAI210     m601(.A0(mai_mai_n623_), .A1(mai_mai_n617_), .B0(i_1_), .Y(mai_mai_n624_));
  AOI210     m602(.A0(mai_mai_n246_), .A1(mai_mai_n89_), .B0(i_1_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n325_), .B(i_2_), .Y(mai_mai_n626_));
  NA2        m604(.A(mai_mai_n626_), .B(mai_mai_n625_), .Y(mai_mai_n627_));
  OAI210     m605(.A0(mai_mai_n593_), .A1(mai_mai_n399_), .B0(mai_mai_n627_), .Y(mai_mai_n628_));
  INV        m606(.A(mai_mai_n628_), .Y(mai_mai_n629_));
  AOI210     m607(.A0(mai_mai_n629_), .A1(mai_mai_n624_), .B0(i_13_), .Y(mai_mai_n630_));
  NA3        m608(.A(i_11_), .B(mai_mai_n98_), .C(mai_mai_n127_), .Y(mai_mai_n631_));
  NA2        m609(.A(mai_mai_n418_), .B(mai_mai_n149_), .Y(mai_mai_n632_));
  OAI210     m610(.A0(mai_mai_n632_), .A1(mai_mai_n44_), .B0(mai_mai_n631_), .Y(mai_mai_n633_));
  NO2        m611(.A(mai_mai_n425_), .B(mai_mai_n24_), .Y(mai_mai_n634_));
  AOI220     m612(.A0(mai_mai_n634_), .A1(mai_mai_n603_), .B0(mai_mai_n224_), .B1(mai_mai_n120_), .Y(mai_mai_n635_));
  NO2        m613(.A(mai_mai_n635_), .B(mai_mai_n40_), .Y(mai_mai_n636_));
  AOI210     m614(.A0(mai_mai_n633_), .A1(mai_mai_n300_), .B0(mai_mai_n636_), .Y(mai_mai_n637_));
  NA2        m615(.A(mai_mai_n343_), .B(mai_mai_n590_), .Y(mai_mai_n638_));
  NO2        m616(.A(mai_mai_n638_), .B(mai_mai_n222_), .Y(mai_mai_n639_));
  AOI210     m617(.A0(mai_mai_n399_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n640_));
  NOi31      m618(.An(mai_mai_n640_), .B(mai_mai_n534_), .C(mai_mai_n44_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n118_), .B(i_13_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n589_), .B(mai_mai_n107_), .Y(mai_mai_n643_));
  INV        m621(.A(mai_mai_n643_), .Y(mai_mai_n644_));
  OAI220     m622(.A0(mai_mai_n644_), .A1(mai_mai_n66_), .B0(mai_mai_n642_), .B1(mai_mai_n625_), .Y(mai_mai_n645_));
  NO3        m623(.A(mai_mai_n66_), .B(mai_mai_n32_), .C(mai_mai_n93_), .Y(mai_mai_n646_));
  NA2        m624(.A(mai_mai_n26_), .B(mai_mai_n178_), .Y(mai_mai_n647_));
  NA2        m625(.A(mai_mai_n647_), .B(i_7_), .Y(mai_mai_n648_));
  NO3        m626(.A(mai_mai_n425_), .B(mai_mai_n218_), .C(mai_mai_n78_), .Y(mai_mai_n649_));
  AOI210     m627(.A0(mai_mai_n649_), .A1(mai_mai_n648_), .B0(mai_mai_n646_), .Y(mai_mai_n650_));
  AOI220     m628(.A0(mai_mai_n343_), .A1(mai_mai_n590_), .B0(mai_mai_n84_), .B1(mai_mai_n94_), .Y(mai_mai_n651_));
  OAI220     m629(.A0(mai_mai_n651_), .A1(mai_mai_n539_), .B0(mai_mai_n650_), .B1(mai_mai_n552_), .Y(mai_mai_n652_));
  NO4        m630(.A(mai_mai_n652_), .B(mai_mai_n645_), .C(mai_mai_n641_), .D(mai_mai_n639_), .Y(mai_mai_n653_));
  OR2        m631(.A(i_11_), .B(i_6_), .Y(mai_mai_n654_));
  NA3        m632(.A(mai_mai_n538_), .B(mai_mai_n647_), .C(i_7_), .Y(mai_mai_n655_));
  AOI210     m633(.A0(mai_mai_n655_), .A1(mai_mai_n644_), .B0(mai_mai_n654_), .Y(mai_mai_n656_));
  NA3        m634(.A(mai_mai_n363_), .B(mai_mai_n542_), .C(mai_mai_n89_), .Y(mai_mai_n657_));
  NA2        m635(.A(mai_mai_n579_), .B(i_13_), .Y(mai_mai_n658_));
  NAi21      m636(.An(i_11_), .B(i_12_), .Y(mai_mai_n659_));
  NOi41      m637(.An(mai_mai_n103_), .B(mai_mai_n659_), .C(i_13_), .D(mai_mai_n78_), .Y(mai_mai_n660_));
  NO3        m638(.A(mai_mai_n425_), .B(mai_mai_n521_), .C(mai_mai_n543_), .Y(mai_mai_n661_));
  AOI210     m639(.A0(mai_mai_n661_), .A1(mai_mai_n282_), .B0(mai_mai_n660_), .Y(mai_mai_n662_));
  NA3        m640(.A(mai_mai_n662_), .B(mai_mai_n658_), .C(mai_mai_n657_), .Y(mai_mai_n663_));
  OAI210     m641(.A0(mai_mai_n663_), .A1(mai_mai_n656_), .B0(mai_mai_n62_), .Y(mai_mai_n664_));
  NO2        m642(.A(i_2_), .B(i_12_), .Y(mai_mai_n665_));
  OAI210     m643(.A0(mai_mai_n546_), .A1(mai_mai_n324_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  OAI210     m644(.A0(mai_mai_n218_), .A1(mai_mai_n326_), .B0(mai_mai_n324_), .Y(mai_mai_n667_));
  NO2        m645(.A(mai_mai_n119_), .B(i_2_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n668_), .B(mai_mai_n573_), .Y(mai_mai_n669_));
  NA3        m647(.A(mai_mai_n669_), .B(mai_mai_n667_), .C(mai_mai_n666_), .Y(mai_mai_n670_));
  NA3        m648(.A(mai_mai_n670_), .B(mai_mai_n45_), .C(mai_mai_n208_), .Y(mai_mai_n671_));
  NA4        m649(.A(mai_mai_n671_), .B(mai_mai_n664_), .C(mai_mai_n653_), .D(mai_mai_n637_), .Y(mai_mai_n672_));
  OR4        m650(.A(mai_mai_n672_), .B(mai_mai_n630_), .C(mai_mai_n615_), .D(mai_mai_n555_), .Y(mai5));
  AOI210     m651(.A0(mai_mai_n600_), .A1(mai_mai_n249_), .B0(mai_mai_n369_), .Y(mai_mai_n674_));
  AO210      m652(.A0(mai_mai_n24_), .A1(i_10_), .B0(mai_mai_n229_), .Y(mai_mai_n675_));
  NA3        m653(.A(mai_mai_n675_), .B(mai_mai_n665_), .C(mai_mai_n100_), .Y(mai_mai_n676_));
  NO2        m654(.A(mai_mai_n539_), .B(i_11_), .Y(mai_mai_n677_));
  OAI210     m655(.A0(mai_mai_n542_), .A1(mai_mai_n81_), .B0(mai_mai_n677_), .Y(mai_mai_n678_));
  NA3        m656(.A(mai_mai_n678_), .B(mai_mai_n676_), .C(mai_mai_n674_), .Y(mai_mai_n679_));
  NO3        m657(.A(i_11_), .B(mai_mai_n218_), .C(i_13_), .Y(mai_mai_n680_));
  NO2        m658(.A(mai_mai_n115_), .B(mai_mai_n23_), .Y(mai_mai_n681_));
  NA2        m659(.A(i_12_), .B(i_8_), .Y(mai_mai_n682_));
  OAI210     m660(.A0(mai_mai_n46_), .A1(i_3_), .B0(mai_mai_n682_), .Y(mai_mai_n683_));
  INV        m661(.A(mai_mai_n398_), .Y(mai_mai_n684_));
  AOI220     m662(.A0(mai_mai_n286_), .A1(mai_mai_n514_), .B0(mai_mai_n683_), .B1(mai_mai_n681_), .Y(mai_mai_n685_));
  INV        m663(.A(mai_mai_n685_), .Y(mai_mai_n686_));
  NO2        m664(.A(mai_mai_n686_), .B(mai_mai_n679_), .Y(mai_mai_n687_));
  INV        m665(.A(mai_mai_n157_), .Y(mai_mai_n688_));
  INV        m666(.A(mai_mai_n224_), .Y(mai_mai_n689_));
  OAI210     m667(.A0(mai_mai_n626_), .A1(mai_mai_n400_), .B0(mai_mai_n103_), .Y(mai_mai_n690_));
  AOI210     m668(.A0(mai_mai_n690_), .A1(mai_mai_n689_), .B0(mai_mai_n688_), .Y(mai_mai_n691_));
  NO2        m669(.A(mai_mai_n407_), .B(mai_mai_n26_), .Y(mai_mai_n692_));
  NO2        m670(.A(mai_mai_n692_), .B(mai_mai_n371_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n693_), .B(i_2_), .Y(mai_mai_n694_));
  INV        m672(.A(mai_mai_n694_), .Y(mai_mai_n695_));
  AOI210     m673(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n368_), .Y(mai_mai_n696_));
  AOI210     m674(.A0(mai_mai_n696_), .A1(mai_mai_n695_), .B0(mai_mai_n691_), .Y(mai_mai_n697_));
  NO2        m675(.A(mai_mai_n175_), .B(mai_mai_n116_), .Y(mai_mai_n698_));
  OAI210     m676(.A0(mai_mai_n698_), .A1(mai_mai_n681_), .B0(i_2_), .Y(mai_mai_n699_));
  INV        m677(.A(mai_mai_n158_), .Y(mai_mai_n700_));
  NO3        m678(.A(mai_mai_n557_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n701_));
  AOI210     m679(.A0(mai_mai_n700_), .A1(mai_mai_n81_), .B0(mai_mai_n701_), .Y(mai_mai_n702_));
  AOI210     m680(.A0(mai_mai_n702_), .A1(mai_mai_n699_), .B0(mai_mai_n178_), .Y(mai_mai_n703_));
  OA210      m681(.A0(mai_mai_n558_), .A1(mai_mai_n117_), .B0(i_13_), .Y(mai_mai_n704_));
  NA2        m682(.A(mai_mai_n184_), .B(mai_mai_n187_), .Y(mai_mai_n705_));
  NA2        m683(.A(mai_mai_n140_), .B(mai_mai_n535_), .Y(mai_mai_n706_));
  AOI210     m684(.A0(mai_mai_n706_), .A1(mai_mai_n705_), .B0(mai_mai_n329_), .Y(mai_mai_n707_));
  NA4        m685(.A(i_2_), .B(mai_mai_n276_), .C(mai_mai_n115_), .D(mai_mai_n42_), .Y(mai_mai_n708_));
  INV        m686(.A(mai_mai_n708_), .Y(mai_mai_n709_));
  NO4        m687(.A(mai_mai_n709_), .B(mai_mai_n707_), .C(mai_mai_n704_), .D(mai_mai_n703_), .Y(mai_mai_n710_));
  NA2        m688(.A(mai_mai_n514_), .B(mai_mai_n28_), .Y(mai_mai_n711_));
  NA2        m689(.A(mai_mai_n680_), .B(mai_mai_n255_), .Y(mai_mai_n712_));
  NA2        m690(.A(mai_mai_n712_), .B(mai_mai_n711_), .Y(mai_mai_n713_));
  NO2        m691(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n714_));
  NO2        m692(.A(mai_mai_n714_), .B(mai_mai_n117_), .Y(mai_mai_n715_));
  NO2        m693(.A(mai_mai_n715_), .B(mai_mai_n535_), .Y(mai_mai_n716_));
  AOI220     m694(.A0(mai_mai_n716_), .A1(mai_mai_n36_), .B0(mai_mai_n713_), .B1(mai_mai_n46_), .Y(mai_mai_n717_));
  NA4        m695(.A(mai_mai_n717_), .B(mai_mai_n710_), .C(mai_mai_n697_), .D(mai_mai_n687_), .Y(mai6));
  OAI210     m696(.A0(mai_mai_n25_), .A1(mai_mai_n959_), .B0(mai_mai_n668_), .Y(mai_mai_n719_));
  NA4        m697(.A(mai_mai_n347_), .B(i_8_), .C(mai_mai_n66_), .D(mai_mai_n93_), .Y(mai_mai_n720_));
  INV        m698(.A(mai_mai_n720_), .Y(mai_mai_n721_));
  NO2        m699(.A(mai_mai_n204_), .B(mai_mai_n432_), .Y(mai_mai_n722_));
  NO2        m700(.A(i_11_), .B(i_9_), .Y(mai_mai_n723_));
  NO3        m701(.A(mai_mai_n722_), .B(mai_mai_n721_), .C(mai_mai_n296_), .Y(mai_mai_n724_));
  AO210      m702(.A0(mai_mai_n724_), .A1(mai_mai_n719_), .B0(i_12_), .Y(mai_mai_n725_));
  NA2        m703(.A(mai_mai_n330_), .B(mai_mai_n302_), .Y(mai_mai_n726_));
  NA2        m704(.A(mai_mai_n521_), .B(mai_mai_n62_), .Y(mai_mai_n727_));
  NA2        m705(.A(mai_mai_n616_), .B(mai_mai_n66_), .Y(mai_mai_n728_));
  NA4        m706(.A(mai_mai_n563_), .B(mai_mai_n728_), .C(mai_mai_n727_), .D(mai_mai_n726_), .Y(mai_mai_n729_));
  INV        m707(.A(mai_mai_n181_), .Y(mai_mai_n730_));
  AOI220     m708(.A0(mai_mai_n730_), .A1(mai_mai_n723_), .B0(mai_mai_n729_), .B1(mai_mai_n68_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n947_), .B(mai_mai_n714_), .Y(mai_mai_n732_));
  AOI210     m710(.A0(mai_mai_n732_), .A1(mai_mai_n462_), .B0(mai_mai_n170_), .Y(mai_mai_n733_));
  NO2        m711(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n734_));
  NA3        m712(.A(mai_mai_n734_), .B(mai_mai_n422_), .C(mai_mai_n347_), .Y(mai_mai_n735_));
  OAI210     m713(.A0(mai_mai_n616_), .A1(mai_mai_n503_), .B0(mai_mai_n502_), .Y(mai_mai_n736_));
  NA2        m714(.A(mai_mai_n736_), .B(mai_mai_n735_), .Y(mai_mai_n737_));
  OR2        m715(.A(mai_mai_n737_), .B(mai_mai_n733_), .Y(mai_mai_n738_));
  NO2        m716(.A(i_11_), .B(i_2_), .Y(mai_mai_n739_));
  NA2        m717(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n740_));
  OAI210     m718(.A0(mai_mai_n740_), .A1(mai_mai_n362_), .B0(mai_mai_n315_), .Y(mai_mai_n741_));
  NA2        m719(.A(mai_mai_n741_), .B(mai_mai_n739_), .Y(mai_mai_n742_));
  NA3        m720(.A(mai_mai_n308_), .B(mai_mai_n234_), .C(i_7_), .Y(mai_mai_n743_));
  NA2        m721(.A(mai_mai_n400_), .B(mai_mai_n136_), .Y(mai_mai_n744_));
  AO210      m722(.A0(mai_mai_n437_), .A1(mai_mai_n684_), .B0(mai_mai_n36_), .Y(mai_mai_n745_));
  NA4        m723(.A(mai_mai_n745_), .B(mai_mai_n744_), .C(mai_mai_n743_), .D(mai_mai_n742_), .Y(mai_mai_n746_));
  AOI220     m724(.A0(mai_mai_n952_), .A1(mai_mai_n502_), .B0(mai_mai_n722_), .B1(mai_mai_n648_), .Y(mai_mai_n747_));
  NA3        m725(.A(mai_mai_n329_), .B(mai_mai_n219_), .C(mai_mai_n136_), .Y(mai_mai_n748_));
  NA3        m726(.A(mai_mai_n748_), .B(mai_mai_n747_), .C(mai_mai_n541_), .Y(mai_mai_n749_));
  AO210      m727(.A0(i_4_), .A1(mai_mai_n46_), .B0(mai_mai_n80_), .Y(mai_mai_n750_));
  NA3        m728(.A(mai_mai_n750_), .B(mai_mai_n428_), .C(mai_mai_n202_), .Y(mai_mai_n751_));
  AOI210     m729(.A0(mai_mai_n400_), .A1(mai_mai_n398_), .B0(mai_mai_n501_), .Y(mai_mai_n752_));
  OAI210     m730(.A0(mai_mai_n954_), .A1(mai_mai_n104_), .B0(mai_mai_n361_), .Y(mai_mai_n753_));
  NA2        m731(.A(i_0_), .B(mai_mai_n526_), .Y(mai_mai_n754_));
  NA3        m732(.A(mai_mai_n754_), .B(mai_mai_n295_), .C(i_7_), .Y(mai_mai_n755_));
  NA4        m733(.A(mai_mai_n755_), .B(mai_mai_n753_), .C(mai_mai_n752_), .D(mai_mai_n751_), .Y(mai_mai_n756_));
  NO4        m734(.A(mai_mai_n756_), .B(mai_mai_n749_), .C(mai_mai_n746_), .D(mai_mai_n738_), .Y(mai_mai_n757_));
  NA4        m735(.A(mai_mai_n757_), .B(mai_mai_n731_), .C(mai_mai_n725_), .D(mai_mai_n337_), .Y(mai3));
  NA2        m736(.A(i_6_), .B(i_7_), .Y(mai_mai_n759_));
  NO2        m737(.A(mai_mai_n759_), .B(i_0_), .Y(mai_mai_n760_));
  NO2        m738(.A(i_11_), .B(mai_mai_n218_), .Y(mai_mai_n761_));
  OAI210     m739(.A0(mai_mai_n760_), .A1(mai_mai_n266_), .B0(mai_mai_n761_), .Y(mai_mai_n762_));
  NO2        m740(.A(mai_mai_n762_), .B(mai_mai_n178_), .Y(mai_mai_n763_));
  AN2        m741(.A(mai_mai_n763_), .B(mai_mai_n160_), .Y(mai_mai_n764_));
  NA3        m742(.A(mai_mai_n748_), .B(mai_mai_n541_), .C(mai_mai_n328_), .Y(mai_mai_n765_));
  NA2        m743(.A(mai_mai_n765_), .B(mai_mai_n39_), .Y(mai_mai_n766_));
  NO3        m744(.A(mai_mai_n568_), .B(mai_mai_n407_), .C(mai_mai_n120_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n363_), .B(mai_mai_n45_), .Y(mai_mai_n768_));
  AN2        m746(.A(mai_mai_n405_), .B(mai_mai_n54_), .Y(mai_mai_n769_));
  NO2        m747(.A(mai_mai_n769_), .B(mai_mai_n767_), .Y(mai_mai_n770_));
  AOI210     m748(.A0(mai_mai_n770_), .A1(mai_mai_n766_), .B0(mai_mai_n48_), .Y(mai_mai_n771_));
  NO4        m749(.A(mai_mai_n333_), .B(mai_mai_n340_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n772_));
  NA2        m750(.A(mai_mai_n640_), .B(mai_mai_n609_), .Y(mai_mai_n773_));
  NA2        m751(.A(i_0_), .B(i_5_), .Y(mai_mai_n774_));
  OAI220     m752(.A0(mai_mai_n774_), .A1(mai_mai_n773_), .B0(mai_mai_n948_), .B1(mai_mai_n62_), .Y(mai_mai_n775_));
  NOi21      m753(.An(i_5_), .B(i_9_), .Y(mai_mai_n776_));
  NA2        m754(.A(mai_mai_n776_), .B(mai_mai_n396_), .Y(mai_mai_n777_));
  NO3        m755(.A(mai_mai_n364_), .B(mai_mai_n246_), .C(mai_mai_n68_), .Y(mai_mai_n778_));
  NO2        m756(.A(mai_mai_n161_), .B(mai_mai_n137_), .Y(mai_mai_n779_));
  AOI210     m757(.A0(mai_mai_n779_), .A1(mai_mai_n223_), .B0(mai_mai_n778_), .Y(mai_mai_n780_));
  OAI220     m758(.A0(mai_mai_n780_), .A1(mai_mai_n166_), .B0(mai_mai_n543_), .B1(mai_mai_n777_), .Y(mai_mai_n781_));
  NO4        m759(.A(mai_mai_n781_), .B(mai_mai_n775_), .C(mai_mai_n771_), .D(mai_mai_n764_), .Y(mai_mai_n782_));
  INV        m760(.A(mai_mai_n282_), .Y(mai_mai_n783_));
  NAi21      m761(.An(mai_mai_n150_), .B(i_5_), .Y(mai_mai_n784_));
  OAI220     m762(.A0(mai_mai_n784_), .A1(i_0_), .B0(mai_mai_n783_), .B1(mai_mai_n355_), .Y(mai_mai_n785_));
  INV        m763(.A(mai_mai_n785_), .Y(mai_mai_n786_));
  NA2        m764(.A(mai_mai_n511_), .B(i_0_), .Y(mai_mai_n787_));
  NO3        m765(.A(mai_mai_n787_), .B(mai_mai_n342_), .C(mai_mai_n81_), .Y(mai_mai_n788_));
  NO4        m766(.A(i_5_), .B(i_12_), .C(mai_mai_n368_), .D(mai_mai_n362_), .Y(mai_mai_n789_));
  AOI210     m767(.A0(mai_mai_n789_), .A1(i_11_), .B0(mai_mai_n788_), .Y(mai_mai_n790_));
  NA2        m768(.A(mai_mai_n680_), .B(mai_mai_n296_), .Y(mai_mai_n791_));
  NO2        m769(.A(mai_mai_n428_), .B(mai_mai_n57_), .Y(mai_mai_n792_));
  NO2        m770(.A(mai_mai_n792_), .B(mai_mai_n791_), .Y(mai_mai_n793_));
  NO2        m771(.A(mai_mai_n232_), .B(mai_mai_n141_), .Y(mai_mai_n794_));
  INV        m772(.A(mai_mai_n478_), .Y(mai_mai_n795_));
  NO4        m773(.A(mai_mai_n107_), .B(mai_mai_n57_), .C(mai_mai_n605_), .D(i_5_), .Y(mai_mai_n796_));
  AO220      m774(.A0(mai_mai_n796_), .A1(mai_mai_n795_), .B0(mai_mai_n794_), .B1(i_6_), .Y(mai_mai_n797_));
  AOI210     m775(.A0(i_0_), .A1(mai_mai_n90_), .B0(mai_mai_n170_), .Y(mai_mai_n798_));
  NA2        m776(.A(mai_mai_n506_), .B(i_4_), .Y(mai_mai_n799_));
  NA2        m777(.A(mai_mai_n173_), .B(mai_mai_n187_), .Y(mai_mai_n800_));
  OAI220     m778(.A0(mai_mai_n800_), .A1(mai_mai_n791_), .B0(mai_mai_n799_), .B1(mai_mai_n798_), .Y(mai_mai_n801_));
  NO3        m779(.A(mai_mai_n801_), .B(mai_mai_n797_), .C(mai_mai_n793_), .Y(mai_mai_n802_));
  NA3        m780(.A(mai_mai_n802_), .B(mai_mai_n790_), .C(mai_mai_n786_), .Y(mai_mai_n803_));
  NA2        m781(.A(i_11_), .B(i_9_), .Y(mai_mai_n804_));
  NO2        m782(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n805_));
  NA2        m783(.A(mai_mai_n351_), .B(mai_mai_n165_), .Y(mai_mai_n806_));
  NAi31      m784(.An(mai_mai_n243_), .B(mai_mai_n806_), .C(mai_mai_n148_), .Y(mai_mai_n807_));
  NO2        m785(.A(mai_mai_n161_), .B(i_0_), .Y(mai_mai_n808_));
  NA2        m786(.A(mai_mai_n422_), .B(mai_mai_n214_), .Y(mai_mai_n809_));
  OAI220     m787(.A0(i_12_), .A1(mai_mai_n777_), .B0(mai_mai_n809_), .B1(mai_mai_n161_), .Y(mai_mai_n810_));
  NO2        m788(.A(mai_mai_n810_), .B(mai_mai_n807_), .Y(mai_mai_n811_));
  AOI210     m789(.A0(mai_mai_n399_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n812_));
  NA2        m790(.A(mai_mai_n157_), .B(mai_mai_n95_), .Y(mai_mai_n813_));
  NOi32      m791(.An(mai_mai_n812_), .Bn(mai_mai_n173_), .C(mai_mai_n813_), .Y(mai_mai_n814_));
  NO2        m792(.A(mai_mai_n955_), .B(mai_mai_n768_), .Y(mai_mai_n815_));
  NO2        m793(.A(mai_mai_n815_), .B(mai_mai_n814_), .Y(mai_mai_n816_));
  NOi21      m794(.An(i_7_), .B(i_5_), .Y(mai_mai_n817_));
  NOi21      m795(.An(mai_mai_n817_), .B(mai_mai_n659_), .Y(mai_mai_n818_));
  NA3        m796(.A(mai_mai_n818_), .B(mai_mai_n341_), .C(i_6_), .Y(mai_mai_n819_));
  OA210      m797(.A0(mai_mai_n813_), .A1(mai_mai_n462_), .B0(mai_mai_n819_), .Y(mai_mai_n820_));
  NO3        m798(.A(mai_mai_n357_), .B(mai_mai_n317_), .C(mai_mai_n313_), .Y(mai_mai_n821_));
  NO2        m799(.A(mai_mai_n240_), .B(mai_mai_n287_), .Y(mai_mai_n822_));
  INV        m800(.A(mai_mai_n821_), .Y(mai_mai_n823_));
  NA4        m801(.A(mai_mai_n823_), .B(mai_mai_n820_), .C(mai_mai_n816_), .D(mai_mai_n811_), .Y(mai_mai_n824_));
  AN2        m802(.A(mai_mai_n300_), .B(mai_mai_n296_), .Y(mai_mai_n825_));
  AN2        m803(.A(mai_mai_n825_), .B(mai_mai_n779_), .Y(mai_mai_n826_));
  NA2        m804(.A(mai_mai_n826_), .B(i_10_), .Y(mai_mai_n827_));
  OA210      m805(.A0(mai_mai_n422_), .A1(mai_mai_n206_), .B0(mai_mai_n421_), .Y(mai_mai_n828_));
  NA3        m806(.A(mai_mai_n421_), .B(mai_mai_n363_), .C(mai_mai_n45_), .Y(mai_mai_n829_));
  OAI210     m807(.A0(mai_mai_n784_), .A1(mai_mai_n422_), .B0(mai_mai_n829_), .Y(mai_mai_n830_));
  INV        m808(.A(mai_mai_n172_), .Y(mai_mai_n831_));
  AOI220     m809(.A0(mai_mai_n831_), .A1(mai_mai_n422_), .B0(mai_mai_n830_), .B1(mai_mai_n68_), .Y(mai_mai_n832_));
  NA3        m810(.A(mai_mai_n740_), .B(mai_mai_n339_), .C(mai_mai_n578_), .Y(mai_mai_n833_));
  NA2        m811(.A(mai_mai_n85_), .B(mai_mai_n44_), .Y(mai_mai_n834_));
  NO2        m812(.A(mai_mai_n70_), .B(mai_mai_n682_), .Y(mai_mai_n835_));
  NA2        m813(.A(mai_mai_n835_), .B(mai_mai_n834_), .Y(mai_mai_n836_));
  AOI210     m814(.A0(mai_mai_n836_), .A1(mai_mai_n833_), .B0(mai_mai_n47_), .Y(mai_mai_n837_));
  NO3        m815(.A(i_5_), .B(i_0_), .C(mai_mai_n24_), .Y(mai_mai_n838_));
  NO2        m816(.A(mai_mai_n485_), .B(mai_mai_n838_), .Y(mai_mai_n839_));
  NAi21      m817(.An(i_9_), .B(i_5_), .Y(mai_mai_n840_));
  NO2        m818(.A(mai_mai_n840_), .B(mai_mai_n357_), .Y(mai_mai_n841_));
  NO2        m819(.A(mai_mai_n537_), .B(mai_mai_n97_), .Y(mai_mai_n842_));
  AOI220     m820(.A0(mai_mai_n842_), .A1(i_0_), .B0(mai_mai_n841_), .B1(mai_mai_n558_), .Y(mai_mai_n843_));
  OAI220     m821(.A0(mai_mai_n843_), .A1(mai_mai_n78_), .B0(mai_mai_n839_), .B1(mai_mai_n158_), .Y(mai_mai_n844_));
  NO3        m822(.A(mai_mai_n844_), .B(mai_mai_n837_), .C(mai_mai_n464_), .Y(mai_mai_n845_));
  NA3        m823(.A(mai_mai_n845_), .B(mai_mai_n832_), .C(mai_mai_n827_), .Y(mai_mai_n846_));
  NO3        m824(.A(mai_mai_n846_), .B(mai_mai_n824_), .C(mai_mai_n803_), .Y(mai_mai_n847_));
  INV        m825(.A(mai_mai_n659_), .Y(mai_mai_n848_));
  NO3        m826(.A(mai_mai_n97_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n849_));
  AO220      m827(.A0(mai_mai_n849_), .A1(mai_mai_n44_), .B0(mai_mai_n848_), .B1(mai_mai_n160_), .Y(mai_mai_n850_));
  AOI210     m828(.A0(mai_mai_n727_), .A1(mai_mai_n618_), .B0(mai_mai_n813_), .Y(mai_mai_n851_));
  AOI210     m829(.A0(mai_mai_n850_), .A1(mai_mai_n307_), .B0(mai_mai_n851_), .Y(mai_mai_n852_));
  NA3        m830(.A(mai_mai_n135_), .B(mai_mai_n609_), .C(mai_mai_n68_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n736_), .B(mai_mai_n357_), .Y(mai_mai_n854_));
  NA3        m832(.A(mai_mai_n760_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n855_));
  NA2        m833(.A(mai_mai_n761_), .B(i_9_), .Y(mai_mai_n856_));
  AOI210     m834(.A0(mai_mai_n855_), .A1(mai_mai_n441_), .B0(mai_mai_n856_), .Y(mai_mai_n857_));
  NO2        m835(.A(mai_mai_n857_), .B(mai_mai_n854_), .Y(mai_mai_n858_));
  NA3        m836(.A(mai_mai_n858_), .B(mai_mai_n853_), .C(mai_mai_n852_), .Y(mai_mai_n859_));
  AOI210     m837(.A0(mai_mai_n274_), .A1(mai_mai_n150_), .B0(mai_mai_n957_), .Y(mai_mai_n860_));
  NA3        m838(.A(mai_mai_n39_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n861_));
  NA2        m839(.A(mai_mai_n805_), .B(mai_mai_n433_), .Y(mai_mai_n862_));
  AOI210     m840(.A0(mai_mai_n861_), .A1(mai_mai_n150_), .B0(mai_mai_n862_), .Y(mai_mai_n863_));
  NO2        m841(.A(mai_mai_n863_), .B(mai_mai_n860_), .Y(mai_mai_n864_));
  NO3        m842(.A(mai_mai_n194_), .B(mai_mai_n340_), .C(i_0_), .Y(mai_mai_n865_));
  OAI210     m843(.A0(mai_mai_n865_), .A1(mai_mai_n71_), .B0(i_13_), .Y(mai_mai_n866_));
  INV        m844(.A(mai_mai_n202_), .Y(mai_mai_n867_));
  OAI220     m845(.A0(mai_mai_n473_), .A1(mai_mai_n128_), .B0(i_12_), .B1(mai_mai_n552_), .Y(mai_mai_n868_));
  NA3        m846(.A(mai_mai_n868_), .B(i_7_), .C(mai_mai_n867_), .Y(mai_mai_n869_));
  NA3        m847(.A(mai_mai_n869_), .B(mai_mai_n866_), .C(mai_mai_n864_), .Y(mai_mai_n870_));
  NO2        m848(.A(mai_mai_n222_), .B(mai_mai_n85_), .Y(mai_mai_n871_));
  AOI210     m849(.A0(mai_mai_n871_), .A1(mai_mai_n848_), .B0(mai_mai_n101_), .Y(mai_mai_n872_));
  AOI220     m850(.A0(mai_mai_n817_), .A1(mai_mai_n433_), .B0(mai_mai_n760_), .B1(mai_mai_n151_), .Y(mai_mai_n873_));
  NA2        m851(.A(mai_mai_n308_), .B(mai_mai_n162_), .Y(mai_mai_n874_));
  OA220      m852(.A0(mai_mai_n874_), .A1(mai_mai_n873_), .B0(mai_mai_n872_), .B1(i_5_), .Y(mai_mai_n875_));
  AOI210     m853(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n161_), .Y(mai_mai_n876_));
  NA2        m854(.A(mai_mai_n876_), .B(mai_mai_n828_), .Y(mai_mai_n877_));
  NA2        m855(.A(mai_mai_n549_), .B(mai_mai_n170_), .Y(mai_mai_n878_));
  NA2        m856(.A(mai_mai_n878_), .B(mai_mai_n484_), .Y(mai_mai_n879_));
  NO3        m857(.A(mai_mai_n768_), .B(mai_mai_n53_), .C(mai_mai_n48_), .Y(mai_mai_n880_));
  NA2        m858(.A(mai_mai_n431_), .B(mai_mai_n419_), .Y(mai_mai_n881_));
  NO3        m859(.A(mai_mai_n881_), .B(mai_mai_n880_), .C(mai_mai_n879_), .Y(mai_mai_n882_));
  NA3        m860(.A(mai_mai_n347_), .B(mai_mai_n301_), .C(mai_mai_n205_), .Y(mai_mai_n883_));
  INV        m861(.A(mai_mai_n883_), .Y(mai_mai_n884_));
  NOi31      m862(.An(mai_mai_n346_), .B(i_11_), .C(mai_mai_n220_), .Y(mai_mai_n885_));
  NO3        m863(.A(mai_mai_n804_), .B(mai_mai_n202_), .C(mai_mai_n175_), .Y(mai_mai_n886_));
  NO3        m864(.A(mai_mai_n886_), .B(mai_mai_n885_), .C(mai_mai_n884_), .Y(mai_mai_n887_));
  NA4        m865(.A(mai_mai_n887_), .B(mai_mai_n882_), .C(mai_mai_n877_), .D(mai_mai_n875_), .Y(mai_mai_n888_));
  INV        m866(.A(mai_mai_n551_), .Y(mai_mai_n889_));
  NO3        m867(.A(mai_mai_n889_), .B(mai_mai_n497_), .C(i_7_), .Y(mai_mai_n890_));
  NO2        m868(.A(mai_mai_n78_), .B(i_5_), .Y(mai_mai_n891_));
  NA3        m869(.A(mai_mai_n761_), .B(mai_mai_n102_), .C(mai_mai_n115_), .Y(mai_mai_n892_));
  INV        m870(.A(mai_mai_n892_), .Y(mai_mai_n893_));
  AOI210     m871(.A0(mai_mai_n893_), .A1(mai_mai_n891_), .B0(mai_mai_n890_), .Y(mai_mai_n894_));
  NA3        m872(.A(mai_mai_n276_), .B(i_5_), .C(mai_mai_n178_), .Y(mai_mai_n895_));
  NO4        m873(.A(mai_mai_n220_), .B(mai_mai_n194_), .C(i_0_), .D(i_12_), .Y(mai_mai_n896_));
  AOI220     m874(.A0(mai_mai_n896_), .A1(mai_mai_n945_), .B0(mai_mai_n721_), .B1(mai_mai_n162_), .Y(mai_mai_n897_));
  BUFFER     m875(.A(mai_mai_n141_), .Y(mai_mai_n898_));
  NO4        m876(.A(mai_mai_n898_), .B(i_12_), .C(mai_mai_n586_), .D(mai_mai_n120_), .Y(mai_mai_n899_));
  NA2        m877(.A(mai_mai_n899_), .B(mai_mai_n202_), .Y(mai_mai_n900_));
  NA2        m878(.A(mai_mai_n817_), .B(mai_mai_n418_), .Y(mai_mai_n901_));
  OAI210     m879(.A0(i_6_), .A1(mai_mai_n895_), .B0(mai_mai_n901_), .Y(mai_mai_n902_));
  NA2        m880(.A(mai_mai_n902_), .B(mai_mai_n808_), .Y(mai_mai_n903_));
  NA4        m881(.A(mai_mai_n903_), .B(mai_mai_n900_), .C(mai_mai_n897_), .D(mai_mai_n894_), .Y(mai_mai_n904_));
  NO4        m882(.A(mai_mai_n904_), .B(mai_mai_n888_), .C(mai_mai_n870_), .D(mai_mai_n859_), .Y(mai_mai_n905_));
  OAI210     m883(.A0(mai_mai_n739_), .A1(mai_mai_n734_), .B0(mai_mai_n37_), .Y(mai_mai_n906_));
  NA3        m884(.A(mai_mai_n812_), .B(mai_mai_n324_), .C(i_5_), .Y(mai_mai_n907_));
  NA3        m885(.A(mai_mai_n907_), .B(mai_mai_n906_), .C(mai_mai_n547_), .Y(mai_mai_n908_));
  NA2        m886(.A(mai_mai_n908_), .B(mai_mai_n191_), .Y(mai_mai_n909_));
  NA2        m887(.A(mai_mai_n171_), .B(mai_mai_n173_), .Y(mai_mai_n910_));
  OAI210     m888(.A0(mai_mai_n551_), .A1(mai_mai_n549_), .B0(mai_mai_n286_), .Y(mai_mai_n911_));
  INV        m889(.A(mai_mai_n583_), .Y(mai_mai_n912_));
  NA3        m890(.A(mai_mai_n912_), .B(mai_mai_n911_), .C(mai_mai_n910_), .Y(mai_mai_n913_));
  NO2        m891(.A(mai_mai_n411_), .B(mai_mai_n246_), .Y(mai_mai_n914_));
  NO2        m892(.A(mai_mai_n914_), .B(mai_mai_n789_), .Y(mai_mai_n915_));
  INV        m893(.A(mai_mai_n915_), .Y(mai_mai_n916_));
  AOI210     m894(.A0(mai_mai_n913_), .A1(mai_mai_n48_), .B0(mai_mai_n916_), .Y(mai_mai_n917_));
  AOI210     m895(.A0(mai_mai_n917_), .A1(mai_mai_n909_), .B0(mai_mai_n68_), .Y(mai_mai_n918_));
  NO2        m896(.A(mai_mai_n504_), .B(mai_mai_n336_), .Y(mai_mai_n919_));
  NO2        m897(.A(mai_mai_n919_), .B(mai_mai_n688_), .Y(mai_mai_n920_));
  AOI210     m898(.A0(mai_mai_n876_), .A1(mai_mai_n805_), .B0(mai_mai_n818_), .Y(mai_mai_n921_));
  NO2        m899(.A(mai_mai_n921_), .B(mai_mai_n610_), .Y(mai_mai_n922_));
  INV        m900(.A(mai_mai_n56_), .Y(mai_mai_n923_));
  NA2        m901(.A(mai_mai_n923_), .B(mai_mai_n71_), .Y(mai_mai_n924_));
  NO2        m902(.A(mai_mai_n924_), .B(mai_mai_n218_), .Y(mai_mai_n925_));
  NO2        m903(.A(mai_mai_n925_), .B(mai_mai_n922_), .Y(mai_mai_n926_));
  OAI210     m904(.A0(mai_mai_n248_), .A1(mai_mai_n146_), .B0(mai_mai_n81_), .Y(mai_mai_n927_));
  NO2        m905(.A(mai_mai_n927_), .B(i_11_), .Y(mai_mai_n928_));
  OAI210     m906(.A0(mai_mai_n946_), .A1(mai_mai_n812_), .B0(mai_mai_n191_), .Y(mai_mai_n929_));
  NA2        m907(.A(i_0_), .B(i_5_), .Y(mai_mai_n930_));
  AOI210     m908(.A0(mai_mai_n929_), .A1(mai_mai_n705_), .B0(mai_mai_n930_), .Y(mai_mai_n931_));
  NO3        m909(.A(mai_mai_n58_), .B(mai_mai_n57_), .C(i_4_), .Y(mai_mai_n932_));
  OAI210     m910(.A0(mai_mai_n822_), .A1(mai_mai_n953_), .B0(mai_mai_n932_), .Y(mai_mai_n933_));
  NO2        m911(.A(mai_mai_n933_), .B(mai_mai_n659_), .Y(mai_mai_n934_));
  NO4        m912(.A(mai_mai_n840_), .B(mai_mai_n424_), .C(mai_mai_n231_), .D(mai_mai_n230_), .Y(mai_mai_n935_));
  NO2        m913(.A(mai_mai_n935_), .B(mai_mai_n501_), .Y(mai_mai_n936_));
  INV        m914(.A(mai_mai_n318_), .Y(mai_mai_n937_));
  AOI210     m915(.A0(mai_mai_n937_), .A1(mai_mai_n936_), .B0(mai_mai_n40_), .Y(mai_mai_n938_));
  NO4        m916(.A(mai_mai_n938_), .B(mai_mai_n934_), .C(mai_mai_n931_), .D(mai_mai_n928_), .Y(mai_mai_n939_));
  OAI210     m917(.A0(mai_mai_n926_), .A1(i_4_), .B0(mai_mai_n939_), .Y(mai_mai_n940_));
  NO3        m918(.A(mai_mai_n940_), .B(mai_mai_n920_), .C(mai_mai_n918_), .Y(mai_mai_n941_));
  NA4        m919(.A(mai_mai_n941_), .B(mai_mai_n905_), .C(mai_mai_n847_), .D(mai_mai_n782_), .Y(mai4));
  INV        m920(.A(mai_mai_n222_), .Y(mai_mai_n945_));
  INV        m921(.A(i_12_), .Y(mai_mai_n946_));
  INV        m922(.A(i_9_), .Y(mai_mai_n947_));
  INV        m923(.A(mai_mai_n772_), .Y(mai_mai_n948_));
  INV        m924(.A(mai_mai_n120_), .Y(mai_mai_n949_));
  INV        m925(.A(i_1_), .Y(mai_mai_n950_));
  INV        m926(.A(mai_mai_n133_), .Y(mai_mai_n951_));
  INV        m927(.A(i_11_), .Y(mai_mai_n952_));
  INV        m928(.A(i_5_), .Y(mai_mai_n953_));
  INV        m929(.A(mai_mai_n548_), .Y(mai_mai_n954_));
  INV        m930(.A(mai_mai_n296_), .Y(mai_mai_n955_));
  INV        m931(.A(mai_mai_n190_), .Y(mai_mai_n956_));
  INV        m932(.A(mai_mai_n296_), .Y(mai_mai_n957_));
  INV        m933(.A(i_1_), .Y(mai_mai_n958_));
  INV        m934(.A(i_9_), .Y(mai_mai_n959_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u0033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  OAI210     u0034(.A0(men_men_n56_), .A1(men_men_n53_), .B0(men_men_n46_), .Y(men_men_n57_));
  NA3        u0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n58_));
  NO2        u0036(.A(i_1_), .B(i_6_), .Y(men_men_n59_));
  NA2        u0037(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  NA2        u0038(.A(i_8_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n51_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(i_3_), .B(i_9_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_7_), .Y(men_men_n83_));
  NO3        u0061(.A(men_men_n83_), .B(men_men_n82_), .C(men_men_n63_), .Y(men_men_n84_));
  INV        u0062(.A(i_6_), .Y(men_men_n85_));
  OR4        u0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n86_));
  INV        u0064(.A(men_men_n86_), .Y(men_men_n87_));
  NO2        u0065(.A(i_2_), .B(i_7_), .Y(men_men_n88_));
  OAI210     u0066(.A0(men_men_n84_), .A1(i_8_), .B0(men_men_n86_), .Y(men_men_n89_));
  NAi21      u0067(.An(i_6_), .B(i_10_), .Y(men_men_n90_));
  NA2        u0068(.A(i_6_), .B(i_9_), .Y(men_men_n91_));
  AOI210     u0069(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n63_), .Y(men_men_n92_));
  NA2        u0070(.A(i_2_), .B(i_6_), .Y(men_men_n93_));
  NO3        u0071(.A(men_men_n93_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n94_));
  NO2        u0072(.A(men_men_n94_), .B(men_men_n92_), .Y(men_men_n95_));
  AOI210     u0073(.A0(men_men_n95_), .A1(men_men_n89_), .B0(men_men_n80_), .Y(men_men_n96_));
  AN3        u0074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n97_));
  NAi21      u0075(.An(i_6_), .B(i_11_), .Y(men_men_n98_));
  NO2        u0076(.A(i_5_), .B(i_8_), .Y(men_men_n99_));
  NOi21      u0077(.An(men_men_n99_), .B(men_men_n98_), .Y(men_men_n100_));
  AOI220     u0078(.A0(men_men_n100_), .A1(men_men_n62_), .B0(men_men_n97_), .B1(men_men_n32_), .Y(men_men_n101_));
  INV        u0079(.A(i_7_), .Y(men_men_n102_));
  NA2        u0080(.A(men_men_n47_), .B(men_men_n102_), .Y(men_men_n103_));
  NO2        u0081(.A(i_0_), .B(i_5_), .Y(men_men_n104_));
  NO2        u0082(.A(men_men_n104_), .B(men_men_n85_), .Y(men_men_n105_));
  NA2        u0083(.A(i_12_), .B(i_3_), .Y(men_men_n106_));
  NAi21      u0084(.An(i_7_), .B(i_11_), .Y(men_men_n107_));
  NO3        u0085(.A(men_men_n107_), .B(men_men_n90_), .C(men_men_n54_), .Y(men_men_n108_));
  AN2        u0086(.A(i_2_), .B(i_10_), .Y(men_men_n109_));
  OR2        u0087(.A(men_men_n80_), .B(men_men_n59_), .Y(men_men_n110_));
  NO2        u0088(.A(i_8_), .B(men_men_n102_), .Y(men_men_n111_));
  NA2        u0089(.A(i_12_), .B(i_7_), .Y(men_men_n112_));
  NO2        u0090(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n113_));
  NA2        u0091(.A(men_men_n113_), .B(i_0_), .Y(men_men_n114_));
  NA2        u0092(.A(i_11_), .B(i_12_), .Y(men_men_n115_));
  OAI210     u0093(.A0(men_men_n114_), .A1(men_men_n112_), .B0(men_men_n115_), .Y(men_men_n116_));
  INV        u0094(.A(men_men_n116_), .Y(men_men_n117_));
  NAi31      u0095(.An(men_men_n108_), .B(men_men_n117_), .C(men_men_n101_), .Y(men_men_n118_));
  NOi21      u0096(.An(i_1_), .B(i_5_), .Y(men_men_n119_));
  NA2        u0097(.A(men_men_n119_), .B(i_11_), .Y(men_men_n120_));
  NA2        u0098(.A(men_men_n102_), .B(men_men_n37_), .Y(men_men_n121_));
  NA2        u0099(.A(i_7_), .B(men_men_n25_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NO2        u0101(.A(men_men_n123_), .B(men_men_n47_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n125_));
  NAi21      u0103(.An(i_3_), .B(i_8_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n126_), .B(men_men_n62_), .Y(men_men_n127_));
  NOi31      u0105(.An(men_men_n127_), .B(men_men_n125_), .C(men_men_n124_), .Y(men_men_n128_));
  NO2        u0106(.A(i_1_), .B(men_men_n85_), .Y(men_men_n129_));
  NO2        u0107(.A(i_6_), .B(i_5_), .Y(men_men_n130_));
  NA2        u0108(.A(men_men_n130_), .B(i_3_), .Y(men_men_n131_));
  AO210      u0109(.A0(men_men_n131_), .A1(men_men_n48_), .B0(men_men_n129_), .Y(men_men_n132_));
  OAI220     u0110(.A0(men_men_n132_), .A1(men_men_n107_), .B0(men_men_n128_), .B1(men_men_n120_), .Y(men_men_n133_));
  NO3        u0111(.A(men_men_n133_), .B(men_men_n118_), .C(men_men_n96_), .Y(men_men_n134_));
  NA3        u0112(.A(men_men_n134_), .B(men_men_n79_), .C(men_men_n57_), .Y(men2));
  NO2        u0113(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n136_));
  NA2        u0114(.A(i_6_), .B(men_men_n25_), .Y(men_men_n137_));
  NA2        u0115(.A(men_men_n137_), .B(men_men_n136_), .Y(men_men_n138_));
  NA4        u0116(.A(men_men_n138_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0117(.A(i_8_), .B(i_7_), .Y(men_men_n140_));
  NA2        u0118(.A(men_men_n140_), .B(i_6_), .Y(men_men_n141_));
  NO2        u0119(.A(i_12_), .B(i_13_), .Y(men_men_n142_));
  NAi21      u0120(.An(i_5_), .B(i_11_), .Y(men_men_n143_));
  NOi21      u0121(.An(men_men_n142_), .B(men_men_n143_), .Y(men_men_n144_));
  NO2        u0122(.A(i_0_), .B(i_1_), .Y(men_men_n145_));
  NA2        u0123(.A(i_2_), .B(i_3_), .Y(men_men_n146_));
  NO2        u0124(.A(men_men_n146_), .B(i_4_), .Y(men_men_n147_));
  NA3        u0125(.A(men_men_n147_), .B(men_men_n145_), .C(men_men_n144_), .Y(men_men_n148_));
  OR2        u0126(.A(men_men_n148_), .B(men_men_n25_), .Y(men_men_n149_));
  AN2        u0127(.A(men_men_n142_), .B(men_men_n82_), .Y(men_men_n150_));
  NO2        u0128(.A(men_men_n150_), .B(men_men_n27_), .Y(men_men_n151_));
  NA2        u0129(.A(i_1_), .B(i_5_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n73_), .B(men_men_n47_), .Y(men_men_n153_));
  NA2        u0131(.A(men_men_n153_), .B(men_men_n36_), .Y(men_men_n154_));
  NO3        u0132(.A(men_men_n154_), .B(men_men_n152_), .C(men_men_n151_), .Y(men_men_n155_));
  OR2        u0133(.A(i_0_), .B(i_1_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n156_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n157_));
  NAi32      u0135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n158_));
  NAi21      u0136(.An(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NOi21      u0137(.An(i_4_), .B(i_10_), .Y(men_men_n160_));
  NA2        u0138(.A(men_men_n160_), .B(men_men_n40_), .Y(men_men_n161_));
  NO2        u0139(.A(i_3_), .B(i_5_), .Y(men_men_n162_));
  NO3        u0140(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n163_));
  NA2        u0141(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  OAI210     u0142(.A0(men_men_n164_), .A1(men_men_n161_), .B0(men_men_n159_), .Y(men_men_n165_));
  NO2        u0143(.A(men_men_n165_), .B(men_men_n155_), .Y(men_men_n166_));
  AOI210     u0144(.A0(men_men_n166_), .A1(men_men_n149_), .B0(men_men_n141_), .Y(men_men_n167_));
  NA3        u0145(.A(men_men_n73_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n168_));
  NA2        u0146(.A(i_3_), .B(men_men_n49_), .Y(men_men_n169_));
  NOi21      u0147(.An(i_4_), .B(i_9_), .Y(men_men_n170_));
  NOi21      u0148(.An(i_11_), .B(i_13_), .Y(men_men_n171_));
  NA2        u0149(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  OR2        u0150(.A(men_men_n172_), .B(men_men_n169_), .Y(men_men_n173_));
  NO2        u0151(.A(i_4_), .B(i_5_), .Y(men_men_n174_));
  NAi21      u0152(.An(i_12_), .B(i_11_), .Y(men_men_n175_));
  NO2        u0153(.A(men_men_n175_), .B(i_13_), .Y(men_men_n176_));
  NA3        u0154(.A(men_men_n176_), .B(men_men_n174_), .C(men_men_n82_), .Y(men_men_n177_));
  AOI210     u0155(.A0(men_men_n177_), .A1(men_men_n173_), .B0(men_men_n168_), .Y(men_men_n178_));
  NO2        u0156(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n179_));
  NA2        u0157(.A(men_men_n179_), .B(men_men_n47_), .Y(men_men_n180_));
  NA2        u0158(.A(men_men_n36_), .B(i_5_), .Y(men_men_n181_));
  NAi31      u0159(.An(men_men_n181_), .B(men_men_n150_), .C(i_11_), .Y(men_men_n182_));
  NA2        u0160(.A(i_3_), .B(i_5_), .Y(men_men_n183_));
  OR2        u0161(.A(men_men_n183_), .B(men_men_n172_), .Y(men_men_n184_));
  AOI210     u0162(.A0(men_men_n184_), .A1(men_men_n182_), .B0(men_men_n180_), .Y(men_men_n185_));
  NO2        u0163(.A(men_men_n73_), .B(i_5_), .Y(men_men_n186_));
  NO2        u0164(.A(i_13_), .B(i_10_), .Y(men_men_n187_));
  NA3        u0165(.A(men_men_n187_), .B(men_men_n186_), .C(men_men_n45_), .Y(men_men_n188_));
  NO2        u0166(.A(i_2_), .B(i_1_), .Y(men_men_n189_));
  NA2        u0167(.A(men_men_n189_), .B(i_3_), .Y(men_men_n190_));
  NAi21      u0168(.An(i_4_), .B(i_12_), .Y(men_men_n191_));
  NO4        u0169(.A(men_men_n191_), .B(men_men_n190_), .C(men_men_n188_), .D(men_men_n25_), .Y(men_men_n192_));
  NO3        u0170(.A(men_men_n192_), .B(men_men_n185_), .C(men_men_n178_), .Y(men_men_n193_));
  INV        u0171(.A(i_8_), .Y(men_men_n194_));
  NO2        u0172(.A(men_men_n194_), .B(i_7_), .Y(men_men_n195_));
  NA2        u0173(.A(men_men_n195_), .B(i_6_), .Y(men_men_n196_));
  NO3        u0174(.A(i_3_), .B(men_men_n85_), .C(men_men_n49_), .Y(men_men_n197_));
  NA2        u0175(.A(men_men_n197_), .B(men_men_n111_), .Y(men_men_n198_));
  NO3        u0176(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n199_));
  NA3        u0177(.A(men_men_n199_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n200_));
  NO3        u0178(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n201_));
  OAI210     u0179(.A0(men_men_n97_), .A1(i_12_), .B0(men_men_n201_), .Y(men_men_n202_));
  AOI210     u0180(.A0(men_men_n202_), .A1(men_men_n200_), .B0(men_men_n198_), .Y(men_men_n203_));
  NO2        u0181(.A(i_3_), .B(i_8_), .Y(men_men_n204_));
  NO3        u0182(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n205_));
  NA3        u0183(.A(men_men_n205_), .B(men_men_n204_), .C(men_men_n40_), .Y(men_men_n206_));
  NO2        u0184(.A(men_men_n104_), .B(men_men_n59_), .Y(men_men_n207_));
  NA2        u0185(.A(men_men_n207_), .B(men_men_n156_), .Y(men_men_n208_));
  NO2        u0186(.A(i_13_), .B(i_9_), .Y(men_men_n209_));
  NA3        u0187(.A(men_men_n209_), .B(i_6_), .C(men_men_n194_), .Y(men_men_n210_));
  NAi21      u0188(.An(i_12_), .B(i_3_), .Y(men_men_n211_));
  OR2        u0189(.A(men_men_n211_), .B(men_men_n210_), .Y(men_men_n212_));
  NO2        u0190(.A(men_men_n45_), .B(i_5_), .Y(men_men_n213_));
  NO3        u0191(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n214_));
  NA3        u0192(.A(men_men_n214_), .B(men_men_n213_), .C(i_10_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(men_men_n212_), .B0(men_men_n208_), .B1(men_men_n206_), .Y(men_men_n216_));
  AOI210     u0194(.A0(men_men_n216_), .A1(i_7_), .B0(men_men_n203_), .Y(men_men_n217_));
  OAI220     u0195(.A0(men_men_n217_), .A1(i_4_), .B0(men_men_n196_), .B1(men_men_n193_), .Y(men_men_n218_));
  NAi21      u0196(.An(i_12_), .B(i_7_), .Y(men_men_n219_));
  NA3        u0197(.A(i_13_), .B(men_men_n194_), .C(i_10_), .Y(men_men_n220_));
  NO2        u0198(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n221_));
  NA2        u0199(.A(i_0_), .B(i_5_), .Y(men_men_n222_));
  NA2        u0200(.A(men_men_n222_), .B(men_men_n105_), .Y(men_men_n223_));
  OAI220     u0201(.A0(men_men_n223_), .A1(men_men_n190_), .B0(men_men_n180_), .B1(men_men_n131_), .Y(men_men_n224_));
  NAi31      u0202(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n36_), .B(i_13_), .Y(men_men_n226_));
  NO2        u0204(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n227_));
  NO2        u0205(.A(men_men_n47_), .B(men_men_n63_), .Y(men_men_n228_));
  NA3        u0206(.A(men_men_n228_), .B(men_men_n227_), .C(men_men_n226_), .Y(men_men_n229_));
  INV        u0207(.A(i_13_), .Y(men_men_n230_));
  NO2        u0208(.A(i_12_), .B(men_men_n230_), .Y(men_men_n231_));
  NA3        u0209(.A(men_men_n231_), .B(men_men_n199_), .C(men_men_n197_), .Y(men_men_n232_));
  OAI210     u0210(.A0(men_men_n229_), .A1(men_men_n225_), .B0(men_men_n232_), .Y(men_men_n233_));
  AOI220     u0211(.A0(men_men_n233_), .A1(men_men_n140_), .B0(men_men_n224_), .B1(men_men_n221_), .Y(men_men_n234_));
  NO2        u0212(.A(i_12_), .B(men_men_n37_), .Y(men_men_n235_));
  NO2        u0213(.A(men_men_n183_), .B(i_4_), .Y(men_men_n236_));
  NA2        u0214(.A(men_men_n236_), .B(men_men_n235_), .Y(men_men_n237_));
  OR2        u0215(.A(i_8_), .B(i_7_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n238_), .B(men_men_n85_), .Y(men_men_n239_));
  NO2        u0217(.A(men_men_n54_), .B(i_1_), .Y(men_men_n240_));
  NA2        u0218(.A(men_men_n240_), .B(men_men_n239_), .Y(men_men_n241_));
  INV        u0219(.A(i_12_), .Y(men_men_n242_));
  NO2        u0220(.A(men_men_n45_), .B(men_men_n242_), .Y(men_men_n243_));
  NO3        u0221(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n244_));
  NA2        u0222(.A(i_2_), .B(i_1_), .Y(men_men_n245_));
  NO2        u0223(.A(men_men_n241_), .B(men_men_n237_), .Y(men_men_n246_));
  NO3        u0224(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n247_));
  NAi21      u0225(.An(i_4_), .B(i_3_), .Y(men_men_n248_));
  NO2        u0226(.A(men_men_n248_), .B(men_men_n75_), .Y(men_men_n249_));
  NO2        u0227(.A(i_0_), .B(i_6_), .Y(men_men_n250_));
  NOi41      u0228(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n251_));
  NA2        u0229(.A(men_men_n251_), .B(men_men_n250_), .Y(men_men_n252_));
  NO2        u0230(.A(men_men_n245_), .B(men_men_n183_), .Y(men_men_n253_));
  NAi21      u0231(.An(men_men_n252_), .B(men_men_n253_), .Y(men_men_n254_));
  INV        u0232(.A(men_men_n254_), .Y(men_men_n255_));
  AOI220     u0233(.A0(men_men_n255_), .A1(men_men_n40_), .B0(men_men_n246_), .B1(men_men_n209_), .Y(men_men_n256_));
  NO2        u0234(.A(i_11_), .B(men_men_n230_), .Y(men_men_n257_));
  NOi21      u0235(.An(i_1_), .B(i_6_), .Y(men_men_n258_));
  NAi21      u0236(.An(i_3_), .B(i_7_), .Y(men_men_n259_));
  NA2        u0237(.A(men_men_n242_), .B(i_9_), .Y(men_men_n260_));
  OR4        u0238(.A(men_men_n260_), .B(men_men_n259_), .C(men_men_n258_), .D(men_men_n186_), .Y(men_men_n261_));
  NO2        u0239(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n262_));
  NO2        u0240(.A(i_12_), .B(i_3_), .Y(men_men_n263_));
  NA2        u0241(.A(men_men_n73_), .B(i_5_), .Y(men_men_n264_));
  NA2        u0242(.A(i_3_), .B(i_9_), .Y(men_men_n265_));
  NAi21      u0243(.An(i_7_), .B(i_10_), .Y(men_men_n266_));
  NO2        u0244(.A(men_men_n266_), .B(men_men_n265_), .Y(men_men_n267_));
  NA3        u0245(.A(men_men_n267_), .B(men_men_n264_), .C(men_men_n64_), .Y(men_men_n268_));
  NA2        u0246(.A(men_men_n268_), .B(men_men_n261_), .Y(men_men_n269_));
  NA3        u0247(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n270_));
  INV        u0248(.A(men_men_n141_), .Y(men_men_n271_));
  NA2        u0249(.A(men_men_n242_), .B(i_13_), .Y(men_men_n272_));
  NO2        u0250(.A(men_men_n272_), .B(men_men_n75_), .Y(men_men_n273_));
  AOI220     u0251(.A0(men_men_n273_), .A1(men_men_n271_), .B0(men_men_n269_), .B1(men_men_n257_), .Y(men_men_n274_));
  NO2        u0252(.A(men_men_n238_), .B(men_men_n37_), .Y(men_men_n275_));
  NA2        u0253(.A(i_12_), .B(i_6_), .Y(men_men_n276_));
  OR2        u0254(.A(i_13_), .B(i_9_), .Y(men_men_n277_));
  NO3        u0255(.A(men_men_n277_), .B(men_men_n276_), .C(men_men_n49_), .Y(men_men_n278_));
  NO2        u0256(.A(men_men_n248_), .B(i_2_), .Y(men_men_n279_));
  NA3        u0257(.A(men_men_n279_), .B(men_men_n278_), .C(men_men_n45_), .Y(men_men_n280_));
  NA2        u0258(.A(men_men_n257_), .B(i_9_), .Y(men_men_n281_));
  OAI210     u0259(.A0(men_men_n73_), .A1(men_men_n281_), .B0(men_men_n280_), .Y(men_men_n282_));
  NA2        u0260(.A(men_men_n153_), .B(men_men_n63_), .Y(men_men_n283_));
  NO3        u0261(.A(i_11_), .B(men_men_n230_), .C(men_men_n25_), .Y(men_men_n284_));
  NO2        u0262(.A(men_men_n259_), .B(i_8_), .Y(men_men_n285_));
  NO2        u0263(.A(i_6_), .B(men_men_n49_), .Y(men_men_n286_));
  NA3        u0264(.A(men_men_n286_), .B(men_men_n285_), .C(men_men_n284_), .Y(men_men_n287_));
  NO3        u0265(.A(men_men_n26_), .B(men_men_n85_), .C(i_5_), .Y(men_men_n288_));
  NA3        u0266(.A(men_men_n288_), .B(men_men_n275_), .C(men_men_n231_), .Y(men_men_n289_));
  AOI210     u0267(.A0(men_men_n289_), .A1(men_men_n287_), .B0(men_men_n283_), .Y(men_men_n290_));
  AOI210     u0268(.A0(men_men_n282_), .A1(men_men_n275_), .B0(men_men_n290_), .Y(men_men_n291_));
  NA4        u0269(.A(men_men_n291_), .B(men_men_n274_), .C(men_men_n256_), .D(men_men_n234_), .Y(men_men_n292_));
  NO3        u0270(.A(i_12_), .B(men_men_n230_), .C(men_men_n37_), .Y(men_men_n293_));
  INV        u0271(.A(men_men_n293_), .Y(men_men_n294_));
  NOi21      u0272(.An(men_men_n162_), .B(men_men_n85_), .Y(men_men_n295_));
  NO3        u0273(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n296_));
  AOI220     u0274(.A0(men_men_n296_), .A1(men_men_n197_), .B0(men_men_n295_), .B1(men_men_n240_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n297_), .B(i_7_), .Y(men_men_n298_));
  NO3        u0276(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n299_));
  NO2        u0277(.A(men_men_n245_), .B(i_0_), .Y(men_men_n300_));
  AOI220     u0278(.A0(men_men_n300_), .A1(men_men_n195_), .B0(men_men_n299_), .B1(men_men_n140_), .Y(men_men_n301_));
  NA2        u0279(.A(men_men_n286_), .B(men_men_n26_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n302_), .B(men_men_n301_), .Y(men_men_n303_));
  NA2        u0281(.A(i_0_), .B(i_1_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n304_), .B(i_2_), .Y(men_men_n305_));
  NO2        u0283(.A(men_men_n60_), .B(i_6_), .Y(men_men_n306_));
  NA3        u0284(.A(men_men_n306_), .B(men_men_n305_), .C(men_men_n162_), .Y(men_men_n307_));
  OAI210     u0285(.A0(men_men_n164_), .A1(men_men_n141_), .B0(men_men_n307_), .Y(men_men_n308_));
  NO3        u0286(.A(men_men_n308_), .B(men_men_n303_), .C(men_men_n298_), .Y(men_men_n309_));
  NO2        u0287(.A(i_3_), .B(i_10_), .Y(men_men_n310_));
  NA3        u0288(.A(men_men_n310_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n311_));
  NO2        u0289(.A(i_2_), .B(men_men_n102_), .Y(men_men_n312_));
  NA2        u0290(.A(i_1_), .B(men_men_n36_), .Y(men_men_n313_));
  NO2        u0291(.A(men_men_n313_), .B(i_8_), .Y(men_men_n314_));
  NOi21      u0292(.An(men_men_n222_), .B(men_men_n104_), .Y(men_men_n315_));
  NA3        u0293(.A(men_men_n315_), .B(men_men_n314_), .C(men_men_n312_), .Y(men_men_n316_));
  AN2        u0294(.A(i_3_), .B(i_10_), .Y(men_men_n317_));
  NA4        u0295(.A(men_men_n317_), .B(men_men_n199_), .C(men_men_n176_), .D(men_men_n174_), .Y(men_men_n318_));
  NO2        u0296(.A(i_5_), .B(men_men_n37_), .Y(men_men_n319_));
  NO2        u0297(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n320_));
  OR2        u0298(.A(men_men_n316_), .B(men_men_n311_), .Y(men_men_n321_));
  OAI220     u0299(.A0(men_men_n321_), .A1(i_6_), .B0(men_men_n309_), .B1(men_men_n294_), .Y(men_men_n322_));
  NO4        u0300(.A(men_men_n322_), .B(men_men_n292_), .C(men_men_n218_), .D(men_men_n167_), .Y(men_men_n323_));
  NO3        u0301(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n324_));
  NO2        u0302(.A(men_men_n60_), .B(men_men_n85_), .Y(men_men_n325_));
  NA2        u0303(.A(men_men_n300_), .B(men_men_n325_), .Y(men_men_n326_));
  NO3        u0304(.A(i_6_), .B(men_men_n194_), .C(i_7_), .Y(men_men_n327_));
  AOI210     u0305(.A0(men_men_n1121_), .A1(men_men_n326_), .B0(men_men_n169_), .Y(men_men_n328_));
  NO2        u0306(.A(i_2_), .B(i_3_), .Y(men_men_n329_));
  OR2        u0307(.A(i_0_), .B(i_5_), .Y(men_men_n330_));
  NA2        u0308(.A(men_men_n222_), .B(men_men_n330_), .Y(men_men_n331_));
  NA4        u0309(.A(men_men_n331_), .B(men_men_n239_), .C(men_men_n329_), .D(i_1_), .Y(men_men_n332_));
  NA3        u0310(.A(men_men_n300_), .B(men_men_n295_), .C(men_men_n111_), .Y(men_men_n333_));
  NAi21      u0311(.An(i_8_), .B(i_7_), .Y(men_men_n334_));
  NO2        u0312(.A(men_men_n334_), .B(i_6_), .Y(men_men_n335_));
  NO2        u0313(.A(men_men_n156_), .B(men_men_n47_), .Y(men_men_n336_));
  NA3        u0314(.A(men_men_n336_), .B(men_men_n335_), .C(men_men_n162_), .Y(men_men_n337_));
  NA3        u0315(.A(men_men_n337_), .B(men_men_n333_), .C(men_men_n332_), .Y(men_men_n338_));
  OAI210     u0316(.A0(men_men_n338_), .A1(men_men_n328_), .B0(i_4_), .Y(men_men_n339_));
  NO2        u0317(.A(i_12_), .B(i_10_), .Y(men_men_n340_));
  NOi21      u0318(.An(i_5_), .B(i_0_), .Y(men_men_n341_));
  AOI210     u0319(.A0(i_2_), .A1(men_men_n49_), .B0(men_men_n102_), .Y(men_men_n342_));
  NO4        u0320(.A(men_men_n342_), .B(men_men_n313_), .C(men_men_n341_), .D(men_men_n126_), .Y(men_men_n343_));
  NA4        u0321(.A(men_men_n83_), .B(men_men_n36_), .C(men_men_n85_), .D(i_8_), .Y(men_men_n344_));
  NA2        u0322(.A(men_men_n343_), .B(men_men_n340_), .Y(men_men_n345_));
  NO2        u0323(.A(i_6_), .B(i_8_), .Y(men_men_n346_));
  NOi21      u0324(.An(i_0_), .B(i_2_), .Y(men_men_n347_));
  AN2        u0325(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NO2        u0326(.A(i_1_), .B(i_7_), .Y(men_men_n349_));
  AO220      u0327(.A0(men_men_n349_), .A1(men_men_n348_), .B0(men_men_n335_), .B1(men_men_n240_), .Y(men_men_n350_));
  NA3        u0328(.A(men_men_n350_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n351_));
  NA3        u0329(.A(men_men_n351_), .B(men_men_n345_), .C(men_men_n339_), .Y(men_men_n352_));
  NO3        u0330(.A(men_men_n238_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n353_));
  NO3        u0331(.A(men_men_n334_), .B(i_2_), .C(i_1_), .Y(men_men_n354_));
  OAI210     u0332(.A0(men_men_n354_), .A1(men_men_n353_), .B0(i_6_), .Y(men_men_n355_));
  NA3        u0333(.A(men_men_n258_), .B(men_men_n312_), .C(men_men_n194_), .Y(men_men_n356_));
  AOI210     u0334(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n331_), .Y(men_men_n357_));
  NOi21      u0335(.An(men_men_n152_), .B(men_men_n105_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n358_), .B(men_men_n122_), .Y(men_men_n359_));
  OAI210     u0337(.A0(men_men_n359_), .A1(men_men_n357_), .B0(i_3_), .Y(men_men_n360_));
  INV        u0338(.A(men_men_n83_), .Y(men_men_n361_));
  NO2        u0339(.A(men_men_n304_), .B(men_men_n81_), .Y(men_men_n362_));
  NA2        u0340(.A(men_men_n362_), .B(men_men_n130_), .Y(men_men_n363_));
  NO2        u0341(.A(men_men_n93_), .B(men_men_n194_), .Y(men_men_n364_));
  NA3        u0342(.A(men_men_n315_), .B(men_men_n364_), .C(men_men_n63_), .Y(men_men_n365_));
  AOI210     u0343(.A0(men_men_n365_), .A1(men_men_n363_), .B0(men_men_n361_), .Y(men_men_n366_));
  NO2        u0344(.A(men_men_n194_), .B(i_9_), .Y(men_men_n367_));
  NA3        u0345(.A(men_men_n367_), .B(men_men_n207_), .C(men_men_n156_), .Y(men_men_n368_));
  NO2        u0346(.A(men_men_n368_), .B(men_men_n47_), .Y(men_men_n369_));
  NO3        u0347(.A(men_men_n369_), .B(men_men_n366_), .C(men_men_n303_), .Y(men_men_n370_));
  AOI210     u0348(.A0(men_men_n370_), .A1(men_men_n360_), .B0(men_men_n161_), .Y(men_men_n371_));
  AOI210     u0349(.A0(men_men_n352_), .A1(men_men_n324_), .B0(men_men_n371_), .Y(men_men_n372_));
  NOi32      u0350(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n373_));
  INV        u0351(.A(men_men_n373_), .Y(men_men_n374_));
  NAi21      u0352(.An(i_0_), .B(i_6_), .Y(men_men_n375_));
  NAi21      u0353(.An(i_1_), .B(i_5_), .Y(men_men_n376_));
  NA2        u0354(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n377_));
  NA2        u0355(.A(men_men_n377_), .B(men_men_n25_), .Y(men_men_n378_));
  OAI210     u0356(.A0(men_men_n378_), .A1(men_men_n158_), .B0(men_men_n252_), .Y(men_men_n379_));
  NAi41      u0357(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n380_));
  OAI220     u0358(.A0(men_men_n380_), .A1(men_men_n376_), .B0(men_men_n225_), .B1(men_men_n158_), .Y(men_men_n381_));
  AOI210     u0359(.A0(men_men_n380_), .A1(men_men_n158_), .B0(men_men_n156_), .Y(men_men_n382_));
  NOi32      u0360(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n383_));
  NAi21      u0361(.An(i_6_), .B(i_1_), .Y(men_men_n384_));
  NA3        u0362(.A(men_men_n384_), .B(men_men_n383_), .C(men_men_n47_), .Y(men_men_n385_));
  NO2        u0363(.A(men_men_n385_), .B(i_0_), .Y(men_men_n386_));
  OR3        u0364(.A(men_men_n386_), .B(men_men_n382_), .C(men_men_n381_), .Y(men_men_n387_));
  NO2        u0365(.A(i_1_), .B(men_men_n102_), .Y(men_men_n388_));
  NAi21      u0366(.An(i_3_), .B(i_4_), .Y(men_men_n389_));
  NO2        u0367(.A(men_men_n389_), .B(i_9_), .Y(men_men_n390_));
  AN2        u0368(.A(i_6_), .B(i_7_), .Y(men_men_n391_));
  OAI210     u0369(.A0(men_men_n391_), .A1(men_men_n388_), .B0(men_men_n390_), .Y(men_men_n392_));
  NA2        u0370(.A(i_2_), .B(i_7_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n389_), .B(i_10_), .Y(men_men_n394_));
  NA3        u0372(.A(men_men_n394_), .B(men_men_n393_), .C(men_men_n250_), .Y(men_men_n395_));
  AOI210     u0373(.A0(men_men_n395_), .A1(men_men_n392_), .B0(men_men_n186_), .Y(men_men_n396_));
  AOI210     u0374(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n397_));
  OAI210     u0375(.A0(men_men_n397_), .A1(men_men_n189_), .B0(men_men_n394_), .Y(men_men_n398_));
  AOI220     u0376(.A0(men_men_n394_), .A1(men_men_n349_), .B0(men_men_n244_), .B1(men_men_n189_), .Y(men_men_n399_));
  AOI210     u0377(.A0(men_men_n399_), .A1(men_men_n398_), .B0(i_5_), .Y(men_men_n400_));
  NO4        u0378(.A(men_men_n400_), .B(men_men_n396_), .C(men_men_n387_), .D(men_men_n379_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n401_), .B(men_men_n374_), .Y(men_men_n402_));
  NO2        u0380(.A(men_men_n60_), .B(men_men_n25_), .Y(men_men_n403_));
  AN2        u0381(.A(i_12_), .B(i_5_), .Y(men_men_n404_));
  NO2        u0382(.A(i_4_), .B(men_men_n26_), .Y(men_men_n405_));
  NA2        u0383(.A(men_men_n405_), .B(men_men_n404_), .Y(men_men_n406_));
  NO2        u0384(.A(i_11_), .B(i_6_), .Y(men_men_n407_));
  NA3        u0385(.A(men_men_n407_), .B(men_men_n336_), .C(men_men_n230_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n408_), .B(men_men_n406_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n248_), .B(i_5_), .Y(men_men_n410_));
  NO2        u0388(.A(i_5_), .B(i_10_), .Y(men_men_n411_));
  AOI220     u0389(.A0(men_men_n411_), .A1(men_men_n279_), .B0(men_men_n410_), .B1(men_men_n199_), .Y(men_men_n412_));
  NA2        u0390(.A(men_men_n142_), .B(men_men_n46_), .Y(men_men_n413_));
  NO2        u0391(.A(men_men_n413_), .B(men_men_n412_), .Y(men_men_n414_));
  OAI210     u0392(.A0(men_men_n414_), .A1(men_men_n409_), .B0(men_men_n403_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n148_), .B(men_men_n85_), .Y(men_men_n417_));
  OAI210     u0395(.A0(men_men_n417_), .A1(men_men_n409_), .B0(men_men_n416_), .Y(men_men_n418_));
  NO3        u0396(.A(men_men_n85_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n419_));
  NO2        u0397(.A(i_3_), .B(men_men_n102_), .Y(men_men_n420_));
  NO2        u0398(.A(i_11_), .B(i_12_), .Y(men_men_n421_));
  NA2        u0399(.A(men_men_n411_), .B(men_men_n242_), .Y(men_men_n422_));
  NA3        u0400(.A(men_men_n111_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n423_));
  OAI220     u0401(.A0(men_men_n423_), .A1(men_men_n225_), .B0(men_men_n422_), .B1(men_men_n344_), .Y(men_men_n424_));
  NAi21      u0402(.An(i_13_), .B(i_0_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n425_), .B(men_men_n245_), .Y(men_men_n426_));
  NA2        u0404(.A(men_men_n424_), .B(men_men_n426_), .Y(men_men_n427_));
  NA3        u0405(.A(men_men_n427_), .B(men_men_n418_), .C(men_men_n415_), .Y(men_men_n428_));
  NA2        u0406(.A(men_men_n45_), .B(men_men_n230_), .Y(men_men_n429_));
  NO3        u0407(.A(i_1_), .B(i_12_), .C(men_men_n85_), .Y(men_men_n430_));
  NO2        u0408(.A(i_0_), .B(i_11_), .Y(men_men_n431_));
  AN2        u0409(.A(i_1_), .B(i_6_), .Y(men_men_n432_));
  NOi21      u0410(.An(i_2_), .B(i_12_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n433_), .B(men_men_n432_), .Y(men_men_n434_));
  NO2        u0412(.A(men_men_n434_), .B(men_men_n1119_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n140_), .B(i_9_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(i_4_), .Y(men_men_n437_));
  NA2        u0415(.A(men_men_n435_), .B(men_men_n437_), .Y(men_men_n438_));
  NAi21      u0416(.An(i_9_), .B(i_4_), .Y(men_men_n439_));
  OR2        u0417(.A(i_13_), .B(i_10_), .Y(men_men_n440_));
  NO3        u0418(.A(men_men_n440_), .B(men_men_n115_), .C(men_men_n439_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n172_), .B(men_men_n121_), .Y(men_men_n442_));
  OR2        u0420(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n443_));
  NO2        u0421(.A(men_men_n102_), .B(men_men_n25_), .Y(men_men_n444_));
  NA2        u0422(.A(men_men_n293_), .B(men_men_n444_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n286_), .B(men_men_n214_), .Y(men_men_n446_));
  OAI220     u0424(.A0(men_men_n446_), .A1(men_men_n443_), .B0(men_men_n445_), .B1(men_men_n358_), .Y(men_men_n447_));
  INV        u0425(.A(men_men_n447_), .Y(men_men_n448_));
  AOI210     u0426(.A0(men_men_n448_), .A1(men_men_n438_), .B0(men_men_n26_), .Y(men_men_n449_));
  NA2        u0427(.A(men_men_n333_), .B(men_men_n332_), .Y(men_men_n450_));
  AOI220     u0428(.A0(men_men_n306_), .A1(men_men_n296_), .B0(men_men_n300_), .B1(men_men_n325_), .Y(men_men_n451_));
  NO2        u0429(.A(men_men_n451_), .B(men_men_n169_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n183_), .B(men_men_n85_), .Y(men_men_n453_));
  AOI220     u0431(.A0(men_men_n453_), .A1(men_men_n305_), .B0(men_men_n288_), .B1(men_men_n214_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n454_), .B(i_7_), .Y(men_men_n455_));
  NO3        u0433(.A(men_men_n455_), .B(men_men_n452_), .C(men_men_n450_), .Y(men_men_n456_));
  NA2        u0434(.A(men_men_n197_), .B(men_men_n97_), .Y(men_men_n457_));
  NA3        u0435(.A(men_men_n336_), .B(men_men_n162_), .C(men_men_n85_), .Y(men_men_n458_));
  AOI210     u0436(.A0(men_men_n458_), .A1(men_men_n457_), .B0(men_men_n334_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n194_), .B(i_10_), .Y(men_men_n460_));
  NA3        u0438(.A(men_men_n264_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n461_));
  NA2        u0439(.A(men_men_n306_), .B(men_men_n240_), .Y(men_men_n462_));
  OAI220     u0440(.A0(men_men_n462_), .A1(men_men_n183_), .B0(men_men_n461_), .B1(men_men_n460_), .Y(men_men_n463_));
  NO2        u0441(.A(i_3_), .B(men_men_n49_), .Y(men_men_n464_));
  NA3        u0442(.A(men_men_n349_), .B(men_men_n348_), .C(men_men_n464_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n327_), .B(men_men_n331_), .Y(men_men_n466_));
  OAI210     u0444(.A0(men_men_n466_), .A1(men_men_n190_), .B0(men_men_n465_), .Y(men_men_n467_));
  NO3        u0445(.A(men_men_n467_), .B(men_men_n463_), .C(men_men_n459_), .Y(men_men_n468_));
  AOI210     u0446(.A0(men_men_n468_), .A1(men_men_n456_), .B0(men_men_n281_), .Y(men_men_n469_));
  NO4        u0447(.A(men_men_n469_), .B(men_men_n449_), .C(men_men_n428_), .D(men_men_n402_), .Y(men_men_n470_));
  NO2        u0448(.A(men_men_n63_), .B(i_4_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n73_), .B(i_13_), .Y(men_men_n472_));
  NA3        u0450(.A(men_men_n472_), .B(men_men_n471_), .C(i_2_), .Y(men_men_n473_));
  NO2        u0451(.A(i_10_), .B(i_9_), .Y(men_men_n474_));
  NAi21      u0452(.An(i_12_), .B(i_8_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n475_), .B(i_3_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n476_), .B(men_men_n474_), .Y(men_men_n477_));
  NO2        u0455(.A(men_men_n47_), .B(i_4_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n478_), .B(men_men_n105_), .Y(men_men_n479_));
  OAI220     u0457(.A0(men_men_n479_), .A1(men_men_n206_), .B0(men_men_n477_), .B1(men_men_n473_), .Y(men_men_n480_));
  NA2        u0458(.A(men_men_n320_), .B(i_0_), .Y(men_men_n481_));
  NO3        u0459(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n276_), .B(men_men_n98_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n483_), .B(men_men_n482_), .Y(men_men_n484_));
  NA2        u0462(.A(i_8_), .B(i_9_), .Y(men_men_n485_));
  AOI210     u0463(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n486_));
  OR2        u0464(.A(men_men_n486_), .B(men_men_n485_), .Y(men_men_n487_));
  NA2        u0465(.A(men_men_n293_), .B(men_men_n207_), .Y(men_men_n488_));
  OAI220     u0466(.A0(men_men_n488_), .A1(men_men_n487_), .B0(men_men_n484_), .B1(men_men_n481_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n257_), .B(men_men_n319_), .Y(men_men_n490_));
  NO3        u0468(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n491_));
  AOI210     u0469(.A0(men_men_n263_), .A1(men_men_n189_), .B0(men_men_n491_), .Y(men_men_n492_));
  NA3        u0470(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n493_));
  NA4        u0471(.A(men_men_n143_), .B(men_men_n113_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n494_));
  OAI220     u0472(.A0(men_men_n494_), .A1(men_men_n493_), .B0(men_men_n492_), .B1(men_men_n490_), .Y(men_men_n495_));
  NO3        u0473(.A(men_men_n495_), .B(men_men_n489_), .C(men_men_n480_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n305_), .B(men_men_n107_), .Y(men_men_n497_));
  OR2        u0475(.A(men_men_n497_), .B(men_men_n210_), .Y(men_men_n498_));
  OA210      u0476(.A0(men_men_n368_), .A1(men_men_n102_), .B0(men_men_n307_), .Y(men_men_n499_));
  OA220      u0477(.A0(men_men_n499_), .A1(men_men_n161_), .B0(men_men_n498_), .B1(men_men_n237_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n97_), .B(i_13_), .Y(men_men_n501_));
  NA2        u0479(.A(men_men_n453_), .B(men_men_n403_), .Y(men_men_n502_));
  NO2        u0480(.A(i_2_), .B(i_13_), .Y(men_men_n503_));
  NA3        u0481(.A(men_men_n503_), .B(men_men_n160_), .C(men_men_n100_), .Y(men_men_n504_));
  OAI220     u0482(.A0(men_men_n504_), .A1(men_men_n242_), .B0(men_men_n502_), .B1(men_men_n501_), .Y(men_men_n505_));
  NO3        u0483(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n506_));
  NO2        u0484(.A(i_6_), .B(i_7_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n507_), .B(men_men_n506_), .Y(men_men_n508_));
  NO2        u0486(.A(i_11_), .B(i_1_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n73_), .B(i_3_), .Y(men_men_n510_));
  OR2        u0488(.A(i_11_), .B(i_8_), .Y(men_men_n511_));
  NOi21      u0489(.An(i_2_), .B(i_7_), .Y(men_men_n512_));
  NAi31      u0490(.An(men_men_n511_), .B(men_men_n512_), .C(men_men_n510_), .Y(men_men_n513_));
  NO2        u0491(.A(men_men_n440_), .B(i_6_), .Y(men_men_n514_));
  NA3        u0492(.A(men_men_n514_), .B(men_men_n471_), .C(men_men_n75_), .Y(men_men_n515_));
  NO2        u0493(.A(men_men_n515_), .B(men_men_n513_), .Y(men_men_n516_));
  NO2        u0494(.A(i_3_), .B(men_men_n194_), .Y(men_men_n517_));
  NO2        u0495(.A(i_6_), .B(i_10_), .Y(men_men_n518_));
  NA4        u0496(.A(men_men_n518_), .B(men_men_n324_), .C(men_men_n517_), .D(men_men_n242_), .Y(men_men_n519_));
  NO2        u0497(.A(men_men_n519_), .B(men_men_n154_), .Y(men_men_n520_));
  NA3        u0498(.A(men_men_n251_), .B(men_men_n171_), .C(men_men_n130_), .Y(men_men_n521_));
  NA2        u0499(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n522_));
  NO2        u0500(.A(men_men_n156_), .B(i_3_), .Y(men_men_n523_));
  NAi31      u0501(.An(men_men_n522_), .B(men_men_n523_), .C(men_men_n231_), .Y(men_men_n524_));
  NA3        u0502(.A(men_men_n416_), .B(men_men_n179_), .C(men_men_n147_), .Y(men_men_n525_));
  NA3        u0503(.A(men_men_n525_), .B(men_men_n524_), .C(men_men_n521_), .Y(men_men_n526_));
  NO4        u0504(.A(men_men_n526_), .B(men_men_n520_), .C(men_men_n516_), .D(men_men_n505_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n491_), .B(men_men_n411_), .Y(men_men_n528_));
  NO2        u0506(.A(men_men_n528_), .B(men_men_n229_), .Y(men_men_n529_));
  NAi21      u0507(.An(men_men_n220_), .B(men_men_n421_), .Y(men_men_n530_));
  NA2        u0508(.A(men_men_n349_), .B(men_men_n222_), .Y(men_men_n531_));
  NO2        u0509(.A(men_men_n26_), .B(i_5_), .Y(men_men_n532_));
  NO2        u0510(.A(i_0_), .B(men_men_n85_), .Y(men_men_n533_));
  NA3        u0511(.A(men_men_n533_), .B(men_men_n532_), .C(men_men_n140_), .Y(men_men_n534_));
  OR3        u0512(.A(men_men_n313_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n535_));
  OAI220     u0513(.A0(men_men_n535_), .A1(men_men_n534_), .B0(men_men_n531_), .B1(men_men_n530_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n27_), .B(i_10_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n324_), .B(men_men_n244_), .Y(men_men_n538_));
  OAI220     u0516(.A0(men_men_n538_), .A1(men_men_n461_), .B0(men_men_n537_), .B1(men_men_n501_), .Y(men_men_n539_));
  NA4        u0517(.A(men_men_n317_), .B(men_men_n228_), .C(men_men_n73_), .D(men_men_n242_), .Y(men_men_n540_));
  NO2        u0518(.A(men_men_n540_), .B(men_men_n508_), .Y(men_men_n541_));
  NO4        u0519(.A(men_men_n541_), .B(men_men_n539_), .C(men_men_n536_), .D(men_men_n529_), .Y(men_men_n542_));
  NA4        u0520(.A(men_men_n542_), .B(men_men_n527_), .C(men_men_n500_), .D(men_men_n496_), .Y(men_men_n543_));
  NA3        u0521(.A(men_men_n317_), .B(men_men_n176_), .C(men_men_n174_), .Y(men_men_n544_));
  OAI210     u0522(.A0(men_men_n311_), .A1(men_men_n181_), .B0(men_men_n544_), .Y(men_men_n545_));
  AN2        u0523(.A(men_men_n296_), .B(men_men_n239_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n546_), .B(men_men_n545_), .Y(men_men_n547_));
  NA2        u0525(.A(men_men_n120_), .B(men_men_n110_), .Y(men_men_n548_));
  AO220      u0526(.A0(men_men_n548_), .A1(men_men_n482_), .B0(men_men_n441_), .B1(i_6_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n324_), .B(men_men_n163_), .Y(men_men_n550_));
  OAI210     u0528(.A0(men_men_n550_), .A1(men_men_n237_), .B0(men_men_n318_), .Y(men_men_n551_));
  AOI220     u0529(.A0(men_men_n551_), .A1(men_men_n335_), .B0(men_men_n549_), .B1(men_men_n320_), .Y(men_men_n552_));
  NA4        u0530(.A(men_men_n472_), .B(men_men_n471_), .C(men_men_n204_), .D(i_2_), .Y(men_men_n553_));
  INV        u0531(.A(men_men_n553_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n404_), .B(men_men_n230_), .Y(men_men_n555_));
  NA2        u0533(.A(men_men_n373_), .B(men_men_n73_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n391_), .B(men_men_n383_), .Y(men_men_n557_));
  AO210      u0535(.A0(men_men_n556_), .A1(men_men_n555_), .B0(men_men_n557_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n36_), .B(i_8_), .Y(men_men_n559_));
  AOI210     u0537(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n441_), .Y(men_men_n560_));
  NA2        u0538(.A(men_men_n560_), .B(men_men_n558_), .Y(men_men_n561_));
  AOI210     u0539(.A0(men_men_n554_), .A1(men_men_n205_), .B0(men_men_n561_), .Y(men_men_n562_));
  NA2        u0540(.A(men_men_n264_), .B(men_men_n64_), .Y(men_men_n563_));
  OAI210     u0541(.A0(i_8_), .A1(men_men_n563_), .B0(men_men_n132_), .Y(men_men_n564_));
  AOI210     u0542(.A0(men_men_n195_), .A1(i_9_), .B0(men_men_n275_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n565_), .B(men_men_n200_), .Y(men_men_n566_));
  OR2        u0544(.A(men_men_n183_), .B(i_4_), .Y(men_men_n567_));
  NO2        u0545(.A(men_men_n567_), .B(men_men_n85_), .Y(men_men_n568_));
  AOI220     u0546(.A0(men_men_n568_), .A1(men_men_n566_), .B0(men_men_n564_), .B1(men_men_n442_), .Y(men_men_n569_));
  NA4        u0547(.A(men_men_n569_), .B(men_men_n562_), .C(men_men_n552_), .D(men_men_n547_), .Y(men_men_n570_));
  NA2        u0548(.A(men_men_n410_), .B(men_men_n305_), .Y(men_men_n571_));
  OAI210     u0549(.A0(men_men_n406_), .A1(men_men_n168_), .B0(men_men_n571_), .Y(men_men_n572_));
  NO2        u0550(.A(i_12_), .B(men_men_n194_), .Y(men_men_n573_));
  NA2        u0551(.A(men_men_n573_), .B(men_men_n230_), .Y(men_men_n574_));
  NA3        u0552(.A(men_men_n518_), .B(men_men_n174_), .C(men_men_n27_), .Y(men_men_n575_));
  NO3        u0553(.A(men_men_n575_), .B(men_men_n574_), .C(men_men_n497_), .Y(men_men_n576_));
  NOi31      u0554(.An(men_men_n327_), .B(men_men_n440_), .C(men_men_n38_), .Y(men_men_n577_));
  OAI210     u0555(.A0(men_men_n577_), .A1(men_men_n576_), .B0(men_men_n572_), .Y(men_men_n578_));
  NO2        u0556(.A(i_8_), .B(i_7_), .Y(men_men_n579_));
  OAI210     u0557(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n580_), .B(men_men_n228_), .Y(men_men_n581_));
  AOI220     u0559(.A0(men_men_n336_), .A1(men_men_n40_), .B0(men_men_n240_), .B1(men_men_n209_), .Y(men_men_n582_));
  OAI220     u0560(.A0(men_men_n582_), .A1(men_men_n567_), .B0(men_men_n581_), .B1(men_men_n248_), .Y(men_men_n583_));
  NA2        u0561(.A(men_men_n45_), .B(i_10_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n584_), .B(i_6_), .Y(men_men_n585_));
  NA3        u0563(.A(men_men_n585_), .B(men_men_n583_), .C(men_men_n579_), .Y(men_men_n586_));
  AOI220     u0564(.A0(men_men_n453_), .A1(men_men_n336_), .B0(men_men_n253_), .B1(men_men_n250_), .Y(men_men_n587_));
  OAI220     u0565(.A0(men_men_n587_), .A1(men_men_n272_), .B0(men_men_n501_), .B1(men_men_n131_), .Y(men_men_n588_));
  NA2        u0566(.A(men_men_n588_), .B(men_men_n275_), .Y(men_men_n589_));
  NOi31      u0567(.An(men_men_n300_), .B(men_men_n311_), .C(men_men_n181_), .Y(men_men_n590_));
  NA3        u0568(.A(men_men_n317_), .B(men_men_n174_), .C(men_men_n97_), .Y(men_men_n591_));
  NO2        u0569(.A(men_men_n226_), .B(men_men_n45_), .Y(men_men_n592_));
  NO2        u0570(.A(men_men_n156_), .B(i_5_), .Y(men_men_n593_));
  NA3        u0571(.A(men_men_n593_), .B(men_men_n429_), .C(men_men_n329_), .Y(men_men_n594_));
  OAI210     u0572(.A0(men_men_n594_), .A1(men_men_n592_), .B0(men_men_n591_), .Y(men_men_n595_));
  OAI210     u0573(.A0(men_men_n595_), .A1(men_men_n590_), .B0(men_men_n491_), .Y(men_men_n596_));
  NA4        u0574(.A(men_men_n596_), .B(men_men_n589_), .C(men_men_n586_), .D(men_men_n578_), .Y(men_men_n597_));
  NA3        u0575(.A(men_men_n222_), .B(men_men_n71_), .C(men_men_n45_), .Y(men_men_n598_));
  NA2        u0576(.A(men_men_n293_), .B(men_men_n83_), .Y(men_men_n599_));
  AOI210     u0577(.A0(men_men_n598_), .A1(men_men_n363_), .B0(men_men_n599_), .Y(men_men_n600_));
  NA2        u0578(.A(men_men_n306_), .B(men_men_n296_), .Y(men_men_n601_));
  NO2        u0579(.A(men_men_n601_), .B(men_men_n173_), .Y(men_men_n602_));
  NA2        u0580(.A(men_men_n228_), .B(men_men_n227_), .Y(men_men_n603_));
  NA2        u0581(.A(men_men_n474_), .B(men_men_n226_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n603_), .B(men_men_n604_), .Y(men_men_n605_));
  AOI210     u0583(.A0(men_men_n384_), .A1(men_men_n47_), .B0(men_men_n388_), .Y(men_men_n606_));
  NA2        u0584(.A(i_0_), .B(men_men_n49_), .Y(men_men_n607_));
  NA3        u0585(.A(men_men_n573_), .B(men_men_n284_), .C(men_men_n607_), .Y(men_men_n608_));
  NO2        u0586(.A(men_men_n606_), .B(men_men_n608_), .Y(men_men_n609_));
  NO4        u0587(.A(men_men_n609_), .B(men_men_n605_), .C(men_men_n602_), .D(men_men_n600_), .Y(men_men_n610_));
  NO4        u0588(.A(men_men_n258_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n611_));
  NO3        u0589(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n612_));
  NO2        u0590(.A(men_men_n238_), .B(men_men_n36_), .Y(men_men_n613_));
  AN2        u0591(.A(men_men_n613_), .B(men_men_n612_), .Y(men_men_n614_));
  OA210      u0592(.A0(men_men_n614_), .A1(men_men_n611_), .B0(men_men_n373_), .Y(men_men_n615_));
  NO2        u0593(.A(men_men_n440_), .B(i_1_), .Y(men_men_n616_));
  NOi31      u0594(.An(men_men_n616_), .B(men_men_n483_), .C(men_men_n73_), .Y(men_men_n617_));
  AN4        u0595(.A(men_men_n617_), .B(men_men_n437_), .C(men_men_n532_), .D(i_2_), .Y(men_men_n618_));
  NO2        u0596(.A(men_men_n451_), .B(men_men_n177_), .Y(men_men_n619_));
  NO3        u0597(.A(men_men_n619_), .B(men_men_n618_), .C(men_men_n615_), .Y(men_men_n620_));
  NOi21      u0598(.An(i_10_), .B(i_6_), .Y(men_men_n621_));
  NO2        u0599(.A(men_men_n85_), .B(men_men_n25_), .Y(men_men_n622_));
  AOI220     u0600(.A0(men_men_n293_), .A1(men_men_n622_), .B0(men_men_n284_), .B1(men_men_n621_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n623_), .B(men_men_n481_), .Y(men_men_n624_));
  NO2        u0602(.A(men_men_n112_), .B(men_men_n23_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n327_), .B(men_men_n163_), .Y(men_men_n626_));
  AOI220     u0604(.A0(men_men_n626_), .A1(men_men_n462_), .B0(men_men_n184_), .B1(men_men_n182_), .Y(men_men_n627_));
  NO2        u0605(.A(men_men_n199_), .B(men_men_n37_), .Y(men_men_n628_));
  NOi31      u0606(.An(men_men_n144_), .B(men_men_n628_), .C(men_men_n344_), .Y(men_men_n629_));
  NO3        u0607(.A(men_men_n629_), .B(men_men_n627_), .C(men_men_n624_), .Y(men_men_n630_));
  NO2        u0608(.A(men_men_n556_), .B(men_men_n399_), .Y(men_men_n631_));
  INV        u0609(.A(men_men_n329_), .Y(men_men_n632_));
  NO2        u0610(.A(i_12_), .B(men_men_n85_), .Y(men_men_n633_));
  NA3        u0611(.A(men_men_n633_), .B(men_men_n284_), .C(men_men_n607_), .Y(men_men_n634_));
  NA3        u0612(.A(men_men_n407_), .B(men_men_n293_), .C(men_men_n222_), .Y(men_men_n635_));
  AOI210     u0613(.A0(men_men_n635_), .A1(men_men_n634_), .B0(men_men_n632_), .Y(men_men_n636_));
  NA2        u0614(.A(men_men_n174_), .B(i_0_), .Y(men_men_n637_));
  NO3        u0615(.A(men_men_n637_), .B(men_men_n355_), .C(men_men_n311_), .Y(men_men_n638_));
  OR2        u0616(.A(i_2_), .B(i_5_), .Y(men_men_n639_));
  OR2        u0617(.A(men_men_n639_), .B(men_men_n432_), .Y(men_men_n640_));
  AOI210     u0618(.A0(men_men_n393_), .A1(men_men_n250_), .B0(men_men_n199_), .Y(men_men_n641_));
  AOI210     u0619(.A0(men_men_n641_), .A1(men_men_n640_), .B0(men_men_n530_), .Y(men_men_n642_));
  NO4        u0620(.A(men_men_n642_), .B(men_men_n638_), .C(men_men_n636_), .D(men_men_n631_), .Y(men_men_n643_));
  NA4        u0621(.A(men_men_n643_), .B(men_men_n630_), .C(men_men_n620_), .D(men_men_n610_), .Y(men_men_n644_));
  NO4        u0622(.A(men_men_n644_), .B(men_men_n597_), .C(men_men_n570_), .D(men_men_n543_), .Y(men_men_n645_));
  NA4        u0623(.A(men_men_n645_), .B(men_men_n470_), .C(men_men_n372_), .D(men_men_n323_), .Y(men7));
  OAI220     u0624(.A0(men_men_n537_), .A1(men_men_n115_), .B0(men_men_n93_), .B1(men_men_n55_), .Y(men_men_n647_));
  NO2        u0625(.A(men_men_n107_), .B(men_men_n90_), .Y(men_men_n648_));
  NA2        u0626(.A(men_men_n405_), .B(men_men_n648_), .Y(men_men_n649_));
  NA2        u0627(.A(men_men_n518_), .B(men_men_n83_), .Y(men_men_n650_));
  NA2        u0628(.A(men_men_n142_), .B(i_8_), .Y(men_men_n651_));
  OAI210     u0629(.A0(men_men_n651_), .A1(men_men_n650_), .B0(men_men_n649_), .Y(men_men_n652_));
  NA3        u0630(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n653_));
  NO2        u0631(.A(men_men_n242_), .B(i_4_), .Y(men_men_n654_));
  NA2        u0632(.A(men_men_n654_), .B(i_8_), .Y(men_men_n655_));
  AOI210     u0633(.A0(men_men_n655_), .A1(men_men_n106_), .B0(men_men_n653_), .Y(men_men_n656_));
  NA2        u0634(.A(i_2_), .B(men_men_n85_), .Y(men_men_n657_));
  OAI210     u0635(.A0(men_men_n88_), .A1(men_men_n204_), .B0(men_men_n205_), .Y(men_men_n658_));
  NO2        u0636(.A(i_7_), .B(men_men_n37_), .Y(men_men_n659_));
  NA2        u0637(.A(i_4_), .B(i_8_), .Y(men_men_n660_));
  AOI210     u0638(.A0(men_men_n660_), .A1(men_men_n317_), .B0(men_men_n659_), .Y(men_men_n661_));
  OAI220     u0639(.A0(men_men_n661_), .A1(men_men_n657_), .B0(men_men_n658_), .B1(i_13_), .Y(men_men_n662_));
  NO4        u0640(.A(men_men_n662_), .B(men_men_n656_), .C(men_men_n652_), .D(men_men_n647_), .Y(men_men_n663_));
  AOI210     u0641(.A0(men_men_n126_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n664_));
  AOI210     u0642(.A0(men_men_n664_), .A1(men_men_n242_), .B0(men_men_n160_), .Y(men_men_n665_));
  NO2        u0643(.A(i_10_), .B(men_men_n23_), .Y(men_men_n666_));
  OR3        u0644(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n667_));
  NO3        u0645(.A(men_men_n667_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n668_));
  INV        u0646(.A(men_men_n201_), .Y(men_men_n669_));
  NO2        u0647(.A(men_men_n668_), .B(men_men_n666_), .Y(men_men_n670_));
  OA220      u0648(.A0(men_men_n670_), .A1(men_men_n632_), .B0(men_men_n665_), .B1(men_men_n277_), .Y(men_men_n671_));
  AOI210     u0649(.A0(men_men_n671_), .A1(men_men_n663_), .B0(men_men_n63_), .Y(men_men_n672_));
  NOi21      u0650(.An(i_11_), .B(i_7_), .Y(men_men_n673_));
  AO210      u0651(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(men_men_n673_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n675_), .B(men_men_n209_), .Y(men_men_n676_));
  NA3        u0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n677_));
  NAi31      u0655(.An(men_men_n677_), .B(men_men_n219_), .C(i_11_), .Y(men_men_n678_));
  AOI210     u0656(.A0(men_men_n678_), .A1(men_men_n676_), .B0(men_men_n63_), .Y(men_men_n679_));
  NA2        u0657(.A(men_men_n87_), .B(men_men_n63_), .Y(men_men_n680_));
  AO210      u0658(.A0(men_men_n680_), .A1(men_men_n399_), .B0(men_men_n41_), .Y(men_men_n681_));
  NO3        u0659(.A(men_men_n266_), .B(men_men_n211_), .C(i_8_), .Y(men_men_n682_));
  OAI210     u0660(.A0(men_men_n682_), .A1(men_men_n231_), .B0(men_men_n63_), .Y(men_men_n683_));
  NA2        u0661(.A(men_men_n433_), .B(men_men_n31_), .Y(men_men_n684_));
  OR2        u0662(.A(men_men_n211_), .B(men_men_n107_), .Y(men_men_n685_));
  INV        u0663(.A(men_men_n684_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n63_), .B(i_9_), .Y(men_men_n687_));
  INV        u0665(.A(i_4_), .Y(men_men_n688_));
  NA2        u0666(.A(men_men_n688_), .B(men_men_n686_), .Y(men_men_n689_));
  NO2        u0667(.A(i_1_), .B(i_12_), .Y(men_men_n690_));
  NA3        u0668(.A(men_men_n690_), .B(men_men_n109_), .C(men_men_n24_), .Y(men_men_n691_));
  NA4        u0669(.A(men_men_n691_), .B(men_men_n689_), .C(men_men_n683_), .D(men_men_n681_), .Y(men_men_n692_));
  OAI210     u0670(.A0(men_men_n692_), .A1(men_men_n679_), .B0(i_6_), .Y(men_men_n693_));
  OAI210     u0671(.A0(men_men_n677_), .A1(men_men_n107_), .B0(men_men_n493_), .Y(men_men_n694_));
  NA2        u0672(.A(men_men_n694_), .B(men_men_n633_), .Y(men_men_n695_));
  NA3        u0673(.A(men_men_n695_), .B(men_men_n560_), .C(men_men_n484_), .Y(men_men_n696_));
  NO4        u0674(.A(men_men_n219_), .B(men_men_n126_), .C(i_13_), .D(men_men_n85_), .Y(men_men_n697_));
  NA2        u0675(.A(men_men_n697_), .B(men_men_n687_), .Y(men_men_n698_));
  NA2        u0676(.A(men_men_n242_), .B(i_6_), .Y(men_men_n699_));
  NO3        u0677(.A(i_10_), .B(men_men_n238_), .C(men_men_n23_), .Y(men_men_n700_));
  AOI210     u0678(.A0(i_1_), .A1(men_men_n267_), .B0(men_men_n700_), .Y(men_men_n701_));
  OAI210     u0679(.A0(men_men_n701_), .A1(men_men_n45_), .B0(men_men_n698_), .Y(men_men_n702_));
  NA3        u0680(.A(men_men_n579_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n703_));
  NA3        u0681(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n704_));
  NA3        u0682(.A(men_men_n1126_), .B(men_men_n276_), .C(men_men_n45_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(men_men_n704_), .Y(men_men_n706_));
  NA3        u0684(.A(men_men_n687_), .B(men_men_n329_), .C(i_6_), .Y(men_men_n707_));
  NO2        u0685(.A(men_men_n707_), .B(men_men_n23_), .Y(men_men_n708_));
  AOI210     u0686(.A0(men_men_n509_), .A1(men_men_n444_), .B0(men_men_n247_), .Y(men_men_n709_));
  NO2        u0687(.A(men_men_n709_), .B(men_men_n657_), .Y(men_men_n710_));
  NAi21      u0688(.An(men_men_n703_), .B(men_men_n92_), .Y(men_men_n711_));
  NO2        u0689(.A(i_11_), .B(men_men_n37_), .Y(men_men_n712_));
  NA2        u0690(.A(men_men_n712_), .B(men_men_n24_), .Y(men_men_n713_));
  OAI210     u0691(.A0(men_men_n713_), .A1(i_6_), .B0(men_men_n711_), .Y(men_men_n714_));
  OR4        u0692(.A(men_men_n714_), .B(men_men_n710_), .C(men_men_n708_), .D(men_men_n706_), .Y(men_men_n715_));
  NO3        u0693(.A(men_men_n715_), .B(men_men_n702_), .C(men_men_n696_), .Y(men_men_n716_));
  NO2        u0694(.A(men_men_n242_), .B(men_men_n102_), .Y(men_men_n717_));
  NO2        u0695(.A(men_men_n717_), .B(men_men_n673_), .Y(men_men_n718_));
  NA2        u0696(.A(men_men_n718_), .B(i_1_), .Y(men_men_n719_));
  NO2        u0697(.A(men_men_n719_), .B(men_men_n667_), .Y(men_men_n720_));
  NO2        u0698(.A(men_men_n439_), .B(men_men_n85_), .Y(men_men_n721_));
  NA2        u0699(.A(men_men_n720_), .B(men_men_n47_), .Y(men_men_n722_));
  NA2        u0700(.A(i_3_), .B(men_men_n194_), .Y(men_men_n723_));
  AOI210     u0701(.A0(men_men_n265_), .A1(men_men_n723_), .B0(men_men_n112_), .Y(men_men_n724_));
  AN2        u0702(.A(men_men_n724_), .B(men_men_n585_), .Y(men_men_n725_));
  NO2        u0703(.A(men_men_n238_), .B(men_men_n45_), .Y(men_men_n726_));
  NO3        u0704(.A(men_men_n726_), .B(men_men_n320_), .C(men_men_n243_), .Y(men_men_n727_));
  NO2        u0705(.A(men_men_n115_), .B(men_men_n37_), .Y(men_men_n728_));
  NO2        u0706(.A(men_men_n728_), .B(i_6_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n85_), .B(i_9_), .Y(men_men_n730_));
  NO2        u0708(.A(men_men_n730_), .B(men_men_n63_), .Y(men_men_n731_));
  NO2        u0709(.A(men_men_n731_), .B(men_men_n690_), .Y(men_men_n732_));
  NO4        u0710(.A(men_men_n732_), .B(men_men_n729_), .C(men_men_n727_), .D(i_4_), .Y(men_men_n733_));
  NA2        u0711(.A(i_1_), .B(i_3_), .Y(men_men_n734_));
  NO2        u0712(.A(men_men_n485_), .B(men_men_n93_), .Y(men_men_n735_));
  AOI210     u0713(.A0(men_men_n726_), .A1(men_men_n621_), .B0(men_men_n735_), .Y(men_men_n736_));
  NO2        u0714(.A(men_men_n736_), .B(men_men_n734_), .Y(men_men_n737_));
  NO3        u0715(.A(men_men_n737_), .B(men_men_n733_), .C(men_men_n725_), .Y(men_men_n738_));
  NA4        u0716(.A(men_men_n738_), .B(men_men_n722_), .C(men_men_n716_), .D(men_men_n693_), .Y(men_men_n739_));
  NO3        u0717(.A(men_men_n511_), .B(i_3_), .C(i_7_), .Y(men_men_n740_));
  NOi21      u0718(.An(men_men_n740_), .B(i_10_), .Y(men_men_n741_));
  OA210      u0719(.A0(men_men_n741_), .A1(men_men_n251_), .B0(men_men_n85_), .Y(men_men_n742_));
  NA2        u0720(.A(men_men_n391_), .B(men_men_n390_), .Y(men_men_n743_));
  NA3        u0721(.A(men_men_n518_), .B(men_men_n559_), .C(men_men_n47_), .Y(men_men_n744_));
  NO3        u0722(.A(men_men_n512_), .B(men_men_n660_), .C(men_men_n85_), .Y(men_men_n745_));
  NA2        u0723(.A(men_men_n745_), .B(men_men_n25_), .Y(men_men_n746_));
  NA3        u0724(.A(men_men_n160_), .B(men_men_n83_), .C(men_men_n85_), .Y(men_men_n747_));
  NA4        u0725(.A(men_men_n747_), .B(men_men_n746_), .C(men_men_n744_), .D(men_men_n743_), .Y(men_men_n748_));
  OAI210     u0726(.A0(men_men_n748_), .A1(men_men_n742_), .B0(i_1_), .Y(men_men_n749_));
  AOI210     u0727(.A0(men_men_n707_), .A1(men_men_n749_), .B0(i_13_), .Y(men_men_n750_));
  OR2        u0728(.A(i_11_), .B(i_7_), .Y(men_men_n751_));
  NA3        u0729(.A(men_men_n751_), .B(i_3_), .C(men_men_n136_), .Y(men_men_n752_));
  AOI220     u0730(.A0(men_men_n503_), .A1(men_men_n160_), .B0(men_men_n478_), .B1(men_men_n136_), .Y(men_men_n753_));
  OAI210     u0731(.A0(men_men_n753_), .A1(men_men_n45_), .B0(men_men_n752_), .Y(men_men_n754_));
  NO2        u0732(.A(men_men_n512_), .B(men_men_n24_), .Y(men_men_n755_));
  AOI220     u0733(.A0(men_men_n755_), .A1(men_men_n721_), .B0(men_men_n251_), .B1(men_men_n129_), .Y(men_men_n756_));
  OAI220     u0734(.A0(men_men_n756_), .A1(men_men_n41_), .B0(men_men_n55_), .B1(men_men_n93_), .Y(men_men_n757_));
  AOI210     u0735(.A0(men_men_n754_), .A1(men_men_n346_), .B0(men_men_n757_), .Y(men_men_n758_));
  AOI220     u0736(.A0(i_7_), .A1(men_men_n72_), .B0(men_men_n407_), .B1(men_men_n1126_), .Y(men_men_n759_));
  NO2        u0737(.A(men_men_n759_), .B(men_men_n248_), .Y(men_men_n760_));
  AOI210     u0738(.A0(men_men_n475_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n761_));
  NOi31      u0739(.An(men_men_n761_), .B(men_men_n650_), .C(men_men_n45_), .Y(men_men_n762_));
  NA2        u0740(.A(men_men_n125_), .B(i_13_), .Y(men_men_n763_));
  NO2        u0741(.A(men_men_n704_), .B(men_men_n112_), .Y(men_men_n764_));
  INV        u0742(.A(men_men_n764_), .Y(men_men_n765_));
  OAI220     u0743(.A0(men_men_n765_), .A1(men_men_n71_), .B0(men_men_n763_), .B1(men_men_n1122_), .Y(men_men_n766_));
  NO3        u0744(.A(men_men_n71_), .B(men_men_n32_), .C(men_men_n102_), .Y(men_men_n767_));
  NA2        u0745(.A(men_men_n26_), .B(men_men_n194_), .Y(men_men_n768_));
  NA2        u0746(.A(men_men_n768_), .B(i_7_), .Y(men_men_n769_));
  NO3        u0747(.A(men_men_n512_), .B(men_men_n242_), .C(men_men_n85_), .Y(men_men_n770_));
  AOI210     u0748(.A0(men_men_n770_), .A1(men_men_n769_), .B0(men_men_n767_), .Y(men_men_n771_));
  OAI220     u0749(.A0(men_men_n1125_), .A1(men_men_n655_), .B0(men_men_n771_), .B1(men_men_n669_), .Y(men_men_n772_));
  NO4        u0750(.A(men_men_n772_), .B(men_men_n766_), .C(men_men_n762_), .D(men_men_n760_), .Y(men_men_n773_));
  OR2        u0751(.A(i_11_), .B(i_6_), .Y(men_men_n774_));
  AOI210     u0752(.A0(men_men_n242_), .A1(men_men_n765_), .B0(men_men_n774_), .Y(men_men_n775_));
  NA2        u0753(.A(men_men_n103_), .B(men_men_n768_), .Y(men_men_n776_));
  NAi21      u0754(.An(i_11_), .B(i_12_), .Y(men_men_n777_));
  NO3        u0755(.A(men_men_n777_), .B(i_13_), .C(men_men_n85_), .Y(men_men_n778_));
  NO3        u0756(.A(men_men_n512_), .B(men_men_n633_), .C(men_men_n660_), .Y(men_men_n779_));
  AOI220     u0757(.A0(men_men_n779_), .A1(men_men_n324_), .B0(men_men_n778_), .B1(men_men_n776_), .Y(men_men_n780_));
  INV        u0758(.A(men_men_n780_), .Y(men_men_n781_));
  OAI210     u0759(.A0(men_men_n781_), .A1(men_men_n775_), .B0(men_men_n63_), .Y(men_men_n782_));
  NO2        u0760(.A(i_2_), .B(i_12_), .Y(men_men_n783_));
  OAI210     u0761(.A0(men_men_n664_), .A1(men_men_n388_), .B0(men_men_n783_), .Y(men_men_n784_));
  NA2        u0762(.A(i_8_), .B(men_men_n25_), .Y(men_men_n785_));
  NO3        u0763(.A(men_men_n785_), .B(men_men_n405_), .C(men_men_n654_), .Y(men_men_n786_));
  OAI210     u0764(.A0(men_men_n786_), .A1(men_men_n390_), .B0(men_men_n388_), .Y(men_men_n787_));
  NO2        u0765(.A(men_men_n126_), .B(i_2_), .Y(men_men_n788_));
  NA2        u0766(.A(men_men_n788_), .B(men_men_n690_), .Y(men_men_n789_));
  NA3        u0767(.A(men_men_n789_), .B(men_men_n787_), .C(men_men_n784_), .Y(men_men_n790_));
  NA3        u0768(.A(men_men_n790_), .B(men_men_n46_), .C(men_men_n230_), .Y(men_men_n791_));
  NA4        u0769(.A(men_men_n791_), .B(men_men_n782_), .C(men_men_n773_), .D(men_men_n758_), .Y(men_men_n792_));
  OR4        u0770(.A(men_men_n792_), .B(men_men_n750_), .C(men_men_n739_), .D(men_men_n672_), .Y(men5));
  NA3        u0771(.A(men_men_n24_), .B(men_men_n783_), .C(men_men_n107_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n655_), .B(i_11_), .Y(men_men_n795_));
  OAI210     u0773(.A0(men_men_n659_), .A1(men_men_n88_), .B0(men_men_n795_), .Y(men_men_n796_));
  NA3        u0774(.A(men_men_n796_), .B(men_men_n794_), .C(men_men_n560_), .Y(men_men_n797_));
  NO3        u0775(.A(i_11_), .B(men_men_n242_), .C(i_13_), .Y(men_men_n798_));
  NO2        u0776(.A(men_men_n122_), .B(men_men_n23_), .Y(men_men_n799_));
  NA2        u0777(.A(i_12_), .B(i_8_), .Y(men_men_n800_));
  OAI210     u0778(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n800_), .Y(men_men_n801_));
  NA2        u0779(.A(men_men_n801_), .B(men_men_n799_), .Y(men_men_n802_));
  INV        u0780(.A(men_men_n802_), .Y(men_men_n803_));
  NO2        u0781(.A(men_men_n803_), .B(men_men_n797_), .Y(men_men_n804_));
  INV        u0782(.A(men_men_n171_), .Y(men_men_n805_));
  INV        u0783(.A(men_men_n251_), .Y(men_men_n806_));
  INV        u0784(.A(men_men_n476_), .Y(men_men_n807_));
  AOI210     u0785(.A0(men_men_n807_), .A1(men_men_n806_), .B0(men_men_n805_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n485_), .B(men_men_n26_), .Y(men_men_n809_));
  NO2        u0787(.A(men_men_n809_), .B(men_men_n444_), .Y(men_men_n810_));
  INV        u0788(.A(men_men_n808_), .Y(men_men_n811_));
  INV        u0789(.A(men_men_n172_), .Y(men_men_n812_));
  NO3        u0790(.A(men_men_n674_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n813_));
  AOI210     u0791(.A0(men_men_n812_), .A1(men_men_n88_), .B0(men_men_n813_), .Y(men_men_n814_));
  NO2        u0792(.A(men_men_n814_), .B(men_men_n194_), .Y(men_men_n815_));
  OA210      u0793(.A0(men_men_n675_), .A1(men_men_n124_), .B0(i_13_), .Y(men_men_n816_));
  NA2        u0794(.A(men_men_n201_), .B(men_men_n204_), .Y(men_men_n817_));
  NA2        u0795(.A(men_men_n150_), .B(i_8_), .Y(men_men_n818_));
  AOI210     u0796(.A0(men_men_n818_), .A1(men_men_n817_), .B0(men_men_n393_), .Y(men_men_n819_));
  AOI210     u0797(.A0(men_men_n211_), .A1(men_men_n146_), .B0(men_men_n559_), .Y(men_men_n820_));
  OAI210     u0798(.A0(men_men_n820_), .A1(men_men_n231_), .B0(men_men_n444_), .Y(men_men_n821_));
  NO2        u0799(.A(men_men_n103_), .B(men_men_n45_), .Y(men_men_n822_));
  NA4        u0800(.A(men_men_n102_), .B(men_men_n317_), .C(men_men_n122_), .D(men_men_n43_), .Y(men_men_n823_));
  OAI210     u0801(.A0(men_men_n823_), .A1(men_men_n822_), .B0(men_men_n821_), .Y(men_men_n824_));
  NO4        u0802(.A(men_men_n824_), .B(men_men_n819_), .C(men_men_n816_), .D(men_men_n815_), .Y(men_men_n825_));
  NA2        u0803(.A(men_men_n625_), .B(men_men_n28_), .Y(men_men_n826_));
  NA2        u0804(.A(men_men_n798_), .B(men_men_n285_), .Y(men_men_n827_));
  NA2        u0805(.A(men_men_n827_), .B(men_men_n826_), .Y(men_men_n828_));
  NO2        u0806(.A(men_men_n62_), .B(i_12_), .Y(men_men_n829_));
  NA2        u0807(.A(men_men_n828_), .B(men_men_n47_), .Y(men_men_n830_));
  NA4        u0808(.A(men_men_n830_), .B(men_men_n825_), .C(men_men_n811_), .D(men_men_n804_), .Y(men6));
  NO3        u0809(.A(men_men_n262_), .B(men_men_n319_), .C(i_1_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n186_), .B(men_men_n137_), .Y(men_men_n833_));
  OAI210     u0811(.A0(men_men_n833_), .A1(men_men_n832_), .B0(men_men_n788_), .Y(men_men_n834_));
  NA4        u0812(.A(men_men_n411_), .B(men_men_n517_), .C(men_men_n71_), .D(men_men_n102_), .Y(men_men_n835_));
  INV        u0813(.A(men_men_n835_), .Y(men_men_n836_));
  NO2        u0814(.A(men_men_n225_), .B(men_men_n522_), .Y(men_men_n837_));
  NO2        u0815(.A(i_11_), .B(i_9_), .Y(men_men_n838_));
  NO3        u0816(.A(men_men_n837_), .B(men_men_n836_), .C(men_men_n341_), .Y(men_men_n839_));
  AO210      u0817(.A0(men_men_n839_), .A1(men_men_n834_), .B0(i_12_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n394_), .B(men_men_n349_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n741_), .B(men_men_n71_), .Y(men_men_n842_));
  NA3        u0820(.A(men_men_n680_), .B(men_men_n842_), .C(men_men_n841_), .Y(men_men_n843_));
  INV        u0821(.A(men_men_n198_), .Y(men_men_n844_));
  AOI220     u0822(.A0(men_men_n844_), .A1(men_men_n838_), .B0(men_men_n843_), .B1(men_men_n73_), .Y(men_men_n845_));
  INV        u0823(.A(men_men_n340_), .Y(men_men_n846_));
  NA2        u0824(.A(men_men_n75_), .B(men_men_n129_), .Y(men_men_n847_));
  OAI210     u0825(.A0(men_men_n774_), .A1(i_5_), .B0(men_men_n122_), .Y(men_men_n848_));
  NA2        u0826(.A(men_men_n848_), .B(men_men_n47_), .Y(men_men_n849_));
  AOI210     u0827(.A0(men_men_n849_), .A1(men_men_n847_), .B0(men_men_n846_), .Y(men_men_n850_));
  NO3        u0828(.A(men_men_n258_), .B(men_men_n130_), .C(i_9_), .Y(men_men_n851_));
  NA2        u0829(.A(men_men_n851_), .B(men_men_n829_), .Y(men_men_n852_));
  AOI210     u0830(.A0(men_men_n852_), .A1(men_men_n557_), .B0(men_men_n186_), .Y(men_men_n853_));
  NO2        u0831(.A(men_men_n32_), .B(i_11_), .Y(men_men_n854_));
  NA3        u0832(.A(men_men_n854_), .B(men_men_n507_), .C(men_men_n411_), .Y(men_men_n855_));
  NAi32      u0833(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n856_));
  AOI210     u0834(.A0(men_men_n774_), .A1(men_men_n86_), .B0(men_men_n856_), .Y(men_men_n857_));
  OAI210     u0835(.A0(men_men_n740_), .A1(men_men_n613_), .B0(men_men_n612_), .Y(men_men_n858_));
  NAi31      u0836(.An(men_men_n857_), .B(men_men_n858_), .C(men_men_n855_), .Y(men_men_n859_));
  OR3        u0837(.A(men_men_n859_), .B(men_men_n853_), .C(men_men_n850_), .Y(men_men_n860_));
  NO2        u0838(.A(men_men_n751_), .B(i_2_), .Y(men_men_n861_));
  NA2        u0839(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n862_));
  NA2        u0840(.A(men_men_n1120_), .B(men_men_n861_), .Y(men_men_n863_));
  AO220      u0841(.A0(men_men_n377_), .A1(men_men_n367_), .B0(men_men_n419_), .B1(i_8_), .Y(men_men_n864_));
  NA3        u0842(.A(men_men_n864_), .B(men_men_n263_), .C(i_7_), .Y(men_men_n865_));
  OR2        u0843(.A(men_men_n675_), .B(men_men_n476_), .Y(men_men_n866_));
  NA3        u0844(.A(men_men_n866_), .B(men_men_n145_), .C(men_men_n69_), .Y(men_men_n867_));
  NA3        u0845(.A(men_men_n867_), .B(men_men_n865_), .C(men_men_n863_), .Y(men_men_n868_));
  AOI220     u0846(.A0(men_men_n1123_), .A1(men_men_n612_), .B0(men_men_n837_), .B1(men_men_n769_), .Y(men_men_n869_));
  NA3        u0847(.A(men_men_n393_), .B(men_men_n244_), .C(men_men_n145_), .Y(men_men_n870_));
  OAI210     u0848(.A0(men_men_n419_), .A1(men_men_n205_), .B0(men_men_n70_), .Y(men_men_n871_));
  NA4        u0849(.A(men_men_n871_), .B(men_men_n870_), .C(men_men_n869_), .D(men_men_n658_), .Y(men_men_n872_));
  AO210      u0850(.A0(men_men_n559_), .A1(men_men_n47_), .B0(men_men_n87_), .Y(men_men_n873_));
  NA3        u0851(.A(men_men_n873_), .B(men_men_n518_), .C(men_men_n222_), .Y(men_men_n874_));
  AOI210     u0852(.A0(men_men_n476_), .A1(men_men_n474_), .B0(men_men_n611_), .Y(men_men_n875_));
  NO2        u0853(.A(i_10_), .B(men_men_n103_), .Y(men_men_n876_));
  OAI210     u0854(.A0(men_men_n876_), .A1(men_men_n110_), .B0(men_men_n431_), .Y(men_men_n877_));
  NA2        u0855(.A(men_men_n250_), .B(men_men_n47_), .Y(men_men_n878_));
  NA2        u0856(.A(men_men_n878_), .B(men_men_n640_), .Y(men_men_n879_));
  NA3        u0857(.A(men_men_n879_), .B(men_men_n340_), .C(i_7_), .Y(men_men_n880_));
  NA4        u0858(.A(men_men_n880_), .B(men_men_n877_), .C(men_men_n875_), .D(men_men_n874_), .Y(men_men_n881_));
  NO4        u0859(.A(men_men_n881_), .B(men_men_n872_), .C(men_men_n868_), .D(men_men_n860_), .Y(men_men_n882_));
  NA4        u0860(.A(men_men_n882_), .B(men_men_n845_), .C(men_men_n840_), .D(men_men_n401_), .Y(men3));
  NA2        u0861(.A(i_12_), .B(i_10_), .Y(men_men_n884_));
  NA2        u0862(.A(i_6_), .B(i_7_), .Y(men_men_n885_));
  NO2        u0863(.A(men_men_n885_), .B(i_0_), .Y(men_men_n886_));
  NO2        u0864(.A(i_11_), .B(men_men_n242_), .Y(men_men_n887_));
  OAI210     u0865(.A0(men_men_n886_), .A1(men_men_n300_), .B0(men_men_n887_), .Y(men_men_n888_));
  NO2        u0866(.A(men_men_n888_), .B(men_men_n194_), .Y(men_men_n889_));
  NO3        u0867(.A(men_men_n481_), .B(men_men_n90_), .C(men_men_n45_), .Y(men_men_n890_));
  OA210      u0868(.A0(men_men_n890_), .A1(men_men_n889_), .B0(men_men_n174_), .Y(men_men_n891_));
  NA3        u0869(.A(men_men_n870_), .B(men_men_n658_), .C(men_men_n392_), .Y(men_men_n892_));
  NA2        u0870(.A(men_men_n892_), .B(men_men_n40_), .Y(men_men_n893_));
  NOi21      u0871(.An(men_men_n97_), .B(men_men_n810_), .Y(men_men_n894_));
  NO3        u0872(.A(men_men_n685_), .B(men_men_n485_), .C(men_men_n129_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n433_), .B(men_men_n46_), .Y(men_men_n896_));
  AN2        u0874(.A(men_men_n483_), .B(men_men_n56_), .Y(men_men_n897_));
  NO3        u0875(.A(men_men_n897_), .B(men_men_n895_), .C(men_men_n894_), .Y(men_men_n898_));
  AOI210     u0876(.A0(men_men_n898_), .A1(men_men_n893_), .B0(men_men_n49_), .Y(men_men_n899_));
  NA2        u0877(.A(men_men_n186_), .B(men_men_n621_), .Y(men_men_n900_));
  NA2        u0878(.A(men_men_n761_), .B(men_men_n730_), .Y(men_men_n901_));
  NA2        u0879(.A(men_men_n347_), .B(men_men_n464_), .Y(men_men_n902_));
  OAI220     u0880(.A0(men_men_n902_), .A1(men_men_n901_), .B0(men_men_n900_), .B1(men_men_n63_), .Y(men_men_n903_));
  NOi21      u0881(.An(i_5_), .B(i_9_), .Y(men_men_n904_));
  NA2        u0882(.A(men_men_n904_), .B(men_men_n472_), .Y(men_men_n905_));
  AOI210     u0883(.A0(men_men_n276_), .A1(men_men_n509_), .B0(men_men_n745_), .Y(men_men_n906_));
  NO3        u0884(.A(men_men_n436_), .B(men_men_n276_), .C(men_men_n73_), .Y(men_men_n907_));
  NO2        u0885(.A(men_men_n175_), .B(men_men_n146_), .Y(men_men_n908_));
  AOI210     u0886(.A0(men_men_n908_), .A1(men_men_n250_), .B0(men_men_n907_), .Y(men_men_n909_));
  OAI220     u0887(.A0(men_men_n909_), .A1(men_men_n181_), .B0(men_men_n906_), .B1(men_men_n905_), .Y(men_men_n910_));
  NO4        u0888(.A(men_men_n910_), .B(men_men_n903_), .C(men_men_n899_), .D(men_men_n891_), .Y(men_men_n911_));
  NOi21      u0889(.An(i_0_), .B(i_10_), .Y(men_men_n912_));
  NA2        u0890(.A(men_men_n186_), .B(men_men_n24_), .Y(men_men_n913_));
  NO2        u0891(.A(men_men_n728_), .B(men_men_n648_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n914_), .B(men_men_n913_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n324_), .B(men_men_n127_), .Y(men_men_n916_));
  NAi21      u0894(.An(men_men_n161_), .B(men_men_n464_), .Y(men_men_n917_));
  OAI220     u0895(.A0(men_men_n917_), .A1(men_men_n878_), .B0(men_men_n916_), .B1(men_men_n422_), .Y(men_men_n918_));
  NO2        u0896(.A(men_men_n918_), .B(men_men_n915_), .Y(men_men_n919_));
  NO2        u0897(.A(men_men_n411_), .B(men_men_n304_), .Y(men_men_n920_));
  NA2        u0898(.A(men_men_n920_), .B(men_men_n764_), .Y(men_men_n921_));
  NA2        u0899(.A(men_men_n622_), .B(i_0_), .Y(men_men_n922_));
  NO3        u0900(.A(men_men_n922_), .B(men_men_n406_), .C(men_men_n88_), .Y(men_men_n923_));
  NO4        u0901(.A(men_men_n639_), .B(men_men_n219_), .C(men_men_n440_), .D(men_men_n432_), .Y(men_men_n924_));
  AOI210     u0902(.A0(men_men_n924_), .A1(i_11_), .B0(men_men_n923_), .Y(men_men_n925_));
  INV        u0903(.A(men_men_n507_), .Y(men_men_n926_));
  AN2        u0904(.A(men_men_n97_), .B(men_men_n249_), .Y(men_men_n927_));
  NA2        u0905(.A(men_men_n798_), .B(men_men_n341_), .Y(men_men_n928_));
  AOI210     u0906(.A0(men_men_n518_), .A1(men_men_n88_), .B0(men_men_n59_), .Y(men_men_n929_));
  OAI220     u0907(.A0(men_men_n929_), .A1(men_men_n928_), .B0(men_men_n713_), .B1(men_men_n581_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n260_), .B(men_men_n152_), .Y(men_men_n931_));
  NA2        u0909(.A(i_0_), .B(i_10_), .Y(men_men_n932_));
  OAI210     u0910(.A0(men_men_n932_), .A1(men_men_n85_), .B0(men_men_n584_), .Y(men_men_n933_));
  NO4        u0911(.A(men_men_n112_), .B(men_men_n59_), .C(men_men_n723_), .D(i_5_), .Y(men_men_n934_));
  AO220      u0912(.A0(men_men_n934_), .A1(men_men_n933_), .B0(men_men_n931_), .B1(i_6_), .Y(men_men_n935_));
  AOI220     u0913(.A0(men_men_n347_), .A1(men_men_n99_), .B0(men_men_n186_), .B1(men_men_n83_), .Y(men_men_n936_));
  NA2        u0914(.A(men_men_n616_), .B(i_4_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n189_), .B(men_men_n204_), .Y(men_men_n938_));
  OAI220     u0916(.A0(men_men_n938_), .A1(men_men_n928_), .B0(men_men_n937_), .B1(men_men_n936_), .Y(men_men_n939_));
  NO4        u0917(.A(men_men_n939_), .B(men_men_n935_), .C(men_men_n930_), .D(men_men_n927_), .Y(men_men_n940_));
  NA4        u0918(.A(men_men_n940_), .B(men_men_n925_), .C(men_men_n921_), .D(men_men_n919_), .Y(men_men_n941_));
  NA2        u0919(.A(i_11_), .B(i_9_), .Y(men_men_n942_));
  NO3        u0920(.A(i_12_), .B(men_men_n942_), .C(men_men_n657_), .Y(men_men_n943_));
  AO220      u0921(.A0(men_men_n943_), .A1(i_10_), .B0(men_men_n278_), .B1(men_men_n87_), .Y(men_men_n944_));
  NO2        u0922(.A(men_men_n49_), .B(i_7_), .Y(men_men_n945_));
  NAi31      u0923(.An(men_men_n273_), .B(men_men_n490_), .C(men_men_n159_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n942_), .B(men_men_n73_), .Y(men_men_n947_));
  NO2        u0925(.A(men_men_n175_), .B(i_0_), .Y(men_men_n948_));
  INV        u0926(.A(men_men_n948_), .Y(men_men_n949_));
  NA2        u0927(.A(men_men_n507_), .B(men_men_n236_), .Y(men_men_n950_));
  AOI210     u0928(.A0(men_men_n391_), .A1(men_men_n42_), .B0(men_men_n430_), .Y(men_men_n951_));
  OAI220     u0929(.A0(men_men_n951_), .A1(men_men_n905_), .B0(men_men_n950_), .B1(men_men_n949_), .Y(men_men_n952_));
  NO3        u0930(.A(men_men_n952_), .B(men_men_n946_), .C(men_men_n944_), .Y(men_men_n953_));
  NA2        u0931(.A(men_men_n712_), .B(men_men_n119_), .Y(men_men_n954_));
  NO2        u0932(.A(i_6_), .B(men_men_n954_), .Y(men_men_n955_));
  AOI210     u0933(.A0(men_men_n475_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n956_));
  NA2        u0934(.A(men_men_n171_), .B(men_men_n104_), .Y(men_men_n957_));
  NOi32      u0935(.An(men_men_n956_), .Bn(men_men_n189_), .C(men_men_n957_), .Y(men_men_n958_));
  AOI210     u0936(.A0(men_men_n659_), .A1(men_men_n341_), .B0(men_men_n249_), .Y(men_men_n959_));
  NO2        u0937(.A(men_men_n959_), .B(men_men_n896_), .Y(men_men_n960_));
  NO3        u0938(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n955_), .Y(men_men_n961_));
  NOi21      u0939(.An(i_7_), .B(i_5_), .Y(men_men_n962_));
  NOi31      u0940(.An(men_men_n962_), .B(men_men_n912_), .C(men_men_n777_), .Y(men_men_n963_));
  NA3        u0941(.A(men_men_n963_), .B(men_men_n405_), .C(i_6_), .Y(men_men_n964_));
  OA210      u0942(.A0(men_men_n957_), .A1(men_men_n557_), .B0(men_men_n964_), .Y(men_men_n965_));
  NO3        u0943(.A(men_men_n425_), .B(men_men_n380_), .C(men_men_n376_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n270_), .B(men_men_n330_), .Y(men_men_n967_));
  NO2        u0945(.A(men_men_n777_), .B(men_men_n265_), .Y(men_men_n968_));
  AOI210     u0946(.A0(men_men_n968_), .A1(men_men_n967_), .B0(men_men_n966_), .Y(men_men_n969_));
  NA4        u0947(.A(men_men_n969_), .B(men_men_n965_), .C(men_men_n961_), .D(men_men_n953_), .Y(men_men_n970_));
  NO2        u0948(.A(men_men_n913_), .B(men_men_n245_), .Y(men_men_n971_));
  AN2        u0949(.A(men_men_n346_), .B(men_men_n341_), .Y(men_men_n972_));
  AO220      u0950(.A0(men_men_n972_), .A1(men_men_n908_), .B0(men_men_n362_), .B1(men_men_n27_), .Y(men_men_n973_));
  OAI210     u0951(.A0(men_men_n973_), .A1(men_men_n971_), .B0(i_10_), .Y(men_men_n974_));
  NO2        u0952(.A(men_men_n884_), .B(men_men_n329_), .Y(men_men_n975_));
  OA210      u0953(.A0(men_men_n507_), .A1(men_men_n228_), .B0(men_men_n506_), .Y(men_men_n976_));
  OAI210     u0954(.A0(men_men_n976_), .A1(men_men_n975_), .B0(men_men_n947_), .Y(men_men_n977_));
  NA3        u0955(.A(men_men_n506_), .B(men_men_n433_), .C(men_men_n46_), .Y(men_men_n978_));
  OAI210     u0956(.A0(men_men_n917_), .A1(men_men_n926_), .B0(men_men_n978_), .Y(men_men_n979_));
  NO2        u0957(.A(men_men_n263_), .B(men_men_n47_), .Y(men_men_n980_));
  NA2        u0958(.A(men_men_n947_), .B(men_men_n317_), .Y(men_men_n981_));
  OAI210     u0959(.A0(men_men_n980_), .A1(men_men_n188_), .B0(men_men_n981_), .Y(men_men_n982_));
  AOI220     u0960(.A0(men_men_n982_), .A1(men_men_n507_), .B0(men_men_n979_), .B1(men_men_n73_), .Y(men_men_n983_));
  NA3        u0961(.A(men_men_n862_), .B(men_men_n403_), .C(i_12_), .Y(men_men_n984_));
  NA2        u0962(.A(men_men_n93_), .B(men_men_n45_), .Y(men_men_n985_));
  NO2        u0963(.A(men_men_n75_), .B(men_men_n800_), .Y(men_men_n986_));
  AOI220     u0964(.A0(men_men_n986_), .A1(men_men_n985_), .B0(men_men_n174_), .B1(men_men_n648_), .Y(men_men_n987_));
  AOI210     u0965(.A0(men_men_n987_), .A1(men_men_n984_), .B0(men_men_n48_), .Y(men_men_n988_));
  NO3        u0966(.A(men_men_n639_), .B(men_men_n375_), .C(men_men_n24_), .Y(men_men_n989_));
  AOI210     u0967(.A0(men_men_n755_), .A1(men_men_n593_), .B0(men_men_n989_), .Y(men_men_n990_));
  NAi21      u0968(.An(i_9_), .B(i_5_), .Y(men_men_n991_));
  NO2        u0969(.A(men_men_n991_), .B(men_men_n425_), .Y(men_men_n992_));
  NO2        u0970(.A(men_men_n653_), .B(men_men_n106_), .Y(men_men_n993_));
  AOI220     u0971(.A0(men_men_n993_), .A1(i_0_), .B0(men_men_n992_), .B1(men_men_n675_), .Y(men_men_n994_));
  OAI220     u0972(.A0(men_men_n994_), .A1(men_men_n85_), .B0(men_men_n990_), .B1(men_men_n172_), .Y(men_men_n995_));
  NO3        u0973(.A(men_men_n995_), .B(men_men_n988_), .C(men_men_n561_), .Y(men_men_n996_));
  NA4        u0974(.A(men_men_n996_), .B(men_men_n983_), .C(men_men_n977_), .D(men_men_n974_), .Y(men_men_n997_));
  NO3        u0975(.A(men_men_n997_), .B(men_men_n970_), .C(men_men_n941_), .Y(men_men_n998_));
  NO2        u0976(.A(men_men_n912_), .B(men_men_n777_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n73_), .B(men_men_n45_), .Y(men_men_n1000_));
  NO3        u0978(.A(men_men_n106_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n1001_));
  AO220      u0979(.A0(men_men_n1001_), .A1(men_men_n73_), .B0(men_men_n999_), .B1(men_men_n174_), .Y(men_men_n1002_));
  NO2        u0980(.A(men_men_n743_), .B(men_men_n957_), .Y(men_men_n1003_));
  AOI210     u0981(.A0(men_men_n1002_), .A1(men_men_n364_), .B0(men_men_n1003_), .Y(men_men_n1004_));
  NA2        u0982(.A(men_men_n788_), .B(men_men_n144_), .Y(men_men_n1005_));
  INV        u0983(.A(men_men_n1005_), .Y(men_men_n1006_));
  NA3        u0984(.A(men_men_n1006_), .B(men_men_n730_), .C(men_men_n73_), .Y(men_men_n1007_));
  NO2        u0985(.A(men_men_n858_), .B(men_men_n425_), .Y(men_men_n1008_));
  NA3        u0986(.A(men_men_n886_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n1009_));
  NA2        u0987(.A(men_men_n887_), .B(i_9_), .Y(men_men_n1010_));
  AOI210     u0988(.A0(men_men_n1009_), .A1(men_men_n534_), .B0(men_men_n1010_), .Y(men_men_n1011_));
  OAI210     u0989(.A0(men_men_n250_), .A1(i_9_), .B0(men_men_n235_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n1012_), .A1(men_men_n922_), .B0(men_men_n152_), .Y(men_men_n1013_));
  NO3        u0991(.A(men_men_n1013_), .B(men_men_n1011_), .C(men_men_n1008_), .Y(men_men_n1014_));
  NA3        u0992(.A(men_men_n1014_), .B(men_men_n1007_), .C(men_men_n1004_), .Y(men_men_n1015_));
  NA2        u0993(.A(men_men_n972_), .B(men_men_n393_), .Y(men_men_n1016_));
  AOI210     u0994(.A0(men_men_n311_), .A1(men_men_n161_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  NA3        u0995(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n1018_));
  NA2        u0996(.A(men_men_n945_), .B(men_men_n523_), .Y(men_men_n1019_));
  AOI210     u0997(.A0(men_men_n1018_), .A1(men_men_n161_), .B0(men_men_n1019_), .Y(men_men_n1020_));
  NO2        u0998(.A(men_men_n1020_), .B(men_men_n1017_), .Y(men_men_n1021_));
  NO3        u0999(.A(men_men_n932_), .B(men_men_n904_), .C(men_men_n191_), .Y(men_men_n1022_));
  AOI220     u1000(.A0(men_men_n1022_), .A1(i_11_), .B0(men_men_n617_), .B1(men_men_n75_), .Y(men_men_n1023_));
  NO3        u1001(.A(men_men_n213_), .B(men_men_n404_), .C(i_0_), .Y(men_men_n1024_));
  OAI210     u1002(.A0(men_men_n1024_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n1025_));
  INV        u1003(.A(men_men_n222_), .Y(men_men_n1026_));
  OAI220     u1004(.A0(men_men_n574_), .A1(men_men_n137_), .B0(men_men_n699_), .B1(men_men_n669_), .Y(men_men_n1027_));
  NA3        u1005(.A(men_men_n1027_), .B(men_men_n420_), .C(men_men_n1026_), .Y(men_men_n1028_));
  NA4        u1006(.A(men_men_n1028_), .B(men_men_n1025_), .C(men_men_n1023_), .D(men_men_n1021_), .Y(men_men_n1029_));
  NO2        u1007(.A(men_men_n248_), .B(men_men_n93_), .Y(men_men_n1030_));
  AOI210     u1008(.A0(men_men_n1030_), .A1(men_men_n999_), .B0(men_men_n108_), .Y(men_men_n1031_));
  AOI220     u1009(.A0(men_men_n962_), .A1(men_men_n523_), .B0(men_men_n886_), .B1(men_men_n162_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n367_), .B(men_men_n176_), .Y(men_men_n1033_));
  OA220      u1011(.A0(men_men_n1033_), .A1(men_men_n1032_), .B0(men_men_n1031_), .B1(i_5_), .Y(men_men_n1034_));
  AOI210     u1012(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n175_), .Y(men_men_n1035_));
  NA2        u1013(.A(men_men_n1035_), .B(men_men_n976_), .Y(men_men_n1036_));
  NA3        u1014(.A(men_men_n666_), .B(men_men_n186_), .C(men_men_n83_), .Y(men_men_n1037_));
  NA2        u1015(.A(men_men_n1037_), .B(men_men_n591_), .Y(men_men_n1038_));
  NO3        u1016(.A(men_men_n896_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n1039_));
  NA2        u1017(.A(men_men_n521_), .B(men_men_n504_), .Y(men_men_n1040_));
  NO3        u1018(.A(men_men_n1040_), .B(men_men_n1039_), .C(men_men_n1038_), .Y(men_men_n1041_));
  NA3        u1019(.A(men_men_n945_), .B(men_men_n300_), .C(men_men_n235_), .Y(men_men_n1042_));
  INV        u1020(.A(men_men_n1042_), .Y(men_men_n1043_));
  NA3        u1021(.A(men_men_n411_), .B(men_men_n348_), .C(men_men_n226_), .Y(men_men_n1044_));
  OAI210     u1022(.A0(men_men_n900_), .A1(men_men_n703_), .B0(men_men_n1044_), .Y(men_men_n1045_));
  NOi31      u1023(.An(men_men_n410_), .B(men_men_n1000_), .C(men_men_n245_), .Y(men_men_n1046_));
  NO3        u1024(.A(men_men_n942_), .B(men_men_n222_), .C(men_men_n191_), .Y(men_men_n1047_));
  NO4        u1025(.A(men_men_n1047_), .B(men_men_n1046_), .C(men_men_n1045_), .D(men_men_n1043_), .Y(men_men_n1048_));
  NA4        u1026(.A(men_men_n1048_), .B(men_men_n1041_), .C(men_men_n1036_), .D(men_men_n1034_), .Y(men_men_n1049_));
  AOI210     u1027(.A0(men_men_n616_), .A1(men_men_n573_), .B0(men_men_n668_), .Y(men_men_n1050_));
  NO3        u1028(.A(men_men_n1050_), .B(men_men_n607_), .C(men_men_n361_), .Y(men_men_n1051_));
  NA3        u1029(.A(men_men_n887_), .B(men_men_n109_), .C(men_men_n122_), .Y(men_men_n1052_));
  INV        u1030(.A(men_men_n1052_), .Y(men_men_n1053_));
  AOI210     u1031(.A0(men_men_n1053_), .A1(men_men_n1124_), .B0(men_men_n1051_), .Y(men_men_n1054_));
  NA3        u1032(.A(men_men_n317_), .B(i_5_), .C(men_men_n194_), .Y(men_men_n1055_));
  NAi31      u1033(.An(men_men_n247_), .B(men_men_n1055_), .C(men_men_n248_), .Y(men_men_n1056_));
  NO4        u1034(.A(men_men_n245_), .B(men_men_n213_), .C(i_0_), .D(i_12_), .Y(men_men_n1057_));
  AOI220     u1035(.A0(men_men_n1057_), .A1(men_men_n1056_), .B0(men_men_n836_), .B1(men_men_n176_), .Y(men_men_n1058_));
  AN2        u1036(.A(men_men_n932_), .B(men_men_n152_), .Y(men_men_n1059_));
  NO4        u1037(.A(men_men_n1059_), .B(i_12_), .C(men_men_n703_), .D(men_men_n129_), .Y(men_men_n1060_));
  NA2        u1038(.A(men_men_n1060_), .B(men_men_n222_), .Y(men_men_n1061_));
  NA3        u1039(.A(men_men_n99_), .B(men_men_n621_), .C(i_11_), .Y(men_men_n1062_));
  NO2        u1040(.A(men_men_n1062_), .B(men_men_n154_), .Y(men_men_n1063_));
  NA2        u1041(.A(men_men_n962_), .B(men_men_n503_), .Y(men_men_n1064_));
  OAI220     u1042(.A0(i_7_), .A1(men_men_n1055_), .B0(men_men_n1064_), .B1(men_men_n731_), .Y(men_men_n1065_));
  AOI210     u1043(.A0(men_men_n1065_), .A1(men_men_n948_), .B0(men_men_n1063_), .Y(men_men_n1066_));
  NA4        u1044(.A(men_men_n1066_), .B(men_men_n1061_), .C(men_men_n1058_), .D(men_men_n1054_), .Y(men_men_n1067_));
  NO4        u1045(.A(men_men_n1067_), .B(men_men_n1049_), .C(men_men_n1029_), .D(men_men_n1015_), .Y(men_men_n1068_));
  OAI210     u1046(.A0(men_men_n861_), .A1(men_men_n854_), .B0(men_men_n37_), .Y(men_men_n1069_));
  NA3        u1047(.A(men_men_n956_), .B(men_men_n388_), .C(i_5_), .Y(men_men_n1070_));
  NA3        u1048(.A(men_men_n1070_), .B(men_men_n1069_), .C(men_men_n665_), .Y(men_men_n1071_));
  NA2        u1049(.A(men_men_n1071_), .B(men_men_n209_), .Y(men_men_n1072_));
  AN2        u1050(.A(men_men_n751_), .B(men_men_n389_), .Y(men_men_n1073_));
  NA2        u1051(.A(men_men_n187_), .B(men_men_n189_), .Y(men_men_n1074_));
  AO210      u1052(.A0(men_men_n1073_), .A1(men_men_n33_), .B0(men_men_n1074_), .Y(men_men_n1075_));
  OAI210     u1053(.A0(men_men_n668_), .A1(men_men_n666_), .B0(men_men_n329_), .Y(men_men_n1076_));
  NAi31      u1054(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1077_));
  AOI210     u1055(.A0(men_men_n115_), .A1(men_men_n70_), .B0(men_men_n1077_), .Y(men_men_n1078_));
  NO2        u1056(.A(men_men_n1078_), .B(men_men_n700_), .Y(men_men_n1079_));
  NA3        u1057(.A(men_men_n1079_), .B(men_men_n1076_), .C(men_men_n1075_), .Y(men_men_n1080_));
  NO2        u1058(.A(men_men_n493_), .B(men_men_n276_), .Y(men_men_n1081_));
  NO4        u1059(.A(men_men_n238_), .B(men_men_n143_), .C(men_men_n734_), .D(men_men_n37_), .Y(men_men_n1082_));
  NO3        u1060(.A(men_men_n1082_), .B(men_men_n1081_), .C(men_men_n924_), .Y(men_men_n1083_));
  OAI210     u1061(.A0(men_men_n1062_), .A1(men_men_n146_), .B0(men_men_n1083_), .Y(men_men_n1084_));
  AOI210     u1062(.A0(men_men_n1080_), .A1(men_men_n49_), .B0(men_men_n1084_), .Y(men_men_n1085_));
  AOI210     u1063(.A0(men_men_n1085_), .A1(men_men_n1072_), .B0(men_men_n73_), .Y(men_men_n1086_));
  NO2        u1064(.A(men_men_n614_), .B(men_men_n400_), .Y(men_men_n1087_));
  NO2        u1065(.A(men_men_n1087_), .B(men_men_n805_), .Y(men_men_n1088_));
  OAI210     u1066(.A0(men_men_n80_), .A1(men_men_n55_), .B0(men_men_n107_), .Y(men_men_n1089_));
  NA2        u1067(.A(men_men_n1089_), .B(men_men_n76_), .Y(men_men_n1090_));
  AOI210     u1068(.A0(men_men_n1035_), .A1(men_men_n945_), .B0(men_men_n963_), .Y(men_men_n1091_));
  AOI210     u1069(.A0(men_men_n1091_), .A1(men_men_n1090_), .B0(men_men_n734_), .Y(men_men_n1092_));
  NA2        u1070(.A(men_men_n270_), .B(men_men_n58_), .Y(men_men_n1093_));
  AOI220     u1071(.A0(men_men_n1093_), .A1(men_men_n76_), .B0(men_men_n362_), .B1(men_men_n262_), .Y(men_men_n1094_));
  NO2        u1072(.A(men_men_n1094_), .B(men_men_n242_), .Y(men_men_n1095_));
  NA3        u1073(.A(men_men_n97_), .B(men_men_n319_), .C(men_men_n31_), .Y(men_men_n1096_));
  INV        u1074(.A(men_men_n1096_), .Y(men_men_n1097_));
  NO3        u1075(.A(men_men_n1097_), .B(men_men_n1095_), .C(men_men_n1092_), .Y(men_men_n1098_));
  OAI210     u1076(.A0(men_men_n278_), .A1(men_men_n157_), .B0(men_men_n88_), .Y(men_men_n1099_));
  NA3        u1077(.A(men_men_n809_), .B(men_men_n300_), .C(men_men_n80_), .Y(men_men_n1100_));
  AOI210     u1078(.A0(men_men_n1100_), .A1(men_men_n1099_), .B0(i_11_), .Y(men_men_n1101_));
  NA2        u1079(.A(men_men_n660_), .B(men_men_n219_), .Y(men_men_n1102_));
  OAI210     u1080(.A0(men_men_n1102_), .A1(men_men_n956_), .B0(men_men_n209_), .Y(men_men_n1103_));
  NA2        u1081(.A(men_men_n163_), .B(i_5_), .Y(men_men_n1104_));
  AOI210     u1082(.A0(men_men_n1103_), .A1(men_men_n817_), .B0(men_men_n1104_), .Y(men_men_n1105_));
  NO3        u1083(.A(men_men_n60_), .B(men_men_n59_), .C(i_4_), .Y(men_men_n1106_));
  OAI210     u1084(.A0(men_men_n967_), .A1(men_men_n319_), .B0(men_men_n1106_), .Y(men_men_n1107_));
  NO2        u1085(.A(men_men_n1107_), .B(men_men_n777_), .Y(men_men_n1108_));
  NO4        u1086(.A(men_men_n991_), .B(men_men_n511_), .C(men_men_n259_), .D(men_men_n258_), .Y(men_men_n1109_));
  NO2        u1087(.A(men_men_n1109_), .B(men_men_n611_), .Y(men_men_n1110_));
  NO2        u1088(.A(men_men_n857_), .B(men_men_n381_), .Y(men_men_n1111_));
  AOI210     u1089(.A0(men_men_n1111_), .A1(men_men_n1110_), .B0(men_men_n41_), .Y(men_men_n1112_));
  NO4        u1090(.A(men_men_n1112_), .B(men_men_n1108_), .C(men_men_n1105_), .D(men_men_n1101_), .Y(men_men_n1113_));
  OAI210     u1091(.A0(men_men_n1098_), .A1(i_4_), .B0(men_men_n1113_), .Y(men_men_n1114_));
  NO3        u1092(.A(men_men_n1114_), .B(men_men_n1088_), .C(men_men_n1086_), .Y(men_men_n1115_));
  NA4        u1093(.A(men_men_n1115_), .B(men_men_n1068_), .C(men_men_n998_), .D(men_men_n911_), .Y(men4));
  INV        u1094(.A(i_5_), .Y(men_men_n1119_));
  INV        u1095(.A(men_men_n862_), .Y(men_men_n1120_));
  INV        u1096(.A(men_men_n199_), .Y(men_men_n1121_));
  INV        u1097(.A(i_1_), .Y(men_men_n1122_));
  INV        u1098(.A(men_men_n86_), .Y(men_men_n1123_));
  INV        u1099(.A(i_5_), .Y(men_men_n1124_));
  INV        u1100(.A(men_men_n407_), .Y(men_men_n1125_));
  INV        u1101(.A(i_1_), .Y(men_men_n1126_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule