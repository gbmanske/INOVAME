// Benchmark "top" written by ABC on Fri Jun 21 17:49:26 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n133_, new_new_n134_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1015_,
    new_new_n1016_, new_new_n1017_, new_new_n1018_, new_new_n1019_,
    new_new_n1020_, new_new_n1021_, new_new_n1022_, new_new_n1023_,
    new_new_n1024_, new_new_n1025_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi21      g0043(.An(new_new_n65_), .B(new_new_n61_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n51_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  INV        g0053(.A(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(new_new_n79_), .B(new_new_n58_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  INV        g0060(.A(i_6_), .Y(new_new_n83_));
  OR4        g0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  NO2        g0062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  NAi21      g0063(.An(i_6_), .B(i_10_), .Y(new_new_n86_));
  NA2        g0064(.A(i_6_), .B(i_9_), .Y(new_new_n87_));
  NA2        g0065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  NO2        g0066(.A(new_new_n1019_), .B(new_new_n78_), .Y(new_new_n89_));
  AN3        g0067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  NO2        g0069(.A(i_5_), .B(i_8_), .Y(new_new_n92_));
  NOi21      g0070(.An(new_new_n92_), .B(new_new_n91_), .Y(new_new_n93_));
  AOI220     g0071(.A0(new_new_n93_), .A1(new_new_n62_), .B0(new_new_n90_), .B1(new_new_n32_), .Y(new_new_n94_));
  INV        g0072(.A(i_7_), .Y(new_new_n95_));
  NA2        g0073(.A(new_new_n47_), .B(new_new_n95_), .Y(new_new_n96_));
  NO2        g0074(.A(i_0_), .B(i_5_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n83_), .Y(new_new_n98_));
  NA2        g0076(.A(i_12_), .B(i_3_), .Y(new_new_n99_));
  INV        g0077(.A(new_new_n99_), .Y(new_new_n100_));
  NA3        g0078(.A(new_new_n100_), .B(new_new_n98_), .C(new_new_n96_), .Y(new_new_n101_));
  NAi21      g0079(.An(i_7_), .B(i_11_), .Y(new_new_n102_));
  AN2        g0080(.A(i_2_), .B(i_10_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(i_7_), .Y(new_new_n104_));
  OR2        g0082(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n105_));
  NO2        g0083(.A(i_8_), .B(new_new_n95_), .Y(new_new_n106_));
  NO3        g0084(.A(new_new_n106_), .B(new_new_n105_), .C(new_new_n104_), .Y(new_new_n107_));
  NA2        g0085(.A(i_12_), .B(i_7_), .Y(new_new_n108_));
  NO2        g0086(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n109_));
  NA2        g0087(.A(new_new_n109_), .B(i_0_), .Y(new_new_n110_));
  NA2        g0088(.A(i_11_), .B(i_12_), .Y(new_new_n111_));
  OAI210     g0089(.A0(new_new_n110_), .A1(new_new_n108_), .B0(new_new_n111_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n112_), .B(new_new_n107_), .Y(new_new_n113_));
  NA3        g0091(.A(new_new_n113_), .B(new_new_n101_), .C(new_new_n94_), .Y(new_new_n114_));
  NOi21      g0092(.An(i_1_), .B(i_5_), .Y(new_new_n115_));
  NA2        g0093(.A(new_new_n115_), .B(i_11_), .Y(new_new_n116_));
  NA2        g0094(.A(new_new_n95_), .B(new_new_n37_), .Y(new_new_n117_));
  NA2        g0095(.A(i_7_), .B(new_new_n25_), .Y(new_new_n118_));
  NA2        g0096(.A(new_new_n118_), .B(new_new_n117_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n119_), .B(new_new_n47_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n87_), .B(new_new_n86_), .Y(new_new_n121_));
  NAi21      g0099(.An(i_3_), .B(i_8_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(new_new_n62_), .Y(new_new_n123_));
  NOi21      g0101(.An(new_new_n123_), .B(new_new_n121_), .Y(new_new_n124_));
  NO2        g0102(.A(i_1_), .B(new_new_n83_), .Y(new_new_n125_));
  NO2        g0103(.A(i_6_), .B(i_5_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(i_3_), .Y(new_new_n127_));
  AO210      g0105(.A0(new_new_n127_), .A1(new_new_n48_), .B0(new_new_n125_), .Y(new_new_n128_));
  OAI220     g0106(.A0(new_new_n128_), .A1(new_new_n102_), .B0(new_new_n124_), .B1(new_new_n116_), .Y(new_new_n129_));
  NO3        g0107(.A(new_new_n129_), .B(new_new_n114_), .C(new_new_n89_), .Y(new_new_n130_));
  NA3        g0108(.A(new_new_n130_), .B(new_new_n77_), .C(new_new_n56_), .Y(men2));
  NO2        g0109(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n132_));
  INV        g0110(.A(i_6_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(new_new_n132_), .Y(new_new_n134_));
  NA4        g0112(.A(new_new_n134_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(men0));
  AN2        g0113(.A(i_8_), .B(i_7_), .Y(new_new_n136_));
  NA2        g0114(.A(new_new_n136_), .B(i_6_), .Y(new_new_n137_));
  NO2        g0115(.A(i_12_), .B(i_13_), .Y(new_new_n138_));
  NAi21      g0116(.An(i_5_), .B(i_11_), .Y(new_new_n139_));
  NOi21      g0117(.An(new_new_n138_), .B(new_new_n139_), .Y(new_new_n140_));
  NO2        g0118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NA2        g0119(.A(i_2_), .B(i_3_), .Y(new_new_n142_));
  NO2        g0120(.A(new_new_n142_), .B(i_4_), .Y(new_new_n143_));
  NA3        g0121(.A(new_new_n143_), .B(new_new_n141_), .C(new_new_n140_), .Y(new_new_n144_));
  OR2        g0122(.A(new_new_n144_), .B(new_new_n25_), .Y(new_new_n145_));
  AN2        g0123(.A(new_new_n138_), .B(new_new_n81_), .Y(new_new_n146_));
  NO2        g0124(.A(new_new_n146_), .B(new_new_n27_), .Y(new_new_n147_));
  NA2        g0125(.A(i_1_), .B(i_5_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n71_), .B(new_new_n47_), .Y(new_new_n149_));
  NA2        g0127(.A(new_new_n149_), .B(new_new_n36_), .Y(new_new_n150_));
  NO3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  OR2        g0129(.A(i_0_), .B(i_1_), .Y(new_new_n152_));
  NO3        g0130(.A(new_new_n152_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n153_));
  NAi32      g0131(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n154_));
  NAi21      g0132(.An(new_new_n154_), .B(new_new_n153_), .Y(new_new_n155_));
  NOi21      g0133(.An(i_4_), .B(i_10_), .Y(new_new_n156_));
  NA2        g0134(.A(new_new_n156_), .B(new_new_n40_), .Y(new_new_n157_));
  NO2        g0135(.A(i_3_), .B(i_5_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n159_));
  NA2        g0137(.A(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  OAI210     g0138(.A0(new_new_n160_), .A1(new_new_n157_), .B0(new_new_n155_), .Y(new_new_n161_));
  NO2        g0139(.A(new_new_n161_), .B(new_new_n151_), .Y(new_new_n162_));
  AOI210     g0140(.A0(new_new_n162_), .A1(new_new_n145_), .B0(new_new_n137_), .Y(new_new_n163_));
  NA3        g0141(.A(new_new_n71_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n164_));
  NOi21      g0142(.An(i_4_), .B(i_9_), .Y(new_new_n165_));
  NOi21      g0143(.An(i_11_), .B(i_13_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  NO2        g0145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g0146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g0147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA3        g0148(.A(new_new_n170_), .B(new_new_n168_), .C(new_new_n81_), .Y(new_new_n171_));
  AOI210     g0149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n164_), .Y(new_new_n172_));
  NO2        g0150(.A(new_new_n71_), .B(new_new_n63_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n36_), .B(i_5_), .Y(new_new_n174_));
  NAi31      g0152(.An(new_new_n174_), .B(new_new_n146_), .C(i_11_), .Y(new_new_n175_));
  NA2        g0153(.A(i_3_), .B(i_5_), .Y(new_new_n176_));
  OR2        g0154(.A(new_new_n176_), .B(new_new_n167_), .Y(new_new_n177_));
  AOI210     g0155(.A0(new_new_n177_), .A1(new_new_n175_), .B0(new_new_n63_), .Y(new_new_n178_));
  NO2        g0156(.A(new_new_n71_), .B(i_5_), .Y(new_new_n179_));
  NO2        g0157(.A(i_13_), .B(i_10_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n179_), .C(new_new_n45_), .Y(new_new_n181_));
  NO2        g0159(.A(i_2_), .B(i_1_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n182_), .B(i_3_), .Y(new_new_n183_));
  NAi21      g0161(.An(i_4_), .B(i_12_), .Y(new_new_n184_));
  NO4        g0162(.A(new_new_n184_), .B(new_new_n183_), .C(new_new_n181_), .D(new_new_n25_), .Y(new_new_n185_));
  NO3        g0163(.A(new_new_n185_), .B(new_new_n178_), .C(new_new_n172_), .Y(new_new_n186_));
  INV        g0164(.A(i_8_), .Y(new_new_n187_));
  NO2        g0165(.A(new_new_n187_), .B(i_7_), .Y(new_new_n188_));
  NA2        g0166(.A(new_new_n188_), .B(i_6_), .Y(new_new_n189_));
  NO3        g0167(.A(i_3_), .B(new_new_n83_), .C(new_new_n49_), .Y(new_new_n190_));
  NA2        g0168(.A(new_new_n190_), .B(new_new_n106_), .Y(new_new_n191_));
  NO3        g0169(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n192_));
  NA3        g0170(.A(new_new_n192_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n193_));
  NO3        g0171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n194_));
  OAI210     g0172(.A0(new_new_n90_), .A1(i_12_), .B0(new_new_n194_), .Y(new_new_n195_));
  AOI210     g0173(.A0(new_new_n195_), .A1(new_new_n193_), .B0(new_new_n191_), .Y(new_new_n196_));
  NO2        g0174(.A(i_3_), .B(i_8_), .Y(new_new_n197_));
  NO3        g0175(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n198_));
  NA3        g0176(.A(new_new_n198_), .B(new_new_n197_), .C(new_new_n40_), .Y(new_new_n199_));
  NO2        g0177(.A(new_new_n97_), .B(new_new_n58_), .Y(new_new_n200_));
  NO2        g0178(.A(i_13_), .B(i_9_), .Y(new_new_n201_));
  NA3        g0179(.A(new_new_n201_), .B(i_6_), .C(new_new_n187_), .Y(new_new_n202_));
  NAi21      g0180(.An(i_12_), .B(i_3_), .Y(new_new_n203_));
  OR2        g0181(.A(new_new_n203_), .B(new_new_n202_), .Y(new_new_n204_));
  NO2        g0182(.A(new_new_n45_), .B(i_5_), .Y(new_new_n205_));
  NO3        g0183(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n206_));
  INV        g0184(.A(new_new_n206_), .Y(new_new_n207_));
  OAI220     g0185(.A0(new_new_n207_), .A1(new_new_n204_), .B0(new_new_n97_), .B1(new_new_n199_), .Y(new_new_n208_));
  AOI210     g0186(.A0(new_new_n208_), .A1(i_7_), .B0(new_new_n196_), .Y(new_new_n209_));
  OAI220     g0187(.A0(new_new_n209_), .A1(i_4_), .B0(new_new_n189_), .B1(new_new_n186_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_7_), .Y(new_new_n211_));
  NA3        g0189(.A(i_13_), .B(new_new_n187_), .C(i_10_), .Y(new_new_n212_));
  NO2        g0190(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n213_));
  NA2        g0191(.A(i_0_), .B(i_5_), .Y(new_new_n214_));
  OAI220     g0192(.A0(new_new_n83_), .A1(new_new_n183_), .B0(new_new_n63_), .B1(new_new_n127_), .Y(new_new_n215_));
  NAi31      g0193(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n36_), .B(i_13_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n218_));
  NA3        g0196(.A(new_new_n218_), .B(i_0_), .C(new_new_n217_), .Y(new_new_n219_));
  INV        g0197(.A(i_13_), .Y(new_new_n220_));
  NO2        g0198(.A(i_12_), .B(new_new_n220_), .Y(new_new_n221_));
  NA3        g0199(.A(new_new_n221_), .B(new_new_n192_), .C(new_new_n190_), .Y(new_new_n222_));
  OAI210     g0200(.A0(new_new_n219_), .A1(new_new_n216_), .B0(new_new_n222_), .Y(new_new_n223_));
  AOI220     g0201(.A0(new_new_n223_), .A1(new_new_n136_), .B0(new_new_n215_), .B1(new_new_n213_), .Y(new_new_n224_));
  NO2        g0202(.A(i_12_), .B(new_new_n37_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n176_), .B(i_4_), .Y(new_new_n226_));
  NA2        g0204(.A(new_new_n226_), .B(new_new_n225_), .Y(new_new_n227_));
  OR2        g0205(.A(i_8_), .B(i_7_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n228_), .B(new_new_n83_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n54_), .B(i_1_), .Y(new_new_n230_));
  NA2        g0208(.A(new_new_n230_), .B(new_new_n229_), .Y(new_new_n231_));
  INV        g0209(.A(i_12_), .Y(new_new_n232_));
  NO3        g0210(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n233_));
  NA2        g0211(.A(i_2_), .B(i_1_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n231_), .B(new_new_n227_), .Y(new_new_n235_));
  NO3        g0213(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n236_));
  NAi21      g0214(.An(i_4_), .B(i_3_), .Y(new_new_n237_));
  NO2        g0215(.A(i_0_), .B(i_6_), .Y(new_new_n238_));
  NOi41      g0216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n234_), .B(new_new_n176_), .Y(new_new_n241_));
  NAi21      g0219(.An(new_new_n240_), .B(new_new_n241_), .Y(new_new_n242_));
  INV        g0220(.A(new_new_n242_), .Y(new_new_n243_));
  AOI220     g0221(.A0(new_new_n243_), .A1(new_new_n40_), .B0(new_new_n235_), .B1(new_new_n201_), .Y(new_new_n244_));
  NO2        g0222(.A(i_11_), .B(new_new_n220_), .Y(new_new_n245_));
  NOi21      g0223(.An(i_1_), .B(i_6_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_3_), .B(i_7_), .Y(new_new_n247_));
  NO2        g0225(.A(i_12_), .B(i_3_), .Y(new_new_n248_));
  NA2        g0226(.A(i_3_), .B(i_9_), .Y(new_new_n249_));
  NA3        g0227(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n250_));
  INV        g0228(.A(new_new_n137_), .Y(new_new_n251_));
  NA2        g0229(.A(new_new_n232_), .B(i_13_), .Y(new_new_n252_));
  NO2        g0230(.A(new_new_n252_), .B(new_new_n73_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n253_), .B(new_new_n251_), .Y(new_new_n254_));
  NO2        g0232(.A(new_new_n228_), .B(new_new_n37_), .Y(new_new_n255_));
  NA2        g0233(.A(i_12_), .B(i_6_), .Y(new_new_n256_));
  OR2        g0234(.A(i_13_), .B(i_9_), .Y(new_new_n257_));
  NO3        g0235(.A(new_new_n257_), .B(new_new_n256_), .C(new_new_n49_), .Y(new_new_n258_));
  NO2        g0236(.A(new_new_n237_), .B(i_2_), .Y(new_new_n259_));
  NA3        g0237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n45_), .Y(new_new_n260_));
  NA2        g0238(.A(new_new_n245_), .B(i_9_), .Y(new_new_n261_));
  OAI210     g0239(.A0(new_new_n63_), .A1(new_new_n261_), .B0(new_new_n260_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n149_), .B(new_new_n63_), .Y(new_new_n263_));
  NO3        g0241(.A(i_11_), .B(new_new_n220_), .C(new_new_n25_), .Y(new_new_n264_));
  NO2        g0242(.A(new_new_n247_), .B(i_8_), .Y(new_new_n265_));
  NO2        g0243(.A(i_6_), .B(new_new_n49_), .Y(new_new_n266_));
  NA2        g0244(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n267_));
  NO3        g0245(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n268_));
  NA3        g0246(.A(new_new_n268_), .B(new_new_n255_), .C(new_new_n221_), .Y(new_new_n269_));
  AOI210     g0247(.A0(new_new_n269_), .A1(new_new_n267_), .B0(new_new_n263_), .Y(new_new_n270_));
  AOI210     g0248(.A0(new_new_n262_), .A1(new_new_n255_), .B0(new_new_n270_), .Y(new_new_n271_));
  NA4        g0249(.A(new_new_n271_), .B(new_new_n254_), .C(new_new_n244_), .D(new_new_n224_), .Y(new_new_n272_));
  NO3        g0250(.A(i_12_), .B(new_new_n220_), .C(new_new_n37_), .Y(new_new_n273_));
  INV        g0251(.A(new_new_n273_), .Y(new_new_n274_));
  NO3        g0252(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n275_));
  AOI220     g0253(.A0(new_new_n275_), .A1(new_new_n190_), .B0(new_new_n158_), .B1(new_new_n230_), .Y(new_new_n276_));
  NO2        g0254(.A(new_new_n276_), .B(new_new_n1025_), .Y(new_new_n277_));
  NO3        g0255(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n234_), .B(i_0_), .Y(new_new_n279_));
  AOI220     g0257(.A0(new_new_n279_), .A1(new_new_n188_), .B0(new_new_n278_), .B1(new_new_n136_), .Y(new_new_n280_));
  NA2        g0258(.A(new_new_n266_), .B(new_new_n26_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n281_), .B(new_new_n280_), .Y(new_new_n282_));
  NA2        g0260(.A(i_0_), .B(i_1_), .Y(new_new_n283_));
  NO2        g0261(.A(new_new_n283_), .B(i_2_), .Y(new_new_n284_));
  NO2        g0262(.A(new_new_n59_), .B(i_6_), .Y(new_new_n285_));
  NA3        g0263(.A(new_new_n285_), .B(new_new_n284_), .C(new_new_n158_), .Y(new_new_n286_));
  OAI210     g0264(.A0(new_new_n160_), .A1(new_new_n137_), .B0(new_new_n286_), .Y(new_new_n287_));
  NO3        g0265(.A(new_new_n287_), .B(new_new_n282_), .C(new_new_n277_), .Y(new_new_n288_));
  NO2        g0266(.A(i_3_), .B(i_10_), .Y(new_new_n289_));
  NA3        g0267(.A(new_new_n289_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n290_));
  NO2        g0268(.A(i_2_), .B(new_new_n95_), .Y(new_new_n291_));
  NA2        g0269(.A(i_1_), .B(new_new_n36_), .Y(new_new_n292_));
  NOi21      g0270(.An(new_new_n214_), .B(new_new_n97_), .Y(new_new_n293_));
  NA3        g0271(.A(new_new_n293_), .B(i_1_), .C(new_new_n291_), .Y(new_new_n294_));
  AN2        g0272(.A(i_3_), .B(i_10_), .Y(new_new_n295_));
  NA4        g0273(.A(new_new_n295_), .B(new_new_n192_), .C(new_new_n170_), .D(new_new_n168_), .Y(new_new_n296_));
  NO2        g0274(.A(i_5_), .B(new_new_n37_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n298_));
  OR2        g0276(.A(new_new_n294_), .B(new_new_n290_), .Y(new_new_n299_));
  OAI220     g0277(.A0(new_new_n299_), .A1(i_6_), .B0(new_new_n288_), .B1(new_new_n274_), .Y(new_new_n300_));
  NO4        g0278(.A(new_new_n300_), .B(new_new_n272_), .C(new_new_n210_), .D(new_new_n163_), .Y(new_new_n301_));
  NO3        g0279(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n59_), .B(new_new_n83_), .Y(new_new_n303_));
  NA2        g0281(.A(new_new_n279_), .B(new_new_n303_), .Y(new_new_n304_));
  NO3        g0282(.A(i_6_), .B(new_new_n187_), .C(i_7_), .Y(new_new_n305_));
  NA2        g0283(.A(new_new_n305_), .B(new_new_n192_), .Y(new_new_n306_));
  AOI210     g0284(.A0(new_new_n306_), .A1(new_new_n304_), .B0(i_5_), .Y(new_new_n307_));
  NO2        g0285(.A(i_2_), .B(i_3_), .Y(new_new_n308_));
  OR2        g0286(.A(i_0_), .B(i_5_), .Y(new_new_n309_));
  NA2        g0287(.A(new_new_n214_), .B(new_new_n309_), .Y(new_new_n310_));
  NA4        g0288(.A(new_new_n310_), .B(new_new_n229_), .C(new_new_n308_), .D(i_1_), .Y(new_new_n311_));
  NA3        g0289(.A(new_new_n279_), .B(new_new_n158_), .C(new_new_n106_), .Y(new_new_n312_));
  NAi21      g0290(.An(i_8_), .B(i_7_), .Y(new_new_n313_));
  NO2        g0291(.A(new_new_n152_), .B(new_new_n47_), .Y(new_new_n314_));
  NA3        g0292(.A(new_new_n314_), .B(i_7_), .C(new_new_n158_), .Y(new_new_n315_));
  NA3        g0293(.A(new_new_n315_), .B(new_new_n312_), .C(new_new_n311_), .Y(new_new_n316_));
  OAI210     g0294(.A0(new_new_n316_), .A1(new_new_n307_), .B0(i_4_), .Y(new_new_n317_));
  NO2        g0295(.A(i_12_), .B(i_10_), .Y(new_new_n318_));
  NOi21      g0296(.An(i_5_), .B(i_0_), .Y(new_new_n319_));
  NO2        g0297(.A(new_new_n292_), .B(new_new_n122_), .Y(new_new_n320_));
  NA4        g0298(.A(new_new_n82_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n320_), .B(new_new_n318_), .Y(new_new_n322_));
  NO2        g0300(.A(i_6_), .B(i_8_), .Y(new_new_n323_));
  AN2        g0301(.A(i_0_), .B(new_new_n323_), .Y(new_new_n324_));
  NO2        g0302(.A(i_1_), .B(i_7_), .Y(new_new_n325_));
  NA2        g0303(.A(new_new_n324_), .B(new_new_n42_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n322_), .C(new_new_n317_), .Y(new_new_n327_));
  NO3        g0305(.A(new_new_n228_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n328_));
  NO3        g0306(.A(new_new_n313_), .B(i_2_), .C(i_1_), .Y(new_new_n329_));
  OAI210     g0307(.A0(new_new_n329_), .A1(new_new_n328_), .B0(i_6_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n246_), .B(new_new_n291_), .C(new_new_n187_), .Y(new_new_n331_));
  NA2        g0309(.A(new_new_n331_), .B(new_new_n330_), .Y(new_new_n332_));
  NA2        g0310(.A(new_new_n332_), .B(i_3_), .Y(new_new_n333_));
  NO2        g0311(.A(new_new_n283_), .B(new_new_n79_), .Y(new_new_n334_));
  NA2        g0312(.A(new_new_n334_), .B(new_new_n126_), .Y(new_new_n335_));
  NO2        g0313(.A(new_new_n88_), .B(new_new_n187_), .Y(new_new_n336_));
  NA2        g0314(.A(new_new_n293_), .B(new_new_n336_), .Y(new_new_n337_));
  AOI210     g0315(.A0(new_new_n337_), .A1(new_new_n335_), .B0(i_3_), .Y(new_new_n338_));
  NO2        g0316(.A(new_new_n187_), .B(i_9_), .Y(new_new_n339_));
  NA2        g0317(.A(new_new_n339_), .B(new_new_n200_), .Y(new_new_n340_));
  NO2        g0318(.A(new_new_n338_), .B(new_new_n282_), .Y(new_new_n341_));
  AOI210     g0319(.A0(new_new_n341_), .A1(new_new_n333_), .B0(new_new_n157_), .Y(new_new_n342_));
  AOI210     g0320(.A0(new_new_n327_), .A1(new_new_n302_), .B0(new_new_n342_), .Y(new_new_n343_));
  NOi32      g0321(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n344_));
  INV        g0322(.A(new_new_n344_), .Y(new_new_n345_));
  NAi21      g0323(.An(i_1_), .B(i_5_), .Y(new_new_n346_));
  INV        g0324(.A(new_new_n240_), .Y(new_new_n347_));
  NAi41      g0325(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n348_));
  OAI220     g0326(.A0(new_new_n348_), .A1(new_new_n346_), .B0(new_new_n216_), .B1(new_new_n154_), .Y(new_new_n349_));
  AOI210     g0327(.A0(new_new_n348_), .A1(new_new_n154_), .B0(new_new_n152_), .Y(new_new_n350_));
  NOi32      g0328(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n351_));
  NAi21      g0329(.An(i_6_), .B(i_1_), .Y(new_new_n352_));
  NA3        g0330(.A(new_new_n352_), .B(new_new_n351_), .C(new_new_n47_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n353_), .B(i_0_), .Y(new_new_n354_));
  OR3        g0332(.A(new_new_n354_), .B(new_new_n350_), .C(new_new_n349_), .Y(new_new_n355_));
  NO2        g0333(.A(i_1_), .B(new_new_n95_), .Y(new_new_n356_));
  NAi21      g0334(.An(i_3_), .B(i_4_), .Y(new_new_n357_));
  NO2        g0335(.A(new_new_n357_), .B(i_9_), .Y(new_new_n358_));
  AN2        g0336(.A(i_6_), .B(i_7_), .Y(new_new_n359_));
  OAI210     g0337(.A0(new_new_n359_), .A1(new_new_n356_), .B0(new_new_n358_), .Y(new_new_n360_));
  NA2        g0338(.A(i_2_), .B(i_7_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n357_), .B(i_10_), .Y(new_new_n362_));
  NA3        g0340(.A(new_new_n362_), .B(new_new_n361_), .C(new_new_n238_), .Y(new_new_n363_));
  AOI210     g0341(.A0(new_new_n363_), .A1(new_new_n360_), .B0(new_new_n179_), .Y(new_new_n364_));
  AOI220     g0342(.A0(new_new_n362_), .A1(new_new_n325_), .B0(new_new_n233_), .B1(new_new_n182_), .Y(new_new_n365_));
  NO2        g0343(.A(new_new_n365_), .B(i_5_), .Y(new_new_n366_));
  NO4        g0344(.A(new_new_n366_), .B(new_new_n364_), .C(new_new_n355_), .D(new_new_n347_), .Y(new_new_n367_));
  NO2        g0345(.A(new_new_n367_), .B(new_new_n345_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n369_));
  AN2        g0347(.A(i_12_), .B(i_5_), .Y(new_new_n370_));
  NO2        g0348(.A(i_4_), .B(new_new_n26_), .Y(new_new_n371_));
  NA2        g0349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  NO2        g0350(.A(i_11_), .B(i_6_), .Y(new_new_n373_));
  NA3        g0351(.A(new_new_n373_), .B(new_new_n314_), .C(new_new_n220_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n374_), .B(new_new_n372_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n237_), .B(i_5_), .Y(new_new_n376_));
  NO2        g0354(.A(i_5_), .B(i_10_), .Y(new_new_n377_));
  AOI220     g0355(.A0(new_new_n377_), .A1(new_new_n259_), .B0(new_new_n376_), .B1(new_new_n192_), .Y(new_new_n378_));
  NO2        g0356(.A(new_new_n1020_), .B(new_new_n378_), .Y(new_new_n379_));
  OAI210     g0357(.A0(new_new_n379_), .A1(new_new_n375_), .B0(new_new_n369_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n382_));
  OAI210     g0360(.A0(new_new_n382_), .A1(new_new_n375_), .B0(new_new_n381_), .Y(new_new_n383_));
  NO3        g0361(.A(new_new_n83_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n384_));
  NA2        g0362(.A(new_new_n289_), .B(new_new_n87_), .Y(new_new_n385_));
  NO2        g0363(.A(i_11_), .B(i_12_), .Y(new_new_n386_));
  NA2        g0364(.A(new_new_n386_), .B(new_new_n36_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n385_), .B(new_new_n387_), .Y(new_new_n388_));
  NA2        g0366(.A(new_new_n377_), .B(new_new_n232_), .Y(new_new_n389_));
  INV        g0367(.A(new_new_n42_), .Y(new_new_n390_));
  NO2        g0368(.A(new_new_n390_), .B(new_new_n216_), .Y(new_new_n391_));
  NAi21      g0369(.An(i_13_), .B(i_0_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n392_), .B(new_new_n234_), .Y(new_new_n393_));
  OAI210     g0371(.A0(new_new_n391_), .A1(new_new_n388_), .B0(new_new_n393_), .Y(new_new_n394_));
  NA3        g0372(.A(new_new_n394_), .B(new_new_n383_), .C(new_new_n380_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n45_), .B(new_new_n220_), .Y(new_new_n396_));
  NO3        g0374(.A(i_1_), .B(i_12_), .C(new_new_n83_), .Y(new_new_n397_));
  NO2        g0375(.A(i_0_), .B(i_11_), .Y(new_new_n398_));
  AN2        g0376(.A(i_1_), .B(i_6_), .Y(new_new_n399_));
  NOi21      g0377(.An(i_2_), .B(i_12_), .Y(new_new_n400_));
  NA2        g0378(.A(new_new_n400_), .B(new_new_n399_), .Y(new_new_n401_));
  INV        g0379(.A(new_new_n401_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n136_), .B(i_9_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(i_4_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n402_), .B(new_new_n404_), .Y(new_new_n405_));
  NAi21      g0383(.An(i_9_), .B(i_4_), .Y(new_new_n406_));
  OR2        g0384(.A(i_13_), .B(i_10_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n167_), .B(new_new_n117_), .Y(new_new_n408_));
  BUFFER     g0386(.A(new_new_n212_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n95_), .B(new_new_n25_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n266_), .B(new_new_n206_), .Y(new_new_n411_));
  NO2        g0389(.A(new_new_n411_), .B(new_new_n409_), .Y(new_new_n412_));
  INV        g0390(.A(new_new_n412_), .Y(new_new_n413_));
  AOI210     g0391(.A0(new_new_n413_), .A1(new_new_n405_), .B0(new_new_n26_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n312_), .B(new_new_n311_), .Y(new_new_n415_));
  AOI220     g0393(.A0(new_new_n285_), .A1(new_new_n275_), .B0(new_new_n279_), .B1(new_new_n303_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n416_), .B(i_5_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n176_), .B(new_new_n83_), .Y(new_new_n418_));
  AOI220     g0396(.A0(new_new_n418_), .A1(new_new_n284_), .B0(new_new_n268_), .B1(new_new_n206_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n1025_), .Y(new_new_n420_));
  NO3        g0398(.A(new_new_n420_), .B(new_new_n417_), .C(new_new_n415_), .Y(new_new_n421_));
  INV        g0399(.A(new_new_n90_), .Y(new_new_n422_));
  NA3        g0400(.A(new_new_n314_), .B(new_new_n158_), .C(new_new_n83_), .Y(new_new_n423_));
  AOI210     g0401(.A0(new_new_n423_), .A1(new_new_n422_), .B0(new_new_n313_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n285_), .B(new_new_n230_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(new_new_n176_), .Y(new_new_n426_));
  NO2        g0404(.A(i_3_), .B(new_new_n49_), .Y(new_new_n427_));
  NA3        g0405(.A(new_new_n325_), .B(new_new_n324_), .C(new_new_n427_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n305_), .B(new_new_n310_), .Y(new_new_n429_));
  OAI210     g0407(.A0(new_new_n429_), .A1(new_new_n183_), .B0(new_new_n428_), .Y(new_new_n430_));
  NO3        g0408(.A(new_new_n430_), .B(new_new_n426_), .C(new_new_n424_), .Y(new_new_n431_));
  AOI210     g0409(.A0(new_new_n431_), .A1(new_new_n421_), .B0(new_new_n261_), .Y(new_new_n432_));
  NO4        g0410(.A(new_new_n432_), .B(new_new_n414_), .C(new_new_n395_), .D(new_new_n368_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n71_), .B(i_13_), .Y(new_new_n434_));
  NO2        g0412(.A(i_10_), .B(i_9_), .Y(new_new_n435_));
  NAi21      g0413(.An(i_12_), .B(i_8_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(i_3_), .Y(new_new_n437_));
  NA2        g0415(.A(i_2_), .B(new_new_n98_), .Y(new_new_n438_));
  NO2        g0416(.A(new_new_n438_), .B(new_new_n199_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n298_), .B(i_0_), .Y(new_new_n440_));
  NO3        g0418(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n256_), .B(new_new_n91_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n442_), .B(new_new_n441_), .Y(new_new_n443_));
  NA2        g0421(.A(i_8_), .B(i_9_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n273_), .B(new_new_n200_), .Y(new_new_n445_));
  OAI220     g0423(.A0(new_new_n445_), .A1(new_new_n444_), .B0(new_new_n443_), .B1(new_new_n440_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n245_), .B(new_new_n297_), .Y(new_new_n447_));
  NO3        g0425(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n448_));
  INV        g0426(.A(new_new_n448_), .Y(new_new_n449_));
  NA3        g0427(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n450_));
  NA4        g0428(.A(new_new_n139_), .B(new_new_n109_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n451_));
  OAI220     g0429(.A0(new_new_n451_), .A1(new_new_n450_), .B0(new_new_n449_), .B1(new_new_n447_), .Y(new_new_n452_));
  NO3        g0430(.A(new_new_n452_), .B(new_new_n446_), .C(new_new_n439_), .Y(new_new_n453_));
  NA2        g0431(.A(new_new_n284_), .B(new_new_n102_), .Y(new_new_n454_));
  OR2        g0432(.A(new_new_n454_), .B(new_new_n202_), .Y(new_new_n455_));
  OR2        g0433(.A(new_new_n340_), .B(new_new_n95_), .Y(new_new_n456_));
  OA220      g0434(.A0(new_new_n456_), .A1(new_new_n157_), .B0(new_new_n455_), .B1(new_new_n227_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n90_), .B(i_13_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n418_), .B(new_new_n369_), .Y(new_new_n459_));
  NO2        g0437(.A(i_2_), .B(i_13_), .Y(new_new_n460_));
  NA3        g0438(.A(new_new_n460_), .B(new_new_n156_), .C(new_new_n93_), .Y(new_new_n461_));
  NO2        g0439(.A(new_new_n459_), .B(new_new_n458_), .Y(new_new_n462_));
  NO3        g0440(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n463_));
  NO2        g0441(.A(i_6_), .B(i_7_), .Y(new_new_n464_));
  NA2        g0442(.A(new_new_n464_), .B(new_new_n463_), .Y(new_new_n465_));
  NO2        g0443(.A(i_11_), .B(i_1_), .Y(new_new_n466_));
  OR2        g0444(.A(i_11_), .B(i_8_), .Y(new_new_n467_));
  NOi21      g0445(.An(i_2_), .B(i_7_), .Y(new_new_n468_));
  NAi31      g0446(.An(new_new_n467_), .B(new_new_n468_), .C(i_0_), .Y(new_new_n469_));
  NO2        g0447(.A(new_new_n407_), .B(i_6_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n470_), .B(i_1_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n471_), .B(new_new_n469_), .Y(new_new_n472_));
  NO2        g0450(.A(i_3_), .B(new_new_n187_), .Y(new_new_n473_));
  NO2        g0451(.A(i_6_), .B(i_10_), .Y(new_new_n474_));
  NA3        g0452(.A(new_new_n474_), .B(new_new_n302_), .C(new_new_n473_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n475_), .B(new_new_n150_), .Y(new_new_n476_));
  NA3        g0454(.A(new_new_n239_), .B(new_new_n166_), .C(new_new_n126_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n152_), .B(i_3_), .Y(new_new_n478_));
  NA3        g0456(.A(new_new_n381_), .B(new_new_n173_), .C(new_new_n143_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n479_), .B(new_new_n477_), .Y(new_new_n480_));
  NO4        g0458(.A(new_new_n480_), .B(new_new_n476_), .C(new_new_n472_), .D(new_new_n462_), .Y(new_new_n481_));
  NA2        g0459(.A(new_new_n441_), .B(new_new_n370_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n448_), .B(new_new_n377_), .Y(new_new_n483_));
  NO2        g0461(.A(new_new_n483_), .B(new_new_n219_), .Y(new_new_n484_));
  NAi21      g0462(.An(new_new_n212_), .B(new_new_n386_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n325_), .B(new_new_n214_), .Y(new_new_n486_));
  NO2        g0464(.A(new_new_n26_), .B(i_5_), .Y(new_new_n487_));
  NA3        g0465(.A(i_6_), .B(new_new_n487_), .C(new_new_n136_), .Y(new_new_n488_));
  OR3        g0466(.A(new_new_n292_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n489_));
  OAI220     g0467(.A0(new_new_n489_), .A1(new_new_n488_), .B0(new_new_n486_), .B1(new_new_n485_), .Y(new_new_n490_));
  NA3        g0468(.A(new_new_n295_), .B(new_new_n218_), .C(new_new_n71_), .Y(new_new_n491_));
  NO2        g0469(.A(new_new_n491_), .B(new_new_n465_), .Y(new_new_n492_));
  NO3        g0470(.A(new_new_n492_), .B(new_new_n490_), .C(new_new_n484_), .Y(new_new_n493_));
  NA4        g0471(.A(new_new_n493_), .B(new_new_n481_), .C(new_new_n457_), .D(new_new_n453_), .Y(new_new_n494_));
  NA3        g0472(.A(new_new_n295_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n495_));
  OAI210     g0473(.A0(new_new_n290_), .A1(new_new_n174_), .B0(new_new_n495_), .Y(new_new_n496_));
  AN2        g0474(.A(new_new_n275_), .B(new_new_n229_), .Y(new_new_n497_));
  NA2        g0475(.A(new_new_n497_), .B(new_new_n496_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n116_), .B(new_new_n105_), .Y(new_new_n499_));
  AN2        g0477(.A(new_new_n499_), .B(new_new_n441_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n302_), .B(new_new_n159_), .Y(new_new_n501_));
  OAI210     g0479(.A0(new_new_n501_), .A1(new_new_n227_), .B0(new_new_n296_), .Y(new_new_n502_));
  AOI220     g0480(.A0(new_new_n502_), .A1(i_7_), .B0(new_new_n500_), .B1(new_new_n298_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n344_), .B(new_new_n71_), .Y(new_new_n504_));
  NA2        g0482(.A(new_new_n359_), .B(new_new_n351_), .Y(new_new_n505_));
  NO2        g0483(.A(new_new_n36_), .B(i_8_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n39_), .B(i_13_), .Y(new_new_n507_));
  OAI210     g0485(.A0(i_8_), .A1(new_new_n63_), .B0(new_new_n128_), .Y(new_new_n508_));
  AOI210     g0486(.A0(new_new_n188_), .A1(i_9_), .B0(new_new_n255_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n509_), .B(new_new_n193_), .Y(new_new_n510_));
  OR2        g0488(.A(new_new_n176_), .B(i_4_), .Y(new_new_n511_));
  INV        g0489(.A(new_new_n511_), .Y(new_new_n512_));
  AOI220     g0490(.A0(new_new_n512_), .A1(new_new_n510_), .B0(new_new_n508_), .B1(new_new_n408_), .Y(new_new_n513_));
  NA4        g0491(.A(new_new_n513_), .B(new_new_n507_), .C(new_new_n503_), .D(new_new_n498_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n376_), .B(new_new_n284_), .Y(new_new_n515_));
  OAI210     g0493(.A0(new_new_n372_), .A1(new_new_n164_), .B0(new_new_n515_), .Y(new_new_n516_));
  NO2        g0494(.A(i_12_), .B(new_new_n187_), .Y(new_new_n517_));
  NOi31      g0495(.An(new_new_n305_), .B(new_new_n407_), .C(new_new_n38_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n518_), .B(new_new_n516_), .Y(new_new_n519_));
  NO2        g0497(.A(i_8_), .B(i_7_), .Y(new_new_n520_));
  OAI210     g0498(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n521_), .B(new_new_n218_), .Y(new_new_n522_));
  NA2        g0500(.A(new_new_n45_), .B(i_10_), .Y(new_new_n523_));
  NO2        g0501(.A(new_new_n523_), .B(i_6_), .Y(new_new_n524_));
  NA3        g0502(.A(new_new_n524_), .B(new_new_n1024_), .C(new_new_n520_), .Y(new_new_n525_));
  AOI220     g0503(.A0(new_new_n418_), .A1(new_new_n314_), .B0(new_new_n241_), .B1(new_new_n238_), .Y(new_new_n526_));
  OAI220     g0504(.A0(new_new_n526_), .A1(new_new_n252_), .B0(new_new_n458_), .B1(new_new_n127_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n527_), .B(new_new_n255_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n290_), .B(new_new_n174_), .Y(new_new_n529_));
  NA3        g0507(.A(new_new_n295_), .B(new_new_n168_), .C(new_new_n90_), .Y(new_new_n530_));
  NO2        g0508(.A(new_new_n152_), .B(i_5_), .Y(new_new_n531_));
  NA3        g0509(.A(new_new_n531_), .B(new_new_n396_), .C(new_new_n308_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n532_), .B(new_new_n530_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n533_), .A1(new_new_n529_), .B0(new_new_n448_), .Y(new_new_n534_));
  NA4        g0512(.A(new_new_n534_), .B(new_new_n528_), .C(new_new_n525_), .D(new_new_n519_), .Y(new_new_n535_));
  NA3        g0513(.A(new_new_n214_), .B(new_new_n69_), .C(new_new_n45_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n273_), .B(new_new_n82_), .Y(new_new_n537_));
  AOI210     g0515(.A0(new_new_n536_), .A1(new_new_n335_), .B0(new_new_n537_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n285_), .B(new_new_n275_), .Y(new_new_n539_));
  NO2        g0517(.A(new_new_n539_), .B(new_new_n167_), .Y(new_new_n540_));
  NA2        g0518(.A(i_0_), .B(new_new_n49_), .Y(new_new_n541_));
  NA3        g0519(.A(new_new_n517_), .B(new_new_n264_), .C(new_new_n541_), .Y(new_new_n542_));
  NO2        g0520(.A(i_1_), .B(new_new_n542_), .Y(new_new_n543_));
  NO3        g0521(.A(new_new_n543_), .B(new_new_n540_), .C(new_new_n538_), .Y(new_new_n544_));
  NO4        g0522(.A(new_new_n246_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n545_));
  NO3        g0523(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n546_));
  NO2        g0524(.A(new_new_n228_), .B(new_new_n36_), .Y(new_new_n547_));
  AN2        g0525(.A(new_new_n547_), .B(new_new_n546_), .Y(new_new_n548_));
  OA210      g0526(.A0(new_new_n548_), .A1(new_new_n545_), .B0(new_new_n344_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n407_), .B(i_1_), .Y(new_new_n550_));
  NOi31      g0528(.An(new_new_n550_), .B(new_new_n442_), .C(new_new_n71_), .Y(new_new_n551_));
  AN3        g0529(.A(new_new_n551_), .B(new_new_n404_), .C(new_new_n487_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n416_), .B(new_new_n171_), .Y(new_new_n553_));
  NO3        g0531(.A(new_new_n553_), .B(new_new_n552_), .C(new_new_n549_), .Y(new_new_n554_));
  NOi21      g0532(.An(i_10_), .B(i_6_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n556_));
  AOI220     g0534(.A0(new_new_n273_), .A1(new_new_n556_), .B0(new_new_n264_), .B1(new_new_n555_), .Y(new_new_n557_));
  NO2        g0535(.A(new_new_n557_), .B(new_new_n440_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n108_), .B(new_new_n23_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n305_), .B(new_new_n159_), .Y(new_new_n560_));
  AOI220     g0538(.A0(new_new_n560_), .A1(new_new_n425_), .B0(new_new_n177_), .B1(new_new_n175_), .Y(new_new_n561_));
  NOi21      g0539(.An(new_new_n140_), .B(new_new_n321_), .Y(new_new_n562_));
  NO3        g0540(.A(new_new_n562_), .B(new_new_n561_), .C(new_new_n558_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n504_), .B(new_new_n365_), .Y(new_new_n564_));
  INV        g0542(.A(new_new_n308_), .Y(new_new_n565_));
  NO2        g0543(.A(i_12_), .B(new_new_n83_), .Y(new_new_n566_));
  NA3        g0544(.A(new_new_n566_), .B(new_new_n264_), .C(new_new_n541_), .Y(new_new_n567_));
  NA3        g0545(.A(new_new_n373_), .B(new_new_n273_), .C(new_new_n214_), .Y(new_new_n568_));
  AOI210     g0546(.A0(new_new_n568_), .A1(new_new_n567_), .B0(new_new_n565_), .Y(new_new_n569_));
  NA2        g0547(.A(new_new_n168_), .B(i_0_), .Y(new_new_n570_));
  NO3        g0548(.A(new_new_n570_), .B(new_new_n330_), .C(new_new_n290_), .Y(new_new_n571_));
  OR2        g0549(.A(i_2_), .B(i_5_), .Y(new_new_n572_));
  OR2        g0550(.A(new_new_n572_), .B(new_new_n399_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n573_), .B(new_new_n485_), .Y(new_new_n574_));
  NO4        g0552(.A(new_new_n574_), .B(new_new_n571_), .C(new_new_n569_), .D(new_new_n564_), .Y(new_new_n575_));
  NA4        g0553(.A(new_new_n575_), .B(new_new_n563_), .C(new_new_n554_), .D(new_new_n544_), .Y(new_new_n576_));
  NO4        g0554(.A(new_new_n576_), .B(new_new_n535_), .C(new_new_n514_), .D(new_new_n494_), .Y(new_new_n577_));
  NA4        g0555(.A(new_new_n577_), .B(new_new_n433_), .C(new_new_n343_), .D(new_new_n301_), .Y(men7));
  NO2        g0556(.A(new_new_n102_), .B(new_new_n86_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n371_), .B(new_new_n579_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n474_), .B(new_new_n82_), .Y(new_new_n581_));
  NA2        g0559(.A(i_11_), .B(new_new_n187_), .Y(new_new_n582_));
  OAI210     g0560(.A0(new_new_n1023_), .A1(new_new_n581_), .B0(new_new_n580_), .Y(new_new_n583_));
  NA3        g0561(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n232_), .B(i_4_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n99_), .B(new_new_n584_), .Y(new_new_n586_));
  NA2        g0564(.A(i_2_), .B(new_new_n83_), .Y(new_new_n587_));
  OAI210     g0565(.A0(new_new_n85_), .A1(new_new_n197_), .B0(new_new_n198_), .Y(new_new_n588_));
  NO2        g0566(.A(i_7_), .B(new_new_n37_), .Y(new_new_n589_));
  NA2        g0567(.A(i_4_), .B(i_8_), .Y(new_new_n590_));
  AOI210     g0568(.A0(new_new_n590_), .A1(new_new_n295_), .B0(new_new_n589_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n591_), .B(new_new_n587_), .Y(new_new_n592_));
  NO3        g0570(.A(new_new_n592_), .B(new_new_n586_), .C(new_new_n583_), .Y(new_new_n593_));
  INV        g0571(.A(new_new_n156_), .Y(new_new_n594_));
  OR2        g0572(.A(i_6_), .B(i_10_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n595_), .B(new_new_n23_), .Y(new_new_n596_));
  OR3        g0574(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n597_));
  NO3        g0575(.A(new_new_n597_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n598_));
  INV        g0576(.A(new_new_n194_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n598_), .B(new_new_n596_), .Y(new_new_n600_));
  OA220      g0578(.A0(new_new_n600_), .A1(new_new_n565_), .B0(new_new_n594_), .B1(new_new_n257_), .Y(new_new_n601_));
  AOI210     g0579(.A0(new_new_n601_), .A1(new_new_n593_), .B0(new_new_n63_), .Y(new_new_n602_));
  NOi21      g0580(.An(i_11_), .B(i_7_), .Y(new_new_n603_));
  AO210      g0581(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n604_), .B(new_new_n603_), .Y(new_new_n605_));
  NA2        g0583(.A(new_new_n605_), .B(new_new_n201_), .Y(new_new_n606_));
  NA3        g0584(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n607_));
  AOI210     g0585(.A0(new_new_n607_), .A1(new_new_n606_), .B0(new_new_n63_), .Y(new_new_n608_));
  AO210      g0586(.A0(new_new_n84_), .A1(new_new_n365_), .B0(new_new_n41_), .Y(new_new_n609_));
  NA2        g0587(.A(new_new_n221_), .B(new_new_n63_), .Y(new_new_n610_));
  NA2        g0588(.A(new_new_n400_), .B(new_new_n31_), .Y(new_new_n611_));
  OR2        g0589(.A(new_new_n203_), .B(new_new_n102_), .Y(new_new_n612_));
  NA2        g0590(.A(new_new_n612_), .B(new_new_n611_), .Y(new_new_n613_));
  NO2        g0591(.A(new_new_n63_), .B(i_9_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n614_), .B(i_4_), .Y(new_new_n615_));
  NA2        g0593(.A(new_new_n615_), .B(new_new_n613_), .Y(new_new_n616_));
  NO2        g0594(.A(i_1_), .B(i_12_), .Y(new_new_n617_));
  NA3        g0595(.A(new_new_n617_), .B(new_new_n103_), .C(new_new_n24_), .Y(new_new_n618_));
  NA4        g0596(.A(new_new_n618_), .B(new_new_n616_), .C(new_new_n610_), .D(new_new_n609_), .Y(new_new_n619_));
  OAI210     g0597(.A0(new_new_n619_), .A1(new_new_n608_), .B0(i_6_), .Y(new_new_n620_));
  NO2        g0598(.A(i_6_), .B(i_11_), .Y(new_new_n621_));
  INV        g0599(.A(new_new_n443_), .Y(new_new_n622_));
  NO4        g0600(.A(new_new_n211_), .B(new_new_n122_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n623_));
  NA2        g0601(.A(new_new_n623_), .B(new_new_n614_), .Y(new_new_n624_));
  INV        g0602(.A(new_new_n624_), .Y(new_new_n625_));
  NA3        g0603(.A(new_new_n520_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n132_), .B(i_9_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n47_), .B(i_1_), .Y(new_new_n628_));
  NO2        g0606(.A(new_new_n627_), .B(new_new_n1016_), .Y(new_new_n629_));
  NA3        g0607(.A(new_new_n614_), .B(new_new_n308_), .C(i_6_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n630_), .B(new_new_n23_), .Y(new_new_n631_));
  AOI210     g0609(.A0(new_new_n466_), .A1(new_new_n410_), .B0(new_new_n236_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n632_), .B(new_new_n587_), .Y(new_new_n633_));
  NA2        g0611(.A(new_new_n628_), .B(new_new_n256_), .Y(new_new_n634_));
  NO2        g0612(.A(i_11_), .B(new_new_n37_), .Y(new_new_n635_));
  NA2        g0613(.A(new_new_n635_), .B(new_new_n24_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n636_), .B(new_new_n634_), .Y(new_new_n637_));
  OR4        g0615(.A(new_new_n637_), .B(new_new_n633_), .C(new_new_n631_), .D(new_new_n629_), .Y(new_new_n638_));
  NO3        g0616(.A(new_new_n638_), .B(new_new_n625_), .C(new_new_n622_), .Y(new_new_n639_));
  NO2        g0617(.A(new_new_n232_), .B(new_new_n95_), .Y(new_new_n640_));
  NO2        g0618(.A(new_new_n640_), .B(new_new_n603_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n641_), .B(i_1_), .Y(new_new_n642_));
  NO2        g0620(.A(new_new_n642_), .B(new_new_n597_), .Y(new_new_n643_));
  NO2        g0621(.A(new_new_n406_), .B(new_new_n83_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n643_), .B(new_new_n47_), .Y(new_new_n645_));
  NA2        g0623(.A(i_3_), .B(new_new_n187_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n228_), .B(new_new_n45_), .Y(new_new_n647_));
  NO3        g0625(.A(new_new_n647_), .B(new_new_n298_), .C(i_12_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n111_), .B(new_new_n37_), .Y(new_new_n649_));
  NO2        g0627(.A(new_new_n649_), .B(i_6_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n83_), .B(i_9_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n651_), .B(new_new_n63_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n617_), .Y(new_new_n653_));
  NO4        g0631(.A(new_new_n653_), .B(new_new_n650_), .C(new_new_n648_), .D(i_4_), .Y(new_new_n654_));
  NA2        g0632(.A(i_1_), .B(i_3_), .Y(new_new_n655_));
  INV        g0633(.A(new_new_n654_), .Y(new_new_n656_));
  NA4        g0634(.A(new_new_n656_), .B(new_new_n645_), .C(new_new_n639_), .D(new_new_n620_), .Y(new_new_n657_));
  NO3        g0635(.A(new_new_n467_), .B(i_3_), .C(i_7_), .Y(new_new_n658_));
  NOi21      g0636(.An(new_new_n658_), .B(i_10_), .Y(new_new_n659_));
  OA210      g0637(.A0(new_new_n659_), .A1(new_new_n239_), .B0(new_new_n83_), .Y(new_new_n660_));
  NA3        g0638(.A(new_new_n474_), .B(new_new_n506_), .C(new_new_n47_), .Y(new_new_n661_));
  NO3        g0639(.A(new_new_n468_), .B(new_new_n590_), .C(new_new_n83_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(new_new_n25_), .Y(new_new_n663_));
  NA3        g0641(.A(new_new_n156_), .B(new_new_n82_), .C(new_new_n83_), .Y(new_new_n664_));
  NA3        g0642(.A(new_new_n664_), .B(new_new_n663_), .C(new_new_n661_), .Y(new_new_n665_));
  OAI210     g0643(.A0(new_new_n665_), .A1(new_new_n660_), .B0(i_1_), .Y(new_new_n666_));
  AOI210     g0644(.A0(new_new_n256_), .A1(new_new_n91_), .B0(i_1_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n357_), .B(i_2_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n668_), .B(new_new_n667_), .Y(new_new_n669_));
  OAI210     g0647(.A0(new_new_n630_), .A1(new_new_n436_), .B0(new_new_n669_), .Y(new_new_n670_));
  INV        g0648(.A(new_new_n670_), .Y(new_new_n671_));
  AOI210     g0649(.A0(new_new_n671_), .A1(new_new_n666_), .B0(i_13_), .Y(new_new_n672_));
  NA3        g0650(.A(i_11_), .B(new_new_n100_), .C(new_new_n132_), .Y(new_new_n673_));
  AOI220     g0651(.A0(new_new_n460_), .A1(new_new_n156_), .B0(i_2_), .B1(new_new_n132_), .Y(new_new_n674_));
  OAI210     g0652(.A0(new_new_n674_), .A1(new_new_n45_), .B0(new_new_n673_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n55_), .B(i_12_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n468_), .B(new_new_n24_), .Y(new_new_n677_));
  AOI220     g0655(.A0(new_new_n677_), .A1(new_new_n644_), .B0(new_new_n239_), .B1(new_new_n125_), .Y(new_new_n678_));
  OAI220     g0656(.A0(new_new_n678_), .A1(new_new_n41_), .B0(new_new_n1015_), .B1(new_new_n88_), .Y(new_new_n679_));
  AOI210     g0657(.A0(new_new_n675_), .A1(new_new_n323_), .B0(new_new_n679_), .Y(new_new_n680_));
  AOI220     g0658(.A0(i_12_), .A1(new_new_n70_), .B0(new_new_n373_), .B1(new_new_n628_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n681_), .B(new_new_n237_), .Y(new_new_n682_));
  AOI210     g0660(.A0(new_new_n436_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n683_));
  NOi31      g0661(.An(new_new_n683_), .B(new_new_n581_), .C(new_new_n45_), .Y(new_new_n684_));
  NA2        g0662(.A(new_new_n121_), .B(i_13_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n685_), .B(new_new_n667_), .Y(new_new_n686_));
  NO3        g0664(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n95_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n26_), .B(new_new_n187_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n1017_), .B(new_new_n599_), .Y(new_new_n689_));
  NO4        g0667(.A(new_new_n689_), .B(new_new_n686_), .C(new_new_n684_), .D(new_new_n682_), .Y(new_new_n690_));
  OR2        g0668(.A(i_11_), .B(i_6_), .Y(new_new_n691_));
  NA3        g0669(.A(new_new_n585_), .B(new_new_n688_), .C(i_7_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n692_), .B(new_new_n691_), .Y(new_new_n693_));
  NA3        g0671(.A(new_new_n400_), .B(new_new_n589_), .C(new_new_n91_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n621_), .B(i_13_), .Y(new_new_n695_));
  NA2        g0673(.A(new_new_n96_), .B(new_new_n688_), .Y(new_new_n696_));
  NAi21      g0674(.An(i_11_), .B(i_12_), .Y(new_new_n697_));
  NOi41      g0675(.An(new_new_n104_), .B(new_new_n697_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n698_));
  NO3        g0676(.A(new_new_n468_), .B(new_new_n566_), .C(new_new_n590_), .Y(new_new_n699_));
  AOI220     g0677(.A0(new_new_n699_), .A1(new_new_n302_), .B0(new_new_n698_), .B1(new_new_n696_), .Y(new_new_n700_));
  NA3        g0678(.A(new_new_n700_), .B(new_new_n695_), .C(new_new_n694_), .Y(new_new_n701_));
  OAI210     g0679(.A0(new_new_n701_), .A1(new_new_n693_), .B0(new_new_n63_), .Y(new_new_n702_));
  NO2        g0680(.A(i_2_), .B(i_12_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n356_), .B(new_new_n703_), .Y(new_new_n704_));
  NA2        g0682(.A(i_8_), .B(new_new_n25_), .Y(new_new_n705_));
  NO3        g0683(.A(new_new_n705_), .B(new_new_n371_), .C(new_new_n585_), .Y(new_new_n706_));
  OAI210     g0684(.A0(new_new_n706_), .A1(new_new_n358_), .B0(new_new_n356_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n122_), .B(i_2_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n707_), .B(new_new_n704_), .Y(new_new_n709_));
  NA3        g0687(.A(new_new_n709_), .B(new_new_n46_), .C(new_new_n220_), .Y(new_new_n710_));
  NA4        g0688(.A(new_new_n710_), .B(new_new_n702_), .C(new_new_n690_), .D(new_new_n680_), .Y(new_new_n711_));
  OR4        g0689(.A(new_new_n711_), .B(new_new_n672_), .C(new_new_n657_), .D(new_new_n602_), .Y(men5));
  AOI210     g0690(.A0(new_new_n641_), .A1(new_new_n259_), .B0(new_new_n408_), .Y(new_new_n713_));
  AN2        g0691(.A(new_new_n24_), .B(i_10_), .Y(new_new_n714_));
  NA3        g0692(.A(new_new_n714_), .B(new_new_n703_), .C(new_new_n102_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n715_), .B(new_new_n713_), .Y(new_new_n716_));
  NO3        g0694(.A(i_11_), .B(new_new_n232_), .C(i_13_), .Y(new_new_n717_));
  NO2        g0695(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n718_));
  NA2        g0696(.A(i_12_), .B(i_8_), .Y(new_new_n719_));
  OAI210     g0697(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n719_), .Y(new_new_n720_));
  INV        g0698(.A(new_new_n435_), .Y(new_new_n721_));
  AOI220     g0699(.A0(new_new_n308_), .A1(new_new_n559_), .B0(new_new_n720_), .B1(new_new_n718_), .Y(new_new_n722_));
  INV        g0700(.A(new_new_n722_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n723_), .B(new_new_n716_), .Y(new_new_n724_));
  INV        g0702(.A(new_new_n166_), .Y(new_new_n725_));
  INV        g0703(.A(new_new_n239_), .Y(new_new_n726_));
  OAI210     g0704(.A0(new_new_n668_), .A1(new_new_n437_), .B0(new_new_n104_), .Y(new_new_n727_));
  AOI210     g0705(.A0(new_new_n727_), .A1(new_new_n726_), .B0(new_new_n725_), .Y(new_new_n728_));
  NO2        g0706(.A(new_new_n444_), .B(new_new_n26_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n729_), .B(new_new_n410_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n730_), .B(i_2_), .Y(new_new_n731_));
  INV        g0709(.A(new_new_n731_), .Y(new_new_n732_));
  AOI210     g0710(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n407_), .Y(new_new_n733_));
  AOI210     g0711(.A0(new_new_n733_), .A1(new_new_n732_), .B0(new_new_n728_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n184_), .B(new_new_n119_), .Y(new_new_n735_));
  OAI210     g0713(.A0(new_new_n735_), .A1(new_new_n718_), .B0(i_2_), .Y(new_new_n736_));
  NO2        g0714(.A(new_new_n736_), .B(new_new_n187_), .Y(new_new_n737_));
  OA210      g0715(.A0(new_new_n605_), .A1(new_new_n120_), .B0(i_13_), .Y(new_new_n738_));
  NA2        g0716(.A(new_new_n194_), .B(new_new_n197_), .Y(new_new_n739_));
  NA2        g0717(.A(new_new_n146_), .B(new_new_n582_), .Y(new_new_n740_));
  AOI210     g0718(.A0(new_new_n740_), .A1(new_new_n739_), .B0(new_new_n361_), .Y(new_new_n741_));
  AOI210     g0719(.A0(new_new_n203_), .A1(new_new_n142_), .B0(new_new_n506_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n742_), .B(new_new_n410_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n96_), .B(new_new_n45_), .Y(new_new_n744_));
  INV        g0722(.A(new_new_n291_), .Y(new_new_n745_));
  NA4        g0723(.A(new_new_n745_), .B(new_new_n295_), .C(new_new_n118_), .D(new_new_n43_), .Y(new_new_n746_));
  OAI210     g0724(.A0(new_new_n746_), .A1(new_new_n744_), .B0(new_new_n743_), .Y(new_new_n747_));
  NO4        g0725(.A(new_new_n747_), .B(new_new_n741_), .C(new_new_n738_), .D(new_new_n737_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n559_), .B(new_new_n28_), .Y(new_new_n749_));
  NA2        g0727(.A(new_new_n717_), .B(new_new_n265_), .Y(new_new_n750_));
  NA2        g0728(.A(new_new_n750_), .B(new_new_n749_), .Y(new_new_n751_));
  NO2        g0729(.A(new_new_n62_), .B(i_12_), .Y(new_new_n752_));
  NO2        g0730(.A(new_new_n752_), .B(new_new_n120_), .Y(new_new_n753_));
  NO2        g0731(.A(new_new_n753_), .B(new_new_n582_), .Y(new_new_n754_));
  AOI220     g0732(.A0(new_new_n754_), .A1(new_new_n36_), .B0(new_new_n751_), .B1(new_new_n47_), .Y(new_new_n755_));
  NA4        g0733(.A(new_new_n755_), .B(new_new_n748_), .C(new_new_n734_), .D(new_new_n724_), .Y(men6));
  NA2        g0734(.A(new_new_n25_), .B(new_new_n708_), .Y(new_new_n757_));
  NA4        g0735(.A(new_new_n377_), .B(new_new_n473_), .C(new_new_n69_), .D(new_new_n95_), .Y(new_new_n758_));
  INV        g0736(.A(new_new_n758_), .Y(new_new_n759_));
  NO2        g0737(.A(i_11_), .B(i_9_), .Y(new_new_n760_));
  NO2        g0738(.A(new_new_n759_), .B(new_new_n319_), .Y(new_new_n761_));
  AO210      g0739(.A0(new_new_n761_), .A1(new_new_n757_), .B0(i_12_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n362_), .B(new_new_n325_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n566_), .B(new_new_n63_), .Y(new_new_n764_));
  INV        g0742(.A(new_new_n659_), .Y(new_new_n765_));
  NA4        g0743(.A(new_new_n84_), .B(new_new_n765_), .C(new_new_n764_), .D(new_new_n763_), .Y(new_new_n766_));
  INV        g0744(.A(new_new_n191_), .Y(new_new_n767_));
  AOI220     g0745(.A0(new_new_n767_), .A1(new_new_n760_), .B0(new_new_n766_), .B1(new_new_n71_), .Y(new_new_n768_));
  NO2        g0746(.A(new_new_n246_), .B(i_9_), .Y(new_new_n769_));
  NA2        g0747(.A(new_new_n769_), .B(new_new_n752_), .Y(new_new_n770_));
  AOI210     g0748(.A0(new_new_n770_), .A1(new_new_n505_), .B0(new_new_n179_), .Y(new_new_n771_));
  NA3        g0749(.A(new_new_n1022_), .B(new_new_n464_), .C(new_new_n377_), .Y(new_new_n772_));
  NAi32      g0750(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n691_), .A1(new_new_n84_), .B0(new_new_n773_), .Y(new_new_n774_));
  OAI210     g0752(.A0(new_new_n658_), .A1(new_new_n547_), .B0(new_new_n546_), .Y(new_new_n775_));
  NAi31      g0753(.An(new_new_n774_), .B(new_new_n775_), .C(new_new_n772_), .Y(new_new_n776_));
  OR2        g0754(.A(new_new_n776_), .B(new_new_n771_), .Y(new_new_n777_));
  NO2        g0755(.A(i_11_), .B(i_2_), .Y(new_new_n778_));
  NA2        g0756(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n779_), .B(new_new_n399_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n780_), .B(new_new_n778_), .Y(new_new_n781_));
  NA3        g0759(.A(new_new_n339_), .B(new_new_n248_), .C(i_7_), .Y(new_new_n782_));
  BUFFER     g0760(.A(new_new_n605_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(new_new_n141_), .Y(new_new_n784_));
  OR2        g0762(.A(new_new_n721_), .B(new_new_n36_), .Y(new_new_n785_));
  NA4        g0763(.A(new_new_n785_), .B(new_new_n784_), .C(new_new_n782_), .D(new_new_n781_), .Y(new_new_n786_));
  NA2        g0764(.A(new_new_n384_), .B(new_new_n68_), .Y(new_new_n787_));
  NA2        g0765(.A(new_new_n787_), .B(new_new_n588_), .Y(new_new_n788_));
  NA3        g0766(.A(new_new_n506_), .B(new_new_n474_), .C(new_new_n214_), .Y(new_new_n789_));
  INV        g0767(.A(new_new_n545_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n105_), .B(new_new_n398_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n238_), .B(new_new_n47_), .Y(new_new_n792_));
  INV        g0770(.A(new_new_n573_), .Y(new_new_n793_));
  NA3        g0771(.A(new_new_n793_), .B(new_new_n318_), .C(i_7_), .Y(new_new_n794_));
  NA4        g0772(.A(new_new_n794_), .B(new_new_n791_), .C(new_new_n790_), .D(new_new_n789_), .Y(new_new_n795_));
  NO4        g0773(.A(new_new_n795_), .B(new_new_n788_), .C(new_new_n786_), .D(new_new_n777_), .Y(new_new_n796_));
  NA4        g0774(.A(new_new_n796_), .B(new_new_n768_), .C(new_new_n762_), .D(new_new_n367_), .Y(men3));
  NA2        g0775(.A(i_12_), .B(i_10_), .Y(new_new_n798_));
  NA2        g0776(.A(i_6_), .B(i_7_), .Y(new_new_n799_));
  NO2        g0777(.A(new_new_n799_), .B(i_0_), .Y(new_new_n800_));
  NO2        g0778(.A(i_11_), .B(new_new_n232_), .Y(new_new_n801_));
  OAI210     g0779(.A0(new_new_n800_), .A1(new_new_n279_), .B0(new_new_n801_), .Y(new_new_n802_));
  NO2        g0780(.A(new_new_n802_), .B(new_new_n187_), .Y(new_new_n803_));
  NO3        g0781(.A(new_new_n440_), .B(new_new_n86_), .C(new_new_n45_), .Y(new_new_n804_));
  OA210      g0782(.A0(new_new_n804_), .A1(new_new_n803_), .B0(new_new_n168_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n588_), .B(new_new_n360_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n806_), .B(new_new_n40_), .Y(new_new_n807_));
  NO3        g0785(.A(new_new_n612_), .B(new_new_n444_), .C(new_new_n125_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n400_), .B(new_new_n46_), .Y(new_new_n809_));
  AOI210     g0787(.A0(new_new_n1018_), .A1(new_new_n807_), .B0(new_new_n49_), .Y(new_new_n810_));
  NA2        g0788(.A(new_new_n179_), .B(new_new_n555_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n683_), .B(new_new_n651_), .Y(new_new_n812_));
  NA2        g0790(.A(i_0_), .B(new_new_n427_), .Y(new_new_n813_));
  OAI220     g0791(.A0(new_new_n813_), .A1(new_new_n812_), .B0(new_new_n811_), .B1(new_new_n63_), .Y(new_new_n814_));
  NOi21      g0792(.An(i_5_), .B(i_9_), .Y(new_new_n815_));
  NA2        g0793(.A(new_new_n815_), .B(new_new_n434_), .Y(new_new_n816_));
  AOI210     g0794(.A0(new_new_n256_), .A1(new_new_n466_), .B0(new_new_n662_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n169_), .B(new_new_n142_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n818_), .B(new_new_n238_), .Y(new_new_n819_));
  OAI220     g0797(.A0(new_new_n819_), .A1(new_new_n174_), .B0(new_new_n817_), .B1(new_new_n816_), .Y(new_new_n820_));
  NO4        g0798(.A(new_new_n820_), .B(new_new_n814_), .C(new_new_n810_), .D(new_new_n805_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n179_), .B(new_new_n24_), .Y(new_new_n822_));
  NO2        g0800(.A(new_new_n649_), .B(new_new_n579_), .Y(new_new_n823_));
  NO2        g0801(.A(new_new_n823_), .B(new_new_n822_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n302_), .B(new_new_n123_), .Y(new_new_n825_));
  NAi21      g0803(.An(new_new_n157_), .B(new_new_n427_), .Y(new_new_n826_));
  OAI220     g0804(.A0(new_new_n826_), .A1(new_new_n792_), .B0(new_new_n825_), .B1(new_new_n389_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n827_), .B(new_new_n824_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n556_), .B(i_0_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n829_), .B(new_new_n372_), .Y(new_new_n830_));
  NO4        g0808(.A(new_new_n572_), .B(new_new_n211_), .C(new_new_n407_), .D(new_new_n399_), .Y(new_new_n831_));
  AOI210     g0809(.A0(new_new_n831_), .A1(i_11_), .B0(new_new_n830_), .Y(new_new_n832_));
  NA2        g0810(.A(new_new_n717_), .B(new_new_n319_), .Y(new_new_n833_));
  INV        g0811(.A(new_new_n58_), .Y(new_new_n834_));
  OAI220     g0812(.A0(new_new_n834_), .A1(new_new_n833_), .B0(new_new_n636_), .B1(new_new_n522_), .Y(new_new_n835_));
  NA2        g0813(.A(i_0_), .B(i_10_), .Y(new_new_n836_));
  OAI210     g0814(.A0(new_new_n836_), .A1(new_new_n83_), .B0(new_new_n523_), .Y(new_new_n837_));
  NO4        g0815(.A(new_new_n108_), .B(new_new_n58_), .C(new_new_n646_), .D(i_5_), .Y(new_new_n838_));
  AN2        g0816(.A(new_new_n838_), .B(new_new_n837_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n179_), .B(new_new_n82_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n550_), .B(i_4_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n182_), .B(new_new_n197_), .Y(new_new_n842_));
  OAI220     g0820(.A0(new_new_n842_), .A1(new_new_n833_), .B0(new_new_n841_), .B1(new_new_n840_), .Y(new_new_n843_));
  NO3        g0821(.A(new_new_n843_), .B(new_new_n839_), .C(new_new_n835_), .Y(new_new_n844_));
  NA3        g0822(.A(new_new_n844_), .B(new_new_n832_), .C(new_new_n828_), .Y(new_new_n845_));
  NO2        g0823(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n846_));
  NA2        g0824(.A(i_11_), .B(i_9_), .Y(new_new_n847_));
  NO3        g0825(.A(i_12_), .B(new_new_n847_), .C(new_new_n587_), .Y(new_new_n848_));
  AN2        g0826(.A(new_new_n848_), .B(new_new_n846_), .Y(new_new_n849_));
  NO2        g0827(.A(new_new_n49_), .B(i_7_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n381_), .B(new_new_n173_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n851_), .B(new_new_n155_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n847_), .B(new_new_n71_), .Y(new_new_n853_));
  NO2        g0831(.A(new_new_n169_), .B(i_0_), .Y(new_new_n854_));
  INV        g0832(.A(new_new_n854_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n464_), .B(new_new_n226_), .Y(new_new_n856_));
  AOI210     g0834(.A0(new_new_n359_), .A1(new_new_n42_), .B0(new_new_n397_), .Y(new_new_n857_));
  OAI220     g0835(.A0(new_new_n857_), .A1(new_new_n816_), .B0(new_new_n856_), .B1(new_new_n855_), .Y(new_new_n858_));
  NO3        g0836(.A(new_new_n858_), .B(new_new_n852_), .C(new_new_n849_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n635_), .B(new_new_n115_), .Y(new_new_n860_));
  NO2        g0838(.A(i_6_), .B(new_new_n860_), .Y(new_new_n861_));
  AOI210     g0839(.A0(new_new_n436_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n166_), .B(new_new_n97_), .Y(new_new_n863_));
  NOi32      g0841(.An(new_new_n862_), .Bn(new_new_n182_), .C(new_new_n863_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n589_), .B(new_new_n319_), .Y(new_new_n865_));
  NO2        g0843(.A(new_new_n865_), .B(new_new_n809_), .Y(new_new_n866_));
  NO3        g0844(.A(new_new_n866_), .B(new_new_n864_), .C(new_new_n861_), .Y(new_new_n867_));
  NOi21      g0845(.An(i_7_), .B(i_5_), .Y(new_new_n868_));
  NOi31      g0846(.An(new_new_n868_), .B(i_0_), .C(new_new_n697_), .Y(new_new_n869_));
  NA3        g0847(.A(new_new_n869_), .B(new_new_n371_), .C(i_6_), .Y(new_new_n870_));
  OA210      g0848(.A0(new_new_n863_), .A1(new_new_n505_), .B0(new_new_n870_), .Y(new_new_n871_));
  NO3        g0849(.A(new_new_n392_), .B(new_new_n348_), .C(new_new_n346_), .Y(new_new_n872_));
  NO2        g0850(.A(new_new_n250_), .B(new_new_n309_), .Y(new_new_n873_));
  NO2        g0851(.A(new_new_n697_), .B(new_new_n249_), .Y(new_new_n874_));
  AOI210     g0852(.A0(new_new_n874_), .A1(new_new_n873_), .B0(new_new_n872_), .Y(new_new_n875_));
  NA4        g0853(.A(new_new_n875_), .B(new_new_n871_), .C(new_new_n867_), .D(new_new_n859_), .Y(new_new_n876_));
  NO2        g0854(.A(new_new_n822_), .B(new_new_n234_), .Y(new_new_n877_));
  AN2        g0855(.A(new_new_n323_), .B(new_new_n319_), .Y(new_new_n878_));
  AN2        g0856(.A(new_new_n878_), .B(new_new_n818_), .Y(new_new_n879_));
  OAI210     g0857(.A0(new_new_n879_), .A1(new_new_n877_), .B0(i_10_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n798_), .B(new_new_n308_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n881_), .B(new_new_n853_), .Y(new_new_n882_));
  NA3        g0860(.A(new_new_n463_), .B(new_new_n400_), .C(new_new_n46_), .Y(new_new_n883_));
  OAI210     g0861(.A0(new_new_n826_), .A1(i_7_), .B0(new_new_n883_), .Y(new_new_n884_));
  NO2        g0862(.A(new_new_n248_), .B(new_new_n47_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n853_), .B(new_new_n295_), .Y(new_new_n886_));
  OAI210     g0864(.A0(new_new_n885_), .A1(new_new_n181_), .B0(new_new_n886_), .Y(new_new_n887_));
  AOI220     g0865(.A0(new_new_n887_), .A1(new_new_n464_), .B0(new_new_n884_), .B1(new_new_n71_), .Y(new_new_n888_));
  NO2        g0866(.A(new_new_n73_), .B(new_new_n719_), .Y(new_new_n889_));
  AOI210     g0867(.A0(new_new_n168_), .A1(new_new_n579_), .B0(new_new_n889_), .Y(new_new_n890_));
  NO2        g0868(.A(new_new_n890_), .B(new_new_n48_), .Y(new_new_n891_));
  NO3        g0869(.A(new_new_n572_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n892_));
  AOI210     g0870(.A0(new_new_n677_), .A1(new_new_n531_), .B0(new_new_n892_), .Y(new_new_n893_));
  NAi21      g0871(.An(i_9_), .B(i_5_), .Y(new_new_n894_));
  NO2        g0872(.A(new_new_n894_), .B(new_new_n392_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n584_), .B(new_new_n99_), .Y(new_new_n896_));
  AOI220     g0874(.A0(new_new_n896_), .A1(i_0_), .B0(new_new_n895_), .B1(new_new_n605_), .Y(new_new_n897_));
  OAI220     g0875(.A0(new_new_n897_), .A1(new_new_n83_), .B0(new_new_n893_), .B1(new_new_n167_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n898_), .B(new_new_n891_), .Y(new_new_n899_));
  NA4        g0877(.A(new_new_n899_), .B(new_new_n888_), .C(new_new_n882_), .D(new_new_n880_), .Y(new_new_n900_));
  NO3        g0878(.A(new_new_n900_), .B(new_new_n876_), .C(new_new_n845_), .Y(new_new_n901_));
  NO2        g0879(.A(i_0_), .B(new_new_n697_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n71_), .B(new_new_n45_), .Y(new_new_n903_));
  NO3        g0881(.A(new_new_n99_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n904_));
  AO220      g0882(.A0(new_new_n904_), .A1(new_new_n45_), .B0(new_new_n902_), .B1(new_new_n168_), .Y(new_new_n905_));
  NO2        g0883(.A(new_new_n764_), .B(new_new_n863_), .Y(new_new_n906_));
  AOI210     g0884(.A0(new_new_n905_), .A1(new_new_n336_), .B0(new_new_n906_), .Y(new_new_n907_));
  NA2        g0885(.A(new_new_n708_), .B(new_new_n140_), .Y(new_new_n908_));
  INV        g0886(.A(new_new_n908_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n909_), .B(new_new_n651_), .Y(new_new_n910_));
  NO2        g0888(.A(new_new_n775_), .B(new_new_n392_), .Y(new_new_n911_));
  NA3        g0889(.A(new_new_n800_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n912_));
  NA2        g0890(.A(new_new_n801_), .B(i_9_), .Y(new_new_n913_));
  AOI210     g0891(.A0(new_new_n912_), .A1(new_new_n488_), .B0(new_new_n913_), .Y(new_new_n914_));
  OAI210     g0892(.A0(new_new_n238_), .A1(i_9_), .B0(new_new_n225_), .Y(new_new_n915_));
  AOI210     g0893(.A0(new_new_n915_), .A1(new_new_n829_), .B0(new_new_n148_), .Y(new_new_n916_));
  NO3        g0894(.A(new_new_n916_), .B(new_new_n914_), .C(new_new_n911_), .Y(new_new_n917_));
  NA3        g0895(.A(new_new_n917_), .B(new_new_n910_), .C(new_new_n907_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n878_), .B(new_new_n361_), .Y(new_new_n919_));
  AOI210     g0897(.A0(new_new_n290_), .A1(new_new_n157_), .B0(new_new_n919_), .Y(new_new_n920_));
  NA3        g0898(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n850_), .B(new_new_n478_), .Y(new_new_n922_));
  AOI210     g0900(.A0(new_new_n921_), .A1(new_new_n157_), .B0(new_new_n922_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n923_), .B(new_new_n920_), .Y(new_new_n924_));
  NO3        g0902(.A(new_new_n836_), .B(new_new_n815_), .C(new_new_n184_), .Y(new_new_n925_));
  AOI220     g0903(.A0(new_new_n925_), .A1(i_11_), .B0(new_new_n551_), .B1(new_new_n73_), .Y(new_new_n926_));
  NO3        g0904(.A(new_new_n205_), .B(new_new_n370_), .C(i_0_), .Y(new_new_n927_));
  OAI210     g0905(.A0(new_new_n927_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n928_));
  INV        g0906(.A(new_new_n214_), .Y(new_new_n929_));
  NO2        g0907(.A(i_12_), .B(new_new_n599_), .Y(new_new_n930_));
  NA3        g0908(.A(new_new_n930_), .B(new_new_n1021_), .C(new_new_n929_), .Y(new_new_n931_));
  NA4        g0909(.A(new_new_n931_), .B(new_new_n928_), .C(new_new_n926_), .D(new_new_n924_), .Y(new_new_n932_));
  NO2        g0910(.A(new_new_n237_), .B(new_new_n88_), .Y(new_new_n933_));
  NA2        g0911(.A(new_new_n933_), .B(new_new_n902_), .Y(new_new_n934_));
  AOI220     g0912(.A0(new_new_n868_), .A1(new_new_n478_), .B0(new_new_n800_), .B1(new_new_n158_), .Y(new_new_n935_));
  NA2        g0913(.A(new_new_n339_), .B(new_new_n170_), .Y(new_new_n936_));
  OA220      g0914(.A0(new_new_n936_), .A1(new_new_n935_), .B0(new_new_n934_), .B1(i_5_), .Y(new_new_n937_));
  AOI210     g0915(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n938_));
  NA3        g0916(.A(new_new_n596_), .B(new_new_n179_), .C(new_new_n82_), .Y(new_new_n939_));
  NA2        g0917(.A(new_new_n939_), .B(new_new_n530_), .Y(new_new_n940_));
  NO3        g0918(.A(new_new_n809_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n941_));
  NA3        g0919(.A(new_new_n482_), .B(new_new_n477_), .C(new_new_n461_), .Y(new_new_n942_));
  NO3        g0920(.A(new_new_n942_), .B(new_new_n941_), .C(new_new_n940_), .Y(new_new_n943_));
  NA3        g0921(.A(new_new_n377_), .B(new_new_n166_), .C(new_new_n165_), .Y(new_new_n944_));
  NA3        g0922(.A(new_new_n850_), .B(new_new_n279_), .C(new_new_n225_), .Y(new_new_n945_));
  NA2        g0923(.A(new_new_n945_), .B(new_new_n944_), .Y(new_new_n946_));
  NA3        g0924(.A(new_new_n377_), .B(new_new_n324_), .C(new_new_n217_), .Y(new_new_n947_));
  INV        g0925(.A(new_new_n947_), .Y(new_new_n948_));
  NOi31      g0926(.An(new_new_n376_), .B(new_new_n903_), .C(new_new_n234_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n847_), .B(new_new_n214_), .C(new_new_n184_), .Y(new_new_n950_));
  NO4        g0928(.A(new_new_n950_), .B(new_new_n949_), .C(new_new_n948_), .D(new_new_n946_), .Y(new_new_n951_));
  NA3        g0929(.A(new_new_n951_), .B(new_new_n943_), .C(new_new_n937_), .Y(new_new_n952_));
  INV        g0930(.A(new_new_n598_), .Y(new_new_n953_));
  NO3        g0931(.A(new_new_n953_), .B(new_new_n541_), .C(i_3_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n83_), .B(i_5_), .Y(new_new_n955_));
  NA3        g0933(.A(new_new_n801_), .B(new_new_n103_), .C(new_new_n118_), .Y(new_new_n956_));
  INV        g0934(.A(new_new_n956_), .Y(new_new_n957_));
  AOI210     g0935(.A0(new_new_n957_), .A1(new_new_n955_), .B0(new_new_n954_), .Y(new_new_n958_));
  NA3        g0936(.A(new_new_n295_), .B(i_5_), .C(new_new_n187_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n959_), .B(new_new_n237_), .Y(new_new_n960_));
  NO4        g0938(.A(new_new_n234_), .B(new_new_n205_), .C(i_0_), .D(i_12_), .Y(new_new_n961_));
  AOI220     g0939(.A0(new_new_n961_), .A1(new_new_n960_), .B0(new_new_n759_), .B1(new_new_n170_), .Y(new_new_n962_));
  AN2        g0940(.A(new_new_n836_), .B(new_new_n148_), .Y(new_new_n963_));
  NO4        g0941(.A(new_new_n963_), .B(i_12_), .C(new_new_n626_), .D(new_new_n125_), .Y(new_new_n964_));
  NA2        g0942(.A(new_new_n964_), .B(new_new_n214_), .Y(new_new_n965_));
  NA3        g0943(.A(new_new_n92_), .B(new_new_n555_), .C(i_11_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n966_), .B(new_new_n150_), .Y(new_new_n967_));
  NA2        g0945(.A(new_new_n868_), .B(new_new_n460_), .Y(new_new_n968_));
  OAI220     g0946(.A0(i_7_), .A1(new_new_n959_), .B0(new_new_n968_), .B1(new_new_n652_), .Y(new_new_n969_));
  AOI210     g0947(.A0(new_new_n969_), .A1(new_new_n854_), .B0(new_new_n967_), .Y(new_new_n970_));
  NA4        g0948(.A(new_new_n970_), .B(new_new_n965_), .C(new_new_n962_), .D(new_new_n958_), .Y(new_new_n971_));
  NO4        g0949(.A(new_new_n971_), .B(new_new_n952_), .C(new_new_n932_), .D(new_new_n918_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n862_), .B(new_new_n356_), .C(i_5_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n973_), .B(new_new_n594_), .Y(new_new_n974_));
  NA2        g0952(.A(new_new_n974_), .B(new_new_n201_), .Y(new_new_n975_));
  NA2        g0953(.A(new_new_n180_), .B(new_new_n182_), .Y(new_new_n976_));
  AO210      g0954(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n976_), .Y(new_new_n977_));
  OAI210     g0955(.A0(new_new_n598_), .A1(new_new_n596_), .B0(new_new_n308_), .Y(new_new_n978_));
  NA2        g0956(.A(new_new_n978_), .B(new_new_n977_), .Y(new_new_n979_));
  NO4        g0957(.A(new_new_n228_), .B(new_new_n139_), .C(new_new_n655_), .D(new_new_n37_), .Y(new_new_n980_));
  NO2        g0958(.A(new_new_n980_), .B(new_new_n831_), .Y(new_new_n981_));
  OAI210     g0959(.A0(new_new_n966_), .A1(new_new_n142_), .B0(new_new_n981_), .Y(new_new_n982_));
  AOI210     g0960(.A0(new_new_n979_), .A1(new_new_n49_), .B0(new_new_n982_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n983_), .A1(new_new_n975_), .B0(new_new_n71_), .Y(new_new_n984_));
  NO2        g0962(.A(new_new_n548_), .B(new_new_n366_), .Y(new_new_n985_));
  NO2        g0963(.A(new_new_n985_), .B(new_new_n725_), .Y(new_new_n986_));
  INV        g0964(.A(new_new_n74_), .Y(new_new_n987_));
  AOI210     g0965(.A0(new_new_n938_), .A1(new_new_n850_), .B0(new_new_n869_), .Y(new_new_n988_));
  AOI210     g0966(.A0(new_new_n988_), .A1(new_new_n987_), .B0(new_new_n655_), .Y(new_new_n989_));
  NA2        g0967(.A(i_8_), .B(new_new_n74_), .Y(new_new_n990_));
  NO2        g0968(.A(new_new_n990_), .B(new_new_n232_), .Y(new_new_n991_));
  NA3        g0969(.A(new_new_n90_), .B(new_new_n297_), .C(new_new_n31_), .Y(new_new_n992_));
  INV        g0970(.A(new_new_n992_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n993_), .B(new_new_n991_), .C(new_new_n989_), .Y(new_new_n994_));
  OAI210     g0972(.A0(new_new_n258_), .A1(new_new_n153_), .B0(new_new_n85_), .Y(new_new_n995_));
  NA3        g0973(.A(new_new_n729_), .B(new_new_n279_), .C(new_new_n78_), .Y(new_new_n996_));
  AOI210     g0974(.A0(new_new_n996_), .A1(new_new_n995_), .B0(i_11_), .Y(new_new_n997_));
  NA2        g0975(.A(new_new_n590_), .B(new_new_n211_), .Y(new_new_n998_));
  OAI210     g0976(.A0(new_new_n998_), .A1(new_new_n862_), .B0(new_new_n201_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n159_), .B(i_5_), .Y(new_new_n1000_));
  NO2        g0978(.A(new_new_n999_), .B(new_new_n1000_), .Y(new_new_n1001_));
  NO3        g0979(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1002_));
  OAI210     g0980(.A0(new_new_n873_), .A1(new_new_n297_), .B0(new_new_n1002_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n1003_), .B(new_new_n697_), .Y(new_new_n1004_));
  NO3        g0982(.A(new_new_n894_), .B(new_new_n467_), .C(new_new_n247_), .Y(new_new_n1005_));
  NO2        g0983(.A(new_new_n1005_), .B(new_new_n545_), .Y(new_new_n1006_));
  INV        g0984(.A(new_new_n349_), .Y(new_new_n1007_));
  AOI210     g0985(.A0(new_new_n1007_), .A1(new_new_n1006_), .B0(new_new_n41_), .Y(new_new_n1008_));
  NO4        g0986(.A(new_new_n1008_), .B(new_new_n1004_), .C(new_new_n1001_), .D(new_new_n997_), .Y(new_new_n1009_));
  OAI210     g0987(.A0(new_new_n994_), .A1(i_4_), .B0(new_new_n1009_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n1010_), .B(new_new_n986_), .C(new_new_n984_), .Y(new_new_n1011_));
  NA4        g0989(.A(new_new_n1011_), .B(new_new_n972_), .C(new_new_n901_), .D(new_new_n821_), .Y(men4));
  INV        g0990(.A(new_new_n676_), .Y(new_new_n1015_));
  INV        g0991(.A(i_2_), .Y(new_new_n1016_));
  INV        g0992(.A(new_new_n687_), .Y(new_new_n1017_));
  INV        g0993(.A(new_new_n808_), .Y(new_new_n1018_));
  INV        g0994(.A(new_new_n80_), .Y(new_new_n1019_));
  INV        g0995(.A(new_new_n138_), .Y(new_new_n1020_));
  INV        g0996(.A(i_3_), .Y(new_new_n1021_));
  INV        g0997(.A(i_11_), .Y(new_new_n1022_));
  INV        g0998(.A(new_new_n138_), .Y(new_new_n1023_));
  INV        g0999(.A(new_new_n237_), .Y(new_new_n1024_));
  INV        g1000(.A(i_8_), .Y(new_new_n1025_));
endmodule


