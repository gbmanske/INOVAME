// Benchmark "top" written by ABC on Thu Jun 20 14:59:10 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n137_, new_new_n138_, new_new_n139_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1107_, new_new_n1108_,
    new_new_n1109_, new_new_n1113_, new_new_n1114_, new_new_n1115_,
    new_new_n1116_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g0028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g0029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g0030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA3        g0031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g0032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g0033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  INV        g0034(.A(new_new_n54_), .Y(new_new_n57_));
  NA2        g0035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g0036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g0037(.A(i_1_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g0039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g0040(.A(new_new_n62_), .B(new_new_n58_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n50_), .B(i_2_), .Y(new_new_n64_));
  AOI210     g0042(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_6_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(new_new_n25_), .Y(new_new_n67_));
  INV        g0045(.A(i_0_), .Y(new_new_n68_));
  NAi21      g0046(.An(i_5_), .B(i_10_), .Y(new_new_n69_));
  NA2        g0047(.A(i_5_), .B(i_9_), .Y(new_new_n70_));
  AOI210     g0048(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n68_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n67_), .Y(new_new_n72_));
  OAI210     g0050(.A0(new_new_n65_), .A1(new_new_n64_), .B0(new_new_n72_), .Y(new_new_n73_));
  OAI210     g0051(.A0(new_new_n73_), .A1(new_new_n63_), .B0(i_0_), .Y(new_new_n74_));
  NA2        g0052(.A(i_12_), .B(i_5_), .Y(new_new_n75_));
  NA2        g0053(.A(i_2_), .B(i_8_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n55_), .Y(new_new_n77_));
  NO2        g0055(.A(i_3_), .B(i_9_), .Y(new_new_n78_));
  NO2        g0056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  NO3        g0057(.A(new_new_n79_), .B(new_new_n78_), .C(new_new_n60_), .Y(new_new_n80_));
  INV        g0058(.A(i_6_), .Y(new_new_n81_));
  OR4        g0059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n82_));
  INV        g0060(.A(new_new_n82_), .Y(new_new_n83_));
  NO2        g0061(.A(i_2_), .B(i_7_), .Y(new_new_n84_));
  AOI210     g0062(.A0(new_new_n83_), .A1(new_new_n81_), .B0(new_new_n84_), .Y(new_new_n85_));
  OAI210     g0063(.A0(new_new_n80_), .A1(new_new_n77_), .B0(new_new_n85_), .Y(new_new_n86_));
  NAi21      g0064(.An(i_6_), .B(i_10_), .Y(new_new_n87_));
  NA2        g0065(.A(i_6_), .B(i_9_), .Y(new_new_n88_));
  AOI210     g0066(.A0(new_new_n88_), .A1(new_new_n87_), .B0(new_new_n60_), .Y(new_new_n89_));
  NA2        g0067(.A(i_2_), .B(i_6_), .Y(new_new_n90_));
  NO3        g0068(.A(new_new_n90_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n91_));
  NO2        g0069(.A(new_new_n91_), .B(new_new_n89_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n86_), .B0(new_new_n75_), .Y(new_new_n93_));
  AN3        g0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g0072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NO2        g0073(.A(i_5_), .B(i_8_), .Y(new_new_n96_));
  NOi21      g0074(.An(new_new_n96_), .B(new_new_n95_), .Y(new_new_n97_));
  AOI220     g0075(.A0(new_new_n97_), .A1(new_new_n59_), .B0(new_new_n94_), .B1(new_new_n32_), .Y(new_new_n98_));
  INV        g0076(.A(i_7_), .Y(new_new_n99_));
  NA2        g0077(.A(new_new_n46_), .B(new_new_n99_), .Y(new_new_n100_));
  NO2        g0078(.A(i_0_), .B(i_5_), .Y(new_new_n101_));
  NO2        g0079(.A(new_new_n101_), .B(new_new_n81_), .Y(new_new_n102_));
  NA2        g0080(.A(i_12_), .B(i_3_), .Y(new_new_n103_));
  INV        g0081(.A(new_new_n103_), .Y(new_new_n104_));
  NA3        g0082(.A(new_new_n104_), .B(new_new_n102_), .C(new_new_n100_), .Y(new_new_n105_));
  NAi21      g0083(.An(i_7_), .B(i_11_), .Y(new_new_n106_));
  NO3        g0084(.A(new_new_n106_), .B(new_new_n87_), .C(new_new_n51_), .Y(new_new_n107_));
  AN2        g0085(.A(i_2_), .B(i_10_), .Y(new_new_n108_));
  NO2        g0086(.A(new_new_n108_), .B(i_7_), .Y(new_new_n109_));
  OR2        g0087(.A(new_new_n75_), .B(new_new_n55_), .Y(new_new_n110_));
  NO2        g0088(.A(i_8_), .B(new_new_n99_), .Y(new_new_n111_));
  NO3        g0089(.A(new_new_n111_), .B(new_new_n110_), .C(new_new_n109_), .Y(new_new_n112_));
  NA2        g0090(.A(i_12_), .B(i_7_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n60_), .B(new_new_n26_), .Y(new_new_n114_));
  NA2        g0092(.A(new_new_n114_), .B(i_0_), .Y(new_new_n115_));
  NA2        g0093(.A(i_11_), .B(i_12_), .Y(new_new_n116_));
  OAI210     g0094(.A0(new_new_n115_), .A1(new_new_n113_), .B0(new_new_n116_), .Y(new_new_n117_));
  NO2        g0095(.A(new_new_n117_), .B(new_new_n112_), .Y(new_new_n118_));
  NAi41      g0096(.An(new_new_n107_), .B(new_new_n118_), .C(new_new_n105_), .D(new_new_n98_), .Y(new_new_n119_));
  NOi21      g0097(.An(i_1_), .B(i_5_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n120_), .B(i_11_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n122_));
  NA2        g0100(.A(i_7_), .B(new_new_n25_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(new_new_n122_), .Y(new_new_n124_));
  NO2        g0102(.A(new_new_n124_), .B(new_new_n46_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n88_), .B(new_new_n87_), .Y(new_new_n126_));
  NAi21      g0104(.An(i_3_), .B(i_8_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n59_), .Y(new_new_n128_));
  NOi21      g0106(.An(new_new_n128_), .B(new_new_n126_), .Y(new_new_n129_));
  NO2        g0107(.A(i_1_), .B(new_new_n81_), .Y(new_new_n130_));
  NO2        g0108(.A(i_6_), .B(i_5_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(i_3_), .Y(new_new_n132_));
  AO210      g0110(.A0(new_new_n132_), .A1(new_new_n47_), .B0(new_new_n130_), .Y(new_new_n133_));
  OAI220     g0111(.A0(new_new_n133_), .A1(new_new_n106_), .B0(new_new_n129_), .B1(new_new_n121_), .Y(new_new_n134_));
  NO3        g0112(.A(new_new_n134_), .B(new_new_n119_), .C(new_new_n93_), .Y(new_new_n135_));
  NA2        g0113(.A(new_new_n135_), .B(new_new_n74_), .Y(men2));
  NO2        g0114(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n137_));
  NA2        g0115(.A(i_6_), .B(new_new_n25_), .Y(new_new_n138_));
  NA2        g0116(.A(new_new_n138_), .B(new_new_n137_), .Y(new_new_n139_));
  NA4        g0117(.A(new_new_n139_), .B(new_new_n72_), .C(new_new_n64_), .D(new_new_n30_), .Y(men0));
  AN2        g0118(.A(i_8_), .B(i_7_), .Y(new_new_n141_));
  NA2        g0119(.A(new_new_n141_), .B(i_6_), .Y(new_new_n142_));
  NO2        g0120(.A(i_12_), .B(i_13_), .Y(new_new_n143_));
  NAi21      g0121(.An(i_5_), .B(i_11_), .Y(new_new_n144_));
  NOi21      g0122(.An(new_new_n143_), .B(new_new_n144_), .Y(new_new_n145_));
  NO2        g0123(.A(i_0_), .B(i_1_), .Y(new_new_n146_));
  NA2        g0124(.A(i_2_), .B(i_3_), .Y(new_new_n147_));
  NO2        g0125(.A(new_new_n147_), .B(i_4_), .Y(new_new_n148_));
  NA3        g0126(.A(new_new_n148_), .B(new_new_n146_), .C(new_new_n145_), .Y(new_new_n149_));
  OR2        g0127(.A(new_new_n149_), .B(new_new_n25_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n143_), .B(new_new_n78_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(new_new_n27_), .Y(new_new_n152_));
  NA2        g0130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n68_), .B(new_new_n46_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n36_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n75_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n39_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n68_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  NO2        g0144(.A(new_new_n166_), .B(new_new_n156_), .Y(new_new_n167_));
  AOI210     g0145(.A0(new_new_n167_), .A1(new_new_n150_), .B0(new_new_n142_), .Y(new_new_n168_));
  NA3        g0146(.A(new_new_n68_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n169_));
  NOi21      g0147(.An(i_4_), .B(i_9_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_11_), .B(i_13_), .Y(new_new_n171_));
  NA2        g0149(.A(new_new_n171_), .B(new_new_n170_), .Y(new_new_n172_));
  NO2        g0150(.A(i_4_), .B(i_5_), .Y(new_new_n173_));
  NAi21      g0151(.An(i_12_), .B(i_11_), .Y(new_new_n174_));
  NO2        g0152(.A(new_new_n174_), .B(i_13_), .Y(new_new_n175_));
  NA3        g0153(.A(new_new_n175_), .B(new_new_n173_), .C(new_new_n78_), .Y(new_new_n176_));
  AOI210     g0154(.A0(new_new_n176_), .A1(new_new_n172_), .B0(new_new_n169_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n68_), .B(new_new_n60_), .Y(new_new_n178_));
  NA2        g0156(.A(new_new_n178_), .B(new_new_n46_), .Y(new_new_n179_));
  NA2        g0157(.A(new_new_n36_), .B(i_5_), .Y(new_new_n180_));
  NAi31      g0158(.An(new_new_n180_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n181_));
  NA2        g0159(.A(i_3_), .B(i_5_), .Y(new_new_n182_));
  OR2        g0160(.A(new_new_n182_), .B(new_new_n172_), .Y(new_new_n183_));
  AOI210     g0161(.A0(new_new_n183_), .A1(new_new_n181_), .B0(new_new_n179_), .Y(new_new_n184_));
  NO2        g0162(.A(new_new_n68_), .B(i_5_), .Y(new_new_n185_));
  NO2        g0163(.A(i_13_), .B(i_10_), .Y(new_new_n186_));
  NA3        g0164(.A(new_new_n186_), .B(new_new_n185_), .C(new_new_n44_), .Y(new_new_n187_));
  NO2        g0165(.A(i_2_), .B(i_1_), .Y(new_new_n188_));
  NA2        g0166(.A(new_new_n188_), .B(i_3_), .Y(new_new_n189_));
  NAi21      g0167(.An(i_4_), .B(i_12_), .Y(new_new_n190_));
  NO4        g0168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n187_), .D(new_new_n25_), .Y(new_new_n191_));
  NO3        g0169(.A(new_new_n191_), .B(new_new_n184_), .C(new_new_n177_), .Y(new_new_n192_));
  INV        g0170(.A(i_8_), .Y(new_new_n193_));
  NO2        g0171(.A(new_new_n193_), .B(i_7_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(i_6_), .Y(new_new_n195_));
  NO3        g0173(.A(i_3_), .B(new_new_n81_), .C(new_new_n48_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(new_new_n111_), .Y(new_new_n197_));
  NO3        g0175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n198_));
  NA3        g0176(.A(new_new_n198_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n199_));
  NO3        g0177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n200_));
  OAI210     g0178(.A0(new_new_n94_), .A1(i_12_), .B0(new_new_n200_), .Y(new_new_n201_));
  AOI210     g0179(.A0(new_new_n201_), .A1(new_new_n199_), .B0(new_new_n197_), .Y(new_new_n202_));
  NO2        g0180(.A(i_3_), .B(i_8_), .Y(new_new_n203_));
  NO3        g0181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(new_new_n203_), .C(new_new_n39_), .Y(new_new_n205_));
  NO2        g0183(.A(new_new_n101_), .B(new_new_n55_), .Y(new_new_n206_));
  NO2        g0184(.A(i_13_), .B(i_9_), .Y(new_new_n207_));
  NAi21      g0185(.An(i_12_), .B(i_3_), .Y(new_new_n208_));
  NO2        g0186(.A(new_new_n44_), .B(i_5_), .Y(new_new_n209_));
  NO3        g0187(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n210_));
  NA2        g0188(.A(new_new_n210_), .B(i_10_), .Y(new_new_n211_));
  OAI220     g0189(.A0(new_new_n211_), .A1(new_new_n208_), .B0(new_new_n101_), .B1(new_new_n205_), .Y(new_new_n212_));
  AOI210     g0190(.A0(new_new_n212_), .A1(i_7_), .B0(new_new_n202_), .Y(new_new_n213_));
  OAI220     g0191(.A0(new_new_n213_), .A1(i_4_), .B0(new_new_n195_), .B1(new_new_n192_), .Y(new_new_n214_));
  NAi21      g0192(.An(i_12_), .B(i_7_), .Y(new_new_n215_));
  NA3        g0193(.A(i_13_), .B(new_new_n193_), .C(i_10_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NA2        g0195(.A(i_0_), .B(i_5_), .Y(new_new_n218_));
  NA2        g0196(.A(new_new_n218_), .B(new_new_n102_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n219_), .A1(new_new_n189_), .B0(new_new_n179_), .B1(new_new_n132_), .Y(new_new_n220_));
  NAi31      g0198(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n36_), .B(i_13_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n68_), .B(new_new_n26_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n46_), .B(new_new_n60_), .Y(new_new_n224_));
  NA3        g0202(.A(new_new_n224_), .B(new_new_n223_), .C(new_new_n222_), .Y(new_new_n225_));
  INV        g0203(.A(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n226_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n198_), .C(new_new_n196_), .Y(new_new_n228_));
  OAI210     g0206(.A0(new_new_n225_), .A1(new_new_n221_), .B0(new_new_n228_), .Y(new_new_n229_));
  AOI220     g0207(.A0(new_new_n229_), .A1(new_new_n141_), .B0(new_new_n220_), .B1(new_new_n217_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n37_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n182_), .B(i_4_), .Y(new_new_n232_));
  NA2        g0210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  OR2        g0211(.A(i_8_), .B(i_7_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n234_), .B(new_new_n81_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n51_), .B(i_1_), .Y(new_new_n236_));
  NA2        g0214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  INV        g0215(.A(i_12_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n44_), .B(new_new_n238_), .Y(new_new_n239_));
  NO3        g0217(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n240_));
  NA2        g0218(.A(i_2_), .B(i_1_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n237_), .B(new_new_n233_), .Y(new_new_n242_));
  NO3        g0220(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n243_));
  NAi21      g0221(.An(i_4_), .B(i_3_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n244_), .B(new_new_n70_), .Y(new_new_n245_));
  NO2        g0223(.A(i_0_), .B(i_6_), .Y(new_new_n246_));
  NOi41      g0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n247_), .B(new_new_n246_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n241_), .B(new_new_n182_), .Y(new_new_n249_));
  NAi21      g0227(.An(new_new_n248_), .B(new_new_n249_), .Y(new_new_n250_));
  INV        g0228(.A(new_new_n250_), .Y(new_new_n251_));
  AOI220     g0229(.A0(new_new_n251_), .A1(new_new_n39_), .B0(new_new_n242_), .B1(new_new_n207_), .Y(new_new_n252_));
  NO2        g0230(.A(i_11_), .B(new_new_n226_), .Y(new_new_n253_));
  NOi21      g0231(.An(i_1_), .B(i_6_), .Y(new_new_n254_));
  NAi21      g0232(.An(i_3_), .B(i_7_), .Y(new_new_n255_));
  NA2        g0233(.A(new_new_n238_), .B(i_9_), .Y(new_new_n256_));
  OR4        g0234(.A(new_new_n256_), .B(new_new_n255_), .C(new_new_n254_), .D(new_new_n185_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n258_));
  NO2        g0236(.A(i_12_), .B(i_3_), .Y(new_new_n259_));
  NA2        g0237(.A(new_new_n68_), .B(i_5_), .Y(new_new_n260_));
  NA2        g0238(.A(i_3_), .B(i_9_), .Y(new_new_n261_));
  NAi21      g0239(.An(i_7_), .B(i_10_), .Y(new_new_n262_));
  NO2        g0240(.A(new_new_n262_), .B(new_new_n261_), .Y(new_new_n263_));
  NA3        g0241(.A(new_new_n263_), .B(new_new_n260_), .C(new_new_n61_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n264_), .B(new_new_n257_), .Y(new_new_n265_));
  NA3        g0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n266_));
  NA2        g0244(.A(new_new_n238_), .B(i_13_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n265_), .B(new_new_n253_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n234_), .B(new_new_n37_), .Y(new_new_n269_));
  NA2        g0247(.A(i_12_), .B(i_6_), .Y(new_new_n270_));
  OR2        g0248(.A(i_13_), .B(i_9_), .Y(new_new_n271_));
  NO3        g0249(.A(new_new_n271_), .B(new_new_n270_), .C(new_new_n48_), .Y(new_new_n272_));
  NO2        g0250(.A(new_new_n244_), .B(i_2_), .Y(new_new_n273_));
  NA3        g0251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n44_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n253_), .B(i_9_), .Y(new_new_n275_));
  OAI210     g0253(.A0(new_new_n68_), .A1(new_new_n275_), .B0(new_new_n274_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n154_), .B(new_new_n60_), .Y(new_new_n277_));
  NO3        g0255(.A(i_11_), .B(new_new_n226_), .C(new_new_n25_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n255_), .B(i_8_), .Y(new_new_n279_));
  NO2        g0257(.A(i_6_), .B(new_new_n48_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n278_), .Y(new_new_n281_));
  NO3        g0259(.A(new_new_n26_), .B(new_new_n81_), .C(i_5_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n269_), .C(new_new_n227_), .Y(new_new_n283_));
  AOI210     g0261(.A0(new_new_n283_), .A1(new_new_n281_), .B0(new_new_n277_), .Y(new_new_n284_));
  AOI210     g0262(.A0(new_new_n276_), .A1(new_new_n269_), .B0(new_new_n284_), .Y(new_new_n285_));
  NA4        g0263(.A(new_new_n285_), .B(new_new_n268_), .C(new_new_n252_), .D(new_new_n230_), .Y(new_new_n286_));
  NO3        g0264(.A(i_12_), .B(new_new_n226_), .C(new_new_n37_), .Y(new_new_n287_));
  INV        g0265(.A(new_new_n287_), .Y(new_new_n288_));
  NA2        g0266(.A(i_8_), .B(new_new_n99_), .Y(new_new_n289_));
  NOi21      g0267(.An(new_new_n163_), .B(new_new_n81_), .Y(new_new_n290_));
  NO3        g0268(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n291_));
  AOI220     g0269(.A0(new_new_n291_), .A1(new_new_n196_), .B0(new_new_n290_), .B1(new_new_n236_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n292_), .B(new_new_n289_), .Y(new_new_n293_));
  NO3        g0271(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n241_), .B(i_0_), .Y(new_new_n295_));
  AOI220     g0273(.A0(new_new_n295_), .A1(new_new_n194_), .B0(new_new_n294_), .B1(new_new_n141_), .Y(new_new_n296_));
  NA2        g0274(.A(new_new_n280_), .B(new_new_n26_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(new_new_n296_), .Y(new_new_n298_));
  NA2        g0276(.A(i_0_), .B(i_1_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(i_2_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n56_), .B(i_6_), .Y(new_new_n301_));
  NA3        g0279(.A(new_new_n301_), .B(new_new_n300_), .C(new_new_n163_), .Y(new_new_n302_));
  OAI210     g0280(.A0(new_new_n165_), .A1(new_new_n142_), .B0(new_new_n302_), .Y(new_new_n303_));
  NO3        g0281(.A(new_new_n303_), .B(new_new_n298_), .C(new_new_n293_), .Y(new_new_n304_));
  NO2        g0282(.A(i_3_), .B(i_10_), .Y(new_new_n305_));
  NA3        g0283(.A(new_new_n305_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n306_));
  NO2        g0284(.A(i_2_), .B(new_new_n99_), .Y(new_new_n307_));
  NOi21      g0285(.An(new_new_n218_), .B(new_new_n101_), .Y(new_new_n308_));
  NA3        g0286(.A(new_new_n308_), .B(i_1_), .C(new_new_n307_), .Y(new_new_n309_));
  AN2        g0287(.A(i_3_), .B(i_10_), .Y(new_new_n310_));
  NA4        g0288(.A(new_new_n310_), .B(new_new_n198_), .C(new_new_n175_), .D(new_new_n173_), .Y(new_new_n311_));
  NO2        g0289(.A(i_5_), .B(new_new_n37_), .Y(new_new_n312_));
  NO2        g0290(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n313_));
  OR2        g0291(.A(new_new_n309_), .B(new_new_n306_), .Y(new_new_n314_));
  OAI220     g0292(.A0(new_new_n314_), .A1(i_6_), .B0(new_new_n304_), .B1(new_new_n288_), .Y(new_new_n315_));
  NO4        g0293(.A(new_new_n315_), .B(new_new_n286_), .C(new_new_n214_), .D(new_new_n168_), .Y(new_new_n316_));
  NO3        g0294(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n317_));
  NO2        g0295(.A(new_new_n56_), .B(new_new_n81_), .Y(new_new_n318_));
  NA2        g0296(.A(new_new_n295_), .B(new_new_n318_), .Y(new_new_n319_));
  NO3        g0297(.A(i_6_), .B(new_new_n193_), .C(i_7_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n320_), .B(new_new_n198_), .Y(new_new_n321_));
  AOI210     g0299(.A0(new_new_n321_), .A1(new_new_n319_), .B0(i_5_), .Y(new_new_n322_));
  NO2        g0300(.A(i_2_), .B(i_3_), .Y(new_new_n323_));
  OR2        g0301(.A(i_0_), .B(i_5_), .Y(new_new_n324_));
  NA2        g0302(.A(new_new_n218_), .B(new_new_n324_), .Y(new_new_n325_));
  NA4        g0303(.A(new_new_n325_), .B(new_new_n235_), .C(new_new_n323_), .D(i_1_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n295_), .B(new_new_n290_), .C(new_new_n111_), .Y(new_new_n327_));
  NAi21      g0305(.An(i_8_), .B(i_7_), .Y(new_new_n328_));
  NO2        g0306(.A(new_new_n157_), .B(new_new_n46_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n329_), .B(i_7_), .C(new_new_n163_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n330_), .B(new_new_n327_), .C(new_new_n326_), .Y(new_new_n331_));
  OAI210     g0309(.A0(new_new_n331_), .A1(new_new_n322_), .B0(i_4_), .Y(new_new_n332_));
  NO2        g0310(.A(i_12_), .B(i_10_), .Y(new_new_n333_));
  NOi21      g0311(.An(i_5_), .B(i_0_), .Y(new_new_n334_));
  AOI210     g0312(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n99_), .Y(new_new_n335_));
  NO4        g0313(.A(new_new_n335_), .B(i_4_), .C(new_new_n334_), .D(new_new_n127_), .Y(new_new_n336_));
  NA4        g0314(.A(new_new_n79_), .B(new_new_n36_), .C(new_new_n81_), .D(i_8_), .Y(new_new_n337_));
  NA2        g0315(.A(new_new_n336_), .B(new_new_n333_), .Y(new_new_n338_));
  NO2        g0316(.A(i_6_), .B(i_8_), .Y(new_new_n339_));
  NOi21      g0317(.An(i_0_), .B(i_2_), .Y(new_new_n340_));
  AN2        g0318(.A(new_new_n340_), .B(new_new_n339_), .Y(new_new_n341_));
  NO2        g0319(.A(i_1_), .B(i_7_), .Y(new_new_n342_));
  NA3        g0320(.A(new_new_n339_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n343_));
  NA3        g0321(.A(new_new_n343_), .B(new_new_n338_), .C(new_new_n332_), .Y(new_new_n344_));
  NO3        g0322(.A(new_new_n234_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n345_));
  NO3        g0323(.A(new_new_n328_), .B(i_2_), .C(i_1_), .Y(new_new_n346_));
  OAI210     g0324(.A0(new_new_n346_), .A1(new_new_n345_), .B0(i_6_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n254_), .B(new_new_n307_), .C(new_new_n193_), .Y(new_new_n348_));
  AOI210     g0326(.A0(new_new_n348_), .A1(new_new_n347_), .B0(new_new_n325_), .Y(new_new_n349_));
  NOi21      g0327(.An(new_new_n153_), .B(new_new_n102_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n350_), .B(new_new_n123_), .Y(new_new_n351_));
  OAI210     g0329(.A0(new_new_n351_), .A1(new_new_n349_), .B0(i_3_), .Y(new_new_n352_));
  INV        g0330(.A(new_new_n79_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n299_), .B(new_new_n76_), .Y(new_new_n354_));
  NA2        g0332(.A(new_new_n354_), .B(new_new_n131_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n90_), .B(new_new_n193_), .Y(new_new_n356_));
  NA3        g0334(.A(new_new_n308_), .B(new_new_n356_), .C(new_new_n60_), .Y(new_new_n357_));
  AOI210     g0335(.A0(new_new_n357_), .A1(new_new_n355_), .B0(new_new_n353_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n193_), .B(i_9_), .Y(new_new_n359_));
  NA3        g0337(.A(new_new_n359_), .B(new_new_n206_), .C(new_new_n157_), .Y(new_new_n360_));
  NO2        g0338(.A(new_new_n360_), .B(new_new_n46_), .Y(new_new_n361_));
  NO3        g0339(.A(new_new_n361_), .B(new_new_n358_), .C(new_new_n298_), .Y(new_new_n362_));
  AOI210     g0340(.A0(new_new_n362_), .A1(new_new_n352_), .B0(new_new_n162_), .Y(new_new_n363_));
  AOI210     g0341(.A0(new_new_n344_), .A1(new_new_n317_), .B0(new_new_n363_), .Y(new_new_n364_));
  NOi32      g0342(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n365_));
  INV        g0343(.A(new_new_n365_), .Y(new_new_n366_));
  NAi21      g0344(.An(i_0_), .B(i_6_), .Y(new_new_n367_));
  NAi21      g0345(.An(i_1_), .B(i_5_), .Y(new_new_n368_));
  NA2        g0346(.A(new_new_n368_), .B(new_new_n367_), .Y(new_new_n369_));
  NA2        g0347(.A(new_new_n369_), .B(new_new_n25_), .Y(new_new_n370_));
  OAI210     g0348(.A0(new_new_n370_), .A1(new_new_n159_), .B0(new_new_n248_), .Y(new_new_n371_));
  NAi41      g0349(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n372_));
  OAI220     g0350(.A0(new_new_n372_), .A1(new_new_n368_), .B0(new_new_n221_), .B1(new_new_n159_), .Y(new_new_n373_));
  AOI210     g0351(.A0(new_new_n372_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n374_));
  NOi32      g0352(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n375_));
  NAi21      g0353(.An(i_6_), .B(i_1_), .Y(new_new_n376_));
  NA3        g0354(.A(new_new_n376_), .B(new_new_n375_), .C(new_new_n46_), .Y(new_new_n377_));
  NO2        g0355(.A(new_new_n377_), .B(i_0_), .Y(new_new_n378_));
  OR3        g0356(.A(new_new_n378_), .B(new_new_n374_), .C(new_new_n373_), .Y(new_new_n379_));
  NO2        g0357(.A(i_1_), .B(new_new_n99_), .Y(new_new_n380_));
  NAi21      g0358(.An(i_3_), .B(i_4_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n381_), .B(i_9_), .Y(new_new_n382_));
  AN2        g0360(.A(i_6_), .B(i_7_), .Y(new_new_n383_));
  OAI210     g0361(.A0(new_new_n383_), .A1(new_new_n380_), .B0(new_new_n382_), .Y(new_new_n384_));
  NA2        g0362(.A(i_2_), .B(i_7_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n381_), .B(i_10_), .Y(new_new_n386_));
  NA3        g0364(.A(new_new_n386_), .B(new_new_n385_), .C(new_new_n246_), .Y(new_new_n387_));
  AOI210     g0365(.A0(new_new_n387_), .A1(new_new_n384_), .B0(new_new_n185_), .Y(new_new_n388_));
  AOI210     g0366(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n389_));
  AOI220     g0367(.A0(new_new_n386_), .A1(new_new_n342_), .B0(new_new_n240_), .B1(new_new_n188_), .Y(new_new_n390_));
  NO3        g0368(.A(new_new_n388_), .B(new_new_n379_), .C(new_new_n371_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n366_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n393_));
  AN2        g0371(.A(i_12_), .B(i_5_), .Y(new_new_n394_));
  NO2        g0372(.A(i_4_), .B(new_new_n26_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n395_), .B(new_new_n394_), .Y(new_new_n396_));
  NO2        g0374(.A(i_11_), .B(i_6_), .Y(new_new_n397_));
  NA3        g0375(.A(new_new_n397_), .B(new_new_n329_), .C(new_new_n226_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n396_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n244_), .B(i_5_), .Y(new_new_n400_));
  NO2        g0378(.A(i_5_), .B(i_10_), .Y(new_new_n401_));
  NA2        g0379(.A(new_new_n143_), .B(new_new_n45_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n402_), .B(new_new_n244_), .Y(new_new_n403_));
  OAI210     g0381(.A0(new_new_n403_), .A1(new_new_n399_), .B0(new_new_n393_), .Y(new_new_n404_));
  NO2        g0382(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n149_), .B(new_new_n81_), .Y(new_new_n406_));
  OAI210     g0384(.A0(new_new_n406_), .A1(new_new_n399_), .B0(new_new_n405_), .Y(new_new_n407_));
  NO3        g0385(.A(new_new_n81_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n408_));
  NO2        g0386(.A(i_3_), .B(new_new_n99_), .Y(new_new_n409_));
  NO2        g0387(.A(i_11_), .B(i_12_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n401_), .B(new_new_n238_), .Y(new_new_n411_));
  NA3        g0389(.A(new_new_n111_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n412_));
  OAI220     g0390(.A0(new_new_n412_), .A1(new_new_n221_), .B0(new_new_n411_), .B1(new_new_n337_), .Y(new_new_n413_));
  NAi21      g0391(.An(i_13_), .B(i_0_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n414_), .B(new_new_n241_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n413_), .B(new_new_n415_), .Y(new_new_n416_));
  NA3        g0394(.A(new_new_n416_), .B(new_new_n407_), .C(new_new_n404_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n44_), .B(new_new_n226_), .Y(new_new_n418_));
  NO3        g0396(.A(i_1_), .B(i_12_), .C(new_new_n81_), .Y(new_new_n419_));
  NO2        g0397(.A(i_0_), .B(i_11_), .Y(new_new_n420_));
  NOi21      g0398(.An(i_2_), .B(i_12_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n421_), .B(i_6_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n422_), .B(new_new_n1114_), .Y(new_new_n423_));
  NA2        g0401(.A(new_new_n141_), .B(i_9_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(i_4_), .Y(new_new_n425_));
  NA2        g0403(.A(new_new_n423_), .B(new_new_n425_), .Y(new_new_n426_));
  NAi21      g0404(.An(i_9_), .B(i_4_), .Y(new_new_n427_));
  OR2        g0405(.A(i_13_), .B(i_10_), .Y(new_new_n428_));
  NO3        g0406(.A(new_new_n428_), .B(new_new_n116_), .C(new_new_n427_), .Y(new_new_n429_));
  NO2        g0407(.A(new_new_n172_), .B(new_new_n122_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n99_), .B(new_new_n25_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n287_), .B(new_new_n431_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n280_), .B(new_new_n210_), .Y(new_new_n433_));
  OAI220     g0411(.A0(new_new_n433_), .A1(new_new_n216_), .B0(new_new_n432_), .B1(new_new_n350_), .Y(new_new_n434_));
  INV        g0412(.A(new_new_n434_), .Y(new_new_n435_));
  AOI210     g0413(.A0(new_new_n435_), .A1(new_new_n426_), .B0(new_new_n26_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n327_), .B(new_new_n326_), .Y(new_new_n437_));
  AOI220     g0415(.A0(new_new_n301_), .A1(new_new_n291_), .B0(new_new_n295_), .B1(new_new_n318_), .Y(new_new_n438_));
  NO2        g0416(.A(new_new_n438_), .B(i_5_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n182_), .B(new_new_n81_), .Y(new_new_n440_));
  AOI220     g0418(.A0(new_new_n440_), .A1(new_new_n300_), .B0(new_new_n282_), .B1(new_new_n210_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n441_), .B(new_new_n289_), .Y(new_new_n442_));
  NO3        g0420(.A(new_new_n442_), .B(new_new_n439_), .C(new_new_n437_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n196_), .B(new_new_n94_), .Y(new_new_n444_));
  NA3        g0422(.A(new_new_n329_), .B(new_new_n163_), .C(new_new_n81_), .Y(new_new_n445_));
  AOI210     g0423(.A0(new_new_n445_), .A1(new_new_n444_), .B0(new_new_n328_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n193_), .B(i_10_), .Y(new_new_n447_));
  NA3        g0425(.A(new_new_n260_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n301_), .B(new_new_n236_), .Y(new_new_n449_));
  OAI220     g0427(.A0(new_new_n449_), .A1(new_new_n182_), .B0(new_new_n448_), .B1(new_new_n447_), .Y(new_new_n450_));
  NO2        g0428(.A(i_3_), .B(new_new_n48_), .Y(new_new_n451_));
  NA3        g0429(.A(new_new_n342_), .B(new_new_n341_), .C(new_new_n451_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n320_), .B(new_new_n325_), .Y(new_new_n453_));
  OAI210     g0431(.A0(new_new_n453_), .A1(new_new_n189_), .B0(new_new_n452_), .Y(new_new_n454_));
  NO3        g0432(.A(new_new_n454_), .B(new_new_n450_), .C(new_new_n446_), .Y(new_new_n455_));
  AOI210     g0433(.A0(new_new_n455_), .A1(new_new_n443_), .B0(new_new_n275_), .Y(new_new_n456_));
  NO4        g0434(.A(new_new_n456_), .B(new_new_n436_), .C(new_new_n417_), .D(new_new_n392_), .Y(new_new_n457_));
  NO2        g0435(.A(new_new_n60_), .B(i_4_), .Y(new_new_n458_));
  NO2        g0436(.A(new_new_n68_), .B(i_13_), .Y(new_new_n459_));
  NA3        g0437(.A(new_new_n459_), .B(new_new_n458_), .C(i_2_), .Y(new_new_n460_));
  NO2        g0438(.A(i_10_), .B(i_9_), .Y(new_new_n461_));
  NAi21      g0439(.An(i_12_), .B(i_8_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n462_), .B(i_3_), .Y(new_new_n463_));
  NA2        g0441(.A(new_new_n463_), .B(new_new_n461_), .Y(new_new_n464_));
  NA2        g0442(.A(i_2_), .B(new_new_n102_), .Y(new_new_n465_));
  OAI220     g0443(.A0(new_new_n465_), .A1(new_new_n205_), .B0(new_new_n464_), .B1(new_new_n460_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n313_), .B(i_0_), .Y(new_new_n467_));
  NO3        g0445(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n270_), .B(new_new_n95_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n470_));
  NA2        g0448(.A(i_8_), .B(i_9_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n287_), .B(new_new_n206_), .Y(new_new_n472_));
  OAI220     g0450(.A0(new_new_n472_), .A1(new_new_n471_), .B0(new_new_n470_), .B1(new_new_n467_), .Y(new_new_n473_));
  NO3        g0451(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n474_));
  NA3        g0452(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n473_), .B(new_new_n466_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n300_), .B(new_new_n106_), .Y(new_new_n477_));
  OA210      g0455(.A0(new_new_n360_), .A1(new_new_n99_), .B0(new_new_n302_), .Y(new_new_n478_));
  OA220      g0456(.A0(new_new_n478_), .A1(new_new_n162_), .B0(new_new_n477_), .B1(new_new_n233_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n94_), .B(i_13_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n440_), .B(new_new_n393_), .Y(new_new_n481_));
  NO2        g0459(.A(i_2_), .B(i_13_), .Y(new_new_n482_));
  NO2        g0460(.A(new_new_n481_), .B(new_new_n480_), .Y(new_new_n483_));
  NO3        g0461(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n484_));
  NO2        g0462(.A(i_6_), .B(i_7_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n485_), .B(new_new_n484_), .Y(new_new_n486_));
  NO2        g0464(.A(i_11_), .B(i_1_), .Y(new_new_n487_));
  OR2        g0465(.A(i_11_), .B(i_8_), .Y(new_new_n488_));
  NOi21      g0466(.An(i_2_), .B(i_7_), .Y(new_new_n489_));
  NAi31      g0467(.An(new_new_n488_), .B(new_new_n489_), .C(new_new_n1115_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n428_), .B(i_6_), .Y(new_new_n491_));
  NA3        g0469(.A(new_new_n491_), .B(new_new_n458_), .C(new_new_n70_), .Y(new_new_n492_));
  NO2        g0470(.A(new_new_n492_), .B(new_new_n490_), .Y(new_new_n493_));
  NO2        g0471(.A(i_3_), .B(new_new_n193_), .Y(new_new_n494_));
  NO2        g0472(.A(i_6_), .B(i_10_), .Y(new_new_n495_));
  NA4        g0473(.A(new_new_n495_), .B(new_new_n317_), .C(new_new_n494_), .D(new_new_n238_), .Y(new_new_n496_));
  NO2        g0474(.A(new_new_n496_), .B(new_new_n155_), .Y(new_new_n497_));
  NA3        g0475(.A(new_new_n247_), .B(new_new_n171_), .C(new_new_n131_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n157_), .B(i_3_), .Y(new_new_n500_));
  NA3        g0478(.A(new_new_n405_), .B(new_new_n178_), .C(new_new_n148_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n501_), .B(new_new_n498_), .Y(new_new_n502_));
  NO4        g0480(.A(new_new_n502_), .B(new_new_n497_), .C(new_new_n493_), .D(new_new_n483_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n468_), .B(new_new_n394_), .Y(new_new_n504_));
  NA2        g0482(.A(new_new_n474_), .B(new_new_n401_), .Y(new_new_n505_));
  OAI220     g0483(.A0(new_new_n505_), .A1(new_new_n225_), .B0(new_new_n504_), .B1(new_new_n54_), .Y(new_new_n506_));
  NAi21      g0484(.An(new_new_n216_), .B(new_new_n410_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n342_), .B(new_new_n218_), .Y(new_new_n508_));
  NO2        g0486(.A(new_new_n26_), .B(i_5_), .Y(new_new_n509_));
  NO2        g0487(.A(i_0_), .B(new_new_n81_), .Y(new_new_n510_));
  NA3        g0488(.A(new_new_n510_), .B(new_new_n509_), .C(new_new_n141_), .Y(new_new_n511_));
  OR3        g0489(.A(i_4_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n512_));
  OAI220     g0490(.A0(new_new_n512_), .A1(new_new_n511_), .B0(new_new_n508_), .B1(new_new_n507_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n27_), .B(i_10_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n317_), .B(new_new_n240_), .Y(new_new_n515_));
  OAI220     g0493(.A0(new_new_n515_), .A1(new_new_n448_), .B0(new_new_n514_), .B1(new_new_n480_), .Y(new_new_n516_));
  NA4        g0494(.A(new_new_n310_), .B(new_new_n224_), .C(new_new_n68_), .D(new_new_n238_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n517_), .B(new_new_n486_), .Y(new_new_n518_));
  NO4        g0496(.A(new_new_n518_), .B(new_new_n516_), .C(new_new_n513_), .D(new_new_n506_), .Y(new_new_n519_));
  NA4        g0497(.A(new_new_n519_), .B(new_new_n503_), .C(new_new_n479_), .D(new_new_n476_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n310_), .B(new_new_n175_), .C(new_new_n173_), .Y(new_new_n521_));
  OAI210     g0499(.A0(new_new_n306_), .A1(new_new_n180_), .B0(new_new_n521_), .Y(new_new_n522_));
  AN2        g0500(.A(new_new_n291_), .B(new_new_n235_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n523_), .B(new_new_n522_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n121_), .B(new_new_n110_), .Y(new_new_n525_));
  AO220      g0503(.A0(new_new_n525_), .A1(new_new_n468_), .B0(new_new_n429_), .B1(i_6_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n317_), .B(new_new_n164_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n527_), .A1(new_new_n233_), .B0(new_new_n311_), .Y(new_new_n528_));
  AOI220     g0506(.A0(new_new_n528_), .A1(i_7_), .B0(new_new_n526_), .B1(new_new_n313_), .Y(new_new_n529_));
  NA4        g0507(.A(new_new_n459_), .B(new_new_n458_), .C(new_new_n203_), .D(i_2_), .Y(new_new_n530_));
  INV        g0508(.A(new_new_n530_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n394_), .B(new_new_n226_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n365_), .B(new_new_n68_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n383_), .B(new_new_n375_), .Y(new_new_n534_));
  AO210      g0512(.A0(new_new_n533_), .A1(new_new_n532_), .B0(new_new_n534_), .Y(new_new_n535_));
  NO2        g0513(.A(new_new_n36_), .B(i_8_), .Y(new_new_n536_));
  NAi41      g0514(.An(new_new_n533_), .B(new_new_n495_), .C(new_new_n536_), .D(new_new_n46_), .Y(new_new_n537_));
  INV        g0515(.A(new_new_n429_), .Y(new_new_n538_));
  NA3        g0516(.A(new_new_n538_), .B(new_new_n537_), .C(new_new_n535_), .Y(new_new_n539_));
  AOI210     g0517(.A0(new_new_n531_), .A1(new_new_n204_), .B0(new_new_n539_), .Y(new_new_n540_));
  OAI210     g0518(.A0(i_8_), .A1(new_new_n60_), .B0(new_new_n133_), .Y(new_new_n541_));
  AOI210     g0519(.A0(new_new_n194_), .A1(i_9_), .B0(new_new_n269_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n542_), .B(new_new_n199_), .Y(new_new_n543_));
  NO2        g0521(.A(new_new_n182_), .B(new_new_n81_), .Y(new_new_n544_));
  AOI220     g0522(.A0(new_new_n544_), .A1(new_new_n543_), .B0(new_new_n541_), .B1(new_new_n430_), .Y(new_new_n545_));
  NA4        g0523(.A(new_new_n545_), .B(new_new_n540_), .C(new_new_n529_), .D(new_new_n524_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n400_), .B(new_new_n300_), .Y(new_new_n547_));
  OAI210     g0525(.A0(new_new_n396_), .A1(new_new_n169_), .B0(new_new_n547_), .Y(new_new_n548_));
  NO2        g0526(.A(i_12_), .B(new_new_n193_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n549_), .B(new_new_n226_), .Y(new_new_n550_));
  NO3        g0528(.A(i_10_), .B(new_new_n550_), .C(new_new_n477_), .Y(new_new_n551_));
  NOi31      g0529(.An(new_new_n320_), .B(new_new_n428_), .C(new_new_n38_), .Y(new_new_n552_));
  OAI210     g0530(.A0(new_new_n552_), .A1(new_new_n551_), .B0(new_new_n548_), .Y(new_new_n553_));
  NO2        g0531(.A(i_8_), .B(i_7_), .Y(new_new_n554_));
  OAI210     g0532(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n555_), .B(new_new_n224_), .Y(new_new_n556_));
  AOI220     g0534(.A0(new_new_n329_), .A1(new_new_n39_), .B0(new_new_n236_), .B1(new_new_n207_), .Y(new_new_n557_));
  OAI220     g0535(.A0(new_new_n557_), .A1(new_new_n182_), .B0(new_new_n556_), .B1(new_new_n244_), .Y(new_new_n558_));
  NA2        g0536(.A(new_new_n44_), .B(i_10_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n559_), .B(i_6_), .Y(new_new_n560_));
  NA3        g0538(.A(new_new_n560_), .B(new_new_n558_), .C(new_new_n554_), .Y(new_new_n561_));
  AOI220     g0539(.A0(new_new_n440_), .A1(new_new_n329_), .B0(new_new_n249_), .B1(new_new_n246_), .Y(new_new_n562_));
  OAI220     g0540(.A0(new_new_n562_), .A1(new_new_n267_), .B0(new_new_n480_), .B1(new_new_n132_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n563_), .B(new_new_n269_), .Y(new_new_n564_));
  NOi31      g0542(.An(new_new_n295_), .B(new_new_n306_), .C(new_new_n180_), .Y(new_new_n565_));
  NA3        g0543(.A(new_new_n310_), .B(new_new_n173_), .C(new_new_n94_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n222_), .B(new_new_n44_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n157_), .B(i_5_), .Y(new_new_n568_));
  NA3        g0546(.A(new_new_n568_), .B(new_new_n418_), .C(new_new_n323_), .Y(new_new_n569_));
  OAI210     g0547(.A0(new_new_n569_), .A1(new_new_n567_), .B0(new_new_n566_), .Y(new_new_n570_));
  OAI210     g0548(.A0(new_new_n570_), .A1(new_new_n565_), .B0(new_new_n474_), .Y(new_new_n571_));
  NA4        g0549(.A(new_new_n571_), .B(new_new_n564_), .C(new_new_n561_), .D(new_new_n553_), .Y(new_new_n572_));
  NA3        g0550(.A(new_new_n218_), .B(new_new_n66_), .C(new_new_n44_), .Y(new_new_n573_));
  NA2        g0551(.A(new_new_n287_), .B(new_new_n79_), .Y(new_new_n574_));
  AOI210     g0552(.A0(new_new_n573_), .A1(new_new_n355_), .B0(new_new_n574_), .Y(new_new_n575_));
  NA2        g0553(.A(new_new_n301_), .B(new_new_n291_), .Y(new_new_n576_));
  NO2        g0554(.A(new_new_n576_), .B(new_new_n172_), .Y(new_new_n577_));
  NA2        g0555(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n578_));
  NA2        g0556(.A(new_new_n461_), .B(new_new_n222_), .Y(new_new_n579_));
  NO2        g0557(.A(new_new_n578_), .B(new_new_n579_), .Y(new_new_n580_));
  AOI210     g0558(.A0(new_new_n376_), .A1(new_new_n46_), .B0(new_new_n380_), .Y(new_new_n581_));
  NA2        g0559(.A(i_0_), .B(new_new_n48_), .Y(new_new_n582_));
  NA3        g0560(.A(new_new_n549_), .B(new_new_n278_), .C(new_new_n582_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n581_), .B(new_new_n583_), .Y(new_new_n584_));
  NO4        g0562(.A(new_new_n584_), .B(new_new_n580_), .C(new_new_n577_), .D(new_new_n575_), .Y(new_new_n585_));
  NO4        g0563(.A(new_new_n254_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n586_));
  NO3        g0564(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n234_), .B(new_new_n36_), .Y(new_new_n588_));
  AN2        g0566(.A(new_new_n588_), .B(new_new_n587_), .Y(new_new_n589_));
  OA210      g0567(.A0(new_new_n589_), .A1(new_new_n586_), .B0(new_new_n365_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n428_), .B(i_1_), .Y(new_new_n591_));
  NOi31      g0569(.An(new_new_n591_), .B(new_new_n469_), .C(new_new_n68_), .Y(new_new_n592_));
  AN4        g0570(.A(new_new_n592_), .B(new_new_n425_), .C(new_new_n509_), .D(i_2_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n438_), .B(new_new_n176_), .Y(new_new_n594_));
  NO3        g0572(.A(new_new_n594_), .B(new_new_n593_), .C(new_new_n590_), .Y(new_new_n595_));
  NOi21      g0573(.An(i_10_), .B(i_6_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n81_), .B(new_new_n25_), .Y(new_new_n597_));
  AOI220     g0575(.A0(new_new_n287_), .A1(new_new_n597_), .B0(new_new_n278_), .B1(new_new_n596_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n598_), .B(new_new_n467_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n113_), .B(new_new_n23_), .Y(new_new_n600_));
  NA2        g0578(.A(new_new_n320_), .B(new_new_n164_), .Y(new_new_n601_));
  AOI220     g0579(.A0(new_new_n601_), .A1(new_new_n449_), .B0(new_new_n183_), .B1(new_new_n181_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n198_), .B(new_new_n37_), .Y(new_new_n603_));
  NOi31      g0581(.An(new_new_n145_), .B(new_new_n603_), .C(new_new_n337_), .Y(new_new_n604_));
  NO3        g0582(.A(new_new_n604_), .B(new_new_n602_), .C(new_new_n599_), .Y(new_new_n605_));
  NO2        g0583(.A(new_new_n533_), .B(new_new_n390_), .Y(new_new_n606_));
  INV        g0584(.A(new_new_n323_), .Y(new_new_n607_));
  NO2        g0585(.A(i_12_), .B(new_new_n81_), .Y(new_new_n608_));
  NA3        g0586(.A(new_new_n608_), .B(new_new_n278_), .C(new_new_n582_), .Y(new_new_n609_));
  NA3        g0587(.A(new_new_n397_), .B(new_new_n287_), .C(new_new_n218_), .Y(new_new_n610_));
  AOI210     g0588(.A0(new_new_n610_), .A1(new_new_n609_), .B0(new_new_n607_), .Y(new_new_n611_));
  NA2        g0589(.A(new_new_n173_), .B(i_0_), .Y(new_new_n612_));
  NO3        g0590(.A(new_new_n612_), .B(new_new_n347_), .C(new_new_n306_), .Y(new_new_n613_));
  OR2        g0591(.A(i_2_), .B(i_5_), .Y(new_new_n614_));
  OR2        g0592(.A(new_new_n614_), .B(i_6_), .Y(new_new_n615_));
  AOI210     g0593(.A0(new_new_n385_), .A1(new_new_n246_), .B0(new_new_n198_), .Y(new_new_n616_));
  AOI210     g0594(.A0(new_new_n616_), .A1(new_new_n615_), .B0(new_new_n507_), .Y(new_new_n617_));
  NO4        g0595(.A(new_new_n617_), .B(new_new_n613_), .C(new_new_n611_), .D(new_new_n606_), .Y(new_new_n618_));
  NA4        g0596(.A(new_new_n618_), .B(new_new_n605_), .C(new_new_n595_), .D(new_new_n585_), .Y(new_new_n619_));
  NO4        g0597(.A(new_new_n619_), .B(new_new_n572_), .C(new_new_n546_), .D(new_new_n520_), .Y(new_new_n620_));
  NA4        g0598(.A(new_new_n620_), .B(new_new_n457_), .C(new_new_n364_), .D(new_new_n316_), .Y(men7));
  NO2        g0599(.A(new_new_n106_), .B(new_new_n87_), .Y(new_new_n622_));
  NA2        g0600(.A(new_new_n395_), .B(new_new_n622_), .Y(new_new_n623_));
  NA2        g0601(.A(new_new_n495_), .B(new_new_n79_), .Y(new_new_n624_));
  NA2        g0602(.A(i_11_), .B(new_new_n193_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n143_), .B(new_new_n625_), .Y(new_new_n626_));
  OAI210     g0604(.A0(new_new_n626_), .A1(new_new_n624_), .B0(new_new_n623_), .Y(new_new_n627_));
  NA3        g0605(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n628_));
  NO2        g0606(.A(new_new_n238_), .B(i_4_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n629_), .B(i_8_), .Y(new_new_n630_));
  NA2        g0608(.A(i_2_), .B(new_new_n81_), .Y(new_new_n631_));
  OAI210     g0609(.A0(new_new_n84_), .A1(new_new_n203_), .B0(new_new_n204_), .Y(new_new_n632_));
  NO2        g0610(.A(i_7_), .B(new_new_n37_), .Y(new_new_n633_));
  NA2        g0611(.A(i_4_), .B(i_8_), .Y(new_new_n634_));
  INV        g0612(.A(new_new_n627_), .Y(new_new_n635_));
  INV        g0613(.A(new_new_n161_), .Y(new_new_n636_));
  OR2        g0614(.A(i_6_), .B(i_10_), .Y(new_new_n637_));
  NO2        g0615(.A(new_new_n637_), .B(new_new_n23_), .Y(new_new_n638_));
  OR3        g0616(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n639_));
  NO3        g0617(.A(new_new_n639_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n640_));
  INV        g0618(.A(new_new_n200_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n640_), .B(new_new_n638_), .Y(new_new_n642_));
  OA220      g0620(.A0(new_new_n642_), .A1(new_new_n607_), .B0(new_new_n636_), .B1(new_new_n271_), .Y(new_new_n643_));
  AOI210     g0621(.A0(new_new_n643_), .A1(new_new_n635_), .B0(new_new_n60_), .Y(new_new_n644_));
  NOi21      g0622(.An(i_11_), .B(i_7_), .Y(new_new_n645_));
  AO210      g0623(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n647_), .B(new_new_n207_), .Y(new_new_n648_));
  NA3        g0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n649_));
  NAi31      g0627(.An(new_new_n649_), .B(new_new_n215_), .C(i_11_), .Y(new_new_n650_));
  AOI210     g0628(.A0(new_new_n650_), .A1(new_new_n648_), .B0(new_new_n60_), .Y(new_new_n651_));
  NA2        g0629(.A(new_new_n83_), .B(new_new_n60_), .Y(new_new_n652_));
  AO210      g0630(.A0(new_new_n652_), .A1(new_new_n390_), .B0(new_new_n40_), .Y(new_new_n653_));
  NO3        g0631(.A(new_new_n262_), .B(new_new_n208_), .C(new_new_n625_), .Y(new_new_n654_));
  OAI210     g0632(.A0(new_new_n654_), .A1(new_new_n227_), .B0(new_new_n60_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n421_), .B(new_new_n31_), .Y(new_new_n656_));
  OR2        g0634(.A(new_new_n208_), .B(new_new_n106_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(new_new_n656_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n60_), .B(i_9_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n659_), .B(i_4_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n660_), .B(new_new_n658_), .Y(new_new_n661_));
  NO2        g0639(.A(i_1_), .B(i_12_), .Y(new_new_n662_));
  NA3        g0640(.A(new_new_n662_), .B(new_new_n108_), .C(new_new_n24_), .Y(new_new_n663_));
  NA4        g0641(.A(new_new_n663_), .B(new_new_n661_), .C(new_new_n655_), .D(new_new_n653_), .Y(new_new_n664_));
  OAI210     g0642(.A0(new_new_n664_), .A1(new_new_n651_), .B0(i_6_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n649_), .B(new_new_n106_), .Y(new_new_n666_));
  NA2        g0644(.A(new_new_n666_), .B(new_new_n608_), .Y(new_new_n667_));
  NO2        g0645(.A(i_6_), .B(i_11_), .Y(new_new_n668_));
  NA3        g0646(.A(new_new_n667_), .B(new_new_n538_), .C(new_new_n470_), .Y(new_new_n669_));
  NO4        g0647(.A(new_new_n215_), .B(new_new_n127_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n670_));
  NA2        g0648(.A(new_new_n670_), .B(new_new_n659_), .Y(new_new_n671_));
  NO3        g0649(.A(new_new_n637_), .B(new_new_n234_), .C(new_new_n23_), .Y(new_new_n672_));
  AOI210     g0650(.A0(i_1_), .A1(new_new_n263_), .B0(new_new_n672_), .Y(new_new_n673_));
  OAI210     g0651(.A0(new_new_n673_), .A1(new_new_n44_), .B0(new_new_n671_), .Y(new_new_n674_));
  NA3        g0652(.A(new_new_n554_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n137_), .B(i_9_), .Y(new_new_n676_));
  NA3        g0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n46_), .B(i_1_), .Y(new_new_n678_));
  NA3        g0656(.A(new_new_n678_), .B(new_new_n270_), .C(new_new_n44_), .Y(new_new_n679_));
  OAI220     g0657(.A0(new_new_n679_), .A1(new_new_n677_), .B0(new_new_n676_), .B1(new_new_n1113_), .Y(new_new_n680_));
  NA3        g0658(.A(new_new_n659_), .B(new_new_n323_), .C(i_6_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n681_), .B(new_new_n23_), .Y(new_new_n682_));
  AOI210     g0660(.A0(new_new_n487_), .A1(new_new_n431_), .B0(new_new_n243_), .Y(new_new_n683_));
  NO2        g0661(.A(new_new_n683_), .B(new_new_n631_), .Y(new_new_n684_));
  NAi21      g0662(.An(new_new_n675_), .B(new_new_n89_), .Y(new_new_n685_));
  NA2        g0663(.A(new_new_n678_), .B(new_new_n270_), .Y(new_new_n686_));
  NO2        g0664(.A(i_11_), .B(new_new_n37_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n687_), .B(new_new_n24_), .Y(new_new_n688_));
  OAI210     g0666(.A0(new_new_n688_), .A1(new_new_n686_), .B0(new_new_n685_), .Y(new_new_n689_));
  OR4        g0667(.A(new_new_n689_), .B(new_new_n684_), .C(new_new_n682_), .D(new_new_n680_), .Y(new_new_n690_));
  NO3        g0668(.A(new_new_n690_), .B(new_new_n674_), .C(new_new_n669_), .Y(new_new_n691_));
  NO2        g0669(.A(new_new_n238_), .B(new_new_n99_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n692_), .B(new_new_n645_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n693_), .B(i_1_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n694_), .B(new_new_n639_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n427_), .B(new_new_n81_), .Y(new_new_n696_));
  NA2        g0674(.A(new_new_n695_), .B(new_new_n46_), .Y(new_new_n697_));
  NA2        g0675(.A(i_3_), .B(new_new_n193_), .Y(new_new_n698_));
  AOI210     g0676(.A0(new_new_n261_), .A1(new_new_n698_), .B0(new_new_n113_), .Y(new_new_n699_));
  AN2        g0677(.A(new_new_n699_), .B(new_new_n560_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n234_), .B(new_new_n44_), .Y(new_new_n701_));
  NO3        g0679(.A(new_new_n701_), .B(new_new_n313_), .C(new_new_n239_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n116_), .B(new_new_n37_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n703_), .B(i_6_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n81_), .B(i_9_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n60_), .Y(new_new_n706_));
  NO2        g0684(.A(new_new_n706_), .B(new_new_n662_), .Y(new_new_n707_));
  NO4        g0685(.A(new_new_n707_), .B(new_new_n704_), .C(new_new_n702_), .D(i_4_), .Y(new_new_n708_));
  NA2        g0686(.A(i_1_), .B(i_3_), .Y(new_new_n709_));
  NO2        g0687(.A(new_new_n471_), .B(new_new_n90_), .Y(new_new_n710_));
  AOI210     g0688(.A0(new_new_n701_), .A1(new_new_n596_), .B0(new_new_n710_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n711_), .B(new_new_n709_), .Y(new_new_n712_));
  NO3        g0690(.A(new_new_n712_), .B(new_new_n708_), .C(new_new_n700_), .Y(new_new_n713_));
  NA4        g0691(.A(new_new_n713_), .B(new_new_n697_), .C(new_new_n691_), .D(new_new_n665_), .Y(new_new_n714_));
  NO3        g0692(.A(new_new_n488_), .B(i_3_), .C(i_7_), .Y(new_new_n715_));
  NOi21      g0693(.An(new_new_n715_), .B(i_10_), .Y(new_new_n716_));
  OA210      g0694(.A0(new_new_n716_), .A1(new_new_n247_), .B0(new_new_n81_), .Y(new_new_n717_));
  NA2        g0695(.A(new_new_n383_), .B(new_new_n382_), .Y(new_new_n718_));
  NA3        g0696(.A(new_new_n495_), .B(new_new_n536_), .C(new_new_n46_), .Y(new_new_n719_));
  NO3        g0697(.A(new_new_n489_), .B(new_new_n634_), .C(new_new_n81_), .Y(new_new_n720_));
  NA2        g0698(.A(new_new_n720_), .B(new_new_n25_), .Y(new_new_n721_));
  NA3        g0699(.A(new_new_n161_), .B(new_new_n79_), .C(new_new_n81_), .Y(new_new_n722_));
  NA4        g0700(.A(new_new_n722_), .B(new_new_n721_), .C(new_new_n719_), .D(new_new_n718_), .Y(new_new_n723_));
  OAI210     g0701(.A0(new_new_n723_), .A1(new_new_n717_), .B0(i_1_), .Y(new_new_n724_));
  AOI210     g0702(.A0(new_new_n270_), .A1(new_new_n95_), .B0(i_1_), .Y(new_new_n725_));
  NO2        g0703(.A(new_new_n381_), .B(i_2_), .Y(new_new_n726_));
  NA2        g0704(.A(new_new_n726_), .B(new_new_n725_), .Y(new_new_n727_));
  OAI210     g0705(.A0(new_new_n681_), .A1(new_new_n462_), .B0(new_new_n727_), .Y(new_new_n728_));
  INV        g0706(.A(new_new_n728_), .Y(new_new_n729_));
  AOI210     g0707(.A0(new_new_n729_), .A1(new_new_n724_), .B0(i_13_), .Y(new_new_n730_));
  OR2        g0708(.A(i_11_), .B(i_7_), .Y(new_new_n731_));
  NA3        g0709(.A(new_new_n731_), .B(new_new_n104_), .C(new_new_n137_), .Y(new_new_n732_));
  AOI220     g0710(.A0(new_new_n482_), .A1(new_new_n161_), .B0(i_2_), .B1(new_new_n137_), .Y(new_new_n733_));
  OAI210     g0711(.A0(new_new_n733_), .A1(new_new_n44_), .B0(new_new_n732_), .Y(new_new_n734_));
  AOI210     g0712(.A0(new_new_n677_), .A1(new_new_n52_), .B0(i_12_), .Y(new_new_n735_));
  INV        g0713(.A(new_new_n735_), .Y(new_new_n736_));
  NO2        g0714(.A(new_new_n489_), .B(new_new_n24_), .Y(new_new_n737_));
  AOI220     g0715(.A0(new_new_n737_), .A1(new_new_n696_), .B0(new_new_n247_), .B1(new_new_n130_), .Y(new_new_n738_));
  OAI220     g0716(.A0(new_new_n738_), .A1(new_new_n40_), .B0(new_new_n736_), .B1(new_new_n90_), .Y(new_new_n739_));
  AOI210     g0717(.A0(new_new_n734_), .A1(new_new_n339_), .B0(new_new_n739_), .Y(new_new_n740_));
  NA2        g0718(.A(new_new_n113_), .B(new_new_n106_), .Y(new_new_n741_));
  AOI220     g0719(.A0(new_new_n741_), .A1(new_new_n67_), .B0(new_new_n397_), .B1(new_new_n678_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n742_), .B(new_new_n244_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n462_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n744_));
  NOi31      g0722(.An(new_new_n744_), .B(new_new_n624_), .C(new_new_n44_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n126_), .B(i_13_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n677_), .B(new_new_n113_), .Y(new_new_n747_));
  INV        g0725(.A(new_new_n747_), .Y(new_new_n748_));
  OAI220     g0726(.A0(new_new_n748_), .A1(new_new_n66_), .B0(new_new_n746_), .B1(new_new_n725_), .Y(new_new_n749_));
  NO3        g0727(.A(new_new_n66_), .B(new_new_n32_), .C(new_new_n99_), .Y(new_new_n750_));
  NA2        g0728(.A(new_new_n26_), .B(new_new_n193_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n751_), .B(i_7_), .Y(new_new_n752_));
  NO3        g0730(.A(new_new_n489_), .B(new_new_n238_), .C(new_new_n81_), .Y(new_new_n753_));
  AOI210     g0731(.A0(new_new_n753_), .A1(new_new_n752_), .B0(new_new_n750_), .Y(new_new_n754_));
  AOI220     g0732(.A0(new_new_n397_), .A1(new_new_n678_), .B0(new_new_n89_), .B1(new_new_n100_), .Y(new_new_n755_));
  OAI220     g0733(.A0(new_new_n755_), .A1(new_new_n630_), .B0(new_new_n754_), .B1(new_new_n641_), .Y(new_new_n756_));
  NO4        g0734(.A(new_new_n756_), .B(new_new_n749_), .C(new_new_n745_), .D(new_new_n743_), .Y(new_new_n757_));
  OR2        g0735(.A(i_11_), .B(i_6_), .Y(new_new_n758_));
  NA3        g0736(.A(new_new_n629_), .B(new_new_n751_), .C(i_7_), .Y(new_new_n759_));
  AOI210     g0737(.A0(new_new_n759_), .A1(new_new_n748_), .B0(new_new_n758_), .Y(new_new_n760_));
  NA3        g0738(.A(new_new_n421_), .B(new_new_n633_), .C(new_new_n95_), .Y(new_new_n761_));
  NA2        g0739(.A(new_new_n668_), .B(i_13_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n100_), .B(new_new_n751_), .Y(new_new_n763_));
  NAi21      g0741(.An(i_11_), .B(i_12_), .Y(new_new_n764_));
  NOi41      g0742(.An(new_new_n109_), .B(new_new_n764_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n765_));
  NO3        g0743(.A(new_new_n489_), .B(new_new_n608_), .C(new_new_n634_), .Y(new_new_n766_));
  AOI220     g0744(.A0(new_new_n766_), .A1(new_new_n317_), .B0(new_new_n765_), .B1(new_new_n763_), .Y(new_new_n767_));
  NA3        g0745(.A(new_new_n767_), .B(new_new_n762_), .C(new_new_n761_), .Y(new_new_n768_));
  OAI210     g0746(.A0(new_new_n768_), .A1(new_new_n760_), .B0(new_new_n60_), .Y(new_new_n769_));
  NO2        g0747(.A(i_2_), .B(i_12_), .Y(new_new_n770_));
  NA2        g0748(.A(new_new_n380_), .B(new_new_n770_), .Y(new_new_n771_));
  NA2        g0749(.A(i_8_), .B(new_new_n25_), .Y(new_new_n772_));
  NO3        g0750(.A(new_new_n772_), .B(new_new_n395_), .C(new_new_n629_), .Y(new_new_n773_));
  OAI210     g0751(.A0(new_new_n773_), .A1(new_new_n382_), .B0(new_new_n380_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n127_), .B(i_2_), .Y(new_new_n775_));
  NA2        g0753(.A(new_new_n775_), .B(new_new_n662_), .Y(new_new_n776_));
  NA3        g0754(.A(new_new_n776_), .B(new_new_n774_), .C(new_new_n771_), .Y(new_new_n777_));
  NA3        g0755(.A(new_new_n777_), .B(new_new_n45_), .C(new_new_n226_), .Y(new_new_n778_));
  NA4        g0756(.A(new_new_n778_), .B(new_new_n769_), .C(new_new_n757_), .D(new_new_n740_), .Y(new_new_n779_));
  OR4        g0757(.A(new_new_n779_), .B(new_new_n730_), .C(new_new_n714_), .D(new_new_n644_), .Y(men5));
  AOI210     g0758(.A0(new_new_n693_), .A1(new_new_n273_), .B0(new_new_n430_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n630_), .B(i_11_), .Y(new_new_n782_));
  OAI210     g0760(.A0(new_new_n633_), .A1(new_new_n84_), .B0(new_new_n782_), .Y(new_new_n783_));
  NA3        g0761(.A(new_new_n783_), .B(new_new_n781_), .C(new_new_n538_), .Y(new_new_n784_));
  NO3        g0762(.A(i_11_), .B(new_new_n238_), .C(i_13_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n123_), .B(new_new_n23_), .Y(new_new_n786_));
  NA2        g0764(.A(i_12_), .B(i_8_), .Y(new_new_n787_));
  OAI210     g0765(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n787_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n461_), .Y(new_new_n789_));
  AOI220     g0767(.A0(new_new_n323_), .A1(new_new_n600_), .B0(new_new_n788_), .B1(new_new_n786_), .Y(new_new_n790_));
  INV        g0768(.A(new_new_n790_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n791_), .B(new_new_n784_), .Y(new_new_n792_));
  INV        g0770(.A(new_new_n171_), .Y(new_new_n793_));
  INV        g0771(.A(new_new_n247_), .Y(new_new_n794_));
  OAI210     g0772(.A0(new_new_n726_), .A1(new_new_n463_), .B0(new_new_n109_), .Y(new_new_n795_));
  AOI210     g0773(.A0(new_new_n795_), .A1(new_new_n794_), .B0(new_new_n793_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n471_), .B(new_new_n26_), .Y(new_new_n797_));
  NO2        g0775(.A(new_new_n797_), .B(new_new_n431_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n798_), .B(i_2_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n799_), .Y(new_new_n800_));
  AOI210     g0778(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n428_), .Y(new_new_n801_));
  AOI210     g0779(.A0(new_new_n801_), .A1(new_new_n800_), .B0(new_new_n796_), .Y(new_new_n802_));
  NO2        g0780(.A(new_new_n190_), .B(new_new_n124_), .Y(new_new_n803_));
  OAI210     g0781(.A0(new_new_n803_), .A1(new_new_n786_), .B0(i_2_), .Y(new_new_n804_));
  INV        g0782(.A(new_new_n172_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n805_), .B(new_new_n84_), .Y(new_new_n806_));
  AOI210     g0784(.A0(new_new_n806_), .A1(new_new_n804_), .B0(new_new_n193_), .Y(new_new_n807_));
  OA210      g0785(.A0(new_new_n647_), .A1(new_new_n125_), .B0(i_13_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n200_), .B(new_new_n203_), .Y(new_new_n809_));
  NA2        g0787(.A(new_new_n151_), .B(new_new_n625_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n810_), .A1(new_new_n809_), .B0(new_new_n385_), .Y(new_new_n811_));
  AOI210     g0789(.A0(new_new_n208_), .A1(new_new_n147_), .B0(new_new_n536_), .Y(new_new_n812_));
  OAI210     g0790(.A0(new_new_n812_), .A1(new_new_n227_), .B0(new_new_n431_), .Y(new_new_n813_));
  NO2        g0791(.A(new_new_n100_), .B(new_new_n44_), .Y(new_new_n814_));
  INV        g0792(.A(new_new_n307_), .Y(new_new_n815_));
  NA4        g0793(.A(new_new_n815_), .B(new_new_n310_), .C(new_new_n123_), .D(new_new_n42_), .Y(new_new_n816_));
  OAI210     g0794(.A0(new_new_n816_), .A1(new_new_n814_), .B0(new_new_n813_), .Y(new_new_n817_));
  NO4        g0795(.A(new_new_n817_), .B(new_new_n811_), .C(new_new_n808_), .D(new_new_n807_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n600_), .B(new_new_n28_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n785_), .B(new_new_n279_), .Y(new_new_n820_));
  NA2        g0798(.A(new_new_n820_), .B(new_new_n819_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n59_), .B(i_12_), .Y(new_new_n822_));
  NO2        g0800(.A(new_new_n822_), .B(new_new_n125_), .Y(new_new_n823_));
  NO2        g0801(.A(new_new_n823_), .B(new_new_n625_), .Y(new_new_n824_));
  AOI220     g0802(.A0(new_new_n824_), .A1(new_new_n36_), .B0(new_new_n821_), .B1(new_new_n46_), .Y(new_new_n825_));
  NA4        g0803(.A(new_new_n825_), .B(new_new_n818_), .C(new_new_n802_), .D(new_new_n792_), .Y(men6));
  NO3        g0804(.A(new_new_n258_), .B(new_new_n312_), .C(i_1_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n185_), .B(new_new_n138_), .Y(new_new_n828_));
  OAI210     g0806(.A0(new_new_n828_), .A1(new_new_n827_), .B0(new_new_n775_), .Y(new_new_n829_));
  NA4        g0807(.A(new_new_n401_), .B(new_new_n494_), .C(new_new_n66_), .D(new_new_n99_), .Y(new_new_n830_));
  INV        g0808(.A(new_new_n830_), .Y(new_new_n831_));
  NO2        g0809(.A(new_new_n221_), .B(new_new_n499_), .Y(new_new_n832_));
  NO2        g0810(.A(i_11_), .B(i_9_), .Y(new_new_n833_));
  NO3        g0811(.A(new_new_n832_), .B(new_new_n831_), .C(new_new_n334_), .Y(new_new_n834_));
  AO210      g0812(.A0(new_new_n834_), .A1(new_new_n829_), .B0(i_12_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n386_), .B(new_new_n342_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n608_), .B(new_new_n60_), .Y(new_new_n837_));
  NA2        g0815(.A(new_new_n716_), .B(new_new_n66_), .Y(new_new_n838_));
  NA4        g0816(.A(new_new_n652_), .B(new_new_n838_), .C(new_new_n837_), .D(new_new_n836_), .Y(new_new_n839_));
  INV        g0817(.A(new_new_n197_), .Y(new_new_n840_));
  AOI220     g0818(.A0(new_new_n840_), .A1(new_new_n833_), .B0(new_new_n839_), .B1(new_new_n68_), .Y(new_new_n841_));
  INV        g0819(.A(new_new_n333_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n70_), .B(new_new_n130_), .Y(new_new_n843_));
  INV        g0821(.A(new_new_n123_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n844_), .B(new_new_n46_), .Y(new_new_n845_));
  AOI210     g0823(.A0(new_new_n845_), .A1(new_new_n843_), .B0(new_new_n842_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n32_), .B(i_11_), .Y(new_new_n847_));
  NA3        g0825(.A(new_new_n847_), .B(new_new_n485_), .C(new_new_n401_), .Y(new_new_n848_));
  NAi32      g0826(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n849_));
  AOI210     g0827(.A0(new_new_n758_), .A1(new_new_n82_), .B0(new_new_n849_), .Y(new_new_n850_));
  OAI210     g0828(.A0(new_new_n715_), .A1(new_new_n588_), .B0(new_new_n587_), .Y(new_new_n851_));
  NAi31      g0829(.An(new_new_n850_), .B(new_new_n851_), .C(new_new_n848_), .Y(new_new_n852_));
  OR2        g0830(.A(new_new_n852_), .B(new_new_n846_), .Y(new_new_n853_));
  AO220      g0831(.A0(new_new_n369_), .A1(new_new_n359_), .B0(new_new_n408_), .B1(new_new_n625_), .Y(new_new_n854_));
  NA3        g0832(.A(new_new_n854_), .B(new_new_n259_), .C(i_7_), .Y(new_new_n855_));
  OR2        g0833(.A(new_new_n647_), .B(new_new_n463_), .Y(new_new_n856_));
  NA3        g0834(.A(new_new_n856_), .B(new_new_n146_), .C(new_new_n64_), .Y(new_new_n857_));
  AO210      g0835(.A0(new_new_n505_), .A1(new_new_n789_), .B0(new_new_n36_), .Y(new_new_n858_));
  NA3        g0836(.A(new_new_n858_), .B(new_new_n857_), .C(new_new_n855_), .Y(new_new_n859_));
  OAI210     g0837(.A0(i_6_), .A1(i_11_), .B0(new_new_n82_), .Y(new_new_n860_));
  AOI220     g0838(.A0(new_new_n860_), .A1(new_new_n587_), .B0(new_new_n832_), .B1(new_new_n752_), .Y(new_new_n861_));
  NA3        g0839(.A(new_new_n385_), .B(new_new_n240_), .C(new_new_n146_), .Y(new_new_n862_));
  OAI210     g0840(.A0(new_new_n408_), .A1(new_new_n204_), .B0(new_new_n65_), .Y(new_new_n863_));
  NA4        g0841(.A(new_new_n863_), .B(new_new_n862_), .C(new_new_n861_), .D(new_new_n632_), .Y(new_new_n864_));
  AO210      g0842(.A0(new_new_n536_), .A1(new_new_n46_), .B0(new_new_n83_), .Y(new_new_n865_));
  NA3        g0843(.A(new_new_n865_), .B(new_new_n495_), .C(new_new_n218_), .Y(new_new_n866_));
  AOI210     g0844(.A0(new_new_n463_), .A1(new_new_n461_), .B0(new_new_n586_), .Y(new_new_n867_));
  NO2        g0845(.A(new_new_n637_), .B(new_new_n100_), .Y(new_new_n868_));
  OAI210     g0846(.A0(new_new_n868_), .A1(new_new_n110_), .B0(new_new_n420_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n246_), .B(new_new_n46_), .Y(new_new_n870_));
  NA2        g0848(.A(new_new_n870_), .B(new_new_n615_), .Y(new_new_n871_));
  NA3        g0849(.A(new_new_n871_), .B(new_new_n333_), .C(i_7_), .Y(new_new_n872_));
  NA4        g0850(.A(new_new_n872_), .B(new_new_n869_), .C(new_new_n867_), .D(new_new_n866_), .Y(new_new_n873_));
  NO4        g0851(.A(new_new_n873_), .B(new_new_n864_), .C(new_new_n859_), .D(new_new_n853_), .Y(new_new_n874_));
  NA4        g0852(.A(new_new_n874_), .B(new_new_n841_), .C(new_new_n835_), .D(new_new_n391_), .Y(men3));
  NA2        g0853(.A(i_12_), .B(i_10_), .Y(new_new_n876_));
  NA2        g0854(.A(i_6_), .B(i_7_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n877_), .B(i_0_), .Y(new_new_n878_));
  NO2        g0856(.A(i_11_), .B(new_new_n238_), .Y(new_new_n879_));
  OAI210     g0857(.A0(new_new_n878_), .A1(new_new_n295_), .B0(new_new_n879_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n880_), .B(new_new_n193_), .Y(new_new_n881_));
  NO3        g0859(.A(new_new_n467_), .B(new_new_n87_), .C(new_new_n44_), .Y(new_new_n882_));
  OA210      g0860(.A0(new_new_n882_), .A1(new_new_n881_), .B0(new_new_n173_), .Y(new_new_n883_));
  NA3        g0861(.A(new_new_n862_), .B(new_new_n632_), .C(new_new_n384_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n884_), .B(new_new_n39_), .Y(new_new_n885_));
  NOi21      g0863(.An(new_new_n94_), .B(new_new_n798_), .Y(new_new_n886_));
  NO3        g0864(.A(new_new_n657_), .B(new_new_n471_), .C(new_new_n130_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n421_), .B(new_new_n45_), .Y(new_new_n888_));
  AN2        g0866(.A(new_new_n469_), .B(new_new_n53_), .Y(new_new_n889_));
  NO3        g0867(.A(new_new_n889_), .B(new_new_n887_), .C(new_new_n886_), .Y(new_new_n890_));
  AOI210     g0868(.A0(new_new_n890_), .A1(new_new_n885_), .B0(new_new_n48_), .Y(new_new_n891_));
  NO4        g0869(.A(new_new_n389_), .B(new_new_n394_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n892_));
  NA2        g0870(.A(new_new_n185_), .B(new_new_n596_), .Y(new_new_n893_));
  NOi21      g0871(.An(new_new_n893_), .B(new_new_n892_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n744_), .B(new_new_n705_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n340_), .B(new_new_n451_), .Y(new_new_n896_));
  OAI220     g0874(.A0(new_new_n896_), .A1(new_new_n895_), .B0(new_new_n894_), .B1(new_new_n60_), .Y(new_new_n897_));
  NOi21      g0875(.An(i_5_), .B(i_9_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n898_), .B(new_new_n459_), .Y(new_new_n899_));
  AOI210     g0877(.A0(new_new_n270_), .A1(new_new_n487_), .B0(new_new_n720_), .Y(new_new_n900_));
  NO3        g0878(.A(new_new_n424_), .B(new_new_n270_), .C(new_new_n68_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n174_), .B(new_new_n147_), .Y(new_new_n902_));
  AOI210     g0880(.A0(new_new_n902_), .A1(new_new_n246_), .B0(new_new_n901_), .Y(new_new_n903_));
  OAI220     g0881(.A0(new_new_n903_), .A1(new_new_n180_), .B0(new_new_n900_), .B1(new_new_n899_), .Y(new_new_n904_));
  NO4        g0882(.A(new_new_n904_), .B(new_new_n897_), .C(new_new_n891_), .D(new_new_n883_), .Y(new_new_n905_));
  NOi21      g0883(.An(i_0_), .B(i_10_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n185_), .B(new_new_n24_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n703_), .B(new_new_n622_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n908_), .B(new_new_n907_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n317_), .B(new_new_n128_), .Y(new_new_n910_));
  NAi21      g0888(.An(new_new_n162_), .B(new_new_n451_), .Y(new_new_n911_));
  OAI220     g0889(.A0(new_new_n911_), .A1(new_new_n870_), .B0(new_new_n910_), .B1(new_new_n411_), .Y(new_new_n912_));
  NO2        g0890(.A(new_new_n912_), .B(new_new_n909_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n401_), .B(new_new_n299_), .Y(new_new_n914_));
  NA2        g0892(.A(new_new_n914_), .B(new_new_n747_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n597_), .B(i_0_), .Y(new_new_n916_));
  NO3        g0894(.A(new_new_n916_), .B(new_new_n396_), .C(new_new_n84_), .Y(new_new_n917_));
  NO4        g0895(.A(new_new_n614_), .B(new_new_n215_), .C(new_new_n428_), .D(i_6_), .Y(new_new_n918_));
  AOI210     g0896(.A0(new_new_n918_), .A1(i_11_), .B0(new_new_n917_), .Y(new_new_n919_));
  INV        g0897(.A(new_new_n485_), .Y(new_new_n920_));
  AN2        g0898(.A(new_new_n94_), .B(new_new_n245_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n785_), .B(new_new_n334_), .Y(new_new_n922_));
  AOI210     g0900(.A0(new_new_n495_), .A1(new_new_n84_), .B0(new_new_n55_), .Y(new_new_n923_));
  OAI220     g0901(.A0(new_new_n923_), .A1(new_new_n922_), .B0(new_new_n688_), .B1(new_new_n556_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n256_), .B(new_new_n153_), .Y(new_new_n925_));
  NA2        g0903(.A(i_0_), .B(i_10_), .Y(new_new_n926_));
  OAI210     g0904(.A0(new_new_n926_), .A1(new_new_n81_), .B0(new_new_n559_), .Y(new_new_n927_));
  NO4        g0905(.A(new_new_n113_), .B(new_new_n55_), .C(new_new_n698_), .D(i_5_), .Y(new_new_n928_));
  AO220      g0906(.A0(new_new_n928_), .A1(new_new_n927_), .B0(new_new_n925_), .B1(i_6_), .Y(new_new_n929_));
  AOI220     g0907(.A0(new_new_n340_), .A1(new_new_n96_), .B0(new_new_n185_), .B1(new_new_n79_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n591_), .B(i_4_), .Y(new_new_n931_));
  NA2        g0909(.A(new_new_n188_), .B(new_new_n203_), .Y(new_new_n932_));
  OAI220     g0910(.A0(new_new_n932_), .A1(new_new_n922_), .B0(new_new_n931_), .B1(new_new_n930_), .Y(new_new_n933_));
  NO4        g0911(.A(new_new_n933_), .B(new_new_n929_), .C(new_new_n924_), .D(new_new_n921_), .Y(new_new_n934_));
  NA4        g0912(.A(new_new_n934_), .B(new_new_n919_), .C(new_new_n915_), .D(new_new_n913_), .Y(new_new_n935_));
  NO2        g0913(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n936_));
  NA2        g0914(.A(i_11_), .B(i_9_), .Y(new_new_n937_));
  NO3        g0915(.A(i_12_), .B(new_new_n937_), .C(new_new_n631_), .Y(new_new_n938_));
  AO220      g0916(.A0(new_new_n938_), .A1(new_new_n936_), .B0(new_new_n272_), .B1(new_new_n83_), .Y(new_new_n939_));
  NO2        g0917(.A(new_new_n48_), .B(i_7_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n405_), .B(new_new_n178_), .Y(new_new_n941_));
  NA2        g0919(.A(new_new_n941_), .B(new_new_n160_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n937_), .B(new_new_n68_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n174_), .B(i_0_), .Y(new_new_n944_));
  INV        g0922(.A(new_new_n944_), .Y(new_new_n945_));
  NA2        g0923(.A(new_new_n485_), .B(new_new_n232_), .Y(new_new_n946_));
  AOI210     g0924(.A0(new_new_n383_), .A1(new_new_n41_), .B0(new_new_n419_), .Y(new_new_n947_));
  OAI220     g0925(.A0(new_new_n947_), .A1(new_new_n899_), .B0(new_new_n946_), .B1(new_new_n945_), .Y(new_new_n948_));
  NO3        g0926(.A(new_new_n948_), .B(new_new_n942_), .C(new_new_n939_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n687_), .B(new_new_n120_), .Y(new_new_n950_));
  NO2        g0928(.A(i_6_), .B(new_new_n950_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n462_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n952_));
  NA2        g0930(.A(new_new_n171_), .B(new_new_n101_), .Y(new_new_n953_));
  NOi32      g0931(.An(new_new_n952_), .Bn(new_new_n188_), .C(new_new_n953_), .Y(new_new_n954_));
  AOI210     g0932(.A0(new_new_n633_), .A1(new_new_n334_), .B0(new_new_n245_), .Y(new_new_n955_));
  NO2        g0933(.A(new_new_n955_), .B(new_new_n888_), .Y(new_new_n956_));
  NO3        g0934(.A(new_new_n956_), .B(new_new_n954_), .C(new_new_n951_), .Y(new_new_n957_));
  NOi21      g0935(.An(i_7_), .B(i_5_), .Y(new_new_n958_));
  NOi31      g0936(.An(new_new_n958_), .B(new_new_n906_), .C(new_new_n764_), .Y(new_new_n959_));
  NA3        g0937(.A(new_new_n959_), .B(new_new_n395_), .C(i_6_), .Y(new_new_n960_));
  OA210      g0938(.A0(new_new_n953_), .A1(new_new_n534_), .B0(new_new_n960_), .Y(new_new_n961_));
  NO3        g0939(.A(new_new_n414_), .B(new_new_n372_), .C(new_new_n368_), .Y(new_new_n962_));
  NO2        g0940(.A(new_new_n266_), .B(new_new_n324_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n764_), .B(new_new_n261_), .Y(new_new_n964_));
  AOI210     g0942(.A0(new_new_n964_), .A1(new_new_n963_), .B0(new_new_n962_), .Y(new_new_n965_));
  NA4        g0943(.A(new_new_n965_), .B(new_new_n961_), .C(new_new_n957_), .D(new_new_n949_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n907_), .B(new_new_n241_), .Y(new_new_n967_));
  AN2        g0945(.A(new_new_n339_), .B(new_new_n334_), .Y(new_new_n968_));
  AO220      g0946(.A0(new_new_n968_), .A1(new_new_n902_), .B0(new_new_n354_), .B1(new_new_n27_), .Y(new_new_n969_));
  OAI210     g0947(.A0(new_new_n969_), .A1(new_new_n967_), .B0(i_10_), .Y(new_new_n970_));
  INV        g0948(.A(new_new_n876_), .Y(new_new_n971_));
  OA210      g0949(.A0(new_new_n485_), .A1(new_new_n224_), .B0(new_new_n484_), .Y(new_new_n972_));
  OAI210     g0950(.A0(new_new_n972_), .A1(new_new_n971_), .B0(new_new_n943_), .Y(new_new_n973_));
  NA3        g0951(.A(new_new_n484_), .B(new_new_n421_), .C(new_new_n45_), .Y(new_new_n974_));
  OAI210     g0952(.A0(new_new_n911_), .A1(new_new_n920_), .B0(new_new_n974_), .Y(new_new_n975_));
  NO2        g0953(.A(new_new_n259_), .B(new_new_n46_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n943_), .B(new_new_n310_), .Y(new_new_n977_));
  OAI210     g0955(.A0(new_new_n976_), .A1(new_new_n187_), .B0(new_new_n977_), .Y(new_new_n978_));
  AOI220     g0956(.A0(new_new_n978_), .A1(new_new_n485_), .B0(new_new_n975_), .B1(new_new_n68_), .Y(new_new_n979_));
  NA3        g0957(.A(i_5_), .B(new_new_n393_), .C(i_6_), .Y(new_new_n980_));
  NA2        g0958(.A(new_new_n90_), .B(new_new_n44_), .Y(new_new_n981_));
  NO2        g0959(.A(new_new_n70_), .B(new_new_n787_), .Y(new_new_n982_));
  AOI220     g0960(.A0(new_new_n982_), .A1(new_new_n981_), .B0(new_new_n173_), .B1(new_new_n622_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n983_), .A1(new_new_n980_), .B0(new_new_n47_), .Y(new_new_n984_));
  NO3        g0962(.A(new_new_n614_), .B(new_new_n367_), .C(new_new_n24_), .Y(new_new_n985_));
  AOI210     g0963(.A0(new_new_n737_), .A1(new_new_n568_), .B0(new_new_n985_), .Y(new_new_n986_));
  NAi21      g0964(.An(i_9_), .B(i_5_), .Y(new_new_n987_));
  NO2        g0965(.A(new_new_n987_), .B(new_new_n414_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n628_), .B(new_new_n103_), .Y(new_new_n989_));
  AOI220     g0967(.A0(new_new_n989_), .A1(i_0_), .B0(new_new_n988_), .B1(new_new_n647_), .Y(new_new_n990_));
  OAI220     g0968(.A0(new_new_n990_), .A1(new_new_n81_), .B0(new_new_n986_), .B1(new_new_n172_), .Y(new_new_n991_));
  NO3        g0969(.A(new_new_n991_), .B(new_new_n984_), .C(new_new_n539_), .Y(new_new_n992_));
  NA4        g0970(.A(new_new_n992_), .B(new_new_n979_), .C(new_new_n973_), .D(new_new_n970_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n993_), .B(new_new_n966_), .C(new_new_n935_), .Y(new_new_n994_));
  NO2        g0972(.A(new_new_n906_), .B(new_new_n764_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n68_), .B(new_new_n44_), .Y(new_new_n996_));
  NO3        g0974(.A(new_new_n103_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n997_));
  AO220      g0975(.A0(new_new_n997_), .A1(new_new_n44_), .B0(new_new_n995_), .B1(new_new_n173_), .Y(new_new_n998_));
  AOI210     g0976(.A0(new_new_n837_), .A1(new_new_n718_), .B0(new_new_n953_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n998_), .A1(new_new_n356_), .B0(new_new_n999_), .Y(new_new_n1000_));
  NA2        g0978(.A(new_new_n775_), .B(new_new_n145_), .Y(new_new_n1001_));
  INV        g0979(.A(new_new_n1001_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n1002_), .B(new_new_n705_), .C(new_new_n68_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n851_), .B(new_new_n414_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n878_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n879_), .B(i_9_), .Y(new_new_n1006_));
  AOI210     g0984(.A0(new_new_n1005_), .A1(new_new_n511_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n246_), .A1(i_9_), .B0(new_new_n231_), .Y(new_new_n1008_));
  AOI210     g0986(.A0(new_new_n1008_), .A1(new_new_n916_), .B0(new_new_n153_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n1009_), .B(new_new_n1007_), .C(new_new_n1004_), .Y(new_new_n1010_));
  NA3        g0988(.A(new_new_n1010_), .B(new_new_n1003_), .C(new_new_n1000_), .Y(new_new_n1011_));
  NA2        g0989(.A(new_new_n968_), .B(new_new_n385_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n306_), .A1(new_new_n162_), .B0(new_new_n1012_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n1014_));
  NA2        g0992(.A(new_new_n940_), .B(new_new_n500_), .Y(new_new_n1015_));
  AOI210     g0993(.A0(new_new_n1014_), .A1(new_new_n162_), .B0(new_new_n1015_), .Y(new_new_n1016_));
  NO2        g0994(.A(new_new_n1016_), .B(new_new_n1013_), .Y(new_new_n1017_));
  NA2        g0995(.A(new_new_n592_), .B(new_new_n70_), .Y(new_new_n1018_));
  NO3        g0996(.A(new_new_n209_), .B(new_new_n394_), .C(i_0_), .Y(new_new_n1019_));
  OAI210     g0997(.A0(new_new_n1019_), .A1(new_new_n71_), .B0(i_13_), .Y(new_new_n1020_));
  INV        g0998(.A(new_new_n218_), .Y(new_new_n1021_));
  OAI220     g0999(.A0(new_new_n550_), .A1(new_new_n138_), .B0(i_12_), .B1(new_new_n641_), .Y(new_new_n1022_));
  NA3        g1000(.A(new_new_n1022_), .B(new_new_n409_), .C(new_new_n1021_), .Y(new_new_n1023_));
  NA4        g1001(.A(new_new_n1023_), .B(new_new_n1020_), .C(new_new_n1018_), .D(new_new_n1017_), .Y(new_new_n1024_));
  NO2        g1002(.A(new_new_n244_), .B(new_new_n90_), .Y(new_new_n1025_));
  AOI210     g1003(.A0(new_new_n1025_), .A1(new_new_n995_), .B0(new_new_n107_), .Y(new_new_n1026_));
  AOI220     g1004(.A0(new_new_n958_), .A1(new_new_n500_), .B0(new_new_n878_), .B1(new_new_n163_), .Y(new_new_n1027_));
  NA2        g1005(.A(new_new_n359_), .B(new_new_n175_), .Y(new_new_n1028_));
  OA220      g1006(.A0(new_new_n1028_), .A1(new_new_n1027_), .B0(new_new_n1026_), .B1(i_5_), .Y(new_new_n1029_));
  AOI210     g1007(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n174_), .Y(new_new_n1030_));
  NA2        g1008(.A(new_new_n1030_), .B(new_new_n972_), .Y(new_new_n1031_));
  NA3        g1009(.A(new_new_n638_), .B(new_new_n185_), .C(new_new_n79_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n1032_), .B(new_new_n566_), .Y(new_new_n1033_));
  NO3        g1011(.A(new_new_n888_), .B(new_new_n52_), .C(new_new_n48_), .Y(new_new_n1034_));
  NA2        g1012(.A(new_new_n504_), .B(new_new_n498_), .Y(new_new_n1035_));
  NO3        g1013(.A(new_new_n1035_), .B(new_new_n1034_), .C(new_new_n1033_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n940_), .B(new_new_n295_), .C(new_new_n231_), .Y(new_new_n1037_));
  INV        g1015(.A(new_new_n1037_), .Y(new_new_n1038_));
  NA3        g1016(.A(new_new_n401_), .B(new_new_n341_), .C(new_new_n222_), .Y(new_new_n1039_));
  OAI210     g1017(.A0(new_new_n893_), .A1(new_new_n675_), .B0(new_new_n1039_), .Y(new_new_n1040_));
  NOi31      g1018(.An(new_new_n400_), .B(new_new_n996_), .C(new_new_n241_), .Y(new_new_n1041_));
  NO3        g1019(.A(new_new_n1041_), .B(new_new_n1040_), .C(new_new_n1038_), .Y(new_new_n1042_));
  NA4        g1020(.A(new_new_n1042_), .B(new_new_n1036_), .C(new_new_n1031_), .D(new_new_n1029_), .Y(new_new_n1043_));
  INV        g1021(.A(new_new_n640_), .Y(new_new_n1044_));
  NO3        g1022(.A(new_new_n1044_), .B(new_new_n582_), .C(new_new_n353_), .Y(new_new_n1045_));
  NO2        g1023(.A(new_new_n81_), .B(i_5_), .Y(new_new_n1046_));
  NA3        g1024(.A(new_new_n879_), .B(new_new_n108_), .C(new_new_n123_), .Y(new_new_n1047_));
  INV        g1025(.A(new_new_n1047_), .Y(new_new_n1048_));
  AOI210     g1026(.A0(new_new_n1048_), .A1(new_new_n1046_), .B0(new_new_n1045_), .Y(new_new_n1049_));
  NA3        g1027(.A(new_new_n310_), .B(i_5_), .C(new_new_n193_), .Y(new_new_n1050_));
  NO4        g1028(.A(new_new_n241_), .B(new_new_n209_), .C(i_0_), .D(i_12_), .Y(new_new_n1051_));
  AOI220     g1029(.A0(new_new_n1051_), .A1(i_10_), .B0(new_new_n831_), .B1(new_new_n175_), .Y(new_new_n1052_));
  AN2        g1030(.A(new_new_n926_), .B(new_new_n153_), .Y(new_new_n1053_));
  NO4        g1031(.A(new_new_n1053_), .B(i_12_), .C(new_new_n675_), .D(new_new_n130_), .Y(new_new_n1054_));
  NA2        g1032(.A(new_new_n1054_), .B(new_new_n218_), .Y(new_new_n1055_));
  NA3        g1033(.A(new_new_n96_), .B(new_new_n596_), .C(i_11_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n1056_), .B(new_new_n155_), .Y(new_new_n1057_));
  NA2        g1035(.A(new_new_n958_), .B(new_new_n482_), .Y(new_new_n1058_));
  NA2        g1036(.A(new_new_n61_), .B(new_new_n99_), .Y(new_new_n1059_));
  OAI220     g1037(.A0(new_new_n1059_), .A1(new_new_n1050_), .B0(new_new_n1058_), .B1(new_new_n706_), .Y(new_new_n1060_));
  AOI210     g1038(.A0(new_new_n1060_), .A1(new_new_n944_), .B0(new_new_n1057_), .Y(new_new_n1061_));
  NA4        g1039(.A(new_new_n1061_), .B(new_new_n1055_), .C(new_new_n1052_), .D(new_new_n1049_), .Y(new_new_n1062_));
  NO4        g1040(.A(new_new_n1062_), .B(new_new_n1043_), .C(new_new_n1024_), .D(new_new_n1011_), .Y(new_new_n1063_));
  NA2        g1041(.A(new_new_n847_), .B(new_new_n37_), .Y(new_new_n1064_));
  NA3        g1042(.A(new_new_n952_), .B(new_new_n380_), .C(i_5_), .Y(new_new_n1065_));
  NA3        g1043(.A(new_new_n1065_), .B(new_new_n1064_), .C(new_new_n636_), .Y(new_new_n1066_));
  NA2        g1044(.A(new_new_n1066_), .B(new_new_n207_), .Y(new_new_n1067_));
  AN2        g1045(.A(new_new_n731_), .B(new_new_n381_), .Y(new_new_n1068_));
  NA2        g1046(.A(new_new_n186_), .B(new_new_n188_), .Y(new_new_n1069_));
  AO210      g1047(.A0(new_new_n1068_), .A1(new_new_n33_), .B0(new_new_n1069_), .Y(new_new_n1070_));
  OAI210     g1048(.A0(new_new_n640_), .A1(new_new_n638_), .B0(new_new_n323_), .Y(new_new_n1071_));
  NAi31      g1049(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1072_));
  AOI210     g1050(.A0(new_new_n116_), .A1(new_new_n65_), .B0(new_new_n1072_), .Y(new_new_n1073_));
  NO2        g1051(.A(new_new_n1073_), .B(new_new_n672_), .Y(new_new_n1074_));
  NA3        g1052(.A(new_new_n1074_), .B(new_new_n1071_), .C(new_new_n1070_), .Y(new_new_n1075_));
  NO2        g1053(.A(new_new_n475_), .B(new_new_n270_), .Y(new_new_n1076_));
  NO4        g1054(.A(new_new_n234_), .B(new_new_n144_), .C(new_new_n709_), .D(new_new_n37_), .Y(new_new_n1077_));
  NO3        g1055(.A(new_new_n1077_), .B(new_new_n1076_), .C(new_new_n918_), .Y(new_new_n1078_));
  OAI210     g1056(.A0(new_new_n1056_), .A1(new_new_n147_), .B0(new_new_n1078_), .Y(new_new_n1079_));
  AOI210     g1057(.A0(new_new_n1075_), .A1(new_new_n48_), .B0(new_new_n1079_), .Y(new_new_n1080_));
  AOI210     g1058(.A0(new_new_n1080_), .A1(new_new_n1067_), .B0(new_new_n68_), .Y(new_new_n1081_));
  NO2        g1059(.A(new_new_n1116_), .B(new_new_n793_), .Y(new_new_n1082_));
  OAI210     g1060(.A0(new_new_n75_), .A1(new_new_n52_), .B0(new_new_n106_), .Y(new_new_n1083_));
  NA2        g1061(.A(new_new_n1083_), .B(new_new_n71_), .Y(new_new_n1084_));
  AOI210     g1062(.A0(new_new_n1030_), .A1(new_new_n940_), .B0(new_new_n959_), .Y(new_new_n1085_));
  AOI210     g1063(.A0(new_new_n1085_), .A1(new_new_n1084_), .B0(new_new_n709_), .Y(new_new_n1086_));
  NA2        g1064(.A(new_new_n266_), .B(new_new_n54_), .Y(new_new_n1087_));
  AOI220     g1065(.A0(new_new_n1087_), .A1(new_new_n71_), .B0(new_new_n354_), .B1(new_new_n258_), .Y(new_new_n1088_));
  NO2        g1066(.A(new_new_n1088_), .B(new_new_n238_), .Y(new_new_n1089_));
  NA3        g1067(.A(new_new_n94_), .B(new_new_n312_), .C(new_new_n31_), .Y(new_new_n1090_));
  INV        g1068(.A(new_new_n1090_), .Y(new_new_n1091_));
  NO3        g1069(.A(new_new_n1091_), .B(new_new_n1089_), .C(new_new_n1086_), .Y(new_new_n1092_));
  OAI210     g1070(.A0(new_new_n272_), .A1(new_new_n158_), .B0(new_new_n84_), .Y(new_new_n1093_));
  NA3        g1071(.A(new_new_n797_), .B(new_new_n295_), .C(new_new_n75_), .Y(new_new_n1094_));
  AOI210     g1072(.A0(new_new_n1094_), .A1(new_new_n1093_), .B0(i_11_), .Y(new_new_n1095_));
  NA2        g1073(.A(new_new_n634_), .B(new_new_n215_), .Y(new_new_n1096_));
  OAI210     g1074(.A0(new_new_n1096_), .A1(new_new_n952_), .B0(new_new_n207_), .Y(new_new_n1097_));
  NA2        g1075(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1098_));
  AOI210     g1076(.A0(new_new_n1097_), .A1(new_new_n809_), .B0(new_new_n1098_), .Y(new_new_n1099_));
  NO3        g1077(.A(new_new_n56_), .B(new_new_n55_), .C(i_4_), .Y(new_new_n1100_));
  OAI210     g1078(.A0(new_new_n963_), .A1(new_new_n312_), .B0(new_new_n1100_), .Y(new_new_n1101_));
  NO2        g1079(.A(new_new_n1101_), .B(new_new_n764_), .Y(new_new_n1102_));
  NO4        g1080(.A(new_new_n987_), .B(new_new_n488_), .C(new_new_n255_), .D(new_new_n254_), .Y(new_new_n1103_));
  NO2        g1081(.A(new_new_n1103_), .B(new_new_n586_), .Y(new_new_n1104_));
  NO2        g1082(.A(new_new_n850_), .B(new_new_n373_), .Y(new_new_n1105_));
  AOI210     g1083(.A0(new_new_n1105_), .A1(new_new_n1104_), .B0(new_new_n40_), .Y(new_new_n1106_));
  NO4        g1084(.A(new_new_n1106_), .B(new_new_n1102_), .C(new_new_n1099_), .D(new_new_n1095_), .Y(new_new_n1107_));
  OAI210     g1085(.A0(new_new_n1092_), .A1(i_4_), .B0(new_new_n1107_), .Y(new_new_n1108_));
  NO3        g1086(.A(new_new_n1108_), .B(new_new_n1082_), .C(new_new_n1081_), .Y(new_new_n1109_));
  NA4        g1087(.A(new_new_n1109_), .B(new_new_n1063_), .C(new_new_n994_), .D(new_new_n905_), .Y(men4));
  INV        g1088(.A(i_2_), .Y(new_new_n1113_));
  INV        g1089(.A(i_5_), .Y(new_new_n1114_));
  INV        g1090(.A(i_3_), .Y(new_new_n1115_));
  INV        g1091(.A(new_new_n589_), .Y(new_new_n1116_));
endmodule


