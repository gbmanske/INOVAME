//Benchmark atmr_5xp1_76_0.25

module atmr_5xp1(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n57_, ori_ori_n61_, ori_ori_n62_, ori_ori_n64_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n54_, mai_mai_n55_, mai_mai_n57_, mai_mai_n61_, mai_mai_n62_, mai_mai_n64_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n61_, men_men_n62_, men_men_n64_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09;
  INV        o00(.A(i_5_), .Y(ori_ori_n18_));
  NO3        o01(.A(i_4_), .B(i_6_), .C(ori_ori_n18_), .Y(ori_ori_n19_));
  INV        o02(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o03(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n21_));
  INV        o04(.A(i_1_), .Y(ori_ori_n22_));
  AOI210     o05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(ori_ori_n23_));
  NA2        o06(.A(ori_ori_n23_), .B(ori_ori_n22_), .Y(ori_ori_n24_));
  NO2        o07(.A(ori_ori_n24_), .B(ori_ori_n21_), .Y(ori_ori_n25_));
  INV        o08(.A(i_6_), .Y(ori_ori_n26_));
  NO2        o09(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n27_));
  INV        o10(.A(i_0_), .Y(ori_ori_n28_));
  NO2        o11(.A(i_2_), .B(i_1_), .Y(ori_ori_n29_));
  OAI210     o12(.A0(ori_ori_n29_), .A1(ori_ori_n28_), .B0(ori_ori_n20_), .Y(ori_ori_n30_));
  NO2        o13(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n31_));
  NO2        o14(.A(i_2_), .B(i_3_), .Y(ori_ori_n32_));
  NO3        o15(.A(ori_ori_n32_), .B(ori_ori_n28_), .C(ori_ori_n22_), .Y(ori_ori_n33_));
  AO220      o16(.A0(ori_ori_n33_), .A1(ori_ori_n31_), .B0(ori_ori_n30_), .B1(ori_ori_n27_), .Y(ori_ori_n34_));
  NA2        o17(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n35_));
  NA2        o18(.A(i_2_), .B(i_3_), .Y(ori_ori_n36_));
  NO2        o19(.A(ori_ori_n35_), .B(i_0_), .Y(ori_ori_n37_));
  OR4        o20(.A(ori_ori_n37_), .B(ori_ori_n34_), .C(ori_ori_n25_), .D(ori_ori_n19_), .Y(ori01));
  NA2        o21(.A(i_0_), .B(i_1_), .Y(ori_ori_n39_));
  NA2        o22(.A(ori_ori_n28_), .B(ori_ori_n18_), .Y(ori_ori_n40_));
  AOI210     o23(.A0(ori_ori_n23_), .A1(ori_ori_n22_), .B0(ori_ori_n26_), .Y(ori_ori_n41_));
  AOI220     o24(.A0(ori_ori_n41_), .A1(ori_ori_n40_), .B0(ori_ori_n39_), .B1(ori_ori_n26_), .Y(ori_ori_n42_));
  NO2        o25(.A(ori_ori_n35_), .B(ori_ori_n28_), .Y(ori_ori_n43_));
  NO3        o26(.A(ori_ori_n43_), .B(ori_ori_n42_), .C(i_4_), .Y(ori_ori_n44_));
  NA2        o27(.A(i_0_), .B(i_6_), .Y(ori_ori_n45_));
  NOi21      o28(.An(i_6_), .B(ori_ori_n18_), .Y(ori_ori_n46_));
  NO2        o29(.A(ori_ori_n45_), .B(ori_ori_n29_), .Y(ori_ori_n47_));
  NO3        o30(.A(ori_ori_n47_), .B(ori_ori_n46_), .C(ori_ori_n20_), .Y(ori_ori_n48_));
  NA2        o31(.A(ori_ori_n28_), .B(ori_ori_n26_), .Y(ori_ori_n49_));
  NO2        o32(.A(ori_ori_n49_), .B(ori_ori_n20_), .Y(ori_ori_n50_));
  INV        o33(.A(ori_ori_n50_), .Y(ori_ori_n51_));
  OAI210     o34(.A0(ori_ori_n48_), .A1(ori_ori_n44_), .B0(ori_ori_n51_), .Y(ori02));
  NAi21      o35(.An(ori_ori_n21_), .B(ori_ori_n41_), .Y(ori_ori_n53_));
  NA3        o36(.A(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n54_));
  NO2        o37(.A(ori_ori_n50_), .B(ori_ori_n31_), .Y(ori_ori_n55_));
  NA2        o38(.A(ori_ori_n55_), .B(ori_ori_n53_), .Y(ori00));
  NA2        o39(.A(ori_ori_n49_), .B(i_5_), .Y(ori_ori_n57_));
  NO2        o40(.A(ori_ori_n57_), .B(ori_ori_n20_), .Y(ori09));
  NOi21      o41(.An(ori_ori_n36_), .B(ori_ori_n32_), .Y(ori07));
  INV        o42(.A(i_3_), .Y(ori08));
  INV        o43(.A(ori_ori_n29_), .Y(ori_ori_n61_));
  NA2        o44(.A(ori07), .B(ori_ori_n61_), .Y(ori_ori_n62_));
  XO2        o45(.A(ori_ori_n62_), .B(ori_ori_n28_), .Y(ori05));
  NO2        o46(.A(i_2_), .B(ori08), .Y(ori_ori_n64_));
  XO2        o47(.A(ori_ori_n64_), .B(i_1_), .Y(ori06));
  NO2        o48(.A(i_1_), .B(i_6_), .Y(ori_ori_n66_));
  NO3        o49(.A(ori_ori_n66_), .B(ori_ori_n40_), .C(ori_ori_n36_), .Y(ori_ori_n67_));
  NO2        o50(.A(ori_ori_n67_), .B(ori_ori_n37_), .Y(ori_ori_n68_));
  AO210      o51(.A0(ori_ori_n39_), .A1(ori_ori_n24_), .B0(ori_ori_n18_), .Y(ori_ori_n69_));
  NA2        o52(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori03));
  NA2        o53(.A(ori_ori_n28_), .B(ori08), .Y(ori_ori_n71_));
  OAI210     o54(.A0(ori_ori_n71_), .A1(i_1_), .B0(ori_ori_n54_), .Y(ori_ori_n72_));
  OAI210     o55(.A0(ori_ori_n72_), .A1(ori_ori_n33_), .B0(i_6_), .Y(ori_ori_n73_));
  INV        o56(.A(ori_ori_n29_), .Y(ori_ori_n74_));
  OR2        o57(.A(ori_ori_n74_), .B(ori_ori_n66_), .Y(ori_ori_n75_));
  NA3        o58(.A(ori_ori_n71_), .B(ori_ori_n66_), .C(i_2_), .Y(ori_ori_n76_));
  NA3        o59(.A(ori_ori_n23_), .B(i_1_), .C(ori_ori_n26_), .Y(ori_ori_n77_));
  NA4        o60(.A(ori_ori_n77_), .B(ori_ori_n76_), .C(ori_ori_n75_), .D(ori_ori_n73_), .Y(ori04));
  INV        m00(.A(i_5_), .Y(mai_mai_n18_));
  NO3        m01(.A(i_4_), .B(i_6_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m02(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m03(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n21_));
  INV        m04(.A(i_1_), .Y(mai_mai_n22_));
  AOI210     m05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(mai_mai_n23_));
  NA2        m06(.A(mai_mai_n23_), .B(mai_mai_n22_), .Y(mai_mai_n24_));
  NO2        m07(.A(mai_mai_n24_), .B(mai_mai_n21_), .Y(mai_mai_n25_));
  INV        m08(.A(i_6_), .Y(mai_mai_n26_));
  NO2        m09(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n27_));
  INV        m10(.A(i_0_), .Y(mai_mai_n28_));
  NO2        m11(.A(i_2_), .B(i_1_), .Y(mai_mai_n29_));
  NO2        m12(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n30_));
  NO2        m13(.A(i_2_), .B(i_3_), .Y(mai_mai_n31_));
  NO3        m14(.A(mai_mai_n31_), .B(mai_mai_n28_), .C(mai_mai_n22_), .Y(mai_mai_n32_));
  AO210      m15(.A0(mai_mai_n32_), .A1(mai_mai_n30_), .B0(mai_mai_n27_), .Y(mai_mai_n33_));
  NA2        m16(.A(i_2_), .B(i_3_), .Y(mai_mai_n34_));
  OR3        m17(.A(mai_mai_n33_), .B(mai_mai_n25_), .C(mai_mai_n19_), .Y(mai01));
  OR2        m18(.A(i_2_), .B(i_3_), .Y(mai_mai_n36_));
  NA3        m19(.A(mai_mai_n36_), .B(i_0_), .C(i_1_), .Y(mai_mai_n37_));
  AOI210     m20(.A0(mai_mai_n23_), .A1(mai_mai_n22_), .B0(mai_mai_n26_), .Y(mai_mai_n38_));
  AOI210     m21(.A0(mai_mai_n37_), .A1(mai_mai_n26_), .B0(mai_mai_n38_), .Y(mai_mai_n39_));
  NA2        m22(.A(mai_mai_n29_), .B(mai_mai_n18_), .Y(mai_mai_n40_));
  NO2        m23(.A(mai_mai_n40_), .B(mai_mai_n26_), .Y(mai_mai_n41_));
  NO3        m24(.A(mai_mai_n41_), .B(mai_mai_n39_), .C(i_4_), .Y(mai_mai_n42_));
  NA2        m25(.A(i_0_), .B(i_6_), .Y(mai_mai_n43_));
  OAI210     m26(.A0(i_0_), .A1(i_1_), .B0(mai_mai_n43_), .Y(mai_mai_n44_));
  NOi31      m27(.An(mai_mai_n44_), .B(mai_mai_n23_), .C(mai_mai_n18_), .Y(mai_mai_n45_));
  NA3        m28(.A(i_1_), .B(i_6_), .C(i_5_), .Y(mai_mai_n46_));
  AOI210     m29(.A0(mai_mai_n46_), .A1(mai_mai_n43_), .B0(mai_mai_n29_), .Y(mai_mai_n47_));
  NO3        m30(.A(mai_mai_n36_), .B(i_6_), .C(i_5_), .Y(mai_mai_n48_));
  NO4        m31(.A(mai_mai_n48_), .B(mai_mai_n47_), .C(mai_mai_n45_), .D(mai_mai_n20_), .Y(mai_mai_n49_));
  AOI210     m32(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(mai_mai_n50_));
  AO220      m33(.A0(mai_mai_n50_), .A1(mai_mai_n30_), .B0(i_1_), .B1(mai_mai_n19_), .Y(mai_mai_n51_));
  INV        m34(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  OAI210     m35(.A0(mai_mai_n49_), .A1(mai_mai_n42_), .B0(mai_mai_n52_), .Y(mai02));
  NAi21      m36(.An(mai_mai_n21_), .B(mai_mai_n38_), .Y(mai_mai_n54_));
  INV        m37(.A(mai_mai_n30_), .Y(mai_mai_n55_));
  NA2        m38(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai00));
  INV        m39(.A(i_5_), .Y(mai_mai_n57_));
  NO2        m40(.A(mai_mai_n57_), .B(mai_mai_n20_), .Y(mai09));
  NOi21      m41(.An(mai_mai_n34_), .B(mai_mai_n31_), .Y(mai07));
  INV        m42(.A(i_3_), .Y(mai08));
  INV        m43(.A(mai_mai_n29_), .Y(mai_mai_n61_));
  NA2        m44(.A(mai07), .B(mai_mai_n61_), .Y(mai_mai_n62_));
  XO2        m45(.A(mai_mai_n62_), .B(mai_mai_n28_), .Y(mai05));
  NO2        m46(.A(i_2_), .B(mai08), .Y(mai_mai_n64_));
  XO2        m47(.A(mai_mai_n64_), .B(i_1_), .Y(mai06));
  NAi21      m48(.An(mai_mai_n48_), .B(mai_mai_n40_), .Y(mai_mai_n66_));
  NA2        m49(.A(mai_mai_n66_), .B(i_0_), .Y(mai_mai_n67_));
  NO2        m50(.A(i_1_), .B(i_6_), .Y(mai_mai_n68_));
  AO210      m51(.A0(mai_mai_n37_), .A1(mai_mai_n24_), .B0(mai_mai_n18_), .Y(mai_mai_n69_));
  NO2        m52(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n70_));
  NO2        m53(.A(mai_mai_n26_), .B(mai_mai_n18_), .Y(mai_mai_n71_));
  OAI210     m54(.A0(mai_mai_n22_), .A1(i_6_), .B0(mai_mai_n18_), .Y(mai_mai_n72_));
  NO2        m55(.A(mai_mai_n72_), .B(mai_mai_n44_), .Y(mai_mai_n73_));
  AOI210     m56(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n73_), .Y(mai_mai_n74_));
  NA3        m57(.A(mai_mai_n74_), .B(mai_mai_n69_), .C(mai_mai_n67_), .Y(mai03));
  NA2        m58(.A(mai_mai_n28_), .B(mai08), .Y(mai_mai_n76_));
  NO2        m59(.A(mai_mai_n76_), .B(i_1_), .Y(mai_mai_n77_));
  OAI210     m60(.A0(mai_mai_n77_), .A1(mai_mai_n32_), .B0(i_6_), .Y(mai_mai_n78_));
  AOI210     m61(.A0(mai_mai_n31_), .A1(mai_mai_n26_), .B0(mai_mai_n29_), .Y(mai_mai_n79_));
  OR2        m62(.A(mai_mai_n79_), .B(mai_mai_n68_), .Y(mai_mai_n80_));
  NA3        m63(.A(mai_mai_n76_), .B(mai_mai_n68_), .C(i_2_), .Y(mai_mai_n81_));
  NA3        m64(.A(mai_mai_n23_), .B(i_1_), .C(mai_mai_n26_), .Y(mai_mai_n82_));
  NA4        m65(.A(mai_mai_n82_), .B(mai_mai_n81_), .C(mai_mai_n80_), .D(mai_mai_n78_), .Y(mai04));
  INV        u00(.A(i_5_), .Y(men_men_n18_));
  NO3        u01(.A(i_4_), .B(i_6_), .C(men_men_n18_), .Y(men_men_n19_));
  INV        u02(.A(i_4_), .Y(men_men_n20_));
  NA2        u03(.A(men_men_n20_), .B(i_5_), .Y(men_men_n21_));
  INV        u04(.A(i_1_), .Y(men_men_n22_));
  INV        u05(.A(i_6_), .Y(men_men_n23_));
  NO2        u06(.A(men_men_n23_), .B(i_5_), .Y(men_men_n24_));
  INV        u07(.A(i_0_), .Y(men_men_n25_));
  NO2        u08(.A(i_2_), .B(i_1_), .Y(men_men_n26_));
  OAI210     u09(.A0(men_men_n26_), .A1(men_men_n25_), .B0(men_men_n20_), .Y(men_men_n27_));
  NO2        u10(.A(men_men_n20_), .B(i_5_), .Y(men_men_n28_));
  NO2        u11(.A(i_2_), .B(i_3_), .Y(men_men_n29_));
  NO3        u12(.A(men_men_n29_), .B(men_men_n25_), .C(men_men_n22_), .Y(men_men_n30_));
  AN2        u13(.A(men_men_n27_), .B(men_men_n24_), .Y(men_men_n31_));
  NA2        u14(.A(men_men_n23_), .B(i_5_), .Y(men_men_n32_));
  NA2        u15(.A(i_2_), .B(i_3_), .Y(men_men_n33_));
  NO2        u16(.A(men_men_n33_), .B(men_men_n22_), .Y(men_men_n34_));
  NO3        u17(.A(men_men_n34_), .B(men_men_n32_), .C(i_0_), .Y(men_men_n35_));
  OR3        u18(.A(men_men_n35_), .B(men_men_n31_), .C(men_men_n19_), .Y(men01));
  NA2        u19(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n37_));
  AOI210     u20(.A0(i_6_), .A1(men_men_n37_), .B0(men_men_n23_), .Y(men_men_n38_));
  NA2        u21(.A(men_men_n26_), .B(men_men_n18_), .Y(men_men_n39_));
  OAI220     u22(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n32_), .B1(men_men_n25_), .Y(men_men_n40_));
  NO3        u23(.A(men_men_n40_), .B(men_men_n38_), .C(i_4_), .Y(men_men_n41_));
  NA2        u24(.A(i_0_), .B(i_6_), .Y(men_men_n42_));
  OAI210     u25(.A0(i_0_), .A1(i_1_), .B0(men_men_n42_), .Y(men_men_n43_));
  NA3        u26(.A(i_1_), .B(i_6_), .C(i_5_), .Y(men_men_n44_));
  AOI210     u27(.A0(men_men_n44_), .A1(men_men_n42_), .B0(men_men_n26_), .Y(men_men_n45_));
  NO2        u28(.A(i_6_), .B(i_5_), .Y(men_men_n46_));
  NO3        u29(.A(men_men_n46_), .B(men_men_n45_), .C(men_men_n20_), .Y(men_men_n47_));
  NA2        u30(.A(men_men_n25_), .B(men_men_n23_), .Y(men_men_n48_));
  NO2        u31(.A(men_men_n48_), .B(men_men_n20_), .Y(men_men_n49_));
  AN2        u32(.A(men_men_n34_), .B(men_men_n19_), .Y(men_men_n50_));
  AOI210     u33(.A0(men_men_n49_), .A1(men_men_n33_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u34(.A0(men_men_n47_), .A1(men_men_n41_), .B0(men_men_n51_), .Y(men02));
  NAi21      u35(.An(men_men_n21_), .B(i_6_), .Y(men_men_n53_));
  NA3        u36(.A(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n54_));
  AOI210     u37(.A0(men_men_n49_), .A1(men_men_n54_), .B0(men_men_n28_), .Y(men_men_n55_));
  NA2        u38(.A(men_men_n55_), .B(men_men_n53_), .Y(men00));
  OAI210     u39(.A0(men_men_n48_), .A1(men_men_n34_), .B0(i_5_), .Y(men_men_n57_));
  NO2        u40(.A(men_men_n57_), .B(men_men_n20_), .Y(men09));
  NOi21      u41(.An(men_men_n33_), .B(men_men_n29_), .Y(men07));
  INV        u42(.A(i_3_), .Y(men08));
  INV        u43(.A(men_men_n26_), .Y(men_men_n61_));
  NA2        u44(.A(men07), .B(men_men_n61_), .Y(men_men_n62_));
  XO2        u45(.A(men_men_n62_), .B(men_men_n25_), .Y(men05));
  NO2        u46(.A(i_2_), .B(men08), .Y(men_men_n64_));
  XO2        u47(.A(men_men_n64_), .B(i_1_), .Y(men06));
  NAi21      u48(.An(men_men_n46_), .B(men_men_n39_), .Y(men_men_n66_));
  NA2        u49(.A(men_men_n66_), .B(i_0_), .Y(men_men_n67_));
  NO2        u50(.A(i_1_), .B(i_6_), .Y(men_men_n68_));
  NO3        u51(.A(men_men_n68_), .B(men_men_n37_), .C(men_men_n33_), .Y(men_men_n69_));
  NO2        u52(.A(men_men_n69_), .B(men_men_n35_), .Y(men_men_n70_));
  NO2        u53(.A(men_men_n23_), .B(men_men_n18_), .Y(men_men_n71_));
  OAI210     u54(.A0(men_men_n22_), .A1(i_6_), .B0(men_men_n18_), .Y(men_men_n72_));
  NO2        u55(.A(men_men_n72_), .B(men_men_n43_), .Y(men_men_n73_));
  AOI210     u56(.A0(men_men_n71_), .A1(i_0_), .B0(men_men_n73_), .Y(men_men_n74_));
  NA3        u57(.A(men_men_n74_), .B(men_men_n70_), .C(men_men_n67_), .Y(men03));
  NA2        u58(.A(men_men_n25_), .B(men08), .Y(men_men_n76_));
  INV        u59(.A(men_men_n54_), .Y(men_men_n77_));
  OAI210     u60(.A0(men_men_n77_), .A1(men_men_n30_), .B0(i_6_), .Y(men_men_n78_));
  NO2        u61(.A(men_men_n23_), .B(men_men_n26_), .Y(men_men_n79_));
  OR2        u62(.A(men_men_n79_), .B(men_men_n68_), .Y(men_men_n80_));
  NA3        u63(.A(men_men_n76_), .B(men_men_n68_), .C(i_2_), .Y(men_men_n81_));
  NA3        u64(.A(men_men_n81_), .B(men_men_n80_), .C(men_men_n78_), .Y(men04));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
endmodule