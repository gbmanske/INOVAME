module ex3_4(A, B, C, D, sum);
input  [3:0] A, B, C, D;
output [5:0] sum;

assign sum = A+B+C+D;

endmodule
