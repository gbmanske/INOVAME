//Benchmark atmr_5xp1_76_0.5

module atmr_5xp1(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n45_, ori_ori_n46_, ori_ori_n48_, ori_ori_n52_, ori_ori_n53_, ori_ori_n55_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n48_, mai_mai_n52_, mai_mai_n53_, mai_mai_n55_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n75_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n61_, men_men_n65_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09;
  INV        o00(.A(i_5_), .Y(ori_ori_n18_));
  NO3        o01(.A(i_4_), .B(i_6_), .C(ori_ori_n18_), .Y(ori_ori_n19_));
  INV        o02(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o03(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n21_));
  INV        o04(.A(i_1_), .Y(ori_ori_n22_));
  INV        o05(.A(i_0_), .Y(ori_ori_n23_));
  INV        o06(.A(i_6_), .Y(ori_ori_n24_));
  NO2        o07(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n25_));
  INV        o08(.A(i_0_), .Y(ori_ori_n26_));
  NO2        o09(.A(i_2_), .B(i_1_), .Y(ori_ori_n27_));
  NO2        o10(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n28_));
  NO2        o11(.A(i_2_), .B(i_3_), .Y(ori_ori_n29_));
  NO3        o12(.A(ori_ori_n29_), .B(ori_ori_n26_), .C(ori_ori_n22_), .Y(ori_ori_n30_));
  BUFFER     o13(.A(ori_ori_n25_), .Y(ori_ori_n31_));
  NA2        o14(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n32_));
  NA2        o15(.A(i_2_), .B(i_3_), .Y(ori_ori_n33_));
  NO2        o16(.A(ori_ori_n32_), .B(i_0_), .Y(ori_ori_n34_));
  OR3        o17(.A(ori_ori_n34_), .B(ori_ori_n31_), .C(ori_ori_n19_), .Y(ori01));
  NA2        o18(.A(i_0_), .B(i_1_), .Y(ori_ori_n36_));
  NO2        o19(.A(ori_ori_n36_), .B(i_6_), .Y(ori_ori_n37_));
  NO2        o20(.A(ori_ori_n32_), .B(ori_ori_n26_), .Y(ori_ori_n38_));
  NO3        o21(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(i_4_), .Y(ori_ori_n39_));
  NO2        o22(.A(i_6_), .B(ori_ori_n20_), .Y(ori_ori_n40_));
  NA2        o23(.A(ori_ori_n26_), .B(ori_ori_n24_), .Y(ori_ori_n41_));
  NO2        o24(.A(ori_ori_n41_), .B(ori_ori_n20_), .Y(ori_ori_n42_));
  INV        o25(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  OAI210     o26(.A0(ori_ori_n40_), .A1(ori_ori_n39_), .B0(ori_ori_n43_), .Y(ori02));
  NAi21      o27(.An(ori_ori_n21_), .B(i_6_), .Y(ori_ori_n45_));
  NO2        o28(.A(ori_ori_n42_), .B(ori_ori_n28_), .Y(ori_ori_n46_));
  NA2        o29(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori00));
  NA2        o30(.A(ori_ori_n41_), .B(i_5_), .Y(ori_ori_n48_));
  NO2        o31(.A(ori_ori_n48_), .B(ori_ori_n20_), .Y(ori09));
  NOi21      o32(.An(ori_ori_n33_), .B(ori_ori_n29_), .Y(ori07));
  INV        o33(.A(i_3_), .Y(ori08));
  INV        o34(.A(ori_ori_n27_), .Y(ori_ori_n52_));
  NA2        o35(.A(ori07), .B(ori_ori_n52_), .Y(ori_ori_n53_));
  XO2        o36(.A(ori_ori_n53_), .B(ori_ori_n26_), .Y(ori05));
  NO2        o37(.A(i_2_), .B(ori08), .Y(ori_ori_n55_));
  XO2        o38(.A(ori_ori_n55_), .B(i_1_), .Y(ori06));
  INV        o39(.A(ori_ori_n34_), .Y(ori_ori_n57_));
  OR2        o40(.A(ori_ori_n36_), .B(ori_ori_n18_), .Y(ori_ori_n58_));
  NA2        o41(.A(ori_ori_n58_), .B(ori_ori_n57_), .Y(ori03));
  NA2        o42(.A(ori_ori_n30_), .B(i_6_), .Y(ori_ori_n60_));
  NA3        o43(.A(ori_ori_n23_), .B(i_1_), .C(ori_ori_n24_), .Y(ori_ori_n61_));
  NA2        o44(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori04));
  INV        m00(.A(i_5_), .Y(mai_mai_n18_));
  NO3        m01(.A(i_4_), .B(i_6_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m02(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m03(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n21_));
  INV        m04(.A(i_1_), .Y(mai_mai_n22_));
  NO2        m05(.A(i_1_), .B(mai_mai_n21_), .Y(mai_mai_n23_));
  INV        m06(.A(i_6_), .Y(mai_mai_n24_));
  NO2        m07(.A(mai_mai_n24_), .B(i_5_), .Y(mai_mai_n25_));
  INV        m08(.A(i_0_), .Y(mai_mai_n26_));
  NO2        m09(.A(i_2_), .B(i_1_), .Y(mai_mai_n27_));
  OAI210     m10(.A0(mai_mai_n27_), .A1(mai_mai_n26_), .B0(mai_mai_n20_), .Y(mai_mai_n28_));
  NO2        m11(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n29_));
  NO2        m12(.A(i_2_), .B(i_3_), .Y(mai_mai_n30_));
  NO3        m13(.A(mai_mai_n30_), .B(mai_mai_n26_), .C(mai_mai_n22_), .Y(mai_mai_n31_));
  AO220      m14(.A0(mai_mai_n31_), .A1(mai_mai_n29_), .B0(mai_mai_n28_), .B1(mai_mai_n25_), .Y(mai_mai_n32_));
  NA2        m15(.A(i_2_), .B(i_3_), .Y(mai_mai_n33_));
  OR2        m16(.A(mai_mai_n32_), .B(mai_mai_n23_), .Y(mai01));
  NA2        m17(.A(mai_mai_n26_), .B(mai_mai_n18_), .Y(mai_mai_n35_));
  AOI210     m18(.A0(i_1_), .A1(mai_mai_n35_), .B0(mai_mai_n24_), .Y(mai_mai_n36_));
  NO3        m19(.A(mai_mai_n27_), .B(mai_mai_n36_), .C(i_4_), .Y(mai_mai_n37_));
  NA2        m20(.A(i_0_), .B(i_6_), .Y(mai_mai_n38_));
  OAI210     m21(.A0(i_0_), .A1(i_1_), .B0(mai_mai_n38_), .Y(mai_mai_n39_));
  NO2        m22(.A(mai_mai_n38_), .B(mai_mai_n27_), .Y(mai_mai_n40_));
  NO2        m23(.A(i_6_), .B(i_5_), .Y(mai_mai_n41_));
  NO3        m24(.A(mai_mai_n41_), .B(mai_mai_n40_), .C(mai_mai_n20_), .Y(mai_mai_n42_));
  OAI210     m25(.A0(mai_mai_n42_), .A1(mai_mai_n37_), .B0(mai_mai_n75_), .Y(mai02));
  NAi21      m26(.An(mai_mai_n21_), .B(i_1_), .Y(mai_mai_n44_));
  NA3        m27(.A(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n45_));
  INV        m28(.A(mai_mai_n29_), .Y(mai_mai_n46_));
  NA2        m29(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai00));
  INV        m30(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m31(.A(mai_mai_n48_), .B(mai_mai_n20_), .Y(mai09));
  NOi21      m32(.An(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai07));
  INV        m33(.A(i_3_), .Y(mai08));
  INV        m34(.A(mai_mai_n27_), .Y(mai_mai_n52_));
  NA2        m35(.A(mai07), .B(mai_mai_n52_), .Y(mai_mai_n53_));
  XO2        m36(.A(mai_mai_n53_), .B(mai_mai_n26_), .Y(mai05));
  NO2        m37(.A(i_2_), .B(mai08), .Y(mai_mai_n55_));
  XO2        m38(.A(mai_mai_n55_), .B(i_1_), .Y(mai06));
  NA2        m39(.A(mai_mai_n27_), .B(i_0_), .Y(mai_mai_n57_));
  NO2        m40(.A(i_1_), .B(i_6_), .Y(mai_mai_n58_));
  NO3        m41(.A(mai_mai_n58_), .B(mai_mai_n35_), .C(mai_mai_n33_), .Y(mai_mai_n59_));
  INV        m42(.A(mai_mai_n59_), .Y(mai_mai_n60_));
  OR2        m43(.A(i_1_), .B(mai_mai_n18_), .Y(mai_mai_n61_));
  NO2        m44(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n62_));
  NO2        m45(.A(i_5_), .B(mai_mai_n39_), .Y(mai_mai_n63_));
  AOI210     m46(.A0(mai_mai_n62_), .A1(i_0_), .B0(mai_mai_n63_), .Y(mai_mai_n64_));
  NA4        m47(.A(mai_mai_n64_), .B(mai_mai_n61_), .C(mai_mai_n60_), .D(mai_mai_n57_), .Y(mai03));
  NA2        m48(.A(mai_mai_n26_), .B(mai08), .Y(mai_mai_n66_));
  OAI210     m49(.A0(mai_mai_n66_), .A1(i_1_), .B0(mai_mai_n45_), .Y(mai_mai_n67_));
  OAI210     m50(.A0(mai_mai_n67_), .A1(mai_mai_n31_), .B0(i_6_), .Y(mai_mai_n68_));
  AOI210     m51(.A0(mai_mai_n30_), .A1(mai_mai_n24_), .B0(mai_mai_n27_), .Y(mai_mai_n69_));
  BUFFER     m52(.A(mai_mai_n69_), .Y(mai_mai_n70_));
  NA2        m53(.A(mai_mai_n66_), .B(mai_mai_n58_), .Y(mai_mai_n71_));
  NA3        m54(.A(mai_mai_n71_), .B(mai_mai_n70_), .C(mai_mai_n68_), .Y(mai04));
  INV        m55(.A(mai_mai_n19_), .Y(mai_mai_n75_));
  INV        u00(.A(i_5_), .Y(men_men_n18_));
  NO3        u01(.A(i_4_), .B(i_6_), .C(men_men_n18_), .Y(men_men_n19_));
  INV        u02(.A(i_4_), .Y(men_men_n20_));
  NA2        u03(.A(men_men_n20_), .B(i_5_), .Y(men_men_n21_));
  INV        u04(.A(i_1_), .Y(men_men_n22_));
  AOI210     u05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(men_men_n23_));
  NA2        u06(.A(men_men_n23_), .B(men_men_n22_), .Y(men_men_n24_));
  NO2        u07(.A(men_men_n24_), .B(men_men_n21_), .Y(men_men_n25_));
  INV        u08(.A(i_6_), .Y(men_men_n26_));
  INV        u09(.A(i_0_), .Y(men_men_n27_));
  NO2        u10(.A(i_2_), .B(i_1_), .Y(men_men_n28_));
  NO2        u11(.A(men_men_n20_), .B(i_5_), .Y(men_men_n29_));
  NO2        u12(.A(i_2_), .B(i_3_), .Y(men_men_n30_));
  NA2        u13(.A(men_men_n26_), .B(i_5_), .Y(men_men_n31_));
  NA2        u14(.A(i_2_), .B(i_3_), .Y(men_men_n32_));
  NO2        u15(.A(men_men_n32_), .B(men_men_n22_), .Y(men_men_n33_));
  NO3        u16(.A(men_men_n33_), .B(men_men_n31_), .C(i_0_), .Y(men_men_n34_));
  OR4        u17(.A(men_men_n34_), .B(men_men_n29_), .C(men_men_n25_), .D(men_men_n19_), .Y(men01));
  OR2        u18(.A(i_2_), .B(i_3_), .Y(men_men_n36_));
  NA3        u19(.A(men_men_n36_), .B(i_0_), .C(i_1_), .Y(men_men_n37_));
  NA2        u20(.A(men_men_n27_), .B(men_men_n18_), .Y(men_men_n38_));
  AOI210     u21(.A0(men_men_n23_), .A1(men_men_n22_), .B0(men_men_n26_), .Y(men_men_n39_));
  AOI220     u22(.A0(men_men_n39_), .A1(men_men_n38_), .B0(men_men_n37_), .B1(men_men_n26_), .Y(men_men_n40_));
  NA2        u23(.A(men_men_n28_), .B(men_men_n18_), .Y(men_men_n41_));
  NO2        u24(.A(men_men_n41_), .B(men_men_n26_), .Y(men_men_n42_));
  NO3        u25(.A(men_men_n42_), .B(men_men_n40_), .C(i_4_), .Y(men_men_n43_));
  NA2        u26(.A(i_0_), .B(i_6_), .Y(men_men_n44_));
  OAI210     u27(.A0(i_0_), .A1(i_1_), .B0(men_men_n44_), .Y(men_men_n45_));
  NOi31      u28(.An(men_men_n45_), .B(men_men_n23_), .C(men_men_n18_), .Y(men_men_n46_));
  NA3        u29(.A(i_1_), .B(i_6_), .C(i_5_), .Y(men_men_n47_));
  NO2        u30(.A(men_men_n47_), .B(men_men_n28_), .Y(men_men_n48_));
  NO3        u31(.A(men_men_n36_), .B(i_6_), .C(i_5_), .Y(men_men_n49_));
  NO4        u32(.A(men_men_n49_), .B(men_men_n48_), .C(men_men_n46_), .D(men_men_n20_), .Y(men_men_n50_));
  NA2        u33(.A(men_men_n27_), .B(men_men_n26_), .Y(men_men_n51_));
  NO2        u34(.A(men_men_n51_), .B(men_men_n20_), .Y(men_men_n52_));
  AOI210     u35(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(men_men_n53_));
  AO220      u36(.A0(men_men_n53_), .A1(men_men_n29_), .B0(men_men_n33_), .B1(men_men_n19_), .Y(men_men_n54_));
  AOI210     u37(.A0(men_men_n52_), .A1(men_men_n32_), .B0(men_men_n54_), .Y(men_men_n55_));
  OAI210     u38(.A0(men_men_n50_), .A1(men_men_n43_), .B0(men_men_n55_), .Y(men02));
  NAi21      u39(.An(men_men_n21_), .B(men_men_n39_), .Y(men_men_n57_));
  NA3        u40(.A(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n58_));
  AOI210     u41(.A0(men_men_n52_), .A1(men_men_n58_), .B0(men_men_n29_), .Y(men_men_n59_));
  NA2        u42(.A(men_men_n59_), .B(men_men_n57_), .Y(men00));
  OAI210     u43(.A0(men_men_n51_), .A1(men_men_n33_), .B0(i_5_), .Y(men_men_n61_));
  NO2        u44(.A(men_men_n61_), .B(men_men_n20_), .Y(men09));
  NOi21      u45(.An(men_men_n32_), .B(men_men_n30_), .Y(men07));
  INV        u46(.A(i_3_), .Y(men08));
  INV        u47(.A(men07), .Y(men_men_n65_));
  XO2        u48(.A(men_men_n65_), .B(men_men_n27_), .Y(men05));
  NAi21      u49(.An(men_men_n49_), .B(men_men_n41_), .Y(men_men_n67_));
  NA2        u50(.A(men_men_n67_), .B(i_0_), .Y(men_men_n68_));
  NO2        u51(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO3        u52(.A(men_men_n69_), .B(men_men_n38_), .C(men_men_n32_), .Y(men_men_n70_));
  NO2        u53(.A(men_men_n70_), .B(men_men_n34_), .Y(men_men_n71_));
  AO210      u54(.A0(men_men_n37_), .A1(men_men_n24_), .B0(men_men_n18_), .Y(men_men_n72_));
  NO2        u55(.A(men_men_n28_), .B(men_men_n27_), .Y(men_men_n73_));
  OAI210     u56(.A0(men_men_n22_), .A1(i_6_), .B0(men_men_n18_), .Y(men_men_n74_));
  NO2        u57(.A(men_men_n74_), .B(men_men_n45_), .Y(men_men_n75_));
  AOI210     u58(.A0(i_6_), .A1(men_men_n73_), .B0(men_men_n75_), .Y(men_men_n76_));
  NA4        u59(.A(men_men_n76_), .B(men_men_n72_), .C(men_men_n71_), .D(men_men_n68_), .Y(men03));
  NA2        u60(.A(men_men_n27_), .B(men08), .Y(men_men_n78_));
  OAI210     u61(.A0(men_men_n78_), .A1(i_1_), .B0(men_men_n58_), .Y(men_men_n79_));
  NA2        u62(.A(men_men_n79_), .B(i_6_), .Y(men_men_n80_));
  OR2        u63(.A(i_2_), .B(men_men_n69_), .Y(men_men_n81_));
  NA3        u64(.A(men_men_n78_), .B(men_men_n69_), .C(i_2_), .Y(men_men_n82_));
  NA3        u65(.A(men_men_n23_), .B(i_1_), .C(men_men_n26_), .Y(men_men_n83_));
  NA4        u66(.A(men_men_n83_), .B(men_men_n82_), .C(men_men_n81_), .D(men_men_n80_), .Y(men04));
  BUFFER     u67(.A(i_1_), .Y(men06));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
endmodule