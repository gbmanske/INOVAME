//Benchmark atmr_max1024_476_0.25

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n257_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  INV        o004(.A(ori_ori_n19_), .Y(ori_ori_n21_));
  NA2        o005(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n22_));
  INV        o006(.A(x5), .Y(ori_ori_n23_));
  NA2        o007(.A(x4), .B(x2), .Y(ori_ori_n24_));
  INV        o008(.A(ori_ori_n22_), .Y(ori_ori_n25_));
  NO2        o009(.A(x4), .B(x3), .Y(ori_ori_n26_));
  INV        o010(.A(ori_ori_n26_), .Y(ori_ori_n27_));
  NOi21      o011(.An(ori_ori_n21_), .B(ori_ori_n25_), .Y(ori00));
  NO2        o012(.A(x1), .B(x0), .Y(ori_ori_n29_));
  INV        o013(.A(x6), .Y(ori_ori_n30_));
  NA2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  NO2        o015(.A(ori_ori_n21_), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NO2        o016(.A(x2), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x3), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n34_), .B(ori_ori_n18_), .Y(ori_ori_n35_));
  INV        o019(.A(ori_ori_n35_), .Y(ori_ori_n36_));
  INV        o020(.A(x4), .Y(ori_ori_n37_));
  OAI210     o021(.A0(ori_ori_n37_), .A1(ori_ori_n36_), .B0(ori_ori_n33_), .Y(ori_ori_n38_));
  INV        o022(.A(x4), .Y(ori_ori_n39_));
  NO2        o023(.A(ori_ori_n39_), .B(ori_ori_n17_), .Y(ori_ori_n40_));
  NA2        o024(.A(ori_ori_n40_), .B(x2), .Y(ori_ori_n41_));
  OAI210     o025(.A0(ori_ori_n41_), .A1(ori_ori_n20_), .B0(ori_ori_n38_), .Y(ori_ori_n42_));
  INV        o026(.A(ori_ori_n29_), .Y(ori_ori_n43_));
  INV        o027(.A(x2), .Y(ori_ori_n44_));
  NO2        o028(.A(ori_ori_n44_), .B(ori_ori_n17_), .Y(ori_ori_n45_));
  NA2        o029(.A(ori_ori_n34_), .B(ori_ori_n18_), .Y(ori_ori_n46_));
  NA2        o030(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  OAI210     o031(.A0(ori_ori_n43_), .A1(ori_ori_n27_), .B0(ori_ori_n47_), .Y(ori_ori_n48_));
  NO3        o032(.A(ori_ori_n48_), .B(ori_ori_n42_), .C(ori_ori_n32_), .Y(ori01));
  INV        o033(.A(x7), .Y(ori_ori_n50_));
  NA2        o034(.A(ori_ori_n34_), .B(x1), .Y(ori_ori_n51_));
  INV        o035(.A(x6), .Y(ori_ori_n52_));
  NO2        o036(.A(ori_ori_n51_), .B(x5), .Y(ori_ori_n53_));
  OAI210     o037(.A0(ori_ori_n35_), .A1(ori_ori_n23_), .B0(ori_ori_n44_), .Y(ori_ori_n54_));
  OAI210     o038(.A0(ori_ori_n46_), .A1(ori_ori_n20_), .B0(ori_ori_n54_), .Y(ori_ori_n55_));
  INV        o039(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(x4), .Y(ori_ori_n57_));
  NA2        o041(.A(ori_ori_n39_), .B(x2), .Y(ori_ori_n58_));
  OAI210     o042(.A0(ori_ori_n58_), .A1(ori_ori_n46_), .B0(x0), .Y(ori_ori_n59_));
  NA2        o043(.A(x5), .B(x3), .Y(ori_ori_n60_));
  INV        o044(.A(x6), .Y(ori_ori_n61_));
  NO3        o045(.A(ori_ori_n60_), .B(ori_ori_n52_), .C(ori_ori_n44_), .Y(ori_ori_n62_));
  NAi21      o046(.An(x4), .B(x3), .Y(ori_ori_n63_));
  INV        o047(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NO2        o048(.A(x4), .B(x2), .Y(ori_ori_n65_));
  NO2        o049(.A(ori_ori_n63_), .B(ori_ori_n18_), .Y(ori_ori_n66_));
  NO3        o050(.A(ori_ori_n66_), .B(ori_ori_n62_), .C(ori_ori_n59_), .Y(ori_ori_n67_));
  NA2        o051(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n68_));
  NO2        o052(.A(ori_ori_n68_), .B(ori_ori_n23_), .Y(ori_ori_n69_));
  INV        o053(.A(x8), .Y(ori_ori_n70_));
  NA2        o054(.A(x2), .B(x1), .Y(ori_ori_n71_));
  AOI210     o055(.A0(ori_ori_n46_), .A1(ori_ori_n23_), .B0(ori_ori_n44_), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n36_), .B(ori_ori_n39_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NA2        o058(.A(x4), .B(ori_ori_n34_), .Y(ori_ori_n75_));
  NO2        o059(.A(ori_ori_n39_), .B(ori_ori_n44_), .Y(ori_ori_n76_));
  NO2        o060(.A(ori_ori_n75_), .B(x1), .Y(ori_ori_n77_));
  NA2        o061(.A(ori_ori_n44_), .B(x1), .Y(ori_ori_n78_));
  OAI210     o062(.A0(ori_ori_n78_), .A1(ori_ori_n31_), .B0(ori_ori_n17_), .Y(ori_ori_n79_));
  NO3        o063(.A(ori_ori_n79_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n80_));
  AO210      o064(.A0(ori_ori_n67_), .A1(ori_ori_n57_), .B0(ori_ori_n80_), .Y(ori02));
  BUFFER     o065(.A(x0), .Y(ori_ori_n82_));
  INV        o066(.A(ori_ori_n82_), .Y(ori_ori_n83_));
  NO2        o067(.A(x4), .B(x1), .Y(ori_ori_n84_));
  NA2        o068(.A(ori_ori_n84_), .B(x2), .Y(ori_ori_n85_));
  NOi21      o069(.An(x0), .B(x1), .Y(ori_ori_n86_));
  NOi21      o070(.An(x0), .B(x4), .Y(ori_ori_n87_));
  NO2        o071(.A(ori_ori_n85_), .B(ori_ori_n60_), .Y(ori_ori_n88_));
  NO2        o072(.A(x5), .B(ori_ori_n39_), .Y(ori_ori_n89_));
  NA2        o073(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n90_), .A1(ori_ori_n78_), .B0(x3), .Y(ori_ori_n91_));
  OAI210     o075(.A0(ori_ori_n91_), .A1(ori_ori_n29_), .B0(ori_ori_n89_), .Y(ori_ori_n92_));
  NAi21      o076(.An(x0), .B(x4), .Y(ori_ori_n93_));
  NO2        o077(.A(x7), .B(x0), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n65_), .B(ori_ori_n76_), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n95_), .B(x3), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n94_), .B(ori_ori_n96_), .Y(ori_ori_n97_));
  NA2        o081(.A(x5), .B(x0), .Y(ori_ori_n98_));
  NO2        o082(.A(ori_ori_n39_), .B(x2), .Y(ori_ori_n99_));
  NA3        o083(.A(ori_ori_n97_), .B(ori_ori_n92_), .C(ori_ori_n30_), .Y(ori_ori_n100_));
  NO2        o084(.A(ori_ori_n100_), .B(ori_ori_n88_), .Y(ori_ori_n101_));
  NO3        o085(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n22_), .Y(ori_ori_n102_));
  NO2        o086(.A(ori_ori_n24_), .B(ori_ori_n23_), .Y(ori_ori_n103_));
  NO2        o087(.A(ori_ori_n75_), .B(x5), .Y(ori_ori_n104_));
  NO2        o088(.A(ori_ori_n34_), .B(x2), .Y(ori_ori_n105_));
  INV        o089(.A(x7), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n106_), .B(ori_ori_n18_), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n107_), .B(ori_ori_n105_), .Y(ori_ori_n108_));
  NO2        o092(.A(ori_ori_n23_), .B(x4), .Y(ori_ori_n109_));
  INV        o093(.A(ori_ori_n87_), .Y(ori_ori_n110_));
  NO2        o094(.A(ori_ori_n110_), .B(ori_ori_n108_), .Y(ori_ori_n111_));
  NA2        o095(.A(x5), .B(x1), .Y(ori_ori_n112_));
  INV        o096(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  AOI210     o097(.A0(ori_ori_n113_), .A1(ori_ori_n87_), .B0(ori_ori_n30_), .Y(ori_ori_n114_));
  BUFFER     o098(.A(x2), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n115_), .B(ori_ori_n39_), .Y(ori_ori_n116_));
  NA2        o100(.A(ori_ori_n116_), .B(ori_ori_n53_), .Y(ori_ori_n117_));
  NA2        o101(.A(ori_ori_n117_), .B(ori_ori_n114_), .Y(ori_ori_n118_));
  NO3        o102(.A(ori_ori_n118_), .B(ori_ori_n111_), .C(ori_ori_n102_), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n119_), .B(ori_ori_n101_), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n98_), .B(ori_ori_n95_), .Y(ori_ori_n121_));
  NA2        o105(.A(ori_ori_n23_), .B(ori_ori_n18_), .Y(ori_ori_n122_));
  NA2        o106(.A(ori_ori_n23_), .B(ori_ori_n17_), .Y(ori_ori_n123_));
  NA3        o107(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(ori_ori_n22_), .Y(ori_ori_n124_));
  AN2        o108(.A(ori_ori_n124_), .B(ori_ori_n99_), .Y(ori_ori_n125_));
  NO2        o109(.A(ori_ori_n106_), .B(ori_ori_n23_), .Y(ori_ori_n126_));
  NA2        o110(.A(x2), .B(x0), .Y(ori_ori_n127_));
  NA2        o111(.A(x4), .B(x1), .Y(ori_ori_n128_));
  NAi21      o112(.An(ori_ori_n84_), .B(ori_ori_n128_), .Y(ori_ori_n129_));
  NOi31      o113(.An(ori_ori_n129_), .B(ori_ori_n109_), .C(ori_ori_n127_), .Y(ori_ori_n130_));
  NO3        o114(.A(ori_ori_n130_), .B(ori_ori_n125_), .C(ori_ori_n121_), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n131_), .B(ori_ori_n34_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n124_), .B(ori_ori_n58_), .Y(ori_ori_n133_));
  INV        o117(.A(ori_ori_n89_), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n78_), .B(ori_ori_n17_), .Y(ori_ori_n135_));
  NA2        o119(.A(ori_ori_n129_), .B(ori_ori_n33_), .Y(ori_ori_n136_));
  OAI210     o120(.A0(ori_ori_n123_), .A1(ori_ori_n95_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n137_), .B(ori_ori_n133_), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n138_), .B(x3), .Y(ori_ori_n139_));
  NO3        o123(.A(ori_ori_n139_), .B(ori_ori_n132_), .C(ori_ori_n120_), .Y(ori03));
  NO2        o124(.A(ori_ori_n39_), .B(x3), .Y(ori_ori_n141_));
  NA2        o125(.A(x6), .B(ori_ori_n23_), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n142_), .B(x4), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n144_));
  NA2        o128(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n145_));
  NO3        o129(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n146_));
  NO2        o130(.A(x5), .B(x1), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n145_), .B(ori_ori_n122_), .Y(ori_ori_n148_));
  NO3        o132(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n149_));
  NA2        o133(.A(x3), .B(ori_ori_n19_), .Y(ori_ori_n150_));
  NO2        o134(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n151_), .B(x6), .Y(ori_ori_n152_));
  NOi21      o136(.An(ori_ori_n65_), .B(ori_ori_n152_), .Y(ori_ori_n153_));
  NA2        o137(.A(ori_ori_n151_), .B(x6), .Y(ori_ori_n154_));
  AOI210     o138(.A0(ori_ori_n154_), .A1(ori_ori_n153_), .B0(ori_ori_n106_), .Y(ori_ori_n155_));
  OR2        o139(.A(ori_ori_n155_), .B(ori_ori_n126_), .Y(ori_ori_n156_));
  NA2        o140(.A(ori_ori_n34_), .B(ori_ori_n44_), .Y(ori_ori_n157_));
  NA2        o141(.A(ori_ori_n99_), .B(ori_ori_n69_), .Y(ori_ori_n158_));
  NA2        o142(.A(x6), .B(ori_ori_n39_), .Y(ori_ori_n159_));
  OAI210     o143(.A0(ori_ori_n83_), .A1(ori_ori_n61_), .B0(x4), .Y(ori_ori_n160_));
  AOI210     o144(.A0(ori_ori_n160_), .A1(ori_ori_n159_), .B0(ori_ori_n60_), .Y(ori_ori_n161_));
  OAI210     o145(.A0(ori_ori_n53_), .A1(ori_ori_n161_), .B0(x2), .Y(ori_ori_n162_));
  NA3        o146(.A(ori_ori_n162_), .B(ori_ori_n158_), .C(ori_ori_n156_), .Y(ori_ori_n163_));
  INV        o147(.A(ori_ori_n163_), .Y(ori_ori_n164_));
  INV        o148(.A(x3), .Y(ori_ori_n165_));
  NA2        o149(.A(ori_ori_n165_), .B(ori_ori_n143_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n68_), .B(ori_ori_n23_), .Y(ori_ori_n167_));
  AOI210     o151(.A0(ori_ori_n152_), .A1(ori_ori_n109_), .B0(ori_ori_n167_), .Y(ori_ori_n168_));
  AOI210     o152(.A0(ori_ori_n168_), .A1(ori_ori_n166_), .B0(x2), .Y(ori_ori_n169_));
  AOI220     o153(.A0(ori_ori_n143_), .A1(ori_ori_n135_), .B0(x2), .B1(ori_ori_n53_), .Y(ori_ori_n170_));
  NA2        o154(.A(ori_ori_n34_), .B(ori_ori_n17_), .Y(ori_ori_n171_));
  NA2        o155(.A(ori_ori_n145_), .B(x6), .Y(ori_ori_n172_));
  NO2        o156(.A(ori_ori_n145_), .B(x6), .Y(ori_ori_n173_));
  INV        o157(.A(ori_ori_n173_), .Y(ori_ori_n174_));
  NA3        o158(.A(ori_ori_n174_), .B(ori_ori_n172_), .C(ori_ori_n103_), .Y(ori_ori_n175_));
  NA3        o159(.A(ori_ori_n175_), .B(ori_ori_n170_), .C(ori_ori_n106_), .Y(ori_ori_n176_));
  BUFFER     o160(.A(x1), .Y(ori_ori_n177_));
  NA2        o161(.A(x6), .B(x2), .Y(ori_ori_n178_));
  NA2        o162(.A(x4), .B(x0), .Y(ori_ori_n179_));
  NO2        o163(.A(ori_ori_n176_), .B(ori_ori_n169_), .Y(ori_ori_n180_));
  NA2        o164(.A(ori_ori_n173_), .B(x2), .Y(ori_ori_n181_));
  OAI210     o165(.A0(x0), .A1(x6), .B0(ori_ori_n35_), .Y(ori_ori_n182_));
  AOI210     o166(.A0(ori_ori_n182_), .A1(ori_ori_n181_), .B0(ori_ori_n134_), .Y(ori_ori_n183_));
  NOi21      o167(.An(ori_ori_n178_), .B(ori_ori_n17_), .Y(ori_ori_n184_));
  NA3        o168(.A(ori_ori_n184_), .B(ori_ori_n147_), .C(ori_ori_n31_), .Y(ori_ori_n185_));
  AOI210     o169(.A0(ori_ori_n30_), .A1(ori_ori_n44_), .B0(x0), .Y(ori_ori_n186_));
  NA3        o170(.A(ori_ori_n186_), .B(ori_ori_n113_), .C(ori_ori_n27_), .Y(ori_ori_n187_));
  NA2        o171(.A(x3), .B(x2), .Y(ori_ori_n188_));
  AOI220     o172(.A0(ori_ori_n188_), .A1(ori_ori_n157_), .B0(ori_ori_n187_), .B1(ori_ori_n185_), .Y(ori_ori_n189_));
  NAi21      o173(.An(x4), .B(x0), .Y(ori_ori_n190_));
  NO3        o174(.A(ori_ori_n190_), .B(ori_ori_n35_), .C(x2), .Y(ori_ori_n191_));
  OAI210     o175(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n191_), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n186_), .B(ori_ori_n184_), .Y(ori_ori_n193_));
  AOI220     o177(.A0(ori_ori_n193_), .A1(ori_ori_n64_), .B0(ori_ori_n18_), .B1(ori_ori_n26_), .Y(ori_ori_n194_));
  AOI210     o178(.A0(ori_ori_n194_), .A1(ori_ori_n192_), .B0(ori_ori_n23_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n186_), .B(ori_ori_n184_), .Y(ori_ori_n196_));
  INV        o180(.A(ori_ori_n148_), .Y(ori_ori_n197_));
  NA2        o181(.A(ori_ori_n30_), .B(ori_ori_n34_), .Y(ori_ori_n198_));
  OR2        o182(.A(ori_ori_n198_), .B(ori_ori_n179_), .Y(ori_ori_n199_));
  OAI220     o183(.A0(ori_ori_n199_), .A1(ori_ori_n112_), .B0(ori_ori_n159_), .B1(ori_ori_n197_), .Y(ori_ori_n200_));
  AO210      o184(.A0(ori_ori_n196_), .A1(ori_ori_n104_), .B0(ori_ori_n200_), .Y(ori_ori_n201_));
  NO4        o185(.A(ori_ori_n201_), .B(ori_ori_n195_), .C(ori_ori_n189_), .D(ori_ori_n183_), .Y(ori_ori_n202_));
  OAI210     o186(.A0(ori_ori_n180_), .A1(ori_ori_n164_), .B0(ori_ori_n202_), .Y(ori04));
  INV        o187(.A(x2), .Y(ori_ori_n204_));
  OAI210     o188(.A0(ori_ori_n171_), .A1(ori_ori_n204_), .B0(ori_ori_n30_), .Y(ori_ori_n205_));
  INV        o189(.A(ori_ori_n190_), .Y(ori_ori_n206_));
  OAI210     o190(.A0(ori_ori_n44_), .A1(ori_ori_n206_), .B0(ori_ori_n165_), .Y(ori_ori_n207_));
  NO2        o191(.A(ori_ori_n188_), .B(ori_ori_n144_), .Y(ori_ori_n208_));
  INV        o192(.A(ori_ori_n208_), .Y(ori_ori_n209_));
  NA3        o193(.A(ori_ori_n209_), .B(x6), .C(ori_ori_n207_), .Y(ori_ori_n210_));
  NA2        o194(.A(ori_ori_n210_), .B(ori_ori_n205_), .Y(ori_ori_n211_));
  NA2        o195(.A(x3), .B(ori_ori_n191_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n146_), .B(ori_ori_n65_), .Y(ori_ori_n213_));
  NA3        o197(.A(ori_ori_n213_), .B(ori_ori_n212_), .C(ori_ori_n106_), .Y(ori_ori_n214_));
  INV        o198(.A(ori_ori_n214_), .Y(ori_ori_n215_));
  XO2        o199(.A(x4), .B(x0), .Y(ori_ori_n216_));
  NA2        o200(.A(x4), .B(ori_ori_n71_), .Y(ori_ori_n217_));
  NO2        o201(.A(ori_ori_n217_), .B(x3), .Y(ori_ori_n218_));
  INV        o202(.A(ori_ori_n71_), .Y(ori_ori_n219_));
  NA2        o203(.A(ori_ori_n87_), .B(ori_ori_n219_), .Y(ori_ori_n220_));
  NO2        o204(.A(ori_ori_n216_), .B(x2), .Y(ori_ori_n221_));
  INV        o205(.A(ori_ori_n221_), .Y(ori_ori_n222_));
  NA4        o206(.A(ori_ori_n222_), .B(ori_ori_n220_), .C(ori_ori_n150_), .D(x6), .Y(ori_ori_n223_));
  NO2        o207(.A(ori_ori_n127_), .B(ori_ori_n70_), .Y(ori_ori_n224_));
  NA2        o208(.A(ori_ori_n224_), .B(ori_ori_n51_), .Y(ori_ori_n225_));
  NO2        o209(.A(x8), .B(ori_ori_n63_), .Y(ori_ori_n226_));
  NO2        o210(.A(ori_ori_n29_), .B(x2), .Y(ori_ori_n227_));
  NA2        o211(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  NA2        o212(.A(ori_ori_n225_), .B(ori_ori_n228_), .Y(ori_ori_n229_));
  OAI220     o213(.A0(ori_ori_n229_), .A1(x6), .B0(ori_ori_n223_), .B1(ori_ori_n218_), .Y(ori_ori_n230_));
  AO220      o214(.A0(x7), .A1(ori_ori_n230_), .B0(ori_ori_n215_), .B1(ori_ori_n211_), .Y(ori_ori_n231_));
  NA2        o215(.A(ori_ori_n149_), .B(ori_ori_n40_), .Y(ori_ori_n232_));
  NA2        o216(.A(ori_ori_n232_), .B(ori_ori_n231_), .Y(ori_ori_n233_));
  NA3        o217(.A(ori_ori_n17_), .B(ori_ori_n141_), .C(ori_ori_n106_), .Y(ori_ori_n234_));
  NA3        o218(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n235_));
  NA2        o219(.A(x3), .B(x0), .Y(ori_ori_n236_));
  OAI220     o220(.A0(ori_ori_n236_), .A1(x2), .B0(ori_ori_n235_), .B1(ori_ori_n219_), .Y(ori_ori_n237_));
  INV        o221(.A(ori_ori_n237_), .Y(ori_ori_n238_));
  AOI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n234_), .B0(ori_ori_n23_), .Y(ori_ori_n239_));
  NA2        o223(.A(ori_ori_n239_), .B(x6), .Y(ori_ori_n240_));
  INV        o224(.A(ori_ori_n93_), .Y(ori_ori_n241_));
  NO2        o225(.A(ori_ori_n241_), .B(ori_ori_n34_), .Y(ori_ori_n242_));
  AOI210     o226(.A0(ori_ori_n177_), .A1(ori_ori_n50_), .B0(ori_ori_n86_), .Y(ori_ori_n243_));
  NO2        o227(.A(ori_ori_n243_), .B(x3), .Y(ori_ori_n244_));
  NO3        o228(.A(ori_ori_n244_), .B(ori_ori_n242_), .C(x2), .Y(ori_ori_n245_));
  OAI210     o229(.A0(ori_ori_n190_), .A1(ori_ori_n34_), .B0(ori_ori_n216_), .Y(ori_ori_n246_));
  AOI220     o230(.A0(x7), .A1(ori_ori_n70_), .B0(ori_ori_n246_), .B1(ori_ori_n106_), .Y(ori_ori_n247_));
  NO2        o231(.A(ori_ori_n247_), .B(ori_ori_n44_), .Y(ori_ori_n248_));
  NO2        o232(.A(ori_ori_n248_), .B(ori_ori_n245_), .Y(ori_ori_n249_));
  AOI210     o233(.A0(ori_ori_n249_), .A1(ori_ori_n41_), .B0(ori_ori_n23_), .Y(ori_ori_n250_));
  NA2        o234(.A(ori_ori_n250_), .B(ori_ori_n30_), .Y(ori_ori_n251_));
  NO4        o235(.A(x0), .B(ori_ori_n60_), .C(x4), .D(ori_ori_n44_), .Y(ori_ori_n252_));
  NA3        o236(.A(ori_ori_n257_), .B(ori_ori_n251_), .C(ori_ori_n240_), .Y(ori_ori_n253_));
  AOI210     o237(.A0(ori_ori_n233_), .A1(ori_ori_n23_), .B0(ori_ori_n253_), .Y(ori05));
  INV        o238(.A(ori_ori_n252_), .Y(ori_ori_n257_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  INV        m047(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  NO2        m048(.A(mai_mai_n64_), .B(mai_mai_n61_), .Y(mai_mai_n65_));
  NO2        m049(.A(x7), .B(x6), .Y(mai_mai_n66_));
  NO2        m050(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n67_));
  NO2        m051(.A(x8), .B(x2), .Y(mai_mai_n68_));
  OA210      m052(.A0(mai_mai_n68_), .A1(mai_mai_n67_), .B0(mai_mai_n66_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n70_), .Y(mai_mai_n71_));
  NAi31      m055(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n72_));
  NO2        m056(.A(mai_mai_n71_), .B(mai_mai_n69_), .Y(mai_mai_n73_));
  OAI210     m057(.A0(mai_mai_n73_), .A1(mai_mai_n65_), .B0(x4), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n75_));
  OAI210     m059(.A0(mai_mai_n75_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n76_));
  NA2        m060(.A(x5), .B(x3), .Y(mai_mai_n77_));
  NO2        m061(.A(x8), .B(x6), .Y(mai_mai_n78_));
  NO2        m062(.A(mai_mai_n77_), .B(mai_mai_n54_), .Y(mai_mai_n79_));
  NAi21      m063(.An(x4), .B(x3), .Y(mai_mai_n80_));
  INV        m064(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m065(.A(mai_mai_n81_), .B(mai_mai_n22_), .Y(mai_mai_n82_));
  NO2        m066(.A(x4), .B(x2), .Y(mai_mai_n83_));
  NO2        m067(.A(mai_mai_n83_), .B(x3), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n82_), .C(mai_mai_n18_), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n79_), .C(mai_mai_n76_), .Y(mai_mai_n86_));
  NO3        m070(.A(mai_mai_n21_), .B(mai_mai_n43_), .C(x1), .Y(mai_mai_n87_));
  NA2        m071(.A(mai_mai_n87_), .B(mai_mai_n48_), .Y(mai_mai_n88_));
  NA2        m072(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n89_), .B(mai_mai_n25_), .Y(mai_mai_n90_));
  INV        m074(.A(x8), .Y(mai_mai_n91_));
  NA2        m075(.A(x2), .B(x1), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n90_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n26_), .Y(mai_mai_n95_));
  AOI210     m079(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n96_));
  OAI210     m080(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n97_));
  NO3        m081(.A(mai_mai_n97_), .B(mai_mai_n96_), .C(mai_mai_n95_), .Y(mai_mai_n98_));
  NA2        m082(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n99_));
  NO2        m083(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n100_));
  OAI210     m084(.A0(mai_mai_n100_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n101_));
  AOI210     m085(.A0(mai_mai_n99_), .A1(mai_mai_n52_), .B0(mai_mai_n101_), .Y(mai_mai_n102_));
  NO2        m086(.A(x3), .B(x2), .Y(mai_mai_n103_));
  NA2        m087(.A(mai_mai_n103_), .B(mai_mai_n25_), .Y(mai_mai_n104_));
  INV        m088(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NA2        m089(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n106_));
  OAI210     m090(.A0(mai_mai_n106_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n107_));
  NO4        m091(.A(mai_mai_n107_), .B(mai_mai_n105_), .C(mai_mai_n102_), .D(mai_mai_n98_), .Y(mai_mai_n108_));
  AO220      m092(.A0(mai_mai_n108_), .A1(mai_mai_n88_), .B0(mai_mai_n86_), .B1(mai_mai_n74_), .Y(mai02));
  NO2        m093(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n110_));
  NO2        m094(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n111_));
  NO2        m095(.A(x4), .B(x2), .Y(mai_mai_n112_));
  AOI220     m096(.A0(mai_mai_n112_), .A1(mai_mai_n111_), .B0(mai_mai_n110_), .B1(x4), .Y(mai_mai_n113_));
  NO3        m097(.A(mai_mai_n113_), .B(x7), .C(x5), .Y(mai_mai_n114_));
  OR2        m098(.A(x8), .B(x0), .Y(mai_mai_n115_));
  INV        m099(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NAi21      m100(.An(x2), .B(x8), .Y(mai_mai_n117_));
  NO2        m101(.A(x4), .B(x1), .Y(mai_mai_n118_));
  NOi21      m102(.An(x0), .B(x1), .Y(mai_mai_n119_));
  NO3        m103(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n120_));
  NOi21      m104(.An(x0), .B(x4), .Y(mai_mai_n121_));
  AOI220     m105(.A0(mai_mai_n398_), .A1(mai_mai_n121_), .B0(mai_mai_n120_), .B1(mai_mai_n119_), .Y(mai_mai_n122_));
  NO2        m106(.A(mai_mai_n122_), .B(mai_mai_n77_), .Y(mai_mai_n123_));
  NO2        m107(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n124_));
  NA2        m108(.A(mai_mai_n35_), .B(mai_mai_n124_), .Y(mai_mai_n125_));
  NAi21      m109(.An(x0), .B(x4), .Y(mai_mai_n126_));
  NO2        m110(.A(mai_mai_n126_), .B(x1), .Y(mai_mai_n127_));
  NO2        m111(.A(x7), .B(x0), .Y(mai_mai_n128_));
  NO2        m112(.A(mai_mai_n83_), .B(mai_mai_n100_), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n129_), .B(x3), .Y(mai_mai_n130_));
  OAI210     m114(.A0(mai_mai_n128_), .A1(mai_mai_n127_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n132_));
  NA2        m116(.A(x5), .B(x0), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n134_));
  NA3        m118(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n132_), .Y(mai_mai_n135_));
  NA4        m119(.A(mai_mai_n135_), .B(mai_mai_n131_), .C(mai_mai_n125_), .D(mai_mai_n36_), .Y(mai_mai_n136_));
  NO3        m120(.A(mai_mai_n136_), .B(mai_mai_n123_), .C(mai_mai_n114_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n138_));
  AOI220     m122(.A0(mai_mai_n119_), .A1(mai_mai_n138_), .B0(mai_mai_n67_), .B1(mai_mai_n17_), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n139_), .B(mai_mai_n60_), .Y(mai_mai_n140_));
  NA2        m124(.A(x7), .B(x3), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n99_), .B(x5), .Y(mai_mai_n142_));
  NO2        m126(.A(x9), .B(x7), .Y(mai_mai_n143_));
  NOi21      m127(.An(x8), .B(x0), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n145_));
  INV        m129(.A(x7), .Y(mai_mai_n146_));
  NA2        m130(.A(mai_mai_n146_), .B(mai_mai_n18_), .Y(mai_mai_n147_));
  AOI220     m131(.A0(mai_mai_n147_), .A1(mai_mai_n145_), .B0(mai_mai_n110_), .B1(mai_mai_n38_), .Y(mai_mai_n148_));
  NO2        m132(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n149_), .B(mai_mai_n121_), .Y(mai_mai_n150_));
  NO2        m134(.A(mai_mai_n150_), .B(mai_mai_n148_), .Y(mai_mai_n151_));
  INV        m135(.A(mai_mai_n151_), .Y(mai_mai_n152_));
  OAI210     m136(.A0(mai_mai_n141_), .A1(mai_mai_n50_), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  NA2        m137(.A(x5), .B(x1), .Y(mai_mai_n154_));
  INV        m138(.A(mai_mai_n154_), .Y(mai_mai_n155_));
  AOI210     m139(.A0(mai_mai_n155_), .A1(mai_mai_n121_), .B0(mai_mai_n36_), .Y(mai_mai_n156_));
  NO2        m140(.A(mai_mai_n62_), .B(mai_mai_n91_), .Y(mai_mai_n157_));
  NAi31      m141(.An(mai_mai_n77_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n158_));
  NA2        m142(.A(mai_mai_n158_), .B(mai_mai_n156_), .Y(mai_mai_n159_));
  NO3        m143(.A(mai_mai_n159_), .B(mai_mai_n153_), .C(mai_mai_n140_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n137_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n133_), .B(mai_mai_n129_), .Y(mai_mai_n162_));
  NA2        m146(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n163_));
  NA2        m147(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n164_));
  NA3        m148(.A(mai_mai_n164_), .B(mai_mai_n163_), .C(mai_mai_n24_), .Y(mai_mai_n165_));
  AN2        m149(.A(mai_mai_n165_), .B(mai_mai_n134_), .Y(mai_mai_n166_));
  NA2        m150(.A(x8), .B(x0), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n146_), .B(mai_mai_n25_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n119_), .B(x4), .Y(mai_mai_n169_));
  NA2        m153(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NO2        m154(.A(mai_mai_n167_), .B(mai_mai_n170_), .Y(mai_mai_n171_));
  NA2        m155(.A(x2), .B(x0), .Y(mai_mai_n172_));
  NA2        m156(.A(x4), .B(x1), .Y(mai_mai_n173_));
  NAi21      m157(.An(mai_mai_n118_), .B(mai_mai_n173_), .Y(mai_mai_n174_));
  NOi31      m158(.An(mai_mai_n174_), .B(mai_mai_n149_), .C(mai_mai_n172_), .Y(mai_mai_n175_));
  NO4        m159(.A(mai_mai_n175_), .B(mai_mai_n171_), .C(mai_mai_n166_), .D(mai_mai_n162_), .Y(mai_mai_n176_));
  NO2        m160(.A(mai_mai_n176_), .B(mai_mai_n43_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n165_), .B(mai_mai_n75_), .Y(mai_mai_n178_));
  INV        m162(.A(mai_mai_n124_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n106_), .B(mai_mai_n17_), .Y(mai_mai_n180_));
  NO2        m164(.A(mai_mai_n35_), .B(mai_mai_n180_), .Y(mai_mai_n181_));
  NO3        m165(.A(mai_mai_n181_), .B(mai_mai_n179_), .C(x7), .Y(mai_mai_n182_));
  NA3        m166(.A(mai_mai_n174_), .B(mai_mai_n179_), .C(mai_mai_n42_), .Y(mai_mai_n183_));
  OAI210     m167(.A0(mai_mai_n164_), .A1(mai_mai_n129_), .B0(mai_mai_n183_), .Y(mai_mai_n184_));
  NO3        m168(.A(mai_mai_n184_), .B(mai_mai_n182_), .C(mai_mai_n178_), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n185_), .B(x3), .Y(mai_mai_n186_));
  NO3        m170(.A(mai_mai_n186_), .B(mai_mai_n177_), .C(mai_mai_n161_), .Y(mai03));
  NO2        m171(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n188_));
  NO2        m172(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n189_));
  OAI220     m173(.A0(mai_mai_n54_), .A1(mai_mai_n17_), .B0(x6), .B1(mai_mai_n106_), .Y(mai_mai_n190_));
  NA2        m174(.A(mai_mai_n190_), .B(mai_mai_n188_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n77_), .B(x6), .Y(mai_mai_n192_));
  NA2        m176(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n193_), .B(x4), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n195_));
  NA2        m179(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n196_));
  NO2        m180(.A(mai_mai_n196_), .B(mai_mai_n193_), .Y(mai_mai_n197_));
  AOI210     m181(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n172_), .Y(mai_mai_n198_));
  AOI210     m182(.A0(mai_mai_n198_), .A1(mai_mai_n25_), .B0(mai_mai_n197_), .Y(mai_mai_n199_));
  NO2        m183(.A(x5), .B(x1), .Y(mai_mai_n200_));
  AOI220     m184(.A0(mai_mai_n200_), .A1(mai_mai_n17_), .B0(mai_mai_n103_), .B1(x5), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n196_), .B(mai_mai_n163_), .Y(mai_mai_n202_));
  NO3        m186(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  OAI210     m188(.A0(mai_mai_n201_), .A1(mai_mai_n64_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  AOI220     m189(.A0(mai_mai_n205_), .A1(mai_mai_n48_), .B0(x1), .B1(mai_mai_n124_), .Y(mai_mai_n206_));
  NA3        m190(.A(mai_mai_n206_), .B(mai_mai_n199_), .C(mai_mai_n191_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n19_), .Y(mai_mai_n209_));
  NO2        m193(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n210_));
  NO2        m194(.A(mai_mai_n210_), .B(x6), .Y(mai_mai_n211_));
  NOi21      m195(.An(mai_mai_n83_), .B(mai_mai_n211_), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n212_), .B(mai_mai_n146_), .Y(mai_mai_n213_));
  AO210      m197(.A0(mai_mai_n213_), .A1(mai_mai_n209_), .B0(mai_mai_n168_), .Y(mai_mai_n214_));
  NA2        m198(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n215_));
  NO3        m199(.A(mai_mai_n173_), .B(mai_mai_n62_), .C(x6), .Y(mai_mai_n216_));
  AOI220     m200(.A0(mai_mai_n216_), .A1(mai_mai_n17_), .B0(mai_mai_n134_), .B1(mai_mai_n90_), .Y(mai_mai_n217_));
  NA2        m201(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n218_));
  INV        m202(.A(mai_mai_n202_), .Y(mai_mai_n219_));
  NA2        m203(.A(mai_mai_n189_), .B(mai_mai_n127_), .Y(mai_mai_n220_));
  NA2        m204(.A(mai_mai_n124_), .B(x6), .Y(mai_mai_n221_));
  OAI210     m205(.A0(mai_mai_n91_), .A1(mai_mai_n36_), .B0(mai_mai_n67_), .Y(mai_mai_n222_));
  NA4        m206(.A(mai_mai_n222_), .B(mai_mai_n221_), .C(mai_mai_n220_), .D(mai_mai_n219_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n223_), .B(x2), .Y(mai_mai_n224_));
  NA3        m208(.A(mai_mai_n224_), .B(mai_mai_n217_), .C(mai_mai_n214_), .Y(mai_mai_n225_));
  AOI210     m209(.A0(mai_mai_n207_), .A1(x8), .B0(mai_mai_n225_), .Y(mai_mai_n226_));
  NO2        m210(.A(mai_mai_n91_), .B(x3), .Y(mai_mai_n227_));
  NO3        m211(.A(mai_mai_n89_), .B(mai_mai_n78_), .C(mai_mai_n25_), .Y(mai_mai_n228_));
  NO2        m212(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n229_));
  AOI220     m213(.A0(mai_mai_n194_), .A1(mai_mai_n180_), .B0(mai_mai_n229_), .B1(mai_mai_n67_), .Y(mai_mai_n230_));
  NA3        m214(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n231_));
  NO2        m215(.A(mai_mai_n231_), .B(mai_mai_n399_), .Y(mai_mai_n232_));
  NA2        m216(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n233_));
  NA2        m217(.A(mai_mai_n232_), .B(mai_mai_n118_), .Y(mai_mai_n234_));
  INV        m218(.A(x6), .Y(mai_mai_n235_));
  NO2        m219(.A(mai_mai_n196_), .B(x6), .Y(mai_mai_n236_));
  NA2        m220(.A(mai_mai_n235_), .B(mai_mai_n138_), .Y(mai_mai_n237_));
  NA4        m221(.A(mai_mai_n237_), .B(mai_mai_n234_), .C(mai_mai_n230_), .D(mai_mai_n146_), .Y(mai_mai_n238_));
  NA2        m222(.A(mai_mai_n189_), .B(mai_mai_n210_), .Y(mai_mai_n239_));
  NO2        m223(.A(x9), .B(x6), .Y(mai_mai_n240_));
  NO2        m224(.A(mai_mai_n133_), .B(mai_mai_n18_), .Y(mai_mai_n241_));
  NAi21      m225(.An(mai_mai_n241_), .B(mai_mai_n231_), .Y(mai_mai_n242_));
  AOI210     m226(.A0(x3), .A1(x2), .B0(mai_mai_n48_), .Y(mai_mai_n243_));
  OAI210     m227(.A0(mai_mai_n133_), .A1(x3), .B0(mai_mai_n243_), .Y(mai_mai_n244_));
  AOI220     m228(.A0(mai_mai_n244_), .A1(x1), .B0(mai_mai_n242_), .B1(mai_mai_n240_), .Y(mai_mai_n245_));
  NA2        m229(.A(mai_mai_n245_), .B(mai_mai_n239_), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n247_));
  NO3        m231(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n248_));
  NA2        m232(.A(x6), .B(x2), .Y(mai_mai_n249_));
  OAI210     m233(.A0(mai_mai_n400_), .A1(mai_mai_n43_), .B0(mai_mai_n169_), .Y(mai_mai_n250_));
  OAI210     m234(.A0(mai_mai_n250_), .A1(mai_mai_n189_), .B0(mai_mai_n246_), .Y(mai_mai_n251_));
  NA2        m235(.A(x9), .B(mai_mai_n43_), .Y(mai_mai_n252_));
  OR2        m236(.A(mai_mai_n192_), .B(mai_mai_n142_), .Y(mai_mai_n253_));
  NA2        m237(.A(x4), .B(x0), .Y(mai_mai_n254_));
  NA2        m238(.A(mai_mai_n253_), .B(mai_mai_n42_), .Y(mai_mai_n255_));
  AOI210     m239(.A0(mai_mai_n255_), .A1(mai_mai_n251_), .B0(x8), .Y(mai_mai_n256_));
  OAI210     m240(.A0(mai_mai_n241_), .A1(mai_mai_n200_), .B0(x6), .Y(mai_mai_n257_));
  INV        m241(.A(mai_mai_n167_), .Y(mai_mai_n258_));
  OAI210     m242(.A0(mai_mai_n258_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n259_));
  AOI210     m243(.A0(mai_mai_n259_), .A1(mai_mai_n257_), .B0(mai_mai_n215_), .Y(mai_mai_n260_));
  NO4        m244(.A(mai_mai_n260_), .B(mai_mai_n256_), .C(mai_mai_n238_), .D(mai_mai_n228_), .Y(mai_mai_n261_));
  NO2        m245(.A(mai_mai_n157_), .B(x1), .Y(mai_mai_n262_));
  NO3        m246(.A(mai_mai_n262_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n263_));
  OAI210     m247(.A0(mai_mai_n263_), .A1(mai_mai_n236_), .B0(x2), .Y(mai_mai_n264_));
  OAI210     m248(.A0(mai_mai_n258_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n265_));
  AOI210     m249(.A0(mai_mai_n265_), .A1(mai_mai_n264_), .B0(mai_mai_n179_), .Y(mai_mai_n266_));
  NOi21      m250(.An(mai_mai_n249_), .B(mai_mai_n17_), .Y(mai_mai_n267_));
  NA3        m251(.A(mai_mai_n267_), .B(mai_mai_n200_), .C(mai_mai_n40_), .Y(mai_mai_n268_));
  AOI210     m252(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n269_));
  NA3        m253(.A(mai_mai_n269_), .B(mai_mai_n155_), .C(mai_mai_n32_), .Y(mai_mai_n270_));
  NA2        m254(.A(x3), .B(x2), .Y(mai_mai_n271_));
  AOI220     m255(.A0(mai_mai_n271_), .A1(mai_mai_n215_), .B0(mai_mai_n270_), .B1(mai_mai_n268_), .Y(mai_mai_n272_));
  NAi21      m256(.An(x4), .B(x0), .Y(mai_mai_n273_));
  NO3        m257(.A(mai_mai_n273_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n274_));
  OAI210     m258(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  OAI220     m259(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n276_));
  OAI210     m260(.A0(mai_mai_n269_), .A1(mai_mai_n267_), .B0(x6), .Y(mai_mai_n277_));
  AOI220     m261(.A0(mai_mai_n277_), .A1(mai_mai_n81_), .B0(mai_mai_n276_), .B1(mai_mai_n31_), .Y(mai_mai_n278_));
  AOI210     m262(.A0(mai_mai_n278_), .A1(mai_mai_n275_), .B0(mai_mai_n25_), .Y(mai_mai_n279_));
  NA3        m263(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n280_));
  OAI210     m264(.A0(mai_mai_n269_), .A1(mai_mai_n267_), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  NA2        m265(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n282_));
  OR2        m266(.A(mai_mai_n282_), .B(mai_mai_n254_), .Y(mai_mai_n283_));
  NO2        m267(.A(mai_mai_n283_), .B(mai_mai_n154_), .Y(mai_mai_n284_));
  AO210      m268(.A0(mai_mai_n281_), .A1(mai_mai_n142_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  NO4        m269(.A(mai_mai_n285_), .B(mai_mai_n279_), .C(mai_mai_n272_), .D(mai_mai_n266_), .Y(mai_mai_n286_));
  OAI210     m270(.A0(mai_mai_n261_), .A1(mai_mai_n226_), .B0(mai_mai_n286_), .Y(mai04));
  OAI210     m271(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n288_));
  NA3        m272(.A(mai_mai_n288_), .B(mai_mai_n248_), .C(mai_mai_n84_), .Y(mai_mai_n289_));
  NO2        m273(.A(x2), .B(x1), .Y(mai_mai_n290_));
  OAI210     m274(.A0(mai_mai_n233_), .A1(mai_mai_n290_), .B0(mai_mai_n36_), .Y(mai_mai_n291_));
  NO2        m275(.A(mai_mai_n247_), .B(mai_mai_n89_), .Y(mai_mai_n292_));
  NA2        m276(.A(mai_mai_n36_), .B(mai_mai_n291_), .Y(mai_mai_n293_));
  NA2        m277(.A(x6), .B(x3), .Y(mai_mai_n294_));
  OAI210     m278(.A0(mai_mai_n247_), .A1(mai_mai_n280_), .B0(mai_mai_n282_), .Y(mai_mai_n295_));
  AOI210     m279(.A0(mai_mai_n144_), .A1(mai_mai_n63_), .B0(mai_mai_n295_), .Y(mai_mai_n296_));
  NA2        m280(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n297_));
  OAI210     m281(.A0(mai_mai_n106_), .A1(mai_mai_n17_), .B0(mai_mai_n297_), .Y(mai_mai_n298_));
  AOI220     m282(.A0(mai_mai_n298_), .A1(mai_mai_n78_), .B0(mai_mai_n292_), .B1(mai_mai_n91_), .Y(mai_mai_n299_));
  NA3        m283(.A(mai_mai_n299_), .B(mai_mai_n296_), .C(mai_mai_n294_), .Y(mai_mai_n300_));
  OAI210     m284(.A0(mai_mai_n111_), .A1(x3), .B0(mai_mai_n274_), .Y(mai_mai_n301_));
  NA2        m285(.A(mai_mai_n301_), .B(mai_mai_n146_), .Y(mai_mai_n302_));
  AOI210     m286(.A0(mai_mai_n300_), .A1(x4), .B0(mai_mai_n302_), .Y(mai_mai_n303_));
  NA2        m287(.A(mai_mai_n403_), .B(mai_mai_n91_), .Y(mai_mai_n304_));
  NOi21      m288(.An(x4), .B(x0), .Y(mai_mai_n305_));
  NA2        m289(.A(x2), .B(x8), .Y(mai_mai_n306_));
  AOI210     m290(.A0(mai_mai_n306_), .A1(mai_mai_n304_), .B0(x3), .Y(mai_mai_n307_));
  NO2        m291(.A(mai_mai_n91_), .B(x4), .Y(mai_mai_n308_));
  NA2        m292(.A(mai_mai_n308_), .B(mai_mai_n44_), .Y(mai_mai_n309_));
  NO2        m293(.A(mai_mai_n28_), .B(mai_mai_n24_), .Y(mai_mai_n310_));
  INV        m294(.A(mai_mai_n310_), .Y(mai_mai_n311_));
  NA4        m295(.A(mai_mai_n311_), .B(mai_mai_n309_), .C(mai_mai_n209_), .D(x6), .Y(mai_mai_n312_));
  NO2        m296(.A(mai_mai_n144_), .B(mai_mai_n106_), .Y(mai_mai_n313_));
  AOI210     m297(.A0(mai_mai_n401_), .A1(mai_mai_n61_), .B0(mai_mai_n313_), .Y(mai_mai_n314_));
  NO2        m298(.A(mai_mai_n144_), .B(mai_mai_n80_), .Y(mai_mai_n315_));
  NO2        m299(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n316_));
  NOi21      m300(.An(mai_mai_n118_), .B(mai_mai_n27_), .Y(mai_mai_n317_));
  AOI210     m301(.A0(mai_mai_n316_), .A1(mai_mai_n315_), .B0(mai_mai_n317_), .Y(mai_mai_n318_));
  OAI210     m302(.A0(mai_mai_n314_), .A1(mai_mai_n62_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  OAI220     m303(.A0(mai_mai_n319_), .A1(x6), .B0(mai_mai_n312_), .B1(mai_mai_n307_), .Y(mai_mai_n320_));
  OAI210     m304(.A0(mai_mai_n404_), .A1(mai_mai_n91_), .B0(mai_mai_n283_), .Y(mai_mai_n321_));
  AOI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n18_), .B0(mai_mai_n146_), .Y(mai_mai_n322_));
  AO220      m306(.A0(mai_mai_n322_), .A1(mai_mai_n320_), .B0(mai_mai_n303_), .B1(mai_mai_n293_), .Y(mai_mai_n323_));
  NA2        m307(.A(mai_mai_n316_), .B(x6), .Y(mai_mai_n324_));
  INV        m308(.A(mai_mai_n145_), .Y(mai_mai_n325_));
  NA2        m309(.A(mai_mai_n308_), .B(x0), .Y(mai_mai_n326_));
  NA2        m310(.A(mai_mai_n83_), .B(x6), .Y(mai_mai_n327_));
  OAI210     m311(.A0(mai_mai_n326_), .A1(mai_mai_n325_), .B0(mai_mai_n327_), .Y(mai_mai_n328_));
  AOI220     m312(.A0(mai_mai_n328_), .A1(mai_mai_n324_), .B0(mai_mai_n203_), .B1(mai_mai_n49_), .Y(mai_mai_n329_));
  NA3        m313(.A(mai_mai_n329_), .B(mai_mai_n323_), .C(mai_mai_n289_), .Y(mai_mai_n330_));
  AOI210     m314(.A0(x2), .A1(x8), .B0(mai_mai_n111_), .Y(mai_mai_n331_));
  INV        m315(.A(mai_mai_n331_), .Y(mai_mai_n332_));
  NA3        m316(.A(mai_mai_n332_), .B(mai_mai_n188_), .C(mai_mai_n146_), .Y(mai_mai_n333_));
  OAI210     m317(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n215_), .Y(mai_mai_n334_));
  AO220      m318(.A0(mai_mai_n334_), .A1(mai_mai_n143_), .B0(mai_mai_n110_), .B1(x4), .Y(mai_mai_n335_));
  NA2        m319(.A(mai_mai_n335_), .B(mai_mai_n116_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(mai_mai_n336_), .A1(mai_mai_n333_), .B0(mai_mai_n25_), .Y(mai_mai_n337_));
  NA2        m321(.A(mai_mai_n68_), .B(mai_mai_n195_), .Y(mai_mai_n338_));
  NA3        m322(.A(x2), .B(mai_mai_n210_), .C(x8), .Y(mai_mai_n339_));
  AOI210     m323(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n25_), .Y(mai_mai_n340_));
  AOI210     m324(.A0(mai_mai_n117_), .A1(mai_mai_n115_), .B0(mai_mai_n42_), .Y(mai_mai_n341_));
  NOi21      m325(.An(mai_mai_n341_), .B(mai_mai_n173_), .Y(mai_mai_n342_));
  OAI210     m326(.A0(mai_mai_n342_), .A1(mai_mai_n340_), .B0(mai_mai_n143_), .Y(mai_mai_n343_));
  NAi31      m327(.An(mai_mai_n50_), .B(mai_mai_n262_), .C(mai_mai_n168_), .Y(mai_mai_n344_));
  NA2        m328(.A(mai_mai_n344_), .B(mai_mai_n343_), .Y(mai_mai_n345_));
  OAI210     m329(.A0(mai_mai_n345_), .A1(mai_mai_n337_), .B0(x6), .Y(mai_mai_n346_));
  INV        m330(.A(mai_mai_n128_), .Y(mai_mai_n347_));
  NA3        m331(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n348_));
  AOI220     m332(.A0(mai_mai_n348_), .A1(mai_mai_n347_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n349_));
  NA2        m333(.A(mai_mai_n188_), .B(mai_mai_n146_), .Y(mai_mai_n350_));
  INV        m334(.A(x1), .Y(mai_mai_n351_));
  OAI210     m335(.A0(mai_mai_n350_), .A1(x8), .B0(mai_mai_n351_), .Y(mai_mai_n352_));
  NAi31      m336(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n353_));
  NO2        m337(.A(mai_mai_n353_), .B(x4), .Y(mai_mai_n354_));
  NA3        m338(.A(mai_mai_n354_), .B(mai_mai_n141_), .C(x9), .Y(mai_mai_n355_));
  NO3        m339(.A(x8), .B(mai_mai_n273_), .C(x2), .Y(mai_mai_n356_));
  NOi21      m340(.An(mai_mai_n120_), .B(mai_mai_n172_), .Y(mai_mai_n357_));
  NO3        m341(.A(mai_mai_n357_), .B(mai_mai_n356_), .C(mai_mai_n18_), .Y(mai_mai_n358_));
  AOI220     m342(.A0(x7), .A1(mai_mai_n227_), .B0(mai_mai_n315_), .B1(mai_mai_n146_), .Y(mai_mai_n359_));
  NA4        m343(.A(mai_mai_n359_), .B(mai_mai_n358_), .C(mai_mai_n355_), .D(mai_mai_n50_), .Y(mai_mai_n360_));
  OAI210     m344(.A0(mai_mai_n352_), .A1(mai_mai_n349_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  NO2        m345(.A(mai_mai_n120_), .B(mai_mai_n43_), .Y(mai_mai_n362_));
  NOi31      m346(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n363_));
  AOI210     m347(.A0(mai_mai_n121_), .A1(x3), .B0(mai_mai_n305_), .Y(mai_mai_n364_));
  NA2        m348(.A(x3), .B(mai_mai_n364_), .Y(mai_mai_n365_));
  NO3        m349(.A(mai_mai_n365_), .B(mai_mai_n362_), .C(x2), .Y(mai_mai_n366_));
  INV        m350(.A(mai_mai_n366_), .Y(mai_mai_n367_));
  AOI210     m351(.A0(mai_mai_n367_), .A1(mai_mai_n361_), .B0(mai_mai_n25_), .Y(mai_mai_n368_));
  NO3        m352(.A(mai_mai_n68_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n369_));
  AOI220     m353(.A0(mai_mai_n369_), .A1(mai_mai_n243_), .B0(mai_mai_n402_), .B1(mai_mai_n341_), .Y(mai_mai_n370_));
  NO2        m354(.A(mai_mai_n370_), .B(mai_mai_n103_), .Y(mai_mai_n371_));
  NA2        m355(.A(mai_mai_n371_), .B(x7), .Y(mai_mai_n372_));
  NA2        m356(.A(x9), .B(x7), .Y(mai_mai_n373_));
  NA3        m357(.A(mai_mai_n373_), .B(mai_mai_n145_), .C(mai_mai_n127_), .Y(mai_mai_n374_));
  NA2        m358(.A(mai_mai_n374_), .B(mai_mai_n372_), .Y(mai_mai_n375_));
  OAI210     m359(.A0(mai_mai_n375_), .A1(mai_mai_n368_), .B0(mai_mai_n36_), .Y(mai_mai_n376_));
  NA2        m360(.A(mai_mai_n233_), .B(mai_mai_n21_), .Y(mai_mai_n377_));
  NO2        m361(.A(mai_mai_n154_), .B(mai_mai_n128_), .Y(mai_mai_n378_));
  NA2        m362(.A(mai_mai_n378_), .B(mai_mai_n377_), .Y(mai_mai_n379_));
  AOI210     m363(.A0(mai_mai_n379_), .A1(mai_mai_n158_), .B0(mai_mai_n28_), .Y(mai_mai_n380_));
  AOI220     m364(.A0(x3), .A1(mai_mai_n91_), .B0(mai_mai_n144_), .B1(x2), .Y(mai_mai_n381_));
  NA3        m365(.A(mai_mai_n381_), .B(mai_mai_n353_), .C(mai_mai_n89_), .Y(mai_mai_n382_));
  NA2        m366(.A(mai_mai_n382_), .B(mai_mai_n168_), .Y(mai_mai_n383_));
  OAI220     m367(.A0(mai_mai_n252_), .A1(x2), .B0(mai_mai_n154_), .B1(mai_mai_n43_), .Y(mai_mai_n384_));
  INV        m368(.A(mai_mai_n72_), .Y(mai_mai_n385_));
  NO3        m369(.A(mai_mai_n363_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n386_));
  NO2        m370(.A(mai_mai_n386_), .B(mai_mai_n385_), .Y(mai_mai_n387_));
  INV        m371(.A(mai_mai_n387_), .Y(mai_mai_n388_));
  AOI220     m372(.A0(mai_mai_n388_), .A1(x0), .B0(mai_mai_n384_), .B1(mai_mai_n128_), .Y(mai_mai_n389_));
  AOI210     m373(.A0(mai_mai_n389_), .A1(mai_mai_n383_), .B0(mai_mai_n218_), .Y(mai_mai_n390_));
  INV        m374(.A(x5), .Y(mai_mai_n391_));
  NO4        m375(.A(mai_mai_n106_), .B(mai_mai_n391_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n392_));
  NO3        m376(.A(mai_mai_n392_), .B(mai_mai_n390_), .C(mai_mai_n380_), .Y(mai_mai_n393_));
  NA3        m377(.A(mai_mai_n393_), .B(mai_mai_n376_), .C(mai_mai_n346_), .Y(mai_mai_n394_));
  AOI210     m378(.A0(mai_mai_n330_), .A1(mai_mai_n25_), .B0(mai_mai_n394_), .Y(mai05));
  INV        m379(.A(x8), .Y(mai_mai_n398_));
  INV        m380(.A(x6), .Y(mai_mai_n399_));
  INV        m381(.A(mai_mai_n248_), .Y(mai_mai_n400_));
  INV        m382(.A(mai_mai_n172_), .Y(mai_mai_n401_));
  INV        m383(.A(x4), .Y(mai_mai_n402_));
  INV        m384(.A(x2), .Y(mai_mai_n403_));
  INV        m385(.A(mai_mai_n42_), .Y(mai_mai_n404_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  NOi21      u016(.An(men_men_n23_), .B(men_men_n30_), .Y(men00));
  NO2        u017(.A(x1), .B(x0), .Y(men_men_n34_));
  INV        u018(.A(x6), .Y(men_men_n35_));
  NO2        u019(.A(men_men_n35_), .B(men_men_n25_), .Y(men_men_n36_));
  AN2        u020(.A(x8), .B(x7), .Y(men_men_n37_));
  NA3        u021(.A(men_men_n37_), .B(men_men_n36_), .C(men_men_n34_), .Y(men_men_n38_));
  NA2        u022(.A(x4), .B(x3), .Y(men_men_n39_));
  AOI210     u023(.A0(men_men_n38_), .A1(men_men_n23_), .B0(men_men_n39_), .Y(men_men_n40_));
  NO2        u024(.A(x2), .B(x0), .Y(men_men_n41_));
  INV        u025(.A(x3), .Y(men_men_n42_));
  NO2        u026(.A(men_men_n42_), .B(men_men_n18_), .Y(men_men_n43_));
  INV        u027(.A(men_men_n43_), .Y(men_men_n44_));
  NO2        u028(.A(men_men_n36_), .B(x4), .Y(men_men_n45_));
  OAI210     u029(.A0(men_men_n45_), .A1(men_men_n44_), .B0(men_men_n41_), .Y(men_men_n46_));
  INV        u030(.A(x4), .Y(men_men_n47_));
  NO2        u031(.A(men_men_n47_), .B(men_men_n17_), .Y(men_men_n48_));
  NA2        u032(.A(men_men_n48_), .B(x2), .Y(men_men_n49_));
  OAI210     u033(.A0(men_men_n49_), .A1(men_men_n20_), .B0(men_men_n46_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n51_));
  AOI220     u035(.A0(men_men_n51_), .A1(men_men_n34_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n52_));
  INV        u036(.A(x2), .Y(men_men_n53_));
  NO2        u037(.A(men_men_n53_), .B(men_men_n17_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n42_), .B(men_men_n18_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  OAI210     u040(.A0(men_men_n52_), .A1(men_men_n32_), .B0(men_men_n56_), .Y(men_men_n57_));
  NO3        u041(.A(men_men_n57_), .B(men_men_n50_), .C(men_men_n40_), .Y(men01));
  NA2        u042(.A(x8), .B(x7), .Y(men_men_n59_));
  NA2        u043(.A(men_men_n42_), .B(x1), .Y(men_men_n60_));
  INV        u044(.A(x9), .Y(men_men_n61_));
  NO2        u045(.A(men_men_n61_), .B(men_men_n35_), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n60_), .B(men_men_n59_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n60_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NO2        u051(.A(men_men_n67_), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n43_), .A1(men_men_n25_), .B0(men_men_n53_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n55_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n42_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n47_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n55_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO4        u062(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n64_), .D(men_men_n53_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(men_men_n22_), .Y(men_men_n82_));
  NO2        u066(.A(x4), .B(x2), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(x3), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n82_), .C(men_men_n18_), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n86_));
  NO3        u070(.A(x6), .B(men_men_n42_), .C(x1), .Y(men_men_n87_));
  NA2        u071(.A(men_men_n61_), .B(men_men_n47_), .Y(men_men_n88_));
  INV        u072(.A(men_men_n88_), .Y(men_men_n89_));
  OAI210     u073(.A0(men_men_n87_), .A1(men_men_n65_), .B0(men_men_n89_), .Y(men_men_n90_));
  NA2        u074(.A(x3), .B(men_men_n18_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n25_), .Y(men_men_n92_));
  INV        u076(.A(x8), .Y(men_men_n93_));
  NA2        u077(.A(x2), .B(x1), .Y(men_men_n94_));
  NO2        u078(.A(x2), .B(men_men_n92_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n26_), .Y(men_men_n96_));
  AOI210     u080(.A0(men_men_n55_), .A1(men_men_n25_), .B0(men_men_n53_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n44_), .A1(men_men_n36_), .B0(men_men_n47_), .Y(men_men_n98_));
  NO3        u082(.A(men_men_n98_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n99_));
  NA2        u083(.A(x4), .B(men_men_n42_), .Y(men_men_n100_));
  NO2        u084(.A(men_men_n47_), .B(men_men_n53_), .Y(men_men_n101_));
  OAI210     u085(.A0(men_men_n101_), .A1(men_men_n42_), .B0(men_men_n18_), .Y(men_men_n102_));
  AOI210     u086(.A0(men_men_n100_), .A1(men_men_n51_), .B0(men_men_n102_), .Y(men_men_n103_));
  NO2        u087(.A(x3), .B(x2), .Y(men_men_n104_));
  NA3        u088(.A(men_men_n104_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n105_));
  AOI210     u089(.A0(x8), .A1(x6), .B0(men_men_n105_), .Y(men_men_n106_));
  NA2        u090(.A(men_men_n53_), .B(x1), .Y(men_men_n107_));
  OAI210     u091(.A0(men_men_n107_), .A1(men_men_n39_), .B0(men_men_n17_), .Y(men_men_n108_));
  NO4        u092(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n103_), .D(men_men_n99_), .Y(men_men_n109_));
  AO220      u093(.A0(men_men_n109_), .A1(men_men_n90_), .B0(men_men_n86_), .B1(men_men_n74_), .Y(men02));
  NO2        u094(.A(x3), .B(men_men_n53_), .Y(men_men_n111_));
  NO2        u095(.A(x8), .B(men_men_n18_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n53_), .B(men_men_n17_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n42_), .B(x0), .Y(men_men_n114_));
  OAI210     u098(.A0(men_men_n88_), .A1(men_men_n113_), .B0(men_men_n114_), .Y(men_men_n115_));
  AOI220     u099(.A0(men_men_n115_), .A1(men_men_n112_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n116_));
  NO3        u100(.A(men_men_n116_), .B(x7), .C(x5), .Y(men_men_n117_));
  NA2        u101(.A(x9), .B(x2), .Y(men_men_n118_));
  OR2        u102(.A(x8), .B(x0), .Y(men_men_n119_));
  INV        u103(.A(men_men_n119_), .Y(men_men_n120_));
  NAi21      u104(.An(x2), .B(x8), .Y(men_men_n121_));
  INV        u105(.A(men_men_n121_), .Y(men_men_n122_));
  OAI210     u106(.A0(men_men_n118_), .A1(x7), .B0(men_men_n120_), .Y(men_men_n123_));
  NO2        u107(.A(x4), .B(x1), .Y(men_men_n124_));
  NA3        u108(.A(men_men_n124_), .B(men_men_n123_), .C(men_men_n59_), .Y(men_men_n125_));
  NOi21      u109(.An(x0), .B(x1), .Y(men_men_n126_));
  NO3        u110(.A(x9), .B(x8), .C(x7), .Y(men_men_n127_));
  NOi21      u111(.An(x0), .B(x4), .Y(men_men_n128_));
  NAi21      u112(.An(x8), .B(x7), .Y(men_men_n129_));
  NO2        u113(.A(men_men_n129_), .B(men_men_n61_), .Y(men_men_n130_));
  AOI220     u114(.A0(men_men_n130_), .A1(men_men_n128_), .B0(men_men_n127_), .B1(men_men_n126_), .Y(men_men_n131_));
  AOI210     u115(.A0(men_men_n131_), .A1(men_men_n125_), .B0(men_men_n77_), .Y(men_men_n132_));
  NO2        u116(.A(x5), .B(men_men_n47_), .Y(men_men_n133_));
  NA2        u117(.A(x2), .B(men_men_n18_), .Y(men_men_n134_));
  AOI210     u118(.A0(men_men_n134_), .A1(men_men_n107_), .B0(men_men_n114_), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n135_), .A1(men_men_n34_), .B0(men_men_n133_), .Y(men_men_n136_));
  NAi21      u120(.An(x0), .B(x4), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x1), .Y(men_men_n138_));
  NO2        u122(.A(x7), .B(x0), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n83_), .B(men_men_n101_), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n140_), .B(x3), .Y(men_men_n141_));
  OAI210     u125(.A0(men_men_n139_), .A1(men_men_n138_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n21_), .B(men_men_n42_), .Y(men_men_n143_));
  NA2        u127(.A(x5), .B(x0), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n47_), .B(x2), .Y(men_men_n145_));
  NA2        u129(.A(men_men_n145_), .B(men_men_n143_), .Y(men_men_n146_));
  NA4        u130(.A(men_men_n146_), .B(men_men_n142_), .C(men_men_n136_), .D(men_men_n35_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n147_), .B(men_men_n132_), .C(men_men_n117_), .Y(men_men_n148_));
  NO3        u132(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n24_), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n150_));
  AOI220     u134(.A0(men_men_n126_), .A1(men_men_n150_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n151_));
  NO3        u135(.A(men_men_n151_), .B(men_men_n59_), .C(men_men_n61_), .Y(men_men_n152_));
  NA2        u136(.A(x7), .B(x3), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n100_), .B(x5), .Y(men_men_n154_));
  NO2        u138(.A(x9), .B(x7), .Y(men_men_n155_));
  NOi21      u139(.An(x8), .B(x0), .Y(men_men_n156_));
  OA210      u140(.A0(men_men_n155_), .A1(x1), .B0(men_men_n156_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n42_), .B(x2), .Y(men_men_n158_));
  INV        u142(.A(x7), .Y(men_men_n159_));
  NA2        u143(.A(men_men_n159_), .B(men_men_n18_), .Y(men_men_n160_));
  AOI220     u144(.A0(men_men_n160_), .A1(men_men_n158_), .B0(men_men_n111_), .B1(men_men_n37_), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n25_), .B(x4), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n128_), .Y(men_men_n163_));
  NO2        u147(.A(men_men_n163_), .B(men_men_n161_), .Y(men_men_n164_));
  AOI210     u148(.A0(men_men_n157_), .A1(men_men_n154_), .B0(men_men_n164_), .Y(men_men_n165_));
  OAI210     u149(.A0(men_men_n153_), .A1(men_men_n49_), .B0(men_men_n165_), .Y(men_men_n166_));
  NA2        u150(.A(x5), .B(x1), .Y(men_men_n167_));
  NO2        u151(.A(men_men_n61_), .B(men_men_n93_), .Y(men_men_n168_));
  NAi21      u152(.An(x2), .B(x7), .Y(men_men_n169_));
  NO3        u153(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n47_), .Y(men_men_n170_));
  NA2        u154(.A(men_men_n170_), .B(men_men_n65_), .Y(men_men_n171_));
  NAi31      u155(.An(men_men_n77_), .B(men_men_n37_), .C(men_men_n34_), .Y(men_men_n172_));
  NA3        u156(.A(men_men_n172_), .B(men_men_n171_), .C(x6), .Y(men_men_n173_));
  NO4        u157(.A(men_men_n173_), .B(men_men_n166_), .C(men_men_n152_), .D(men_men_n149_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n174_), .B(men_men_n148_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n144_), .B(men_men_n140_), .Y(men_men_n176_));
  NA2        u160(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n178_));
  NA3        u162(.A(men_men_n178_), .B(men_men_n177_), .C(men_men_n24_), .Y(men_men_n179_));
  AN2        u163(.A(men_men_n179_), .B(men_men_n145_), .Y(men_men_n180_));
  NA2        u164(.A(x8), .B(x0), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n159_), .B(men_men_n25_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n126_), .B(x4), .Y(men_men_n183_));
  NA2        u167(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  AOI210     u168(.A0(men_men_n181_), .A1(men_men_n134_), .B0(men_men_n184_), .Y(men_men_n185_));
  NA2        u169(.A(x2), .B(x0), .Y(men_men_n186_));
  NA2        u170(.A(x4), .B(x1), .Y(men_men_n187_));
  NO3        u171(.A(men_men_n185_), .B(men_men_n180_), .C(men_men_n176_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n188_), .B(men_men_n42_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n179_), .B(men_men_n75_), .Y(men_men_n190_));
  INV        u174(.A(men_men_n133_), .Y(men_men_n191_));
  NA2        u175(.A(men_men_n34_), .B(men_men_n93_), .Y(men_men_n192_));
  NO3        u176(.A(men_men_n192_), .B(men_men_n191_), .C(x7), .Y(men_men_n193_));
  NO2        u177(.A(men_men_n178_), .B(men_men_n140_), .Y(men_men_n194_));
  NO3        u178(.A(men_men_n194_), .B(men_men_n193_), .C(men_men_n190_), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n195_), .B(x3), .Y(men_men_n196_));
  NO3        u180(.A(men_men_n196_), .B(men_men_n189_), .C(men_men_n175_), .Y(men03));
  NO2        u181(.A(men_men_n47_), .B(x3), .Y(men_men_n198_));
  NO2        u182(.A(x6), .B(men_men_n25_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n53_), .B(x1), .Y(men_men_n200_));
  OAI210     u184(.A0(men_men_n200_), .A1(men_men_n25_), .B0(men_men_n62_), .Y(men_men_n201_));
  OAI220     u185(.A0(men_men_n201_), .A1(men_men_n17_), .B0(men_men_n25_), .B1(men_men_n107_), .Y(men_men_n202_));
  NA2        u186(.A(men_men_n202_), .B(men_men_n198_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n77_), .B(x6), .Y(men_men_n204_));
  NA2        u188(.A(x6), .B(men_men_n25_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n205_), .B(x4), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n18_), .B(x0), .Y(men_men_n207_));
  AO220      u191(.A0(men_men_n207_), .A1(men_men_n206_), .B0(men_men_n204_), .B1(men_men_n54_), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n208_), .B(men_men_n61_), .Y(men_men_n209_));
  NA2        u193(.A(x3), .B(men_men_n17_), .Y(men_men_n210_));
  NO2        u194(.A(men_men_n210_), .B(men_men_n205_), .Y(men_men_n211_));
  NA2        u195(.A(x9), .B(men_men_n53_), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n212_), .B(x4), .Y(men_men_n213_));
  NA2        u197(.A(men_men_n205_), .B(men_men_n80_), .Y(men_men_n214_));
  AOI210     u198(.A0(men_men_n25_), .A1(x3), .B0(men_men_n186_), .Y(men_men_n215_));
  AOI220     u199(.A0(men_men_n215_), .A1(men_men_n214_), .B0(men_men_n213_), .B1(men_men_n211_), .Y(men_men_n216_));
  NO3        u200(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n217_));
  NO2        u201(.A(x5), .B(x1), .Y(men_men_n218_));
  AOI220     u202(.A0(men_men_n218_), .A1(men_men_n17_), .B0(men_men_n104_), .B1(x5), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n210_), .B(men_men_n177_), .Y(men_men_n220_));
  AOI220     u204(.A0(men_men_n462_), .A1(men_men_n47_), .B0(men_men_n217_), .B1(men_men_n133_), .Y(men_men_n221_));
  NA4        u205(.A(men_men_n221_), .B(men_men_n216_), .C(men_men_n209_), .D(men_men_n203_), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n47_), .B(men_men_n42_), .Y(men_men_n223_));
  NO2        u207(.A(x3), .B(men_men_n17_), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n224_), .B(x6), .Y(men_men_n225_));
  NOi21      u209(.An(men_men_n83_), .B(men_men_n225_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n61_), .B(men_men_n93_), .Y(men_men_n227_));
  NA3        u211(.A(men_men_n227_), .B(men_men_n224_), .C(x6), .Y(men_men_n228_));
  AOI210     u212(.A0(men_men_n228_), .A1(men_men_n226_), .B0(men_men_n159_), .Y(men_men_n229_));
  OR2        u213(.A(men_men_n229_), .B(men_men_n182_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n42_), .B(men_men_n53_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n25_), .B0(men_men_n178_), .Y(men_men_n232_));
  NO3        u216(.A(men_men_n187_), .B(men_men_n61_), .C(x6), .Y(men_men_n233_));
  AOI220     u217(.A0(men_men_n233_), .A1(men_men_n232_), .B0(men_men_n145_), .B1(men_men_n92_), .Y(men_men_n234_));
  NA2        u218(.A(x6), .B(men_men_n47_), .Y(men_men_n235_));
  OAI210     u219(.A0(men_men_n120_), .A1(men_men_n78_), .B0(x4), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n77_), .Y(men_men_n237_));
  NO2        u221(.A(men_men_n61_), .B(x6), .Y(men_men_n238_));
  NO2        u222(.A(men_men_n167_), .B(men_men_n42_), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n239_), .A1(men_men_n220_), .B0(men_men_n238_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n199_), .B(men_men_n138_), .Y(men_men_n241_));
  NA3        u225(.A(men_men_n210_), .B(men_men_n133_), .C(x6), .Y(men_men_n242_));
  OAI210     u226(.A0(men_men_n93_), .A1(men_men_n35_), .B0(men_men_n65_), .Y(men_men_n243_));
  NA4        u227(.A(men_men_n243_), .B(men_men_n242_), .C(men_men_n241_), .D(men_men_n240_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n237_), .B0(x2), .Y(men_men_n245_));
  NA3        u229(.A(men_men_n245_), .B(men_men_n234_), .C(men_men_n230_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n222_), .A1(x8), .B0(men_men_n246_), .Y(men_men_n247_));
  NO2        u231(.A(men_men_n93_), .B(x3), .Y(men_men_n248_));
  NA2        u232(.A(men_men_n248_), .B(men_men_n206_), .Y(men_men_n249_));
  NA2        u233(.A(men_men_n225_), .B(men_men_n162_), .Y(men_men_n250_));
  AOI210     u234(.A0(men_men_n250_), .A1(men_men_n249_), .B0(x2), .Y(men_men_n251_));
  NO2        u235(.A(x4), .B(men_men_n53_), .Y(men_men_n252_));
  NA2        u236(.A(men_men_n252_), .B(men_men_n65_), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n61_), .B(x6), .Y(men_men_n254_));
  NA3        u238(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n255_), .A1(men_men_n144_), .B0(men_men_n254_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n42_), .B(men_men_n17_), .Y(men_men_n257_));
  NO2        u241(.A(men_men_n257_), .B(men_men_n25_), .Y(men_men_n258_));
  OAI210     u242(.A0(men_men_n258_), .A1(men_men_n256_), .B0(men_men_n124_), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n210_), .B(x6), .Y(men_men_n260_));
  NO2        u244(.A(men_men_n210_), .B(x6), .Y(men_men_n261_));
  NAi21      u245(.An(men_men_n168_), .B(men_men_n261_), .Y(men_men_n262_));
  NA3        u246(.A(men_men_n262_), .B(men_men_n260_), .C(men_men_n150_), .Y(men_men_n263_));
  NA4        u247(.A(men_men_n263_), .B(men_men_n259_), .C(men_men_n253_), .D(men_men_n159_), .Y(men_men_n264_));
  NA2        u248(.A(men_men_n199_), .B(men_men_n224_), .Y(men_men_n265_));
  NO2        u249(.A(men_men_n144_), .B(men_men_n18_), .Y(men_men_n266_));
  NAi21      u250(.An(men_men_n266_), .B(men_men_n255_), .Y(men_men_n267_));
  AOI210     u251(.A0(x3), .A1(x2), .B0(men_men_n47_), .Y(men_men_n268_));
  NO2        u252(.A(men_men_n47_), .B(men_men_n267_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n269_), .B(men_men_n265_), .Y(men_men_n270_));
  NA2        u254(.A(men_men_n61_), .B(x2), .Y(men_men_n271_));
  NO2        u255(.A(men_men_n271_), .B(men_men_n265_), .Y(men_men_n272_));
  NO3        u256(.A(x9), .B(x6), .C(x0), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n107_), .B(men_men_n25_), .Y(men_men_n274_));
  NA2        u258(.A(x6), .B(x2), .Y(men_men_n275_));
  NO2        u259(.A(men_men_n275_), .B(men_men_n177_), .Y(men_men_n276_));
  AOI210     u260(.A0(men_men_n274_), .A1(men_men_n273_), .B0(men_men_n276_), .Y(men_men_n277_));
  OAI220     u261(.A0(men_men_n277_), .A1(men_men_n42_), .B0(men_men_n183_), .B1(men_men_n45_), .Y(men_men_n278_));
  OAI210     u262(.A0(men_men_n278_), .A1(men_men_n272_), .B0(men_men_n270_), .Y(men_men_n279_));
  OR3        u263(.A(x9), .B(men_men_n204_), .C(men_men_n154_), .Y(men_men_n280_));
  NA2        u264(.A(x4), .B(x0), .Y(men_men_n281_));
  NO3        u265(.A(men_men_n72_), .B(men_men_n281_), .C(x6), .Y(men_men_n282_));
  AOI210     u266(.A0(men_men_n280_), .A1(men_men_n41_), .B0(men_men_n282_), .Y(men_men_n283_));
  AOI210     u267(.A0(men_men_n283_), .A1(men_men_n279_), .B0(x8), .Y(men_men_n284_));
  INV        u268(.A(men_men_n254_), .Y(men_men_n285_));
  OAI210     u269(.A0(men_men_n266_), .A1(men_men_n218_), .B0(men_men_n285_), .Y(men_men_n286_));
  AOI210     u270(.A0(men_men_n465_), .A1(men_men_n286_), .B0(men_men_n231_), .Y(men_men_n287_));
  NO4        u271(.A(men_men_n287_), .B(men_men_n284_), .C(men_men_n264_), .D(men_men_n251_), .Y(men_men_n288_));
  NO2        u272(.A(x3), .B(men_men_n35_), .Y(men_men_n289_));
  OAI210     u273(.A0(men_men_n289_), .A1(men_men_n261_), .B0(x2), .Y(men_men_n290_));
  NA2        u274(.A(x6), .B(men_men_n43_), .Y(men_men_n291_));
  AOI210     u275(.A0(men_men_n291_), .A1(men_men_n290_), .B0(men_men_n191_), .Y(men_men_n292_));
  NA2        u276(.A(x3), .B(x2), .Y(men_men_n293_));
  NAi21      u277(.An(x4), .B(x0), .Y(men_men_n294_));
  NO3        u278(.A(men_men_n294_), .B(men_men_n43_), .C(x2), .Y(men_men_n295_));
  OAI210     u279(.A0(x6), .A1(men_men_n18_), .B0(men_men_n295_), .Y(men_men_n296_));
  NO2        u280(.A(x9), .B(x8), .Y(men_men_n297_));
  NA3        u281(.A(men_men_n297_), .B(men_men_n35_), .C(men_men_n53_), .Y(men_men_n298_));
  INV        u282(.A(men_men_n298_), .Y(men_men_n299_));
  NA2        u283(.A(men_men_n299_), .B(men_men_n81_), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n300_), .A1(men_men_n296_), .B0(men_men_n25_), .Y(men_men_n301_));
  NA3        u285(.A(men_men_n35_), .B(x1), .C(men_men_n17_), .Y(men_men_n302_));
  INV        u286(.A(men_men_n220_), .Y(men_men_n303_));
  NA2        u287(.A(men_men_n35_), .B(men_men_n42_), .Y(men_men_n304_));
  OR2        u288(.A(men_men_n304_), .B(men_men_n281_), .Y(men_men_n305_));
  NO2        u289(.A(men_men_n235_), .B(men_men_n303_), .Y(men_men_n306_));
  NO3        u290(.A(men_men_n306_), .B(men_men_n301_), .C(men_men_n292_), .Y(men_men_n307_));
  OAI210     u291(.A0(men_men_n288_), .A1(men_men_n247_), .B0(men_men_n307_), .Y(men04));
  OAI210     u292(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n309_));
  NA3        u293(.A(men_men_n309_), .B(men_men_n273_), .C(men_men_n84_), .Y(men_men_n310_));
  NO2        u294(.A(x2), .B(x1), .Y(men_men_n311_));
  NO2        u295(.A(men_men_n311_), .B(men_men_n294_), .Y(men_men_n312_));
  AOI210     u296(.A0(men_men_n61_), .A1(x4), .B0(men_men_n113_), .Y(men_men_n313_));
  OAI210     u297(.A0(men_men_n313_), .A1(men_men_n312_), .B0(men_men_n248_), .Y(men_men_n314_));
  NO2        u298(.A(men_men_n271_), .B(men_men_n91_), .Y(men_men_n315_));
  NO2        u299(.A(men_men_n315_), .B(men_men_n35_), .Y(men_men_n316_));
  NO2        u300(.A(men_men_n293_), .B(men_men_n207_), .Y(men_men_n317_));
  NA2        u301(.A(x9), .B(x0), .Y(men_men_n318_));
  AOI210     u302(.A0(men_men_n91_), .A1(men_men_n75_), .B0(men_men_n318_), .Y(men_men_n319_));
  OAI210     u303(.A0(men_men_n319_), .A1(men_men_n317_), .B0(men_men_n93_), .Y(men_men_n320_));
  NA3        u304(.A(men_men_n320_), .B(men_men_n316_), .C(men_men_n314_), .Y(men_men_n321_));
  NA2        u305(.A(men_men_n321_), .B(x6), .Y(men_men_n322_));
  NO2        u306(.A(men_men_n212_), .B(men_men_n114_), .Y(men_men_n323_));
  NO3        u307(.A(men_men_n254_), .B(men_men_n121_), .C(men_men_n18_), .Y(men_men_n324_));
  NO2        u308(.A(men_men_n324_), .B(men_men_n323_), .Y(men_men_n325_));
  OAI210     u309(.A0(men_men_n119_), .A1(men_men_n107_), .B0(men_men_n181_), .Y(men_men_n326_));
  NA3        u310(.A(men_men_n326_), .B(x6), .C(x3), .Y(men_men_n327_));
  NOi21      u311(.An(men_men_n156_), .B(men_men_n134_), .Y(men_men_n328_));
  AOI210     u312(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n329_));
  OAI220     u313(.A0(men_men_n329_), .A1(men_men_n304_), .B0(men_men_n271_), .B1(men_men_n302_), .Y(men_men_n330_));
  AOI210     u314(.A0(men_men_n328_), .A1(men_men_n62_), .B0(men_men_n330_), .Y(men_men_n331_));
  NA2        u315(.A(x2), .B(men_men_n17_), .Y(men_men_n332_));
  OAI210     u316(.A0(men_men_n107_), .A1(men_men_n17_), .B0(men_men_n332_), .Y(men_men_n333_));
  AOI220     u317(.A0(men_men_n333_), .A1(men_men_n78_), .B0(men_men_n315_), .B1(men_men_n93_), .Y(men_men_n334_));
  NA4        u318(.A(men_men_n334_), .B(men_men_n331_), .C(men_men_n327_), .D(men_men_n325_), .Y(men_men_n335_));
  OAI210     u319(.A0(men_men_n112_), .A1(x3), .B0(men_men_n295_), .Y(men_men_n336_));
  NA3        u320(.A(men_men_n227_), .B(men_men_n217_), .C(men_men_n83_), .Y(men_men_n337_));
  NA3        u321(.A(men_men_n337_), .B(men_men_n336_), .C(men_men_n159_), .Y(men_men_n338_));
  AOI210     u322(.A0(men_men_n335_), .A1(x4), .B0(men_men_n338_), .Y(men_men_n339_));
  NA3        u323(.A(men_men_n312_), .B(men_men_n212_), .C(men_men_n93_), .Y(men_men_n340_));
  NOi21      u324(.An(x4), .B(x0), .Y(men_men_n341_));
  XO2        u325(.A(x4), .B(x0), .Y(men_men_n342_));
  NO2        u326(.A(men_men_n342_), .B(men_men_n118_), .Y(men_men_n343_));
  AOI220     u327(.A0(men_men_n343_), .A1(x8), .B0(men_men_n341_), .B1(men_men_n94_), .Y(men_men_n344_));
  AOI210     u328(.A0(men_men_n344_), .A1(men_men_n340_), .B0(x3), .Y(men_men_n345_));
  INV        u329(.A(men_men_n94_), .Y(men_men_n346_));
  NO2        u330(.A(men_men_n93_), .B(x4), .Y(men_men_n347_));
  AOI220     u331(.A0(men_men_n347_), .A1(men_men_n43_), .B0(men_men_n128_), .B1(men_men_n346_), .Y(men_men_n348_));
  NO3        u332(.A(men_men_n342_), .B(men_men_n168_), .C(x2), .Y(men_men_n349_));
  NO3        u333(.A(men_men_n227_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n350_));
  NO2        u334(.A(men_men_n350_), .B(men_men_n349_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n351_), .B(men_men_n348_), .C(x6), .Y(men_men_n352_));
  NO2        u336(.A(men_men_n294_), .B(men_men_n91_), .Y(men_men_n353_));
  NO2        u337(.A(men_men_n42_), .B(x0), .Y(men_men_n354_));
  OR2        u338(.A(men_men_n347_), .B(men_men_n354_), .Y(men_men_n355_));
  NO2        u339(.A(men_men_n156_), .B(men_men_n107_), .Y(men_men_n356_));
  AOI220     u340(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n353_), .B1(men_men_n60_), .Y(men_men_n357_));
  NO2        u341(.A(men_men_n156_), .B(men_men_n80_), .Y(men_men_n358_));
  NO2        u342(.A(men_men_n34_), .B(x2), .Y(men_men_n359_));
  NOi21      u343(.An(men_men_n124_), .B(men_men_n27_), .Y(men_men_n360_));
  INV        u344(.A(men_men_n360_), .Y(men_men_n361_));
  OAI210     u345(.A0(men_men_n357_), .A1(men_men_n61_), .B0(men_men_n361_), .Y(men_men_n362_));
  OAI220     u346(.A0(men_men_n362_), .A1(x6), .B0(men_men_n352_), .B1(men_men_n345_), .Y(men_men_n363_));
  OAI210     u347(.A0(men_men_n62_), .A1(men_men_n47_), .B0(men_men_n41_), .Y(men_men_n364_));
  OAI210     u348(.A0(men_men_n364_), .A1(men_men_n93_), .B0(men_men_n305_), .Y(men_men_n365_));
  AOI210     u349(.A0(men_men_n365_), .A1(men_men_n18_), .B0(men_men_n159_), .Y(men_men_n366_));
  AO220      u350(.A0(men_men_n366_), .A1(men_men_n363_), .B0(men_men_n339_), .B1(men_men_n322_), .Y(men_men_n367_));
  NA2        u351(.A(men_men_n359_), .B(x6), .Y(men_men_n368_));
  AOI210     u352(.A0(x6), .A1(x1), .B0(men_men_n158_), .Y(men_men_n369_));
  NA2        u353(.A(men_men_n347_), .B(x0), .Y(men_men_n370_));
  NA2        u354(.A(men_men_n83_), .B(x6), .Y(men_men_n371_));
  OAI210     u355(.A0(men_men_n370_), .A1(men_men_n369_), .B0(men_men_n371_), .Y(men_men_n372_));
  NA2        u356(.A(men_men_n372_), .B(men_men_n368_), .Y(men_men_n373_));
  NA3        u357(.A(men_men_n373_), .B(men_men_n367_), .C(men_men_n310_), .Y(men_men_n374_));
  AOI210     u358(.A0(men_men_n200_), .A1(x8), .B0(men_men_n112_), .Y(men_men_n375_));
  INV        u359(.A(men_men_n375_), .Y(men_men_n376_));
  NA3        u360(.A(men_men_n376_), .B(men_men_n198_), .C(men_men_n159_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n28_), .A1(x1), .B0(men_men_n231_), .Y(men_men_n378_));
  AO220      u362(.A0(men_men_n378_), .A1(men_men_n155_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n379_));
  NA3        u363(.A(x7), .B(x3), .C(x0), .Y(men_men_n380_));
  NA2        u364(.A(men_men_n223_), .B(x0), .Y(men_men_n381_));
  OAI220     u365(.A0(men_men_n381_), .A1(men_men_n212_), .B0(men_men_n380_), .B1(men_men_n346_), .Y(men_men_n382_));
  AOI210     u366(.A0(men_men_n379_), .A1(men_men_n120_), .B0(men_men_n382_), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n383_), .A1(men_men_n377_), .B0(men_men_n25_), .Y(men_men_n384_));
  NA3        u368(.A(men_men_n122_), .B(men_men_n223_), .C(x0), .Y(men_men_n385_));
  OAI210     u369(.A0(men_men_n198_), .A1(men_men_n66_), .B0(men_men_n207_), .Y(men_men_n386_));
  NA3        u370(.A(men_men_n200_), .B(men_men_n224_), .C(x8), .Y(men_men_n387_));
  AOI210     u371(.A0(men_men_n387_), .A1(men_men_n386_), .B0(men_men_n25_), .Y(men_men_n388_));
  AOI210     u372(.A0(men_men_n121_), .A1(men_men_n119_), .B0(men_men_n41_), .Y(men_men_n389_));
  NOi31      u373(.An(men_men_n389_), .B(men_men_n354_), .C(men_men_n187_), .Y(men_men_n390_));
  OAI210     u374(.A0(men_men_n390_), .A1(men_men_n388_), .B0(men_men_n155_), .Y(men_men_n391_));
  NAi31      u375(.An(men_men_n49_), .B(men_men_n463_), .C(men_men_n182_), .Y(men_men_n392_));
  NA3        u376(.A(men_men_n392_), .B(men_men_n391_), .C(men_men_n385_), .Y(men_men_n393_));
  OAI210     u377(.A0(men_men_n393_), .A1(men_men_n384_), .B0(x6), .Y(men_men_n394_));
  OAI210     u378(.A0(men_men_n168_), .A1(men_men_n47_), .B0(men_men_n139_), .Y(men_men_n395_));
  NA3        u379(.A(men_men_n54_), .B(men_men_n37_), .C(men_men_n31_), .Y(men_men_n396_));
  AOI220     u380(.A0(men_men_n396_), .A1(men_men_n395_), .B0(men_men_n39_), .B1(men_men_n32_), .Y(men_men_n397_));
  NO2        u381(.A(men_men_n159_), .B(x0), .Y(men_men_n398_));
  AOI220     u382(.A0(men_men_n398_), .A1(men_men_n223_), .B0(men_men_n198_), .B1(men_men_n159_), .Y(men_men_n399_));
  AOI210     u383(.A0(men_men_n130_), .A1(men_men_n252_), .B0(x1), .Y(men_men_n400_));
  OAI210     u384(.A0(men_men_n399_), .A1(x8), .B0(men_men_n400_), .Y(men_men_n401_));
  NAi31      u385(.An(x2), .B(x8), .C(x0), .Y(men_men_n402_));
  OAI210     u386(.A0(men_men_n402_), .A1(x4), .B0(men_men_n169_), .Y(men_men_n403_));
  NA3        u387(.A(men_men_n403_), .B(men_men_n153_), .C(x9), .Y(men_men_n404_));
  NO4        u388(.A(men_men_n129_), .B(men_men_n294_), .C(x9), .D(x2), .Y(men_men_n405_));
  NOi21      u389(.An(men_men_n127_), .B(men_men_n186_), .Y(men_men_n406_));
  NO3        u390(.A(men_men_n406_), .B(men_men_n405_), .C(men_men_n18_), .Y(men_men_n407_));
  NO3        u391(.A(x9), .B(men_men_n159_), .C(x0), .Y(men_men_n408_));
  AOI220     u392(.A0(men_men_n408_), .A1(men_men_n248_), .B0(men_men_n358_), .B1(men_men_n159_), .Y(men_men_n409_));
  NA4        u393(.A(men_men_n409_), .B(men_men_n407_), .C(men_men_n404_), .D(men_men_n49_), .Y(men_men_n410_));
  OAI210     u394(.A0(men_men_n401_), .A1(men_men_n397_), .B0(men_men_n410_), .Y(men_men_n411_));
  NOi31      u395(.An(men_men_n398_), .B(men_men_n32_), .C(x8), .Y(men_men_n412_));
  AOI210     u396(.A0(men_men_n37_), .A1(x9), .B0(men_men_n137_), .Y(men_men_n413_));
  NO3        u397(.A(men_men_n413_), .B(men_men_n127_), .C(men_men_n42_), .Y(men_men_n414_));
  NOi31      u398(.An(x1), .B(x8), .C(x7), .Y(men_men_n415_));
  AOI220     u399(.A0(men_men_n415_), .A1(men_men_n341_), .B0(men_men_n128_), .B1(x3), .Y(men_men_n416_));
  AOI210     u400(.A0(x1), .A1(men_men_n59_), .B0(men_men_n126_), .Y(men_men_n417_));
  OAI210     u401(.A0(men_men_n417_), .A1(x3), .B0(men_men_n416_), .Y(men_men_n418_));
  NO3        u402(.A(men_men_n418_), .B(men_men_n414_), .C(x2), .Y(men_men_n419_));
  OAI220     u403(.A0(men_men_n342_), .A1(men_men_n297_), .B0(men_men_n294_), .B1(men_men_n42_), .Y(men_men_n420_));
  AOI210     u404(.A0(x9), .A1(men_men_n47_), .B0(men_men_n380_), .Y(men_men_n421_));
  AOI220     u405(.A0(men_men_n421_), .A1(men_men_n93_), .B0(men_men_n420_), .B1(men_men_n159_), .Y(men_men_n422_));
  NO2        u406(.A(men_men_n422_), .B(men_men_n53_), .Y(men_men_n423_));
  NO3        u407(.A(men_men_n423_), .B(men_men_n419_), .C(men_men_n412_), .Y(men_men_n424_));
  AOI210     u408(.A0(men_men_n424_), .A1(men_men_n411_), .B0(men_men_n25_), .Y(men_men_n425_));
  NA4        u409(.A(men_men_n31_), .B(men_men_n93_), .C(x2), .D(men_men_n17_), .Y(men_men_n426_));
  NO3        u410(.A(men_men_n61_), .B(x4), .C(x1), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n428_));
  AOI220     u412(.A0(men_men_n428_), .A1(men_men_n268_), .B0(men_men_n427_), .B1(men_men_n389_), .Y(men_men_n429_));
  NO2        u413(.A(men_men_n429_), .B(men_men_n104_), .Y(men_men_n430_));
  NO3        u414(.A(men_men_n271_), .B(men_men_n181_), .C(men_men_n39_), .Y(men_men_n431_));
  OAI210     u415(.A0(men_men_n431_), .A1(men_men_n430_), .B0(x7), .Y(men_men_n432_));
  NA2        u416(.A(men_men_n227_), .B(x7), .Y(men_men_n433_));
  NA3        u417(.A(men_men_n433_), .B(men_men_n158_), .C(men_men_n138_), .Y(men_men_n434_));
  NA3        u418(.A(men_men_n434_), .B(men_men_n432_), .C(men_men_n426_), .Y(men_men_n435_));
  OAI210     u419(.A0(men_men_n435_), .A1(men_men_n425_), .B0(men_men_n35_), .Y(men_men_n436_));
  NO2        u420(.A(men_men_n408_), .B(men_men_n207_), .Y(men_men_n437_));
  NO4        u421(.A(men_men_n437_), .B(men_men_n77_), .C(x4), .D(men_men_n53_), .Y(men_men_n438_));
  NA2        u422(.A(men_men_n257_), .B(men_men_n21_), .Y(men_men_n439_));
  NO2        u423(.A(men_men_n167_), .B(men_men_n139_), .Y(men_men_n440_));
  NA2        u424(.A(men_men_n440_), .B(men_men_n439_), .Y(men_men_n441_));
  AOI210     u425(.A0(men_men_n441_), .A1(men_men_n172_), .B0(men_men_n28_), .Y(men_men_n442_));
  AOI220     u426(.A0(men_men_n354_), .A1(men_men_n93_), .B0(men_men_n156_), .B1(men_men_n200_), .Y(men_men_n443_));
  NA3        u427(.A(men_men_n443_), .B(men_men_n402_), .C(men_men_n91_), .Y(men_men_n444_));
  NA2        u428(.A(men_men_n444_), .B(men_men_n182_), .Y(men_men_n445_));
  OAI220     u429(.A0(men_men_n464_), .A1(men_men_n67_), .B0(men_men_n167_), .B1(men_men_n42_), .Y(men_men_n446_));
  NA2        u430(.A(x3), .B(men_men_n53_), .Y(men_men_n447_));
  AOI210     u431(.A0(men_men_n169_), .A1(men_men_n27_), .B0(men_men_n72_), .Y(men_men_n448_));
  OAI210     u432(.A0(men_men_n155_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n449_));
  NO3        u433(.A(men_men_n415_), .B(x3), .C(men_men_n53_), .Y(men_men_n450_));
  AOI210     u434(.A0(men_men_n450_), .A1(men_men_n449_), .B0(men_men_n448_), .Y(men_men_n451_));
  OAI210     u435(.A0(men_men_n160_), .A1(men_men_n447_), .B0(men_men_n451_), .Y(men_men_n452_));
  AOI220     u436(.A0(men_men_n452_), .A1(x0), .B0(men_men_n446_), .B1(men_men_n139_), .Y(men_men_n453_));
  AOI210     u437(.A0(men_men_n453_), .A1(men_men_n445_), .B0(men_men_n235_), .Y(men_men_n454_));
  NA2        u438(.A(x9), .B(x5), .Y(men_men_n455_));
  NO4        u439(.A(men_men_n107_), .B(men_men_n455_), .C(men_men_n59_), .D(men_men_n32_), .Y(men_men_n456_));
  NO4        u440(.A(men_men_n456_), .B(men_men_n454_), .C(men_men_n442_), .D(men_men_n438_), .Y(men_men_n457_));
  NA3        u441(.A(men_men_n457_), .B(men_men_n436_), .C(men_men_n394_), .Y(men_men_n458_));
  AOI210     u442(.A0(men_men_n374_), .A1(men_men_n25_), .B0(men_men_n458_), .Y(men05));
  INV        u443(.A(men_men_n219_), .Y(men_men_n462_));
  INV        u444(.A(x1), .Y(men_men_n463_));
  INV        u445(.A(x9), .Y(men_men_n464_));
  INV        u446(.A(men_men_n20_), .Y(men_men_n465_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule