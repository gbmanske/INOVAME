// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n142_, new_new_n143_,
    new_new_n144_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1042_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g0068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g0069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g0070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g0071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g0073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g0074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g0076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g0078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g0079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g0080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g0081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g0082(.A(i_7_), .Y(new_new_n105_));
  NA2        g0083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g0084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g0085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g0087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g0088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g0089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  AN2        g0090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g0092(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n115_));
  NO2        g0093(.A(i_8_), .B(new_new_n105_), .Y(new_new_n116_));
  NO3        g0094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g0095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g0097(.A(new_new_n119_), .B(i_0_), .Y(new_new_n120_));
  NA2        g0098(.A(i_11_), .B(i_12_), .Y(new_new_n121_));
  OAI210     g0099(.A0(new_new_n120_), .A1(new_new_n118_), .B0(new_new_n121_), .Y(new_new_n122_));
  NO2        g0100(.A(new_new_n122_), .B(new_new_n117_), .Y(new_new_n123_));
  NA3        g0101(.A(new_new_n123_), .B(new_new_n111_), .C(new_new_n104_), .Y(new_new_n124_));
  NOi21      g0102(.An(i_1_), .B(i_5_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(i_11_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g0105(.A(i_7_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NO2        g0107(.A(new_new_n129_), .B(new_new_n47_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n131_));
  NAi21      g0109(.An(i_3_), .B(i_8_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(new_new_n63_), .Y(new_new_n133_));
  NOi31      g0111(.An(new_new_n133_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n134_));
  NO2        g0112(.A(i_1_), .B(new_new_n87_), .Y(new_new_n135_));
  NO2        g0113(.A(i_6_), .B(i_5_), .Y(new_new_n136_));
  NA2        g0114(.A(new_new_n136_), .B(i_3_), .Y(new_new_n137_));
  AO210      g0115(.A0(new_new_n137_), .A1(new_new_n48_), .B0(new_new_n135_), .Y(new_new_n138_));
  OAI220     g0116(.A0(new_new_n138_), .A1(new_new_n112_), .B0(new_new_n134_), .B1(new_new_n126_), .Y(new_new_n139_));
  NO3        g0117(.A(new_new_n139_), .B(new_new_n124_), .C(new_new_n99_), .Y(new_new_n140_));
  NA3        g0118(.A(new_new_n140_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g0119(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n142_));
  INV        g0120(.A(i_6_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NA4        g0122(.A(new_new_n144_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g0123(.A(i_8_), .B(i_7_), .Y(new_new_n146_));
  NA2        g0124(.A(new_new_n146_), .B(i_6_), .Y(new_new_n147_));
  NO2        g0125(.A(i_12_), .B(i_13_), .Y(new_new_n148_));
  NAi21      g0126(.An(i_5_), .B(i_11_), .Y(new_new_n149_));
  NOi21      g0127(.An(new_new_n148_), .B(new_new_n149_), .Y(new_new_n150_));
  NO2        g0128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NA2        g0129(.A(i_2_), .B(i_3_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(i_4_), .Y(new_new_n153_));
  NA3        g0131(.A(new_new_n153_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n154_));
  AN2        g0132(.A(new_new_n148_), .B(new_new_n84_), .Y(new_new_n155_));
  NA2        g0133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  INV        g0144(.A(new_new_n166_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n147_), .Y(new_new_n168_));
  NA3        g0146(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n169_));
  NA2        g0147(.A(i_3_), .B(new_new_n49_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_4_), .B(i_9_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_11_), .B(i_13_), .Y(new_new_n172_));
  NA2        g0150(.A(new_new_n172_), .B(new_new_n171_), .Y(new_new_n173_));
  OR2        g0151(.A(new_new_n173_), .B(new_new_n170_), .Y(new_new_n174_));
  NO2        g0152(.A(i_4_), .B(i_5_), .Y(new_new_n175_));
  NAi21      g0153(.An(i_12_), .B(i_11_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n176_), .B(i_13_), .Y(new_new_n177_));
  NA3        g0155(.A(new_new_n177_), .B(new_new_n175_), .C(new_new_n84_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(new_new_n169_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n180_));
  NA2        g0158(.A(new_new_n180_), .B(new_new_n47_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n36_), .B(i_5_), .Y(new_new_n182_));
  NA2        g0160(.A(i_3_), .B(i_5_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n74_), .B(i_5_), .Y(new_new_n184_));
  NO2        g0162(.A(i_13_), .B(i_10_), .Y(new_new_n185_));
  NA3        g0163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n45_), .Y(new_new_n186_));
  NO2        g0164(.A(i_2_), .B(i_1_), .Y(new_new_n187_));
  NA2        g0165(.A(new_new_n187_), .B(i_3_), .Y(new_new_n188_));
  NAi21      g0166(.An(i_4_), .B(i_12_), .Y(new_new_n189_));
  NO4        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n186_), .D(new_new_n25_), .Y(new_new_n190_));
  NO2        g0168(.A(new_new_n190_), .B(new_new_n179_), .Y(new_new_n191_));
  INV        g0169(.A(i_8_), .Y(new_new_n192_));
  NO2        g0170(.A(new_new_n192_), .B(i_7_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_6_), .Y(new_new_n194_));
  NO3        g0172(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(new_new_n116_), .Y(new_new_n196_));
  NO3        g0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n197_));
  NO3        g0175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n198_));
  NA2        g0176(.A(i_12_), .B(new_new_n198_), .Y(new_new_n199_));
  NO2        g0177(.A(new_new_n199_), .B(new_new_n196_), .Y(new_new_n200_));
  NO2        g0178(.A(i_3_), .B(i_8_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n202_));
  NO2        g0180(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n203_));
  NO2        g0181(.A(i_13_), .B(i_9_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(i_6_), .C(new_new_n192_), .Y(new_new_n205_));
  NAi21      g0183(.An(i_12_), .B(i_3_), .Y(new_new_n206_));
  NO2        g0184(.A(new_new_n45_), .B(i_5_), .Y(new_new_n207_));
  NO3        g0185(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(new_new_n207_), .C(i_10_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n209_), .B(new_new_n205_), .Y(new_new_n210_));
  AOI210     g0188(.A0(new_new_n210_), .A1(i_7_), .B0(new_new_n200_), .Y(new_new_n211_));
  OAI220     g0189(.A0(new_new_n211_), .A1(i_4_), .B0(new_new_n194_), .B1(new_new_n191_), .Y(new_new_n212_));
  NAi21      g0190(.An(i_12_), .B(i_7_), .Y(new_new_n213_));
  NA3        g0191(.A(i_13_), .B(new_new_n192_), .C(i_10_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n214_), .B(new_new_n213_), .Y(new_new_n215_));
  NA2        g0193(.A(i_0_), .B(i_5_), .Y(new_new_n216_));
  NA2        g0194(.A(new_new_n216_), .B(new_new_n108_), .Y(new_new_n217_));
  OAI220     g0195(.A0(new_new_n217_), .A1(new_new_n188_), .B0(new_new_n181_), .B1(new_new_n137_), .Y(new_new_n218_));
  NAi31      g0196(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n36_), .B(i_13_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n222_));
  NA3        g0200(.A(new_new_n222_), .B(new_new_n221_), .C(new_new_n220_), .Y(new_new_n223_));
  INV        g0201(.A(i_13_), .Y(new_new_n224_));
  NO2        g0202(.A(i_12_), .B(new_new_n224_), .Y(new_new_n225_));
  NA3        g0203(.A(new_new_n225_), .B(new_new_n197_), .C(new_new_n195_), .Y(new_new_n226_));
  OAI210     g0204(.A0(new_new_n223_), .A1(new_new_n219_), .B0(new_new_n226_), .Y(new_new_n227_));
  AOI220     g0205(.A0(new_new_n227_), .A1(new_new_n146_), .B0(new_new_n218_), .B1(new_new_n215_), .Y(new_new_n228_));
  NO2        g0206(.A(i_12_), .B(new_new_n37_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n183_), .B(i_4_), .Y(new_new_n230_));
  NA2        g0208(.A(new_new_n230_), .B(new_new_n229_), .Y(new_new_n231_));
  OR2        g0209(.A(i_8_), .B(i_7_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n232_), .B(new_new_n87_), .Y(new_new_n233_));
  NO2        g0211(.A(new_new_n54_), .B(i_1_), .Y(new_new_n234_));
  NA2        g0212(.A(new_new_n234_), .B(new_new_n233_), .Y(new_new_n235_));
  INV        g0213(.A(i_12_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n45_), .B(new_new_n236_), .Y(new_new_n237_));
  NO3        g0215(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n238_));
  NA2        g0216(.A(i_2_), .B(i_1_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n235_), .B(new_new_n231_), .Y(new_new_n240_));
  NO3        g0218(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n241_));
  NAi21      g0219(.An(i_4_), .B(i_3_), .Y(new_new_n242_));
  NO2        g0220(.A(i_0_), .B(i_6_), .Y(new_new_n243_));
  NOi41      g0221(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n244_));
  NA2        g0222(.A(new_new_n244_), .B(new_new_n243_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n239_), .B(new_new_n183_), .Y(new_new_n246_));
  NAi21      g0224(.An(new_new_n245_), .B(new_new_n246_), .Y(new_new_n247_));
  INV        g0225(.A(new_new_n247_), .Y(new_new_n248_));
  AOI220     g0226(.A0(new_new_n248_), .A1(new_new_n40_), .B0(new_new_n240_), .B1(new_new_n204_), .Y(new_new_n249_));
  NO2        g0227(.A(i_11_), .B(new_new_n224_), .Y(new_new_n250_));
  NOi21      g0228(.An(i_1_), .B(i_6_), .Y(new_new_n251_));
  NAi21      g0229(.An(i_3_), .B(i_7_), .Y(new_new_n252_));
  NA2        g0230(.A(new_new_n236_), .B(i_9_), .Y(new_new_n253_));
  OR4        g0231(.A(new_new_n253_), .B(new_new_n252_), .C(new_new_n251_), .D(new_new_n184_), .Y(new_new_n254_));
  NO2        g0232(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n255_));
  NO2        g0233(.A(i_12_), .B(i_3_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n74_), .B(i_5_), .Y(new_new_n257_));
  NA2        g0235(.A(i_3_), .B(i_9_), .Y(new_new_n258_));
  NAi21      g0236(.An(i_7_), .B(i_10_), .Y(new_new_n259_));
  NO2        g0237(.A(new_new_n259_), .B(new_new_n258_), .Y(new_new_n260_));
  NA3        g0238(.A(new_new_n260_), .B(new_new_n257_), .C(new_new_n65_), .Y(new_new_n261_));
  NA2        g0239(.A(new_new_n261_), .B(new_new_n254_), .Y(new_new_n262_));
  NA3        g0240(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n263_));
  INV        g0241(.A(new_new_n147_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n236_), .B(i_13_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n76_), .Y(new_new_n266_));
  AOI220     g0244(.A0(new_new_n266_), .A1(new_new_n264_), .B0(new_new_n262_), .B1(new_new_n250_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n232_), .B(new_new_n37_), .Y(new_new_n268_));
  NA2        g0246(.A(i_12_), .B(i_6_), .Y(new_new_n269_));
  OR2        g0247(.A(i_13_), .B(i_9_), .Y(new_new_n270_));
  NO3        g0248(.A(new_new_n270_), .B(new_new_n269_), .C(new_new_n49_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n242_), .B(i_2_), .Y(new_new_n272_));
  NA3        g0250(.A(new_new_n272_), .B(new_new_n271_), .C(new_new_n45_), .Y(new_new_n273_));
  NA2        g0251(.A(new_new_n250_), .B(i_9_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n257_), .B(new_new_n65_), .Y(new_new_n275_));
  OAI210     g0253(.A0(new_new_n275_), .A1(new_new_n274_), .B0(new_new_n273_), .Y(new_new_n276_));
  NO3        g0254(.A(i_11_), .B(new_new_n224_), .C(new_new_n25_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n252_), .B(i_8_), .Y(new_new_n278_));
  NO2        g0256(.A(i_6_), .B(new_new_n49_), .Y(new_new_n279_));
  NO3        g0257(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n280_));
  NA2        g0258(.A(new_new_n276_), .B(new_new_n268_), .Y(new_new_n281_));
  NA4        g0259(.A(new_new_n281_), .B(new_new_n267_), .C(new_new_n249_), .D(new_new_n228_), .Y(new_new_n282_));
  NO3        g0260(.A(i_12_), .B(new_new_n224_), .C(new_new_n37_), .Y(new_new_n283_));
  INV        g0261(.A(new_new_n283_), .Y(new_new_n284_));
  NA2        g0262(.A(i_8_), .B(new_new_n105_), .Y(new_new_n285_));
  NOi21      g0263(.An(new_new_n163_), .B(new_new_n87_), .Y(new_new_n286_));
  NO3        g0264(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n287_));
  AOI220     g0265(.A0(new_new_n287_), .A1(new_new_n195_), .B0(new_new_n286_), .B1(new_new_n234_), .Y(new_new_n288_));
  NO2        g0266(.A(new_new_n288_), .B(new_new_n285_), .Y(new_new_n289_));
  NO3        g0267(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n239_), .B(i_0_), .Y(new_new_n291_));
  AOI220     g0269(.A0(new_new_n291_), .A1(new_new_n193_), .B0(new_new_n290_), .B1(new_new_n146_), .Y(new_new_n292_));
  NA2        g0270(.A(new_new_n279_), .B(new_new_n26_), .Y(new_new_n293_));
  NO2        g0271(.A(new_new_n293_), .B(new_new_n292_), .Y(new_new_n294_));
  NA2        g0272(.A(i_0_), .B(i_1_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(i_2_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n60_), .B(i_6_), .Y(new_new_n297_));
  NA3        g0275(.A(new_new_n297_), .B(new_new_n296_), .C(new_new_n163_), .Y(new_new_n298_));
  OAI210     g0276(.A0(new_new_n165_), .A1(new_new_n147_), .B0(new_new_n298_), .Y(new_new_n299_));
  NO3        g0277(.A(new_new_n299_), .B(new_new_n294_), .C(new_new_n289_), .Y(new_new_n300_));
  NO2        g0278(.A(i_3_), .B(i_10_), .Y(new_new_n301_));
  NA3        g0279(.A(new_new_n301_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n302_));
  NO2        g0280(.A(i_2_), .B(new_new_n105_), .Y(new_new_n303_));
  NA2        g0281(.A(i_1_), .B(new_new_n36_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n304_), .B(i_8_), .Y(new_new_n305_));
  NA2        g0283(.A(new_new_n305_), .B(new_new_n303_), .Y(new_new_n306_));
  AN2        g0284(.A(i_3_), .B(i_10_), .Y(new_new_n307_));
  NA4        g0285(.A(new_new_n307_), .B(new_new_n197_), .C(new_new_n177_), .D(new_new_n175_), .Y(new_new_n308_));
  NO2        g0286(.A(i_5_), .B(new_new_n37_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n310_));
  OR2        g0288(.A(new_new_n306_), .B(new_new_n302_), .Y(new_new_n311_));
  OAI220     g0289(.A0(new_new_n311_), .A1(i_6_), .B0(new_new_n300_), .B1(new_new_n284_), .Y(new_new_n312_));
  NO4        g0290(.A(new_new_n312_), .B(new_new_n282_), .C(new_new_n212_), .D(new_new_n168_), .Y(new_new_n313_));
  NO3        g0291(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n314_));
  NO2        g0292(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n315_));
  NA2        g0293(.A(new_new_n291_), .B(new_new_n315_), .Y(new_new_n316_));
  NO3        g0294(.A(i_6_), .B(new_new_n192_), .C(i_7_), .Y(new_new_n317_));
  NA2        g0295(.A(new_new_n317_), .B(new_new_n197_), .Y(new_new_n318_));
  AOI210     g0296(.A0(new_new_n318_), .A1(new_new_n316_), .B0(new_new_n170_), .Y(new_new_n319_));
  NO2        g0297(.A(i_2_), .B(i_3_), .Y(new_new_n320_));
  OR2        g0298(.A(i_0_), .B(i_5_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n216_), .B(new_new_n321_), .Y(new_new_n322_));
  NA3        g0300(.A(new_new_n291_), .B(new_new_n286_), .C(new_new_n116_), .Y(new_new_n323_));
  NAi21      g0301(.An(i_8_), .B(i_7_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n324_), .B(i_6_), .Y(new_new_n325_));
  NO2        g0303(.A(new_new_n157_), .B(new_new_n47_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n325_), .C(new_new_n163_), .Y(new_new_n327_));
  NA2        g0305(.A(new_new_n327_), .B(new_new_n323_), .Y(new_new_n328_));
  OAI210     g0306(.A0(new_new_n328_), .A1(new_new_n319_), .B0(i_4_), .Y(new_new_n329_));
  NO2        g0307(.A(i_12_), .B(i_10_), .Y(new_new_n330_));
  NOi21      g0308(.An(i_5_), .B(i_0_), .Y(new_new_n331_));
  NO3        g0309(.A(new_new_n304_), .B(new_new_n331_), .C(new_new_n132_), .Y(new_new_n332_));
  NA4        g0310(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n333_));
  NA2        g0311(.A(new_new_n332_), .B(new_new_n330_), .Y(new_new_n334_));
  NO2        g0312(.A(i_6_), .B(i_8_), .Y(new_new_n335_));
  NOi21      g0313(.An(i_0_), .B(i_2_), .Y(new_new_n336_));
  AN2        g0314(.A(new_new_n336_), .B(new_new_n335_), .Y(new_new_n337_));
  NO2        g0315(.A(i_1_), .B(i_7_), .Y(new_new_n338_));
  AO220      g0316(.A0(new_new_n338_), .A1(new_new_n337_), .B0(new_new_n325_), .B1(new_new_n234_), .Y(new_new_n339_));
  NA3        g0317(.A(new_new_n339_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n340_), .B(new_new_n334_), .C(new_new_n329_), .Y(new_new_n341_));
  NO3        g0319(.A(new_new_n232_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n342_));
  NO3        g0320(.A(new_new_n324_), .B(i_2_), .C(i_1_), .Y(new_new_n343_));
  OAI210     g0321(.A0(new_new_n343_), .A1(new_new_n342_), .B0(i_6_), .Y(new_new_n344_));
  NA3        g0322(.A(new_new_n251_), .B(new_new_n303_), .C(new_new_n192_), .Y(new_new_n345_));
  AOI210     g0323(.A0(new_new_n345_), .A1(new_new_n344_), .B0(new_new_n322_), .Y(new_new_n346_));
  NOi21      g0324(.An(new_new_n156_), .B(new_new_n108_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n347_), .B(new_new_n128_), .Y(new_new_n348_));
  OAI210     g0326(.A0(new_new_n348_), .A1(new_new_n346_), .B0(i_3_), .Y(new_new_n349_));
  INV        g0327(.A(new_new_n85_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n295_), .B(new_new_n82_), .Y(new_new_n351_));
  NO2        g0329(.A(new_new_n96_), .B(new_new_n192_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n192_), .B(i_9_), .Y(new_new_n353_));
  NA2        g0331(.A(new_new_n353_), .B(new_new_n203_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n354_), .B(new_new_n47_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n355_), .B(new_new_n294_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n356_), .A1(new_new_n349_), .B0(new_new_n162_), .Y(new_new_n357_));
  AOI210     g0335(.A0(new_new_n341_), .A1(new_new_n314_), .B0(new_new_n357_), .Y(new_new_n358_));
  NOi32      g0336(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n359_));
  INV        g0337(.A(new_new_n359_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_1_), .B(i_5_), .Y(new_new_n361_));
  INV        g0339(.A(new_new_n245_), .Y(new_new_n362_));
  NAi41      g0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n363_));
  OAI220     g0341(.A0(new_new_n363_), .A1(new_new_n361_), .B0(new_new_n219_), .B1(new_new_n159_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n363_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n365_));
  NOi32      g0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n366_));
  NAi21      g0344(.An(i_6_), .B(i_1_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n366_), .C(new_new_n47_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n368_), .B(i_0_), .Y(new_new_n369_));
  OR3        g0347(.A(new_new_n369_), .B(new_new_n365_), .C(new_new_n364_), .Y(new_new_n370_));
  NO2        g0348(.A(i_1_), .B(new_new_n105_), .Y(new_new_n371_));
  NAi21      g0349(.An(i_3_), .B(i_4_), .Y(new_new_n372_));
  NO2        g0350(.A(new_new_n372_), .B(i_9_), .Y(new_new_n373_));
  AN2        g0351(.A(i_6_), .B(i_7_), .Y(new_new_n374_));
  OAI210     g0352(.A0(new_new_n374_), .A1(new_new_n371_), .B0(new_new_n373_), .Y(new_new_n375_));
  NA2        g0353(.A(i_2_), .B(i_7_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n372_), .B(i_10_), .Y(new_new_n377_));
  NA3        g0355(.A(new_new_n377_), .B(new_new_n376_), .C(new_new_n243_), .Y(new_new_n378_));
  AOI210     g0356(.A0(new_new_n378_), .A1(new_new_n375_), .B0(new_new_n184_), .Y(new_new_n379_));
  AOI210     g0357(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n380_));
  OAI210     g0358(.A0(new_new_n380_), .A1(new_new_n187_), .B0(new_new_n377_), .Y(new_new_n381_));
  AOI220     g0359(.A0(new_new_n377_), .A1(new_new_n338_), .B0(new_new_n238_), .B1(new_new_n187_), .Y(new_new_n382_));
  AOI210     g0360(.A0(new_new_n382_), .A1(new_new_n381_), .B0(i_5_), .Y(new_new_n383_));
  NO4        g0361(.A(new_new_n383_), .B(new_new_n379_), .C(new_new_n370_), .D(new_new_n362_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n384_), .B(new_new_n360_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n386_));
  AN2        g0364(.A(i_12_), .B(i_5_), .Y(new_new_n387_));
  NO2        g0365(.A(i_4_), .B(new_new_n26_), .Y(new_new_n388_));
  NA2        g0366(.A(new_new_n388_), .B(new_new_n387_), .Y(new_new_n389_));
  NO2        g0367(.A(i_11_), .B(i_6_), .Y(new_new_n390_));
  NA3        g0368(.A(new_new_n390_), .B(new_new_n326_), .C(new_new_n224_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n389_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n242_), .B(i_5_), .Y(new_new_n393_));
  NO2        g0371(.A(i_5_), .B(i_10_), .Y(new_new_n394_));
  AOI220     g0372(.A0(new_new_n394_), .A1(new_new_n272_), .B0(new_new_n393_), .B1(new_new_n197_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n148_), .B(new_new_n46_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n396_), .B(new_new_n395_), .Y(new_new_n397_));
  OAI210     g0375(.A0(new_new_n397_), .A1(new_new_n392_), .B0(new_new_n386_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n154_), .B(new_new_n87_), .Y(new_new_n400_));
  OAI210     g0378(.A0(new_new_n400_), .A1(new_new_n392_), .B0(new_new_n399_), .Y(new_new_n401_));
  NO3        g0379(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n402_));
  NO2        g0380(.A(i_11_), .B(i_12_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n394_), .B(new_new_n236_), .Y(new_new_n404_));
  NA3        g0382(.A(new_new_n116_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n405_));
  OAI220     g0383(.A0(new_new_n405_), .A1(new_new_n219_), .B0(new_new_n404_), .B1(new_new_n333_), .Y(new_new_n406_));
  NAi21      g0384(.An(i_13_), .B(i_0_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n239_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n406_), .B(new_new_n408_), .Y(new_new_n409_));
  NA3        g0387(.A(new_new_n409_), .B(new_new_n401_), .C(new_new_n398_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n45_), .B(new_new_n224_), .Y(new_new_n411_));
  NO3        g0389(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n412_));
  NO2        g0390(.A(i_0_), .B(i_11_), .Y(new_new_n413_));
  AN2        g0391(.A(i_1_), .B(i_6_), .Y(new_new_n414_));
  NOi21      g0392(.An(i_2_), .B(i_12_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n146_), .B(i_9_), .Y(new_new_n416_));
  NAi21      g0394(.An(i_9_), .B(i_4_), .Y(new_new_n417_));
  OR2        g0395(.A(i_13_), .B(i_10_), .Y(new_new_n418_));
  NO3        g0396(.A(new_new_n418_), .B(new_new_n121_), .C(new_new_n417_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n173_), .B(new_new_n127_), .Y(new_new_n420_));
  NO2        g0398(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n283_), .B(new_new_n421_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n422_), .B(new_new_n347_), .Y(new_new_n423_));
  INV        g0401(.A(new_new_n423_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(new_new_n26_), .Y(new_new_n425_));
  INV        g0403(.A(new_new_n323_), .Y(new_new_n426_));
  NO2        g0404(.A(new_new_n183_), .B(new_new_n87_), .Y(new_new_n427_));
  AOI220     g0405(.A0(new_new_n427_), .A1(new_new_n296_), .B0(new_new_n280_), .B1(new_new_n208_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n428_), .B(new_new_n285_), .Y(new_new_n429_));
  NO2        g0407(.A(new_new_n429_), .B(new_new_n426_), .Y(new_new_n430_));
  NA2        g0408(.A(new_new_n195_), .B(new_new_n100_), .Y(new_new_n431_));
  NA3        g0409(.A(new_new_n326_), .B(new_new_n163_), .C(new_new_n87_), .Y(new_new_n432_));
  AOI210     g0410(.A0(new_new_n432_), .A1(new_new_n431_), .B0(new_new_n324_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n192_), .B(i_10_), .Y(new_new_n434_));
  NA3        g0412(.A(new_new_n257_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n435_), .B(new_new_n434_), .Y(new_new_n436_));
  NO2        g0414(.A(i_3_), .B(new_new_n49_), .Y(new_new_n437_));
  NA3        g0415(.A(new_new_n338_), .B(new_new_n337_), .C(new_new_n437_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n317_), .B(new_new_n322_), .Y(new_new_n439_));
  OAI210     g0417(.A0(new_new_n439_), .A1(new_new_n188_), .B0(new_new_n438_), .Y(new_new_n440_));
  NO3        g0418(.A(new_new_n440_), .B(new_new_n436_), .C(new_new_n433_), .Y(new_new_n441_));
  AOI210     g0419(.A0(new_new_n441_), .A1(new_new_n430_), .B0(new_new_n274_), .Y(new_new_n442_));
  NO4        g0420(.A(new_new_n442_), .B(new_new_n425_), .C(new_new_n410_), .D(new_new_n385_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n64_), .B(i_4_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n74_), .B(i_13_), .Y(new_new_n445_));
  NO2        g0423(.A(i_10_), .B(i_9_), .Y(new_new_n446_));
  NAi21      g0424(.An(i_12_), .B(i_8_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(i_3_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n310_), .B(i_0_), .Y(new_new_n449_));
  NO3        g0427(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n269_), .B(new_new_n101_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n451_), .B(new_new_n450_), .Y(new_new_n452_));
  NA2        g0430(.A(i_8_), .B(i_9_), .Y(new_new_n453_));
  AOI210     g0431(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n454_));
  OR2        g0432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n283_), .B(new_new_n203_), .Y(new_new_n456_));
  OAI220     g0434(.A0(new_new_n456_), .A1(new_new_n455_), .B0(new_new_n452_), .B1(new_new_n449_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n250_), .B(new_new_n309_), .Y(new_new_n458_));
  NO3        g0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n459_));
  INV        g0437(.A(new_new_n459_), .Y(new_new_n460_));
  NA3        g0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n461_));
  NA4        g0439(.A(new_new_n149_), .B(new_new_n119_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n461_), .B0(new_new_n460_), .B1(new_new_n458_), .Y(new_new_n463_));
  NO2        g0441(.A(new_new_n463_), .B(new_new_n457_), .Y(new_new_n464_));
  NA2        g0442(.A(new_new_n296_), .B(new_new_n112_), .Y(new_new_n465_));
  OR2        g0443(.A(new_new_n465_), .B(new_new_n205_), .Y(new_new_n466_));
  OA210      g0444(.A0(new_new_n354_), .A1(new_new_n105_), .B0(new_new_n298_), .Y(new_new_n467_));
  OA220      g0445(.A0(new_new_n467_), .A1(new_new_n162_), .B0(new_new_n466_), .B1(new_new_n231_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n100_), .B(i_13_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n427_), .B(new_new_n386_), .Y(new_new_n470_));
  NO2        g0448(.A(i_2_), .B(i_13_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n470_), .B(new_new_n469_), .Y(new_new_n472_));
  NO3        g0450(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n473_));
  NO2        g0451(.A(i_6_), .B(i_7_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NO2        g0453(.A(i_11_), .B(i_1_), .Y(new_new_n476_));
  NO2        g0454(.A(new_new_n74_), .B(i_3_), .Y(new_new_n477_));
  OR2        g0455(.A(i_11_), .B(i_8_), .Y(new_new_n478_));
  NOi21      g0456(.An(i_2_), .B(i_7_), .Y(new_new_n479_));
  NAi31      g0457(.An(new_new_n478_), .B(new_new_n479_), .C(new_new_n477_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n418_), .B(i_6_), .Y(new_new_n481_));
  NA3        g0459(.A(new_new_n481_), .B(new_new_n444_), .C(new_new_n76_), .Y(new_new_n482_));
  NO2        g0460(.A(new_new_n482_), .B(new_new_n480_), .Y(new_new_n483_));
  NO2        g0461(.A(i_6_), .B(i_10_), .Y(new_new_n484_));
  NA3        g0462(.A(new_new_n244_), .B(new_new_n172_), .C(new_new_n136_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n486_));
  NO2        g0464(.A(new_new_n157_), .B(i_3_), .Y(new_new_n487_));
  NAi31      g0465(.An(new_new_n486_), .B(new_new_n487_), .C(new_new_n225_), .Y(new_new_n488_));
  NA3        g0466(.A(new_new_n399_), .B(new_new_n180_), .C(new_new_n153_), .Y(new_new_n489_));
  NA3        g0467(.A(new_new_n489_), .B(new_new_n488_), .C(new_new_n485_), .Y(new_new_n490_));
  NO3        g0468(.A(new_new_n490_), .B(new_new_n483_), .C(new_new_n472_), .Y(new_new_n491_));
  NA2        g0469(.A(new_new_n450_), .B(new_new_n387_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n459_), .B(new_new_n394_), .Y(new_new_n493_));
  NO2        g0471(.A(new_new_n493_), .B(new_new_n223_), .Y(new_new_n494_));
  NAi21      g0472(.An(new_new_n214_), .B(new_new_n403_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n338_), .B(new_new_n216_), .Y(new_new_n496_));
  NO2        g0474(.A(new_new_n496_), .B(new_new_n495_), .Y(new_new_n497_));
  NA2        g0475(.A(new_new_n27_), .B(i_10_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n314_), .B(new_new_n238_), .Y(new_new_n499_));
  OAI220     g0477(.A0(new_new_n499_), .A1(new_new_n435_), .B0(new_new_n498_), .B1(new_new_n469_), .Y(new_new_n500_));
  NA4        g0478(.A(new_new_n307_), .B(new_new_n222_), .C(new_new_n74_), .D(new_new_n236_), .Y(new_new_n501_));
  NO2        g0479(.A(new_new_n501_), .B(new_new_n475_), .Y(new_new_n502_));
  NO4        g0480(.A(new_new_n502_), .B(new_new_n500_), .C(new_new_n497_), .D(new_new_n494_), .Y(new_new_n503_));
  NA4        g0481(.A(new_new_n503_), .B(new_new_n491_), .C(new_new_n468_), .D(new_new_n464_), .Y(new_new_n504_));
  NA3        g0482(.A(new_new_n307_), .B(new_new_n177_), .C(new_new_n175_), .Y(new_new_n505_));
  OAI210     g0483(.A0(new_new_n302_), .A1(new_new_n182_), .B0(new_new_n505_), .Y(new_new_n506_));
  AN2        g0484(.A(new_new_n287_), .B(new_new_n233_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n507_), .B(new_new_n506_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n314_), .B(new_new_n164_), .Y(new_new_n509_));
  OAI210     g0487(.A0(new_new_n509_), .A1(new_new_n231_), .B0(new_new_n308_), .Y(new_new_n510_));
  NA2        g0488(.A(new_new_n510_), .B(new_new_n325_), .Y(new_new_n511_));
  NA4        g0489(.A(new_new_n445_), .B(new_new_n444_), .C(new_new_n201_), .D(i_2_), .Y(new_new_n512_));
  INV        g0490(.A(new_new_n512_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n387_), .B(new_new_n224_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n359_), .B(new_new_n74_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n374_), .B(new_new_n366_), .Y(new_new_n516_));
  OR2        g0494(.A(new_new_n514_), .B(new_new_n516_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n36_), .B(i_8_), .Y(new_new_n518_));
  NAi41      g0496(.An(new_new_n515_), .B(new_new_n484_), .C(new_new_n518_), .D(new_new_n47_), .Y(new_new_n519_));
  AOI210     g0497(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n419_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n520_), .B(new_new_n519_), .C(new_new_n517_), .Y(new_new_n521_));
  AOI210     g0499(.A0(new_new_n513_), .A1(new_new_n202_), .B0(new_new_n521_), .Y(new_new_n522_));
  NA2        g0500(.A(new_new_n257_), .B(new_new_n65_), .Y(new_new_n523_));
  OAI210     g0501(.A0(i_8_), .A1(new_new_n523_), .B0(new_new_n138_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n524_), .B(new_new_n420_), .Y(new_new_n525_));
  NA4        g0503(.A(new_new_n525_), .B(new_new_n522_), .C(new_new_n511_), .D(new_new_n508_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n393_), .B(new_new_n296_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n389_), .A1(new_new_n169_), .B0(new_new_n527_), .Y(new_new_n528_));
  NO2        g0506(.A(i_12_), .B(new_new_n192_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n529_), .B(new_new_n224_), .Y(new_new_n530_));
  NA3        g0508(.A(new_new_n484_), .B(new_new_n175_), .C(new_new_n27_), .Y(new_new_n531_));
  NO2        g0509(.A(new_new_n531_), .B(new_new_n530_), .Y(new_new_n532_));
  NOi31      g0510(.An(new_new_n317_), .B(new_new_n418_), .C(new_new_n38_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n533_), .A1(new_new_n532_), .B0(new_new_n528_), .Y(new_new_n534_));
  NO2        g0512(.A(i_8_), .B(i_7_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n45_), .B(i_10_), .Y(new_new_n536_));
  NO2        g0514(.A(new_new_n536_), .B(i_6_), .Y(new_new_n537_));
  AOI220     g0515(.A0(new_new_n427_), .A1(new_new_n326_), .B0(new_new_n246_), .B1(new_new_n243_), .Y(new_new_n538_));
  NO2        g0516(.A(new_new_n538_), .B(new_new_n265_), .Y(new_new_n539_));
  NA2        g0517(.A(new_new_n539_), .B(new_new_n268_), .Y(new_new_n540_));
  NOi31      g0518(.An(new_new_n291_), .B(new_new_n302_), .C(new_new_n182_), .Y(new_new_n541_));
  NA3        g0519(.A(new_new_n307_), .B(new_new_n175_), .C(new_new_n100_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n220_), .B(new_new_n45_), .Y(new_new_n543_));
  NO2        g0521(.A(new_new_n157_), .B(i_5_), .Y(new_new_n544_));
  NA3        g0522(.A(new_new_n544_), .B(new_new_n411_), .C(new_new_n320_), .Y(new_new_n545_));
  OAI210     g0523(.A0(new_new_n545_), .A1(new_new_n543_), .B0(new_new_n542_), .Y(new_new_n546_));
  OAI210     g0524(.A0(new_new_n546_), .A1(new_new_n541_), .B0(new_new_n459_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n547_), .B(new_new_n540_), .C(new_new_n534_), .Y(new_new_n548_));
  NA3        g0526(.A(new_new_n216_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n283_), .B(new_new_n85_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n549_), .B(new_new_n550_), .Y(new_new_n551_));
  NA2        g0529(.A(new_new_n297_), .B(new_new_n287_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n552_), .B(new_new_n174_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n446_), .B(new_new_n220_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n554_), .B(new_new_n555_), .Y(new_new_n556_));
  AOI210     g0534(.A0(new_new_n367_), .A1(new_new_n47_), .B0(new_new_n371_), .Y(new_new_n557_));
  NA2        g0535(.A(i_0_), .B(new_new_n49_), .Y(new_new_n558_));
  NA3        g0536(.A(new_new_n529_), .B(new_new_n277_), .C(new_new_n558_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n557_), .B(new_new_n559_), .Y(new_new_n560_));
  NO4        g0538(.A(new_new_n560_), .B(new_new_n556_), .C(new_new_n553_), .D(new_new_n551_), .Y(new_new_n561_));
  NO4        g0539(.A(new_new_n251_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n562_));
  NO3        g0540(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n232_), .B(new_new_n36_), .Y(new_new_n564_));
  AN2        g0542(.A(new_new_n564_), .B(new_new_n563_), .Y(new_new_n565_));
  OA210      g0543(.A0(new_new_n565_), .A1(new_new_n562_), .B0(new_new_n359_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n418_), .B(i_1_), .Y(new_new_n567_));
  NOi31      g0545(.An(new_new_n567_), .B(new_new_n451_), .C(new_new_n74_), .Y(new_new_n568_));
  INV        g0546(.A(new_new_n566_), .Y(new_new_n569_));
  NOi21      g0547(.An(i_10_), .B(i_6_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n571_));
  AOI220     g0549(.A0(new_new_n283_), .A1(new_new_n571_), .B0(new_new_n277_), .B1(new_new_n570_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n572_), .B(new_new_n449_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n574_));
  INV        g0552(.A(new_new_n573_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n515_), .B(new_new_n382_), .Y(new_new_n576_));
  INV        g0554(.A(new_new_n320_), .Y(new_new_n577_));
  NO2        g0555(.A(i_12_), .B(new_new_n87_), .Y(new_new_n578_));
  NA3        g0556(.A(new_new_n578_), .B(new_new_n277_), .C(new_new_n558_), .Y(new_new_n579_));
  NA3        g0557(.A(new_new_n390_), .B(new_new_n283_), .C(new_new_n216_), .Y(new_new_n580_));
  AOI210     g0558(.A0(new_new_n580_), .A1(new_new_n579_), .B0(new_new_n577_), .Y(new_new_n581_));
  NA2        g0559(.A(new_new_n175_), .B(i_0_), .Y(new_new_n582_));
  NO3        g0560(.A(new_new_n582_), .B(new_new_n344_), .C(new_new_n302_), .Y(new_new_n583_));
  OR2        g0561(.A(i_2_), .B(i_5_), .Y(new_new_n584_));
  OR2        g0562(.A(new_new_n584_), .B(new_new_n414_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n585_), .B(new_new_n495_), .Y(new_new_n586_));
  NO4        g0564(.A(new_new_n586_), .B(new_new_n583_), .C(new_new_n581_), .D(new_new_n576_), .Y(new_new_n587_));
  NA4        g0565(.A(new_new_n587_), .B(new_new_n575_), .C(new_new_n569_), .D(new_new_n561_), .Y(new_new_n588_));
  NO4        g0566(.A(new_new_n588_), .B(new_new_n548_), .C(new_new_n526_), .D(new_new_n504_), .Y(new_new_n589_));
  NA4        g0567(.A(new_new_n589_), .B(new_new_n443_), .C(new_new_n358_), .D(new_new_n313_), .Y(mai7));
  NO2        g0568(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n112_), .B(new_new_n93_), .Y(new_new_n592_));
  NA2        g0570(.A(new_new_n388_), .B(new_new_n592_), .Y(new_new_n593_));
  NA2        g0571(.A(new_new_n484_), .B(new_new_n85_), .Y(new_new_n594_));
  NA2        g0572(.A(i_11_), .B(new_new_n192_), .Y(new_new_n595_));
  NA2        g0573(.A(new_new_n148_), .B(new_new_n595_), .Y(new_new_n596_));
  OAI210     g0574(.A0(new_new_n596_), .A1(new_new_n594_), .B0(new_new_n593_), .Y(new_new_n597_));
  NA3        g0575(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n236_), .B(i_4_), .Y(new_new_n599_));
  NA2        g0577(.A(new_new_n599_), .B(i_8_), .Y(new_new_n600_));
  NO2        g0578(.A(new_new_n109_), .B(new_new_n598_), .Y(new_new_n601_));
  NA2        g0579(.A(i_2_), .B(new_new_n87_), .Y(new_new_n602_));
  OAI210     g0580(.A0(new_new_n90_), .A1(new_new_n201_), .B0(new_new_n202_), .Y(new_new_n603_));
  NO2        g0581(.A(i_7_), .B(new_new_n37_), .Y(new_new_n604_));
  NA2        g0582(.A(i_4_), .B(i_8_), .Y(new_new_n605_));
  AOI210     g0583(.A0(new_new_n605_), .A1(new_new_n307_), .B0(new_new_n604_), .Y(new_new_n606_));
  OAI220     g0584(.A0(new_new_n606_), .A1(new_new_n602_), .B0(new_new_n603_), .B1(i_13_), .Y(new_new_n607_));
  NO4        g0585(.A(new_new_n607_), .B(new_new_n601_), .C(new_new_n597_), .D(new_new_n591_), .Y(new_new_n608_));
  AOI210     g0586(.A0(new_new_n132_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n609_));
  AOI210     g0587(.A0(new_new_n609_), .A1(new_new_n236_), .B0(new_new_n161_), .Y(new_new_n610_));
  OR2        g0588(.A(i_6_), .B(i_10_), .Y(new_new_n611_));
  NO2        g0589(.A(new_new_n611_), .B(new_new_n23_), .Y(new_new_n612_));
  OR3        g0590(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n613_));
  NO3        g0591(.A(new_new_n613_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n614_));
  INV        g0592(.A(new_new_n198_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n614_), .B(new_new_n612_), .Y(new_new_n616_));
  OA220      g0594(.A0(new_new_n616_), .A1(new_new_n577_), .B0(new_new_n610_), .B1(new_new_n270_), .Y(new_new_n617_));
  AOI210     g0595(.A0(new_new_n617_), .A1(new_new_n608_), .B0(new_new_n64_), .Y(new_new_n618_));
  NOi21      g0596(.An(i_11_), .B(i_7_), .Y(new_new_n619_));
  AO210      g0597(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n620_), .B(new_new_n619_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n621_), .B(new_new_n204_), .Y(new_new_n622_));
  NA3        g0600(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n623_));
  NAi31      g0601(.An(new_new_n623_), .B(new_new_n213_), .C(i_11_), .Y(new_new_n624_));
  AOI210     g0602(.A0(new_new_n624_), .A1(new_new_n622_), .B0(new_new_n64_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n626_));
  AO210      g0604(.A0(new_new_n626_), .A1(new_new_n382_), .B0(new_new_n41_), .Y(new_new_n627_));
  NO3        g0605(.A(new_new_n259_), .B(new_new_n206_), .C(new_new_n595_), .Y(new_new_n628_));
  OAI210     g0606(.A0(new_new_n628_), .A1(new_new_n225_), .B0(new_new_n64_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n415_), .B(new_new_n31_), .Y(new_new_n630_));
  OR2        g0608(.A(new_new_n206_), .B(new_new_n112_), .Y(new_new_n631_));
  NA2        g0609(.A(new_new_n631_), .B(new_new_n630_), .Y(new_new_n632_));
  NO2        g0610(.A(i_1_), .B(i_4_), .Y(new_new_n633_));
  NA2        g0611(.A(new_new_n633_), .B(new_new_n632_), .Y(new_new_n634_));
  NO2        g0612(.A(i_1_), .B(i_12_), .Y(new_new_n635_));
  NA3        g0613(.A(new_new_n635_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n636_));
  BUFFER     g0614(.A(new_new_n636_), .Y(new_new_n637_));
  NA4        g0615(.A(new_new_n637_), .B(new_new_n634_), .C(new_new_n629_), .D(new_new_n627_), .Y(new_new_n638_));
  OAI210     g0616(.A0(new_new_n638_), .A1(new_new_n625_), .B0(i_6_), .Y(new_new_n639_));
  NO2        g0617(.A(new_new_n623_), .B(new_new_n112_), .Y(new_new_n640_));
  NA2        g0618(.A(new_new_n640_), .B(new_new_n578_), .Y(new_new_n641_));
  NO2        g0619(.A(i_6_), .B(i_11_), .Y(new_new_n642_));
  NA2        g0620(.A(new_new_n641_), .B(new_new_n452_), .Y(new_new_n643_));
  NO3        g0621(.A(new_new_n611_), .B(new_new_n232_), .C(new_new_n23_), .Y(new_new_n644_));
  AOI210     g0622(.A0(i_1_), .A1(new_new_n260_), .B0(new_new_n644_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n645_), .B(new_new_n45_), .Y(new_new_n646_));
  NA3        g0624(.A(new_new_n535_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n647_));
  INV        g0625(.A(i_2_), .Y(new_new_n648_));
  NA2        g0626(.A(new_new_n142_), .B(i_9_), .Y(new_new_n649_));
  NA3        g0627(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n47_), .B(i_1_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n649_), .B(new_new_n648_), .Y(new_new_n652_));
  AOI210     g0630(.A0(new_new_n476_), .A1(new_new_n421_), .B0(new_new_n241_), .Y(new_new_n653_));
  NO2        g0631(.A(new_new_n653_), .B(new_new_n602_), .Y(new_new_n654_));
  NAi21      g0632(.An(new_new_n647_), .B(new_new_n95_), .Y(new_new_n655_));
  NO2        g0633(.A(i_11_), .B(new_new_n37_), .Y(new_new_n656_));
  INV        g0634(.A(new_new_n655_), .Y(new_new_n657_));
  OR3        g0635(.A(new_new_n657_), .B(new_new_n654_), .C(new_new_n652_), .Y(new_new_n658_));
  NO3        g0636(.A(new_new_n658_), .B(new_new_n646_), .C(new_new_n643_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n236_), .B(new_new_n105_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n660_), .B(new_new_n619_), .Y(new_new_n661_));
  NA2        g0639(.A(new_new_n661_), .B(i_1_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n662_), .B(new_new_n613_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n417_), .B(new_new_n87_), .Y(new_new_n664_));
  NA2        g0642(.A(new_new_n663_), .B(new_new_n47_), .Y(new_new_n665_));
  NA2        g0643(.A(i_3_), .B(new_new_n192_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n666_), .B(new_new_n118_), .Y(new_new_n667_));
  AN2        g0645(.A(new_new_n667_), .B(new_new_n537_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n232_), .B(new_new_n45_), .Y(new_new_n669_));
  NO3        g0647(.A(new_new_n669_), .B(new_new_n310_), .C(new_new_n237_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n121_), .B(new_new_n37_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n671_), .B(i_6_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n87_), .B(i_9_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n673_), .B(new_new_n64_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n635_), .Y(new_new_n675_));
  NO4        g0653(.A(new_new_n675_), .B(new_new_n672_), .C(new_new_n670_), .D(i_4_), .Y(new_new_n676_));
  NA2        g0654(.A(i_1_), .B(i_3_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n453_), .B(new_new_n96_), .Y(new_new_n678_));
  AOI210     g0656(.A0(new_new_n669_), .A1(new_new_n570_), .B0(new_new_n678_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n679_), .B(new_new_n677_), .Y(new_new_n680_));
  NO3        g0658(.A(new_new_n680_), .B(new_new_n676_), .C(new_new_n668_), .Y(new_new_n681_));
  NA4        g0659(.A(new_new_n681_), .B(new_new_n665_), .C(new_new_n659_), .D(new_new_n639_), .Y(new_new_n682_));
  NO3        g0660(.A(new_new_n478_), .B(i_3_), .C(i_7_), .Y(new_new_n683_));
  NOi21      g0661(.An(new_new_n683_), .B(i_10_), .Y(new_new_n684_));
  OA210      g0662(.A0(new_new_n684_), .A1(new_new_n244_), .B0(new_new_n87_), .Y(new_new_n685_));
  NA2        g0663(.A(new_new_n374_), .B(new_new_n373_), .Y(new_new_n686_));
  NA3        g0664(.A(new_new_n484_), .B(new_new_n518_), .C(new_new_n47_), .Y(new_new_n687_));
  NO3        g0665(.A(new_new_n479_), .B(new_new_n605_), .C(new_new_n87_), .Y(new_new_n688_));
  NA2        g0666(.A(new_new_n688_), .B(new_new_n25_), .Y(new_new_n689_));
  NA3        g0667(.A(new_new_n689_), .B(new_new_n687_), .C(new_new_n686_), .Y(new_new_n690_));
  OAI210     g0668(.A0(new_new_n690_), .A1(new_new_n685_), .B0(i_1_), .Y(new_new_n691_));
  AOI210     g0669(.A0(new_new_n269_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n372_), .B(i_2_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n693_), .B(new_new_n692_), .Y(new_new_n694_));
  AOI210     g0672(.A0(new_new_n694_), .A1(new_new_n691_), .B0(i_13_), .Y(new_new_n695_));
  OR2        g0673(.A(i_11_), .B(i_7_), .Y(new_new_n696_));
  AOI210     g0674(.A0(new_new_n650_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n697_));
  INV        g0675(.A(new_new_n697_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n479_), .B(new_new_n24_), .Y(new_new_n699_));
  AOI220     g0677(.A0(new_new_n699_), .A1(new_new_n664_), .B0(new_new_n244_), .B1(new_new_n135_), .Y(new_new_n700_));
  OAI220     g0678(.A0(new_new_n700_), .A1(new_new_n41_), .B0(new_new_n698_), .B1(new_new_n96_), .Y(new_new_n701_));
  INV        g0679(.A(new_new_n701_), .Y(new_new_n702_));
  NA2        g0680(.A(new_new_n390_), .B(new_new_n651_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n703_), .B(new_new_n242_), .Y(new_new_n704_));
  AOI210     g0682(.A0(new_new_n447_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n705_));
  NOi31      g0683(.An(new_new_n705_), .B(new_new_n594_), .C(new_new_n45_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n131_), .B(i_13_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n650_), .B(new_new_n118_), .Y(new_new_n708_));
  INV        g0686(.A(new_new_n708_), .Y(new_new_n709_));
  OAI220     g0687(.A0(new_new_n709_), .A1(new_new_n72_), .B0(new_new_n707_), .B1(new_new_n692_), .Y(new_new_n710_));
  NO3        g0688(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n105_), .Y(new_new_n711_));
  NA2        g0689(.A(new_new_n26_), .B(new_new_n192_), .Y(new_new_n712_));
  INV        g0690(.A(i_7_), .Y(new_new_n713_));
  INV        g0691(.A(new_new_n711_), .Y(new_new_n714_));
  AOI220     g0692(.A0(new_new_n390_), .A1(new_new_n651_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n715_));
  OAI220     g0693(.A0(new_new_n715_), .A1(new_new_n600_), .B0(new_new_n714_), .B1(new_new_n615_), .Y(new_new_n716_));
  NO4        g0694(.A(new_new_n716_), .B(new_new_n710_), .C(new_new_n706_), .D(new_new_n704_), .Y(new_new_n717_));
  OR2        g0695(.A(i_11_), .B(i_6_), .Y(new_new_n718_));
  NA3        g0696(.A(new_new_n599_), .B(new_new_n712_), .C(i_7_), .Y(new_new_n719_));
  AOI210     g0697(.A0(new_new_n719_), .A1(new_new_n709_), .B0(new_new_n718_), .Y(new_new_n720_));
  NA3        g0698(.A(new_new_n415_), .B(new_new_n604_), .C(new_new_n101_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n642_), .B(i_13_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n106_), .B(new_new_n712_), .Y(new_new_n723_));
  NAi21      g0701(.An(i_11_), .B(i_12_), .Y(new_new_n724_));
  NOi41      g0702(.An(new_new_n114_), .B(new_new_n724_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n725_));
  NO3        g0703(.A(new_new_n479_), .B(new_new_n578_), .C(new_new_n605_), .Y(new_new_n726_));
  AOI220     g0704(.A0(new_new_n726_), .A1(new_new_n314_), .B0(new_new_n725_), .B1(new_new_n723_), .Y(new_new_n727_));
  NA3        g0705(.A(new_new_n727_), .B(new_new_n722_), .C(new_new_n721_), .Y(new_new_n728_));
  OAI210     g0706(.A0(new_new_n728_), .A1(new_new_n720_), .B0(new_new_n64_), .Y(new_new_n729_));
  NO2        g0707(.A(i_2_), .B(i_12_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n371_), .B(new_new_n730_), .Y(new_new_n731_));
  NA2        g0709(.A(new_new_n373_), .B(new_new_n371_), .Y(new_new_n732_));
  NO2        g0710(.A(new_new_n132_), .B(i_2_), .Y(new_new_n733_));
  NA2        g0711(.A(new_new_n733_), .B(new_new_n635_), .Y(new_new_n734_));
  NA3        g0712(.A(new_new_n734_), .B(new_new_n732_), .C(new_new_n731_), .Y(new_new_n735_));
  NA3        g0713(.A(new_new_n735_), .B(new_new_n46_), .C(new_new_n224_), .Y(new_new_n736_));
  NA4        g0714(.A(new_new_n736_), .B(new_new_n729_), .C(new_new_n717_), .D(new_new_n702_), .Y(new_new_n737_));
  OR4        g0715(.A(new_new_n737_), .B(new_new_n695_), .C(new_new_n682_), .D(new_new_n618_), .Y(mai5));
  NA2        g0716(.A(new_new_n661_), .B(new_new_n272_), .Y(new_new_n739_));
  AN2        g0717(.A(new_new_n24_), .B(i_10_), .Y(new_new_n740_));
  NA3        g0718(.A(new_new_n740_), .B(new_new_n730_), .C(new_new_n112_), .Y(new_new_n741_));
  NO2        g0719(.A(new_new_n600_), .B(i_11_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n90_), .B(new_new_n742_), .Y(new_new_n743_));
  NA3        g0721(.A(new_new_n743_), .B(new_new_n741_), .C(new_new_n739_), .Y(new_new_n744_));
  NO3        g0722(.A(i_11_), .B(new_new_n236_), .C(i_13_), .Y(new_new_n745_));
  NO2        g0723(.A(new_new_n128_), .B(new_new_n23_), .Y(new_new_n746_));
  NA2        g0724(.A(i_12_), .B(i_8_), .Y(new_new_n747_));
  OAI210     g0725(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n747_), .Y(new_new_n748_));
  INV        g0726(.A(new_new_n446_), .Y(new_new_n749_));
  AOI220     g0727(.A0(new_new_n320_), .A1(new_new_n574_), .B0(new_new_n748_), .B1(new_new_n746_), .Y(new_new_n750_));
  INV        g0728(.A(new_new_n750_), .Y(new_new_n751_));
  NO2        g0729(.A(new_new_n751_), .B(new_new_n744_), .Y(new_new_n752_));
  INV        g0730(.A(new_new_n172_), .Y(new_new_n753_));
  INV        g0731(.A(new_new_n244_), .Y(new_new_n754_));
  OAI210     g0732(.A0(new_new_n693_), .A1(new_new_n448_), .B0(new_new_n114_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n755_), .A1(new_new_n754_), .B0(new_new_n753_), .Y(new_new_n756_));
  NO2        g0734(.A(new_new_n453_), .B(new_new_n26_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n757_), .B(new_new_n421_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n758_), .B(i_2_), .Y(new_new_n759_));
  INV        g0737(.A(new_new_n759_), .Y(new_new_n760_));
  AOI210     g0738(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n418_), .Y(new_new_n761_));
  AOI210     g0739(.A0(new_new_n761_), .A1(new_new_n760_), .B0(new_new_n756_), .Y(new_new_n762_));
  NO2        g0740(.A(new_new_n189_), .B(new_new_n129_), .Y(new_new_n763_));
  OAI210     g0741(.A0(new_new_n763_), .A1(new_new_n746_), .B0(i_2_), .Y(new_new_n764_));
  INV        g0742(.A(new_new_n173_), .Y(new_new_n765_));
  NO3        g0743(.A(new_new_n620_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n766_));
  AOI210     g0744(.A0(new_new_n765_), .A1(new_new_n90_), .B0(new_new_n766_), .Y(new_new_n767_));
  AOI210     g0745(.A0(new_new_n767_), .A1(new_new_n764_), .B0(new_new_n192_), .Y(new_new_n768_));
  OA210      g0746(.A0(new_new_n621_), .A1(new_new_n130_), .B0(i_13_), .Y(new_new_n769_));
  NA2        g0747(.A(new_new_n198_), .B(new_new_n201_), .Y(new_new_n770_));
  NA2        g0748(.A(new_new_n155_), .B(new_new_n595_), .Y(new_new_n771_));
  AOI210     g0749(.A0(new_new_n771_), .A1(new_new_n770_), .B0(new_new_n376_), .Y(new_new_n772_));
  AOI210     g0750(.A0(new_new_n206_), .A1(new_new_n152_), .B0(new_new_n518_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n773_), .B(new_new_n421_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n775_));
  INV        g0753(.A(new_new_n303_), .Y(new_new_n776_));
  NA4        g0754(.A(new_new_n776_), .B(new_new_n307_), .C(new_new_n128_), .D(new_new_n43_), .Y(new_new_n777_));
  OAI210     g0755(.A0(new_new_n777_), .A1(new_new_n775_), .B0(new_new_n774_), .Y(new_new_n778_));
  NO4        g0756(.A(new_new_n778_), .B(new_new_n772_), .C(new_new_n769_), .D(new_new_n768_), .Y(new_new_n779_));
  NA2        g0757(.A(new_new_n574_), .B(new_new_n28_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n745_), .B(new_new_n278_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n781_), .B(new_new_n780_), .Y(new_new_n782_));
  NO2        g0760(.A(new_new_n63_), .B(i_12_), .Y(new_new_n783_));
  NO2        g0761(.A(new_new_n783_), .B(new_new_n130_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n784_), .B(new_new_n595_), .Y(new_new_n785_));
  AOI220     g0763(.A0(new_new_n785_), .A1(new_new_n36_), .B0(new_new_n782_), .B1(new_new_n47_), .Y(new_new_n786_));
  NA4        g0764(.A(new_new_n786_), .B(new_new_n779_), .C(new_new_n762_), .D(new_new_n752_), .Y(mai6));
  NO2        g0765(.A(new_new_n219_), .B(new_new_n486_), .Y(new_new_n788_));
  NO2        g0766(.A(i_11_), .B(i_9_), .Y(new_new_n789_));
  INV        g0767(.A(new_new_n331_), .Y(new_new_n790_));
  OR2        g0768(.A(new_new_n790_), .B(i_12_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n377_), .B(new_new_n338_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n578_), .B(new_new_n64_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n684_), .B(new_new_n72_), .Y(new_new_n794_));
  BUFFER     g0772(.A(new_new_n626_), .Y(new_new_n795_));
  NA4        g0773(.A(new_new_n795_), .B(new_new_n794_), .C(new_new_n793_), .D(new_new_n792_), .Y(new_new_n796_));
  INV        g0774(.A(new_new_n196_), .Y(new_new_n797_));
  AOI220     g0775(.A0(new_new_n797_), .A1(new_new_n789_), .B0(new_new_n796_), .B1(new_new_n74_), .Y(new_new_n798_));
  INV        g0776(.A(new_new_n330_), .Y(new_new_n799_));
  NA2        g0777(.A(new_new_n76_), .B(new_new_n135_), .Y(new_new_n800_));
  INV        g0778(.A(new_new_n128_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n801_), .B(new_new_n47_), .Y(new_new_n802_));
  AOI210     g0780(.A0(new_new_n802_), .A1(new_new_n800_), .B0(new_new_n799_), .Y(new_new_n803_));
  NO3        g0781(.A(new_new_n251_), .B(new_new_n136_), .C(i_9_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n804_), .B(new_new_n783_), .Y(new_new_n805_));
  AOI210     g0783(.A0(new_new_n805_), .A1(new_new_n516_), .B0(new_new_n184_), .Y(new_new_n806_));
  NO2        g0784(.A(new_new_n32_), .B(i_11_), .Y(new_new_n807_));
  NA3        g0785(.A(new_new_n807_), .B(new_new_n474_), .C(new_new_n394_), .Y(new_new_n808_));
  NAi32      g0786(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n809_));
  NO2        g0787(.A(new_new_n718_), .B(new_new_n809_), .Y(new_new_n810_));
  OAI210     g0788(.A0(new_new_n683_), .A1(new_new_n564_), .B0(new_new_n563_), .Y(new_new_n811_));
  NAi31      g0789(.An(new_new_n810_), .B(new_new_n811_), .C(new_new_n808_), .Y(new_new_n812_));
  OR3        g0790(.A(new_new_n812_), .B(new_new_n806_), .C(new_new_n803_), .Y(new_new_n813_));
  NO2        g0791(.A(new_new_n696_), .B(i_2_), .Y(new_new_n814_));
  NA2        g0792(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n815_));
  NO2        g0793(.A(new_new_n815_), .B(new_new_n414_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n816_), .B(new_new_n814_), .Y(new_new_n817_));
  BUFFER     g0795(.A(new_new_n621_), .Y(new_new_n818_));
  NA3        g0796(.A(new_new_n818_), .B(new_new_n151_), .C(new_new_n70_), .Y(new_new_n819_));
  AO210      g0797(.A0(new_new_n493_), .A1(new_new_n749_), .B0(new_new_n36_), .Y(new_new_n820_));
  NA3        g0798(.A(new_new_n820_), .B(new_new_n819_), .C(new_new_n817_), .Y(new_new_n821_));
  OAI210     g0799(.A0(i_6_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n822_));
  AOI220     g0800(.A0(new_new_n822_), .A1(new_new_n563_), .B0(new_new_n788_), .B1(new_new_n713_), .Y(new_new_n823_));
  NA3        g0801(.A(new_new_n376_), .B(new_new_n238_), .C(new_new_n151_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n402_), .B(new_new_n71_), .Y(new_new_n825_));
  NA4        g0803(.A(new_new_n825_), .B(new_new_n824_), .C(new_new_n823_), .D(new_new_n603_), .Y(new_new_n826_));
  AO210      g0804(.A0(new_new_n518_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n827_));
  NA3        g0805(.A(new_new_n827_), .B(new_new_n484_), .C(new_new_n216_), .Y(new_new_n828_));
  AOI210     g0806(.A0(new_new_n448_), .A1(new_new_n446_), .B0(new_new_n562_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n611_), .B(new_new_n106_), .Y(new_new_n830_));
  OAI210     g0808(.A0(new_new_n830_), .A1(new_new_n115_), .B0(new_new_n413_), .Y(new_new_n831_));
  NA2        g0809(.A(new_new_n243_), .B(new_new_n47_), .Y(new_new_n832_));
  INV        g0810(.A(new_new_n585_), .Y(new_new_n833_));
  NA3        g0811(.A(new_new_n833_), .B(new_new_n330_), .C(i_7_), .Y(new_new_n834_));
  NA4        g0812(.A(new_new_n834_), .B(new_new_n831_), .C(new_new_n829_), .D(new_new_n828_), .Y(new_new_n835_));
  NO4        g0813(.A(new_new_n835_), .B(new_new_n826_), .C(new_new_n821_), .D(new_new_n813_), .Y(new_new_n836_));
  NA4        g0814(.A(new_new_n836_), .B(new_new_n798_), .C(new_new_n791_), .D(new_new_n384_), .Y(mai3));
  NO2        g0815(.A(i_11_), .B(new_new_n236_), .Y(new_new_n838_));
  NA2        g0816(.A(new_new_n291_), .B(new_new_n838_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n839_), .B(new_new_n192_), .Y(new_new_n840_));
  NO3        g0818(.A(new_new_n449_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n841_));
  OA210      g0819(.A0(new_new_n841_), .A1(new_new_n840_), .B0(new_new_n175_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n824_), .B(new_new_n375_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n843_), .B(new_new_n40_), .Y(new_new_n844_));
  NOi21      g0822(.An(new_new_n100_), .B(new_new_n758_), .Y(new_new_n845_));
  NO3        g0823(.A(new_new_n631_), .B(new_new_n453_), .C(new_new_n135_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n415_), .B(new_new_n46_), .Y(new_new_n847_));
  AN2        g0825(.A(new_new_n451_), .B(new_new_n56_), .Y(new_new_n848_));
  NO3        g0826(.A(new_new_n848_), .B(new_new_n846_), .C(new_new_n845_), .Y(new_new_n849_));
  AOI210     g0827(.A0(new_new_n849_), .A1(new_new_n844_), .B0(new_new_n49_), .Y(new_new_n850_));
  NO4        g0828(.A(new_new_n380_), .B(new_new_n387_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n184_), .B(new_new_n570_), .Y(new_new_n852_));
  NOi21      g0830(.An(new_new_n852_), .B(new_new_n851_), .Y(new_new_n853_));
  NO2        g0831(.A(new_new_n853_), .B(new_new_n64_), .Y(new_new_n854_));
  NOi21      g0832(.An(i_5_), .B(i_9_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n855_), .B(new_new_n445_), .Y(new_new_n856_));
  BUFFER     g0834(.A(new_new_n269_), .Y(new_new_n857_));
  AOI210     g0835(.A0(new_new_n857_), .A1(new_new_n476_), .B0(new_new_n688_), .Y(new_new_n858_));
  NO3        g0836(.A(new_new_n416_), .B(new_new_n269_), .C(new_new_n74_), .Y(new_new_n859_));
  NO2        g0837(.A(new_new_n176_), .B(new_new_n152_), .Y(new_new_n860_));
  AOI210     g0838(.A0(new_new_n860_), .A1(new_new_n243_), .B0(new_new_n859_), .Y(new_new_n861_));
  OAI220     g0839(.A0(new_new_n861_), .A1(new_new_n182_), .B0(new_new_n858_), .B1(new_new_n856_), .Y(new_new_n862_));
  NO4        g0840(.A(new_new_n862_), .B(new_new_n854_), .C(new_new_n850_), .D(new_new_n842_), .Y(new_new_n863_));
  NA2        g0841(.A(new_new_n184_), .B(new_new_n24_), .Y(new_new_n864_));
  NO2        g0842(.A(new_new_n671_), .B(new_new_n592_), .Y(new_new_n865_));
  NO2        g0843(.A(new_new_n865_), .B(new_new_n864_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n314_), .B(new_new_n133_), .Y(new_new_n867_));
  NAi21      g0845(.An(new_new_n162_), .B(new_new_n437_), .Y(new_new_n868_));
  OAI220     g0846(.A0(new_new_n868_), .A1(new_new_n832_), .B0(new_new_n867_), .B1(new_new_n404_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n869_), .B(new_new_n866_), .Y(new_new_n870_));
  NO2        g0848(.A(new_new_n394_), .B(new_new_n295_), .Y(new_new_n871_));
  NA2        g0849(.A(new_new_n871_), .B(new_new_n708_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n571_), .B(i_0_), .Y(new_new_n873_));
  NO3        g0851(.A(new_new_n873_), .B(new_new_n389_), .C(new_new_n90_), .Y(new_new_n874_));
  NO4        g0852(.A(new_new_n584_), .B(new_new_n213_), .C(new_new_n418_), .D(new_new_n414_), .Y(new_new_n875_));
  AOI210     g0853(.A0(new_new_n875_), .A1(i_11_), .B0(new_new_n874_), .Y(new_new_n876_));
  INV        g0854(.A(new_new_n474_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n745_), .B(new_new_n331_), .Y(new_new_n878_));
  AOI210     g0856(.A0(new_new_n484_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n879_));
  NO2        g0857(.A(new_new_n879_), .B(new_new_n878_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n253_), .B(new_new_n156_), .Y(new_new_n881_));
  NA2        g0859(.A(i_0_), .B(i_10_), .Y(new_new_n882_));
  INV        g0860(.A(new_new_n536_), .Y(new_new_n883_));
  NO4        g0861(.A(new_new_n118_), .B(new_new_n59_), .C(new_new_n666_), .D(i_5_), .Y(new_new_n884_));
  AO220      g0862(.A0(new_new_n884_), .A1(new_new_n883_), .B0(new_new_n881_), .B1(i_6_), .Y(new_new_n885_));
  NO2        g0863(.A(new_new_n885_), .B(new_new_n880_), .Y(new_new_n886_));
  NA4        g0864(.A(new_new_n886_), .B(new_new_n876_), .C(new_new_n872_), .D(new_new_n870_), .Y(new_new_n887_));
  NO2        g0865(.A(new_new_n107_), .B(new_new_n37_), .Y(new_new_n888_));
  NA2        g0866(.A(i_11_), .B(i_9_), .Y(new_new_n889_));
  NO3        g0867(.A(i_12_), .B(new_new_n889_), .C(new_new_n602_), .Y(new_new_n890_));
  AN2        g0868(.A(new_new_n890_), .B(new_new_n888_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n49_), .B(i_7_), .Y(new_new_n892_));
  NA2        g0870(.A(new_new_n399_), .B(new_new_n180_), .Y(new_new_n893_));
  NA2        g0871(.A(new_new_n893_), .B(new_new_n160_), .Y(new_new_n894_));
  NO2        g0872(.A(new_new_n889_), .B(new_new_n74_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n176_), .B(i_0_), .Y(new_new_n896_));
  INV        g0874(.A(new_new_n896_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n474_), .B(new_new_n230_), .Y(new_new_n898_));
  AOI210     g0876(.A0(new_new_n374_), .A1(new_new_n42_), .B0(new_new_n412_), .Y(new_new_n899_));
  OAI220     g0877(.A0(new_new_n899_), .A1(new_new_n856_), .B0(new_new_n898_), .B1(new_new_n897_), .Y(new_new_n900_));
  NO3        g0878(.A(new_new_n900_), .B(new_new_n894_), .C(new_new_n891_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n656_), .B(new_new_n125_), .Y(new_new_n902_));
  NO2        g0880(.A(i_6_), .B(new_new_n902_), .Y(new_new_n903_));
  AOI210     g0881(.A0(new_new_n447_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n172_), .B(new_new_n107_), .Y(new_new_n905_));
  NOi32      g0883(.An(new_new_n904_), .Bn(new_new_n187_), .C(new_new_n905_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n604_), .B(new_new_n331_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n907_), .B(new_new_n847_), .Y(new_new_n908_));
  NO3        g0886(.A(new_new_n908_), .B(new_new_n906_), .C(new_new_n903_), .Y(new_new_n909_));
  NOi21      g0887(.An(i_7_), .B(i_5_), .Y(new_new_n910_));
  NOi31      g0888(.An(new_new_n910_), .B(i_0_), .C(new_new_n724_), .Y(new_new_n911_));
  NA3        g0889(.A(new_new_n911_), .B(new_new_n388_), .C(i_6_), .Y(new_new_n912_));
  OA210      g0890(.A0(new_new_n905_), .A1(new_new_n516_), .B0(new_new_n912_), .Y(new_new_n913_));
  NO3        g0891(.A(new_new_n407_), .B(new_new_n363_), .C(new_new_n361_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n263_), .B(new_new_n321_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n724_), .B(new_new_n258_), .Y(new_new_n916_));
  AOI210     g0894(.A0(new_new_n916_), .A1(new_new_n915_), .B0(new_new_n914_), .Y(new_new_n917_));
  NA4        g0895(.A(new_new_n917_), .B(new_new_n913_), .C(new_new_n909_), .D(new_new_n901_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n864_), .B(new_new_n239_), .Y(new_new_n919_));
  AN2        g0897(.A(new_new_n335_), .B(new_new_n331_), .Y(new_new_n920_));
  AN2        g0898(.A(new_new_n920_), .B(new_new_n860_), .Y(new_new_n921_));
  OAI210     g0899(.A0(new_new_n921_), .A1(new_new_n919_), .B0(i_10_), .Y(new_new_n922_));
  NA3        g0900(.A(new_new_n473_), .B(new_new_n415_), .C(new_new_n46_), .Y(new_new_n923_));
  OAI210     g0901(.A0(new_new_n868_), .A1(new_new_n877_), .B0(new_new_n923_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n256_), .B(new_new_n47_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n895_), .B(new_new_n307_), .Y(new_new_n926_));
  OAI210     g0904(.A0(new_new_n925_), .A1(new_new_n186_), .B0(new_new_n926_), .Y(new_new_n927_));
  AOI220     g0905(.A0(new_new_n927_), .A1(new_new_n474_), .B0(new_new_n924_), .B1(new_new_n74_), .Y(new_new_n928_));
  NA2        g0906(.A(new_new_n96_), .B(new_new_n45_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n76_), .B(new_new_n747_), .Y(new_new_n930_));
  AOI220     g0908(.A0(new_new_n930_), .A1(new_new_n929_), .B0(new_new_n175_), .B1(new_new_n592_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n931_), .B(new_new_n48_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n699_), .B(new_new_n544_), .Y(new_new_n933_));
  NAi21      g0911(.An(i_9_), .B(i_5_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n934_), .B(new_new_n407_), .Y(new_new_n935_));
  NO2        g0913(.A(new_new_n598_), .B(new_new_n109_), .Y(new_new_n936_));
  AOI220     g0914(.A0(new_new_n936_), .A1(i_0_), .B0(new_new_n935_), .B1(new_new_n621_), .Y(new_new_n937_));
  OAI220     g0915(.A0(new_new_n937_), .A1(new_new_n87_), .B0(new_new_n933_), .B1(new_new_n173_), .Y(new_new_n938_));
  NO3        g0916(.A(new_new_n938_), .B(new_new_n932_), .C(new_new_n521_), .Y(new_new_n939_));
  NA3        g0917(.A(new_new_n939_), .B(new_new_n928_), .C(new_new_n922_), .Y(new_new_n940_));
  NO3        g0918(.A(new_new_n940_), .B(new_new_n918_), .C(new_new_n887_), .Y(new_new_n941_));
  NO2        g0919(.A(i_0_), .B(new_new_n724_), .Y(new_new_n942_));
  NA2        g0920(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n943_));
  INV        g0921(.A(new_new_n943_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n945_));
  AO220      g0923(.A0(new_new_n945_), .A1(new_new_n944_), .B0(new_new_n942_), .B1(new_new_n175_), .Y(new_new_n946_));
  AOI210     g0924(.A0(new_new_n793_), .A1(new_new_n686_), .B0(new_new_n905_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n946_), .A1(new_new_n352_), .B0(new_new_n947_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n733_), .B(new_new_n150_), .Y(new_new_n949_));
  INV        g0927(.A(new_new_n949_), .Y(new_new_n950_));
  NA3        g0928(.A(new_new_n950_), .B(new_new_n673_), .C(new_new_n74_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n811_), .B(new_new_n407_), .Y(new_new_n952_));
  OAI210     g0930(.A0(new_new_n243_), .A1(i_9_), .B0(new_new_n229_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n953_), .A1(new_new_n873_), .B0(new_new_n156_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n954_), .B(new_new_n952_), .Y(new_new_n955_));
  NA3        g0933(.A(new_new_n955_), .B(new_new_n951_), .C(new_new_n948_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n920_), .B(new_new_n376_), .Y(new_new_n957_));
  AOI210     g0935(.A0(new_new_n302_), .A1(new_new_n162_), .B0(new_new_n957_), .Y(new_new_n958_));
  NA3        g0936(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n892_), .B(new_new_n487_), .Y(new_new_n960_));
  AOI210     g0938(.A0(new_new_n959_), .A1(new_new_n162_), .B0(new_new_n960_), .Y(new_new_n961_));
  NO2        g0939(.A(new_new_n961_), .B(new_new_n958_), .Y(new_new_n962_));
  NO3        g0940(.A(new_new_n882_), .B(new_new_n855_), .C(new_new_n189_), .Y(new_new_n963_));
  AOI220     g0941(.A0(new_new_n963_), .A1(i_11_), .B0(new_new_n568_), .B1(new_new_n76_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n207_), .B(new_new_n387_), .C(i_0_), .Y(new_new_n965_));
  OAI210     g0943(.A0(new_new_n965_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n966_));
  NA3        g0944(.A(new_new_n966_), .B(new_new_n964_), .C(new_new_n962_), .Y(new_new_n967_));
  INV        g0945(.A(new_new_n542_), .Y(new_new_n968_));
  NO3        g0946(.A(new_new_n847_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n492_), .B(new_new_n485_), .Y(new_new_n970_));
  NO3        g0948(.A(new_new_n970_), .B(new_new_n969_), .C(new_new_n968_), .Y(new_new_n971_));
  NA3        g0949(.A(new_new_n394_), .B(new_new_n172_), .C(new_new_n171_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n394_), .B(new_new_n337_), .C(new_new_n220_), .Y(new_new_n973_));
  INV        g0951(.A(new_new_n973_), .Y(new_new_n974_));
  NOi31      g0952(.An(new_new_n393_), .B(new_new_n943_), .C(new_new_n239_), .Y(new_new_n975_));
  NO3        g0953(.A(new_new_n889_), .B(new_new_n216_), .C(new_new_n189_), .Y(new_new_n976_));
  NO4        g0954(.A(new_new_n976_), .B(new_new_n975_), .C(new_new_n974_), .D(new_new_n1042_), .Y(new_new_n977_));
  NA2        g0955(.A(new_new_n977_), .B(new_new_n971_), .Y(new_new_n978_));
  INV        g0956(.A(new_new_n614_), .Y(new_new_n979_));
  NO3        g0957(.A(new_new_n979_), .B(new_new_n558_), .C(new_new_n350_), .Y(new_new_n980_));
  NO2        g0958(.A(new_new_n87_), .B(i_5_), .Y(new_new_n981_));
  NA3        g0959(.A(new_new_n838_), .B(new_new_n113_), .C(new_new_n128_), .Y(new_new_n982_));
  INV        g0960(.A(new_new_n982_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n983_), .A1(new_new_n981_), .B0(new_new_n980_), .Y(new_new_n984_));
  NA3        g0962(.A(new_new_n307_), .B(i_5_), .C(new_new_n192_), .Y(new_new_n985_));
  NAi31      g0963(.An(new_new_n241_), .B(new_new_n985_), .C(new_new_n242_), .Y(new_new_n986_));
  NO4        g0964(.A(new_new_n239_), .B(new_new_n207_), .C(i_0_), .D(i_12_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n987_), .B(new_new_n986_), .Y(new_new_n988_));
  AN2        g0966(.A(new_new_n882_), .B(new_new_n156_), .Y(new_new_n989_));
  NO4        g0967(.A(new_new_n989_), .B(i_12_), .C(new_new_n647_), .D(new_new_n135_), .Y(new_new_n990_));
  NA2        g0968(.A(new_new_n990_), .B(new_new_n216_), .Y(new_new_n991_));
  NA2        g0969(.A(new_new_n910_), .B(new_new_n471_), .Y(new_new_n992_));
  NA2        g0970(.A(new_new_n65_), .B(new_new_n105_), .Y(new_new_n993_));
  OAI220     g0971(.A0(new_new_n993_), .A1(new_new_n985_), .B0(new_new_n992_), .B1(new_new_n674_), .Y(new_new_n994_));
  NA2        g0972(.A(new_new_n994_), .B(new_new_n896_), .Y(new_new_n995_));
  NA4        g0973(.A(new_new_n995_), .B(new_new_n991_), .C(new_new_n988_), .D(new_new_n984_), .Y(new_new_n996_));
  NO4        g0974(.A(new_new_n996_), .B(new_new_n978_), .C(new_new_n967_), .D(new_new_n956_), .Y(new_new_n997_));
  OAI210     g0975(.A0(new_new_n814_), .A1(new_new_n807_), .B0(new_new_n37_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n998_), .B(new_new_n610_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n999_), .B(new_new_n204_), .Y(new_new_n1000_));
  AN2        g0978(.A(new_new_n696_), .B(new_new_n372_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n185_), .B(new_new_n187_), .Y(new_new_n1002_));
  AO210      g0980(.A0(new_new_n1001_), .A1(new_new_n33_), .B0(new_new_n1002_), .Y(new_new_n1003_));
  OAI210     g0981(.A0(new_new_n614_), .A1(new_new_n612_), .B0(new_new_n320_), .Y(new_new_n1004_));
  NAi31      g0982(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1005_));
  AOI210     g0983(.A0(new_new_n121_), .A1(new_new_n71_), .B0(new_new_n1005_), .Y(new_new_n1006_));
  NO2        g0984(.A(new_new_n1006_), .B(new_new_n644_), .Y(new_new_n1007_));
  NA3        g0985(.A(new_new_n1007_), .B(new_new_n1004_), .C(new_new_n1003_), .Y(new_new_n1008_));
  NO2        g0986(.A(new_new_n461_), .B(new_new_n269_), .Y(new_new_n1009_));
  NO4        g0987(.A(new_new_n232_), .B(new_new_n149_), .C(new_new_n677_), .D(new_new_n37_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n1010_), .B(new_new_n1009_), .C(new_new_n875_), .Y(new_new_n1011_));
  INV        g0989(.A(new_new_n1011_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1008_), .A1(new_new_n49_), .B0(new_new_n1012_), .Y(new_new_n1013_));
  AOI210     g0991(.A0(new_new_n1013_), .A1(new_new_n1000_), .B0(new_new_n74_), .Y(new_new_n1014_));
  NO2        g0992(.A(new_new_n565_), .B(new_new_n383_), .Y(new_new_n1015_));
  NO2        g0993(.A(new_new_n1015_), .B(new_new_n753_), .Y(new_new_n1016_));
  NA2        g0994(.A(new_new_n263_), .B(new_new_n58_), .Y(new_new_n1017_));
  AOI220     g0995(.A0(new_new_n1017_), .A1(new_new_n77_), .B0(new_new_n351_), .B1(new_new_n255_), .Y(new_new_n1018_));
  NO2        g0996(.A(new_new_n1018_), .B(new_new_n236_), .Y(new_new_n1019_));
  NA3        g0997(.A(new_new_n100_), .B(new_new_n309_), .C(new_new_n31_), .Y(new_new_n1020_));
  INV        g0998(.A(new_new_n1020_), .Y(new_new_n1021_));
  NO2        g0999(.A(new_new_n1021_), .B(new_new_n1019_), .Y(new_new_n1022_));
  OAI210     g1000(.A0(new_new_n271_), .A1(new_new_n158_), .B0(new_new_n90_), .Y(new_new_n1023_));
  NO2        g1001(.A(new_new_n1023_), .B(i_11_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n605_), .B(new_new_n213_), .Y(new_new_n1025_));
  OAI210     g1003(.A0(new_new_n1025_), .A1(new_new_n904_), .B0(new_new_n204_), .Y(new_new_n1026_));
  NA2        g1004(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1027_));
  NO2        g1005(.A(new_new_n1026_), .B(new_new_n1027_), .Y(new_new_n1028_));
  NO3        g1006(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1029_));
  OAI210     g1007(.A0(new_new_n915_), .A1(new_new_n309_), .B0(new_new_n1029_), .Y(new_new_n1030_));
  NO2        g1008(.A(new_new_n1030_), .B(new_new_n724_), .Y(new_new_n1031_));
  NO4        g1009(.A(new_new_n934_), .B(new_new_n478_), .C(new_new_n252_), .D(new_new_n251_), .Y(new_new_n1032_));
  NO2        g1010(.A(new_new_n1032_), .B(new_new_n562_), .Y(new_new_n1033_));
  INV        g1011(.A(new_new_n364_), .Y(new_new_n1034_));
  AOI210     g1012(.A0(new_new_n1034_), .A1(new_new_n1033_), .B0(new_new_n41_), .Y(new_new_n1035_));
  NO4        g1013(.A(new_new_n1035_), .B(new_new_n1031_), .C(new_new_n1028_), .D(new_new_n1024_), .Y(new_new_n1036_));
  OAI210     g1014(.A0(new_new_n1022_), .A1(i_4_), .B0(new_new_n1036_), .Y(new_new_n1037_));
  NO3        g1015(.A(new_new_n1037_), .B(new_new_n1016_), .C(new_new_n1014_), .Y(new_new_n1038_));
  NA4        g1016(.A(new_new_n1038_), .B(new_new_n997_), .C(new_new_n941_), .D(new_new_n863_), .Y(mai4));
  INV        g1017(.A(new_new_n972_), .Y(new_new_n1042_));
endmodule


