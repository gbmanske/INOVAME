//Benchmark atmr_9sym_175_0.125

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n146_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, ori00, mai00, men00;
  INV        o00(.A(i_3_), .Y(ori_ori_n11_));
  INV        o01(.A(i_6_), .Y(ori_ori_n12_));
  INV        o02(.A(i_5_), .Y(ori_ori_n13_));
  NOi21      o03(.An(i_1_), .B(i_3_), .Y(ori_ori_n14_));
  INV        o04(.A(i_2_), .Y(ori_ori_n15_));
  NOi21      o05(.An(i_6_), .B(i_8_), .Y(ori_ori_n16_));
  NOi21      o06(.An(i_5_), .B(i_6_), .Y(ori_ori_n17_));
  NOi21      o07(.An(i_0_), .B(i_4_), .Y(ori_ori_n18_));
  INV        o08(.A(i_1_), .Y(ori_ori_n19_));
  NOi21      o09(.An(i_3_), .B(i_0_), .Y(ori_ori_n20_));
  NOi21      o10(.An(i_2_), .B(i_1_), .Y(ori_ori_n21_));
  NOi21      o11(.An(i_1_), .B(i_4_), .Y(ori_ori_n22_));
  BUFFER     o12(.A(i_7_), .Y(ori_ori_n23_));
  INV        o13(.A(ori_ori_n23_), .Y(ori_ori_n24_));
  NOi21      o14(.An(i_8_), .B(i_7_), .Y(ori_ori_n25_));
  NO2        o15(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n26_));
  NA2        o16(.A(ori_ori_n26_), .B(ori_ori_n15_), .Y(ori_ori_n27_));
  INV        o17(.A(ori_ori_n27_), .Y(ori_ori_n28_));
  INV        o18(.A(i_7_), .Y(ori_ori_n29_));
  NO2        o19(.A(ori_ori_n29_), .B(i_6_), .Y(ori_ori_n30_));
  INV        o20(.A(i_2_), .Y(ori_ori_n31_));
  BUFFER     o21(.A(i_1_), .Y(ori_ori_n32_));
  NO2        o22(.A(ori_ori_n31_), .B(i_7_), .Y(ori_ori_n33_));
  OAI210     o23(.A0(ori_ori_n33_), .A1(ori_ori_n30_), .B0(ori_ori_n13_), .Y(ori_ori_n34_));
  NA2        o24(.A(ori_ori_n14_), .B(i_2_), .Y(ori_ori_n35_));
  NA2        o25(.A(ori_ori_n35_), .B(ori_ori_n34_), .Y(ori_ori_n36_));
  INV        o26(.A(i_6_), .Y(ori_ori_n37_));
  INV        o27(.A(i_8_), .Y(ori_ori_n38_));
  NA2        o28(.A(ori_ori_n38_), .B(ori_ori_n12_), .Y(ori_ori_n39_));
  NO2        o29(.A(ori_ori_n39_), .B(ori_ori_n11_), .Y(ori_ori_n40_));
  NA2        o30(.A(ori_ori_n40_), .B(ori_ori_n32_), .Y(ori_ori_n41_));
  AOI220     o31(.A0(ori_ori_n20_), .A1(ori_ori_n19_), .B0(ori_ori_n14_), .B1(ori_ori_n15_), .Y(ori_ori_n42_));
  INV        o32(.A(i_5_), .Y(ori_ori_n43_));
  NO2        o33(.A(ori_ori_n43_), .B(ori_ori_n42_), .Y(ori_ori_n44_));
  INV        o34(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  INV        o35(.A(i_0_), .Y(ori_ori_n46_));
  NA2        o36(.A(ori_ori_n45_), .B(ori_ori_n41_), .Y(ori_ori_n47_));
  NA2        o37(.A(ori_ori_n16_), .B(ori_ori_n18_), .Y(ori_ori_n48_));
  NA2        o38(.A(ori_ori_n22_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o39(.A(ori_ori_n22_), .B(ori_ori_n20_), .Y(ori_ori_n50_));
  NA2        o40(.A(ori_ori_n50_), .B(ori_ori_n49_), .Y(ori_ori_n51_));
  NO2        o41(.A(ori_ori_n51_), .B(ori_ori_n21_), .Y(ori_ori_n52_));
  INV        o42(.A(i_4_), .Y(ori_ori_n53_));
  AOI210     o43(.A0(ori_ori_n46_), .A1(ori_ori_n37_), .B0(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o44(.A(i_7_), .Y(ori_ori_n55_));
  AN2        o45(.A(ori_ori_n54_), .B(ori_ori_n55_), .Y(ori_ori_n56_));
  INV        o46(.A(ori_ori_n56_), .Y(ori_ori_n57_));
  NA2        o47(.A(ori_ori_n23_), .B(ori_ori_n19_), .Y(ori_ori_n58_));
  INV        o48(.A(ori_ori_n58_), .Y(ori_ori_n59_));
  NO2        o49(.A(ori_ori_n59_), .B(ori_ori_n25_), .Y(ori_ori_n60_));
  NA4        o50(.A(ori_ori_n60_), .B(ori_ori_n57_), .C(ori_ori_n52_), .D(ori_ori_n48_), .Y(ori_ori_n61_));
  OR4        o51(.A(ori_ori_n61_), .B(ori_ori_n47_), .C(ori_ori_n36_), .D(ori_ori_n28_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  INV        m005(.A(i_0_), .Y(mai_mai_n16_));
  NOi21      m006(.An(i_1_), .B(i_3_), .Y(mai_mai_n17_));
  INV        m007(.A(i_4_), .Y(mai_mai_n18_));
  NA2        m008(.A(i_0_), .B(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m009(.A(i_7_), .Y(mai_mai_n20_));
  NA3        m010(.A(i_6_), .B(i_5_), .C(mai_mai_n20_), .Y(mai_mai_n21_));
  NOi21      m011(.An(i_8_), .B(i_6_), .Y(mai_mai_n22_));
  NOi21      m012(.An(i_1_), .B(i_8_), .Y(mai_mai_n23_));
  AOI220     m013(.A0(mai_mai_n23_), .A1(i_2_), .B0(mai_mai_n22_), .B1(i_5_), .Y(mai_mai_n24_));
  AOI210     m014(.A0(mai_mai_n24_), .A1(mai_mai_n21_), .B0(mai_mai_n19_), .Y(mai_mai_n25_));
  NA2        m015(.A(mai_mai_n25_), .B(mai_mai_n11_), .Y(mai_mai_n26_));
  NA2        m016(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n27_));
  NA2        m017(.A(mai_mai_n16_), .B(i_5_), .Y(mai_mai_n28_));
  NO2        m018(.A(i_2_), .B(i_4_), .Y(mai_mai_n29_));
  NA3        m019(.A(mai_mai_n29_), .B(i_6_), .C(i_8_), .Y(mai_mai_n30_));
  AOI210     m020(.A0(mai_mai_n28_), .A1(mai_mai_n27_), .B0(mai_mai_n30_), .Y(mai_mai_n31_));
  INV        m021(.A(i_2_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_5_), .B(i_0_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_6_), .B(i_8_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_7_), .B(i_1_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_5_), .B(i_6_), .Y(mai_mai_n36_));
  NA2        m026(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n37_));
  NO3        m027(.A(mai_mai_n37_), .B(mai_mai_n32_), .C(i_4_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_0_), .B(i_4_), .Y(mai_mai_n39_));
  XO2        m029(.A(i_1_), .B(i_3_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_7_), .B(i_5_), .Y(mai_mai_n41_));
  AN3        m031(.A(mai_mai_n41_), .B(mai_mai_n40_), .C(mai_mai_n39_), .Y(mai_mai_n42_));
  INV        m032(.A(i_1_), .Y(mai_mai_n43_));
  NOi21      m033(.An(i_3_), .B(i_0_), .Y(mai_mai_n44_));
  NO3        m034(.A(mai_mai_n42_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_4_), .B(i_0_), .Y(mai_mai_n46_));
  NA2        m036(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n47_));
  NOi21      m037(.An(i_2_), .B(i_8_), .Y(mai_mai_n48_));
  NO3        m038(.A(mai_mai_n48_), .B(mai_mai_n46_), .C(mai_mai_n39_), .Y(mai_mai_n49_));
  NO3        m039(.A(mai_mai_n49_), .B(mai_mai_n47_), .C(mai_mai_n146_), .Y(mai_mai_n50_));
  INV        m040(.A(mai_mai_n50_), .Y(mai_mai_n51_));
  NOi31      m041(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n52_));
  NA2        m042(.A(mai_mai_n52_), .B(i_0_), .Y(mai_mai_n53_));
  NOi21      m043(.An(i_4_), .B(i_3_), .Y(mai_mai_n54_));
  NOi21      m044(.An(i_1_), .B(i_4_), .Y(mai_mai_n55_));
  OAI210     m045(.A0(mai_mai_n55_), .A1(mai_mai_n54_), .B0(mai_mai_n48_), .Y(mai_mai_n56_));
  NA2        m046(.A(mai_mai_n56_), .B(mai_mai_n53_), .Y(mai_mai_n57_));
  AN2        m047(.A(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  NA2        m048(.A(mai_mai_n58_), .B(mai_mai_n12_), .Y(mai_mai_n59_));
  NOi21      m049(.An(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  NA3        m050(.A(mai_mai_n60_), .B(mai_mai_n54_), .C(i_6_), .Y(mai_mai_n61_));
  OAI210     m051(.A0(mai_mai_n59_), .A1(mai_mai_n47_), .B0(mai_mai_n61_), .Y(mai_mai_n62_));
  AOI220     m052(.A0(mai_mai_n62_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .B1(mai_mai_n36_), .Y(mai_mai_n63_));
  NA4        m053(.A(mai_mai_n63_), .B(mai_mai_n51_), .C(mai_mai_n45_), .D(mai_mai_n26_), .Y(mai_mai_n64_));
  NA2        m054(.A(i_8_), .B(i_7_), .Y(mai_mai_n65_));
  NO3        m055(.A(mai_mai_n65_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n66_));
  NA2        m056(.A(i_8_), .B(mai_mai_n20_), .Y(mai_mai_n67_));
  AOI220     m057(.A0(mai_mai_n44_), .A1(i_1_), .B0(mai_mai_n40_), .B1(i_2_), .Y(mai_mai_n68_));
  NOi21      m058(.An(i_1_), .B(i_2_), .Y(mai_mai_n69_));
  NO2        m059(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n70_));
  OAI210     m060(.A0(mai_mai_n70_), .A1(mai_mai_n66_), .B0(mai_mai_n14_), .Y(mai_mai_n71_));
  NA3        m061(.A(mai_mai_n60_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n72_));
  NA3        m062(.A(mai_mai_n23_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NOi32      m064(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n75_));
  NA2        m065(.A(mai_mai_n75_), .B(i_3_), .Y(mai_mai_n76_));
  NA3        m066(.A(mai_mai_n17_), .B(i_2_), .C(i_6_), .Y(mai_mai_n77_));
  NA2        m067(.A(mai_mai_n77_), .B(mai_mai_n76_), .Y(mai_mai_n78_));
  NO2        m068(.A(i_0_), .B(i_4_), .Y(mai_mai_n79_));
  AOI220     m069(.A0(mai_mai_n79_), .A1(mai_mai_n78_), .B0(mai_mai_n74_), .B1(mai_mai_n54_), .Y(mai_mai_n80_));
  NA2        m070(.A(mai_mai_n80_), .B(mai_mai_n71_), .Y(mai_mai_n81_));
  NAi21      m071(.An(i_3_), .B(i_6_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n83_));
  NOi21      m073(.An(i_7_), .B(i_8_), .Y(mai_mai_n84_));
  NA3        m074(.A(mai_mai_n60_), .B(mai_mai_n32_), .C(i_3_), .Y(mai_mai_n85_));
  NA2        m075(.A(mai_mai_n43_), .B(i_6_), .Y(mai_mai_n86_));
  AOI210     m076(.A0(mai_mai_n86_), .A1(mai_mai_n19_), .B0(mai_mai_n85_), .Y(mai_mai_n87_));
  NAi21      m077(.An(i_6_), .B(i_0_), .Y(mai_mai_n88_));
  NOi21      m078(.An(i_4_), .B(i_6_), .Y(mai_mai_n89_));
  NOi21      m079(.An(i_5_), .B(i_3_), .Y(mai_mai_n90_));
  NA3        m080(.A(mai_mai_n90_), .B(mai_mai_n69_), .C(mai_mai_n89_), .Y(mai_mai_n91_));
  INV        m081(.A(mai_mai_n91_), .Y(mai_mai_n92_));
  NA2        m082(.A(mai_mai_n69_), .B(mai_mai_n34_), .Y(mai_mai_n93_));
  NOi21      m083(.An(mai_mai_n41_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  NO3        m084(.A(mai_mai_n94_), .B(mai_mai_n92_), .C(mai_mai_n87_), .Y(mai_mai_n95_));
  AOI220     m085(.A0(i_6_), .A1(i_7_), .B0(mai_mai_n22_), .B1(i_5_), .Y(mai_mai_n96_));
  NOi31      m086(.An(mai_mai_n46_), .B(mai_mai_n96_), .C(i_2_), .Y(mai_mai_n97_));
  NA2        m087(.A(mai_mai_n60_), .B(mai_mai_n12_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n34_), .B(mai_mai_n14_), .Y(mai_mai_n99_));
  NOi21      m089(.An(i_3_), .B(i_1_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n100_), .B(i_4_), .Y(mai_mai_n101_));
  AOI210     m091(.A0(mai_mai_n99_), .A1(mai_mai_n98_), .B0(mai_mai_n101_), .Y(mai_mai_n102_));
  AOI220     m092(.A0(mai_mai_n84_), .A1(mai_mai_n14_), .B0(mai_mai_n89_), .B1(mai_mai_n20_), .Y(mai_mai_n103_));
  NOi31      m093(.An(mai_mai_n44_), .B(mai_mai_n103_), .C(mai_mai_n32_), .Y(mai_mai_n104_));
  NO3        m094(.A(mai_mai_n104_), .B(mai_mai_n102_), .C(mai_mai_n97_), .Y(mai_mai_n105_));
  NA3        m095(.A(mai_mai_n105_), .B(mai_mai_n95_), .C(mai_mai_n83_), .Y(mai_mai_n106_));
  NA2        m096(.A(mai_mai_n48_), .B(mai_mai_n15_), .Y(mai_mai_n107_));
  NOi31      m097(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n108_));
  NOi31      m098(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n109_));
  OAI210     m099(.A0(mai_mai_n109_), .A1(mai_mai_n108_), .B0(i_7_), .Y(mai_mai_n110_));
  NA3        m100(.A(mai_mai_n110_), .B(mai_mai_n107_), .C(mai_mai_n93_), .Y(mai_mai_n111_));
  NA2        m101(.A(mai_mai_n111_), .B(mai_mai_n39_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n54_), .B(mai_mai_n35_), .Y(mai_mai_n113_));
  AOI210     m103(.A0(mai_mai_n113_), .A1(mai_mai_n72_), .B0(mai_mai_n28_), .Y(mai_mai_n114_));
  NA3        m104(.A(mai_mai_n60_), .B(mai_mai_n52_), .C(i_6_), .Y(mai_mai_n115_));
  INV        m105(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NOi21      m106(.An(i_0_), .B(i_2_), .Y(mai_mai_n117_));
  NA3        m107(.A(mai_mai_n117_), .B(mai_mai_n35_), .C(mai_mai_n89_), .Y(mai_mai_n118_));
  NA3        m108(.A(mai_mai_n46_), .B(mai_mai_n41_), .C(mai_mai_n17_), .Y(mai_mai_n119_));
  NA3        m109(.A(mai_mai_n117_), .B(mai_mai_n54_), .C(mai_mai_n34_), .Y(mai_mai_n120_));
  NA3        m110(.A(mai_mai_n120_), .B(mai_mai_n119_), .C(mai_mai_n118_), .Y(mai_mai_n121_));
  NA4        m111(.A(mai_mai_n52_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n122_));
  NA4        m112(.A(mai_mai_n55_), .B(mai_mai_n36_), .C(mai_mai_n16_), .D(i_8_), .Y(mai_mai_n123_));
  NA2        m113(.A(mai_mai_n123_), .B(mai_mai_n122_), .Y(mai_mai_n124_));
  NO4        m114(.A(mai_mai_n124_), .B(mai_mai_n121_), .C(mai_mai_n116_), .D(mai_mai_n114_), .Y(mai_mai_n125_));
  NA2        m115(.A(mai_mai_n58_), .B(mai_mai_n29_), .Y(mai_mai_n126_));
  AOI210     m116(.A0(mai_mai_n126_), .A1(mai_mai_n107_), .B0(mai_mai_n86_), .Y(mai_mai_n127_));
  NO4        m117(.A(i_2_), .B(mai_mai_n18_), .C(mai_mai_n11_), .D(mai_mai_n14_), .Y(mai_mai_n128_));
  NA2        m118(.A(i_2_), .B(i_4_), .Y(mai_mai_n129_));
  AOI210     m119(.A0(mai_mai_n88_), .A1(mai_mai_n82_), .B0(mai_mai_n129_), .Y(mai_mai_n130_));
  NO2        m120(.A(i_8_), .B(i_7_), .Y(mai_mai_n131_));
  OA210      m121(.A0(mai_mai_n130_), .A1(mai_mai_n128_), .B0(mai_mai_n131_), .Y(mai_mai_n132_));
  NA4        m122(.A(mai_mai_n100_), .B(i_0_), .C(i_5_), .D(mai_mai_n20_), .Y(mai_mai_n133_));
  NO2        m123(.A(mai_mai_n133_), .B(i_4_), .Y(mai_mai_n134_));
  NO3        m124(.A(mai_mai_n134_), .B(mai_mai_n132_), .C(mai_mai_n127_), .Y(mai_mai_n135_));
  NA2        m125(.A(mai_mai_n84_), .B(mai_mai_n12_), .Y(mai_mai_n136_));
  NA2        m126(.A(mai_mai_n46_), .B(i_3_), .Y(mai_mai_n137_));
  NO2        m127(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n138_));
  NA3        m128(.A(mai_mai_n117_), .B(mai_mai_n60_), .C(mai_mai_n89_), .Y(mai_mai_n139_));
  OAI210     m129(.A0(mai_mai_n85_), .A1(mai_mai_n28_), .B0(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m130(.A(mai_mai_n140_), .B(mai_mai_n138_), .Y(mai_mai_n141_));
  NA4        m131(.A(mai_mai_n141_), .B(mai_mai_n135_), .C(mai_mai_n125_), .D(mai_mai_n112_), .Y(mai_mai_n142_));
  OR4        m132(.A(mai_mai_n142_), .B(mai_mai_n106_), .C(mai_mai_n81_), .D(mai_mai_n64_), .Y(mai00));
  INV        m133(.A(i_3_), .Y(mai_mai_n146_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NA3        u013(.A(i_6_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n24_));
  NOi21      u014(.An(i_8_), .B(i_6_), .Y(men_men_n25_));
  NO2        u015(.A(men_men_n24_), .B(men_men_n22_), .Y(men_men_n26_));
  AOI210     u016(.A0(men_men_n26_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n27_));
  NA2        u017(.A(i_0_), .B(men_men_n14_), .Y(men_men_n28_));
  NA2        u018(.A(men_men_n17_), .B(i_5_), .Y(men_men_n29_));
  INV        u019(.A(i_2_), .Y(men_men_n30_));
  NOi21      u020(.An(i_5_), .B(i_0_), .Y(men_men_n31_));
  NOi21      u021(.An(i_6_), .B(i_8_), .Y(men_men_n32_));
  NOi21      u022(.An(i_5_), .B(i_6_), .Y(men_men_n33_));
  NOi21      u023(.An(i_0_), .B(i_4_), .Y(men_men_n34_));
  XO2        u024(.A(i_1_), .B(i_3_), .Y(men_men_n35_));
  INV        u025(.A(i_1_), .Y(men_men_n36_));
  NOi21      u026(.An(i_3_), .B(i_0_), .Y(men_men_n37_));
  NA2        u027(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NA3        u028(.A(i_6_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n39_));
  AOI210     u029(.A0(men_men_n39_), .A1(men_men_n24_), .B0(men_men_n38_), .Y(men_men_n40_));
  INV        u030(.A(men_men_n40_), .Y(men_men_n41_));
  NA2        u031(.A(i_1_), .B(men_men_n11_), .Y(men_men_n42_));
  NO3        u032(.A(men_men_n42_), .B(men_men_n28_), .C(i_2_), .Y(men_men_n43_));
  NOi21      u033(.An(i_4_), .B(i_0_), .Y(men_men_n44_));
  AOI210     u034(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n15_), .Y(men_men_n45_));
  NA2        u035(.A(i_1_), .B(men_men_n14_), .Y(men_men_n46_));
  NOi21      u036(.An(i_2_), .B(i_8_), .Y(men_men_n47_));
  NO2        u037(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NO3        u038(.A(men_men_n48_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n49_));
  NO2        u039(.A(men_men_n49_), .B(men_men_n43_), .Y(men_men_n50_));
  NOi31      u040(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n51_));
  NA2        u041(.A(men_men_n51_), .B(i_0_), .Y(men_men_n52_));
  NOi21      u042(.An(i_4_), .B(i_3_), .Y(men_men_n53_));
  NOi21      u043(.An(i_1_), .B(i_4_), .Y(men_men_n54_));
  OAI210     u044(.A0(men_men_n54_), .A1(men_men_n53_), .B0(men_men_n47_), .Y(men_men_n55_));
  NA2        u045(.A(men_men_n55_), .B(men_men_n52_), .Y(men_men_n56_));
  AN2        u046(.A(i_8_), .B(i_7_), .Y(men_men_n57_));
  NOi21      u047(.An(i_8_), .B(i_7_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n56_), .B(men_men_n33_), .Y(men_men_n59_));
  NA4        u049(.A(men_men_n59_), .B(men_men_n50_), .C(men_men_n41_), .D(men_men_n27_), .Y(men_men_n60_));
  NA2        u050(.A(i_8_), .B(i_7_), .Y(men_men_n61_));
  NO3        u051(.A(men_men_n61_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n62_));
  NA2        u052(.A(i_8_), .B(men_men_n23_), .Y(men_men_n63_));
  AOI220     u053(.A0(men_men_n37_), .A1(i_1_), .B0(men_men_n35_), .B1(i_2_), .Y(men_men_n64_));
  NOi21      u054(.An(i_1_), .B(i_2_), .Y(men_men_n65_));
  NA3        u055(.A(men_men_n65_), .B(men_men_n44_), .C(i_6_), .Y(men_men_n66_));
  OAI210     u056(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n66_), .Y(men_men_n67_));
  OAI210     u057(.A0(men_men_n67_), .A1(men_men_n62_), .B0(men_men_n14_), .Y(men_men_n68_));
  NA3        u058(.A(men_men_n58_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n69_));
  INV        u059(.A(men_men_n69_), .Y(men_men_n70_));
  NOi32      u060(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n71_));
  NA2        u061(.A(men_men_n71_), .B(i_3_), .Y(men_men_n72_));
  NA3        u062(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n73_));
  NA2        u063(.A(men_men_n73_), .B(men_men_n72_), .Y(men_men_n74_));
  NO2        u064(.A(i_0_), .B(i_4_), .Y(men_men_n75_));
  AOI220     u065(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n70_), .B1(men_men_n53_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n76_), .B(men_men_n68_), .Y(men_men_n77_));
  NAi21      u067(.An(i_3_), .B(i_6_), .Y(men_men_n78_));
  NO2        u068(.A(men_men_n78_), .B(i_0_), .Y(men_men_n79_));
  NA2        u069(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n80_));
  NOi21      u070(.An(i_7_), .B(i_8_), .Y(men_men_n81_));
  NOi31      u071(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n82_));
  AOI210     u072(.A0(men_men_n81_), .A1(men_men_n12_), .B0(men_men_n82_), .Y(men_men_n83_));
  OAI210     u073(.A0(men_men_n83_), .A1(men_men_n11_), .B0(men_men_n80_), .Y(men_men_n84_));
  OAI210     u074(.A0(men_men_n84_), .A1(men_men_n79_), .B0(men_men_n65_), .Y(men_men_n85_));
  NA3        u075(.A(men_men_n25_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n86_));
  AOI210     u076(.A0(men_men_n22_), .A1(men_men_n42_), .B0(men_men_n86_), .Y(men_men_n87_));
  AOI220     u077(.A0(men_men_n37_), .A1(men_men_n36_), .B0(men_men_n18_), .B1(men_men_n30_), .Y(men_men_n88_));
  NA3        u078(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n89_));
  OAI210     u079(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n90_));
  NA3        u080(.A(men_men_n61_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n91_));
  OAI220     u081(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n89_), .B1(men_men_n88_), .Y(men_men_n92_));
  NO2        u082(.A(men_men_n92_), .B(men_men_n87_), .Y(men_men_n93_));
  NA3        u083(.A(men_men_n58_), .B(men_men_n30_), .C(i_3_), .Y(men_men_n94_));
  NA2        u084(.A(men_men_n36_), .B(i_6_), .Y(men_men_n95_));
  AOI210     u085(.A0(men_men_n95_), .A1(men_men_n22_), .B0(men_men_n94_), .Y(men_men_n96_));
  NOi21      u086(.An(i_2_), .B(i_1_), .Y(men_men_n97_));
  AN3        u087(.A(men_men_n81_), .B(men_men_n97_), .C(men_men_n44_), .Y(men_men_n98_));
  NAi21      u088(.An(i_6_), .B(i_0_), .Y(men_men_n99_));
  NA3        u089(.A(men_men_n54_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n100_));
  NOi21      u090(.An(i_5_), .B(i_3_), .Y(men_men_n101_));
  NO2        u091(.A(men_men_n100_), .B(men_men_n99_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n65_), .B(men_men_n32_), .Y(men_men_n103_));
  NO3        u093(.A(men_men_n102_), .B(men_men_n98_), .C(men_men_n96_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n25_), .B(i_5_), .Y(men_men_n105_));
  NOi31      u095(.An(men_men_n44_), .B(men_men_n105_), .C(i_2_), .Y(men_men_n106_));
  NOi21      u096(.An(i_3_), .B(i_1_), .Y(men_men_n107_));
  NA2        u097(.A(men_men_n81_), .B(men_men_n14_), .Y(men_men_n108_));
  NOi31      u098(.An(men_men_n37_), .B(men_men_n108_), .C(men_men_n30_), .Y(men_men_n109_));
  NO2        u099(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n110_));
  NA4        u100(.A(men_men_n110_), .B(men_men_n104_), .C(men_men_n93_), .D(men_men_n85_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n47_), .B(men_men_n15_), .Y(men_men_n112_));
  NOi31      u102(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n113_));
  NOi31      u103(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n114_));
  OAI210     u104(.A0(men_men_n114_), .A1(men_men_n113_), .B0(i_7_), .Y(men_men_n115_));
  NA3        u105(.A(men_men_n32_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n116_));
  NA4        u106(.A(men_men_n116_), .B(men_men_n115_), .C(men_men_n112_), .D(men_men_n103_), .Y(men_men_n117_));
  NA2        u107(.A(men_men_n117_), .B(men_men_n34_), .Y(men_men_n118_));
  NO2        u108(.A(men_men_n69_), .B(men_men_n29_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n57_), .B(men_men_n97_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n120_));
  NAi31      u110(.An(men_men_n99_), .B(men_men_n81_), .C(men_men_n97_), .Y(men_men_n121_));
  NA3        u111(.A(men_men_n58_), .B(men_men_n51_), .C(i_6_), .Y(men_men_n122_));
  NA3        u112(.A(men_men_n122_), .B(men_men_n121_), .C(men_men_n120_), .Y(men_men_n123_));
  NOi32      u113(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n124_));
  NA2        u114(.A(men_men_n124_), .B(men_men_n113_), .Y(men_men_n125_));
  INV        u115(.A(men_men_n125_), .Y(men_men_n126_));
  NA4        u116(.A(men_men_n51_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n54_), .B(men_men_n33_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n128_));
  NA4        u118(.A(men_men_n54_), .B(men_men_n37_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n129_));
  NA3        u119(.A(men_men_n129_), .B(men_men_n128_), .C(men_men_n127_), .Y(men_men_n130_));
  NO4        u120(.A(men_men_n130_), .B(men_men_n126_), .C(men_men_n123_), .D(men_men_n119_), .Y(men_men_n131_));
  NOi21      u121(.An(i_5_), .B(i_2_), .Y(men_men_n132_));
  NA2        u122(.A(men_men_n132_), .B(men_men_n81_), .Y(men_men_n133_));
  AOI210     u123(.A0(men_men_n133_), .A1(men_men_n112_), .B0(men_men_n95_), .Y(men_men_n134_));
  NO4        u124(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n135_));
  NA2        u125(.A(i_2_), .B(i_4_), .Y(men_men_n136_));
  AOI210     u126(.A0(men_men_n99_), .A1(men_men_n78_), .B0(men_men_n136_), .Y(men_men_n137_));
  NO2        u127(.A(i_8_), .B(i_7_), .Y(men_men_n138_));
  OA210      u128(.A0(men_men_n137_), .A1(men_men_n135_), .B0(men_men_n138_), .Y(men_men_n139_));
  NA4        u129(.A(men_men_n107_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n140_));
  NO2        u130(.A(men_men_n140_), .B(i_4_), .Y(men_men_n141_));
  NO3        u131(.A(men_men_n141_), .B(men_men_n139_), .C(men_men_n134_), .Y(men_men_n142_));
  NA2        u132(.A(men_men_n81_), .B(men_men_n12_), .Y(men_men_n143_));
  NA3        u133(.A(i_2_), .B(i_1_), .C(men_men_n14_), .Y(men_men_n144_));
  NA2        u134(.A(men_men_n44_), .B(i_3_), .Y(men_men_n145_));
  AOI210     u135(.A0(men_men_n145_), .A1(men_men_n144_), .B0(men_men_n143_), .Y(men_men_n146_));
  NA4        u136(.A(men_men_n101_), .B(men_men_n57_), .C(men_men_n36_), .D(men_men_n21_), .Y(men_men_n147_));
  NA3        u137(.A(men_men_n82_), .B(men_men_n107_), .C(i_0_), .Y(men_men_n148_));
  NA3        u138(.A(men_men_n47_), .B(men_men_n31_), .C(men_men_n15_), .Y(men_men_n149_));
  NOi31      u139(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n150_));
  OAI210     u140(.A0(men_men_n124_), .A1(men_men_n71_), .B0(men_men_n150_), .Y(men_men_n151_));
  NA4        u141(.A(men_men_n151_), .B(men_men_n149_), .C(men_men_n148_), .D(men_men_n147_), .Y(men_men_n152_));
  NO2        u142(.A(men_men_n152_), .B(men_men_n146_), .Y(men_men_n153_));
  NA4        u143(.A(men_men_n153_), .B(men_men_n142_), .C(men_men_n131_), .D(men_men_n118_), .Y(men_men_n154_));
  OR4        u144(.A(men_men_n154_), .B(men_men_n111_), .C(men_men_n77_), .D(men_men_n60_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule