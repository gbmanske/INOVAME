// Benchmark "top" written by ABC on Thu Jun 20 14:59:10 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n127_,
    new_new_n128_, new_new_n129_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n945_, new_new_n946_, new_new_n947_,
    new_new_n948_, new_new_n949_, new_new_n950_, new_new_n951_,
    new_new_n952_, new_new_n953_, new_new_n954_, new_new_n955_,
    new_new_n956_, new_new_n957_, new_new_n958_, new_new_n959_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NO2        g028(.A(new_new_n47_), .B(new_new_n46_), .Y(new_new_n51_));
  NA2        g029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NO2        g031(.A(new_new_n53_), .B(new_new_n52_), .Y(new_new_n54_));
  OAI210     g032(.A0(new_new_n54_), .A1(new_new_n51_), .B0(new_new_n45_), .Y(new_new_n55_));
  NA3        g033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  OAI210     g036(.A0(new_new_n58_), .A1(new_new_n57_), .B0(new_new_n56_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  INV        g041(.A(new_new_n60_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n50_), .B(i_2_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_6_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(new_new_n25_), .Y(new_new_n67_));
  INV        g045(.A(i_0_), .Y(new_new_n68_));
  NAi21      g046(.An(i_5_), .B(i_10_), .Y(new_new_n69_));
  NA2        g047(.A(i_5_), .B(i_9_), .Y(new_new_n70_));
  AOI210     g048(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n68_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n67_), .Y(new_new_n72_));
  INV        g050(.A(new_new_n72_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n73_), .A1(new_new_n64_), .B0(i_0_), .Y(new_new_n74_));
  NA2        g052(.A(i_12_), .B(i_5_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_9_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_7_), .Y(new_new_n77_));
  INV        g055(.A(i_6_), .Y(new_new_n78_));
  OR4        g056(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n79_));
  INV        g057(.A(new_new_n79_), .Y(new_new_n80_));
  NO2        g058(.A(i_2_), .B(i_7_), .Y(new_new_n81_));
  NAi21      g059(.An(i_6_), .B(i_10_), .Y(new_new_n82_));
  NA2        g060(.A(i_6_), .B(i_9_), .Y(new_new_n83_));
  AOI210     g061(.A0(new_new_n83_), .A1(new_new_n82_), .B0(new_new_n62_), .Y(new_new_n84_));
  NA2        g062(.A(i_2_), .B(i_6_), .Y(new_new_n85_));
  INV        g063(.A(new_new_n84_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n86_), .B(new_new_n75_), .Y(new_new_n87_));
  AN3        g065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_11_), .Y(new_new_n89_));
  NO2        g067(.A(i_5_), .B(i_8_), .Y(new_new_n90_));
  NOi21      g068(.An(new_new_n90_), .B(new_new_n89_), .Y(new_new_n91_));
  AOI220     g069(.A0(new_new_n91_), .A1(new_new_n61_), .B0(new_new_n88_), .B1(new_new_n32_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n46_), .B(new_new_n93_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n78_), .Y(new_new_n96_));
  NA2        g074(.A(i_12_), .B(i_3_), .Y(new_new_n97_));
  INV        g075(.A(new_new_n97_), .Y(new_new_n98_));
  NA3        g076(.A(new_new_n98_), .B(new_new_n96_), .C(new_new_n94_), .Y(new_new_n99_));
  NAi21      g077(.An(i_7_), .B(i_11_), .Y(new_new_n100_));
  NO3        g078(.A(new_new_n100_), .B(new_new_n82_), .C(new_new_n52_), .Y(new_new_n101_));
  AN2        g079(.A(i_2_), .B(i_10_), .Y(new_new_n102_));
  NO2        g080(.A(new_new_n102_), .B(i_7_), .Y(new_new_n103_));
  OR2        g081(.A(new_new_n75_), .B(new_new_n57_), .Y(new_new_n104_));
  NO2        g082(.A(i_8_), .B(new_new_n93_), .Y(new_new_n105_));
  NO3        g083(.A(new_new_n105_), .B(new_new_n104_), .C(new_new_n103_), .Y(new_new_n106_));
  NA2        g084(.A(i_12_), .B(i_7_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n108_));
  NA2        g086(.A(new_new_n108_), .B(i_0_), .Y(new_new_n109_));
  NA2        g087(.A(i_11_), .B(i_12_), .Y(new_new_n110_));
  OAI210     g088(.A0(new_new_n109_), .A1(new_new_n107_), .B0(new_new_n110_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(new_new_n106_), .Y(new_new_n112_));
  NAi41      g090(.An(new_new_n101_), .B(new_new_n112_), .C(new_new_n99_), .D(new_new_n92_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n114_));
  NA2        g092(.A(i_7_), .B(new_new_n25_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n115_), .B(new_new_n114_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n116_), .B(new_new_n46_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n83_), .B(new_new_n82_), .Y(new_new_n118_));
  NAi21      g096(.An(i_3_), .B(i_8_), .Y(new_new_n119_));
  NO2        g097(.A(i_1_), .B(new_new_n78_), .Y(new_new_n120_));
  NO2        g098(.A(i_6_), .B(i_5_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(i_3_), .Y(new_new_n122_));
  AO210      g100(.A0(new_new_n122_), .A1(new_new_n47_), .B0(new_new_n120_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n123_), .B(new_new_n100_), .Y(new_new_n124_));
  NO3        g102(.A(new_new_n124_), .B(new_new_n113_), .C(new_new_n87_), .Y(new_new_n125_));
  NA3        g103(.A(new_new_n125_), .B(new_new_n74_), .C(new_new_n55_), .Y(mai2));
  NO2        g104(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g105(.A(i_6_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NA4        g107(.A(new_new_n129_), .B(new_new_n72_), .C(new_new_n65_), .D(new_new_n30_), .Y(mai0));
  AN2        g108(.A(i_8_), .B(i_7_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(i_6_), .Y(new_new_n132_));
  NO2        g110(.A(i_12_), .B(i_13_), .Y(new_new_n133_));
  NAi21      g111(.An(i_5_), .B(i_11_), .Y(new_new_n134_));
  NOi21      g112(.An(new_new_n133_), .B(new_new_n134_), .Y(new_new_n135_));
  NO2        g113(.A(i_0_), .B(i_1_), .Y(new_new_n136_));
  NA2        g114(.A(i_2_), .B(i_3_), .Y(new_new_n137_));
  NO2        g115(.A(new_new_n137_), .B(i_4_), .Y(new_new_n138_));
  NA3        g116(.A(new_new_n138_), .B(new_new_n136_), .C(new_new_n135_), .Y(new_new_n139_));
  AN2        g117(.A(new_new_n133_), .B(new_new_n76_), .Y(new_new_n140_));
  NA2        g118(.A(i_1_), .B(i_5_), .Y(new_new_n141_));
  NO2        g119(.A(new_new_n68_), .B(new_new_n46_), .Y(new_new_n142_));
  NA2        g120(.A(new_new_n142_), .B(new_new_n36_), .Y(new_new_n143_));
  NO3        g121(.A(new_new_n143_), .B(new_new_n141_), .C(i_13_), .Y(new_new_n144_));
  OR2        g122(.A(i_0_), .B(i_1_), .Y(new_new_n145_));
  NO3        g123(.A(new_new_n145_), .B(new_new_n75_), .C(i_13_), .Y(new_new_n146_));
  NAi32      g124(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n147_));
  NAi21      g125(.An(new_new_n147_), .B(new_new_n146_), .Y(new_new_n148_));
  NOi21      g126(.An(i_4_), .B(i_10_), .Y(new_new_n149_));
  NA2        g127(.A(new_new_n149_), .B(new_new_n39_), .Y(new_new_n150_));
  NO2        g128(.A(i_3_), .B(i_5_), .Y(new_new_n151_));
  NA2        g129(.A(i_0_), .B(new_new_n151_), .Y(new_new_n152_));
  OAI210     g130(.A0(new_new_n152_), .A1(new_new_n150_), .B0(new_new_n148_), .Y(new_new_n153_));
  NO2        g131(.A(new_new_n153_), .B(new_new_n144_), .Y(new_new_n154_));
  AOI210     g132(.A0(new_new_n154_), .A1(new_new_n139_), .B0(new_new_n132_), .Y(new_new_n155_));
  NOi21      g133(.An(i_4_), .B(i_9_), .Y(new_new_n156_));
  NOi21      g134(.An(i_11_), .B(i_13_), .Y(new_new_n157_));
  NA2        g135(.A(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  BUFFER     g136(.A(new_new_n158_), .Y(new_new_n159_));
  NO2        g137(.A(i_4_), .B(i_5_), .Y(new_new_n160_));
  NAi21      g138(.An(i_12_), .B(i_11_), .Y(new_new_n161_));
  NO2        g139(.A(new_new_n161_), .B(i_13_), .Y(new_new_n162_));
  NA3        g140(.A(new_new_n162_), .B(new_new_n160_), .C(new_new_n76_), .Y(new_new_n163_));
  AOI210     g141(.A0(new_new_n163_), .A1(new_new_n159_), .B0(new_new_n950_), .Y(new_new_n164_));
  NO2        g142(.A(new_new_n68_), .B(new_new_n62_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n36_), .B(i_5_), .Y(new_new_n166_));
  NAi31      g144(.An(new_new_n166_), .B(new_new_n140_), .C(i_11_), .Y(new_new_n167_));
  NA2        g145(.A(i_3_), .B(i_5_), .Y(new_new_n168_));
  AOI210     g146(.A0(new_new_n158_), .A1(new_new_n167_), .B0(new_new_n62_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n68_), .B(i_5_), .Y(new_new_n170_));
  NO2        g148(.A(i_13_), .B(i_10_), .Y(new_new_n171_));
  NA3        g149(.A(new_new_n171_), .B(new_new_n170_), .C(new_new_n44_), .Y(new_new_n172_));
  NO2        g150(.A(i_2_), .B(i_1_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(i_3_), .Y(new_new_n174_));
  NAi21      g152(.An(i_4_), .B(i_12_), .Y(new_new_n175_));
  NO4        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n172_), .D(new_new_n25_), .Y(new_new_n176_));
  NO3        g154(.A(new_new_n176_), .B(new_new_n169_), .C(new_new_n164_), .Y(new_new_n177_));
  INV        g155(.A(i_8_), .Y(new_new_n178_));
  NA2        g156(.A(i_8_), .B(i_6_), .Y(new_new_n179_));
  NO3        g157(.A(i_3_), .B(new_new_n78_), .C(new_new_n48_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(new_new_n105_), .Y(new_new_n181_));
  NO3        g159(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n182_));
  NA3        g160(.A(new_new_n182_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n183_));
  NO3        g161(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n184_));
  OAI210     g162(.A0(new_new_n88_), .A1(i_12_), .B0(new_new_n184_), .Y(new_new_n185_));
  AOI210     g163(.A0(new_new_n185_), .A1(new_new_n183_), .B0(new_new_n181_), .Y(new_new_n186_));
  NO2        g164(.A(i_3_), .B(i_8_), .Y(new_new_n187_));
  NO3        g165(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n188_));
  NA3        g166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n39_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n95_), .B(new_new_n57_), .Y(new_new_n190_));
  NO2        g168(.A(i_13_), .B(i_9_), .Y(new_new_n191_));
  NA3        g169(.A(new_new_n191_), .B(i_6_), .C(new_new_n178_), .Y(new_new_n192_));
  NAi21      g170(.An(i_12_), .B(i_3_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n44_), .B(i_5_), .Y(new_new_n194_));
  NO3        g172(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n195_));
  NA2        g173(.A(new_new_n195_), .B(i_10_), .Y(new_new_n196_));
  OAI220     g174(.A0(new_new_n196_), .A1(new_new_n192_), .B0(new_new_n57_), .B1(new_new_n189_), .Y(new_new_n197_));
  AOI210     g175(.A0(new_new_n197_), .A1(i_7_), .B0(new_new_n186_), .Y(new_new_n198_));
  OAI220     g176(.A0(new_new_n198_), .A1(i_4_), .B0(new_new_n179_), .B1(new_new_n177_), .Y(new_new_n199_));
  NA3        g177(.A(i_13_), .B(new_new_n178_), .C(i_10_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n200_), .B(i_12_), .Y(new_new_n201_));
  NA2        g179(.A(i_0_), .B(i_5_), .Y(new_new_n202_));
  OAI220     g180(.A0(new_new_n78_), .A1(new_new_n174_), .B0(new_new_n62_), .B1(new_new_n122_), .Y(new_new_n203_));
  NAi31      g181(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n36_), .B(i_13_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n206_));
  NA3        g184(.A(new_new_n206_), .B(i_0_), .C(new_new_n205_), .Y(new_new_n207_));
  INV        g185(.A(i_13_), .Y(new_new_n208_));
  NO2        g186(.A(i_12_), .B(new_new_n208_), .Y(new_new_n209_));
  NA3        g187(.A(new_new_n209_), .B(new_new_n182_), .C(new_new_n180_), .Y(new_new_n210_));
  OAI210     g188(.A0(new_new_n207_), .A1(new_new_n204_), .B0(new_new_n210_), .Y(new_new_n211_));
  AOI220     g189(.A0(new_new_n211_), .A1(new_new_n131_), .B0(new_new_n203_), .B1(new_new_n201_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(new_new_n37_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n168_), .B(i_4_), .Y(new_new_n214_));
  NA2        g192(.A(new_new_n214_), .B(new_new_n213_), .Y(new_new_n215_));
  OR2        g193(.A(i_8_), .B(i_7_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n216_), .B(new_new_n78_), .Y(new_new_n217_));
  INV        g195(.A(i_12_), .Y(new_new_n218_));
  NO3        g196(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n219_));
  NA2        g197(.A(i_2_), .B(i_1_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n221_));
  NAi21      g199(.An(i_4_), .B(i_3_), .Y(new_new_n222_));
  NO2        g200(.A(i_0_), .B(i_6_), .Y(new_new_n223_));
  NOi41      g201(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  BUFFER     g203(.A(new_new_n225_), .Y(new_new_n226_));
  INV        g204(.A(new_new_n226_), .Y(new_new_n227_));
  AOI220     g205(.A0(new_new_n227_), .A1(new_new_n39_), .B0(new_new_n221_), .B1(new_new_n191_), .Y(new_new_n228_));
  NO2        g206(.A(i_11_), .B(new_new_n208_), .Y(new_new_n229_));
  NOi21      g207(.An(i_1_), .B(i_6_), .Y(new_new_n230_));
  NAi21      g208(.An(i_3_), .B(i_7_), .Y(new_new_n231_));
  NA2        g209(.A(new_new_n218_), .B(i_9_), .Y(new_new_n232_));
  OR4        g210(.A(new_new_n232_), .B(new_new_n231_), .C(new_new_n230_), .D(new_new_n170_), .Y(new_new_n233_));
  NO2        g211(.A(i_12_), .B(i_3_), .Y(new_new_n234_));
  NA2        g212(.A(i_3_), .B(i_9_), .Y(new_new_n235_));
  NAi21      g213(.An(i_7_), .B(i_10_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n237_), .B(new_new_n63_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n233_), .Y(new_new_n239_));
  NA3        g217(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n240_));
  INV        g218(.A(new_new_n132_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n218_), .B(i_13_), .Y(new_new_n242_));
  NO2        g220(.A(new_new_n242_), .B(new_new_n70_), .Y(new_new_n243_));
  AOI220     g221(.A0(new_new_n243_), .A1(new_new_n241_), .B0(new_new_n239_), .B1(new_new_n229_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n216_), .B(new_new_n37_), .Y(new_new_n245_));
  NA2        g223(.A(i_12_), .B(i_6_), .Y(new_new_n246_));
  OR2        g224(.A(i_13_), .B(i_9_), .Y(new_new_n247_));
  NO3        g225(.A(new_new_n247_), .B(new_new_n246_), .C(new_new_n48_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n222_), .B(i_2_), .Y(new_new_n249_));
  NA3        g227(.A(new_new_n249_), .B(new_new_n248_), .C(new_new_n44_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n229_), .B(i_9_), .Y(new_new_n251_));
  OAI210     g229(.A0(new_new_n62_), .A1(new_new_n251_), .B0(new_new_n250_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n142_), .B(new_new_n62_), .Y(new_new_n253_));
  NO3        g231(.A(i_11_), .B(new_new_n208_), .C(new_new_n25_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n231_), .B(i_8_), .Y(new_new_n255_));
  NO2        g233(.A(i_6_), .B(new_new_n48_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n255_), .B(new_new_n254_), .Y(new_new_n257_));
  NA3        g235(.A(i_3_), .B(new_new_n245_), .C(new_new_n209_), .Y(new_new_n258_));
  AOI210     g236(.A0(new_new_n258_), .A1(new_new_n257_), .B0(new_new_n253_), .Y(new_new_n259_));
  AOI210     g237(.A0(new_new_n252_), .A1(new_new_n245_), .B0(new_new_n259_), .Y(new_new_n260_));
  NA4        g238(.A(new_new_n260_), .B(new_new_n244_), .C(new_new_n228_), .D(new_new_n212_), .Y(new_new_n261_));
  NO3        g239(.A(i_12_), .B(new_new_n208_), .C(new_new_n37_), .Y(new_new_n262_));
  INV        g240(.A(new_new_n262_), .Y(new_new_n263_));
  NA2        g241(.A(i_8_), .B(new_new_n93_), .Y(new_new_n264_));
  NO2        g242(.A(i_3_), .B(new_new_n264_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n220_), .B(i_0_), .Y(new_new_n266_));
  NA2        g244(.A(new_new_n256_), .B(new_new_n26_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n267_), .B(new_new_n958_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n58_), .B(i_6_), .Y(new_new_n269_));
  NA3        g247(.A(new_new_n269_), .B(i_1_), .C(new_new_n151_), .Y(new_new_n270_));
  OAI210     g248(.A0(new_new_n152_), .A1(new_new_n132_), .B0(new_new_n270_), .Y(new_new_n271_));
  NO3        g249(.A(new_new_n271_), .B(new_new_n268_), .C(new_new_n265_), .Y(new_new_n272_));
  NO2        g250(.A(i_3_), .B(i_10_), .Y(new_new_n273_));
  NA3        g251(.A(new_new_n273_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n274_));
  NA2        g252(.A(i_1_), .B(new_new_n36_), .Y(new_new_n275_));
  AN2        g253(.A(i_3_), .B(i_10_), .Y(new_new_n276_));
  NA4        g254(.A(new_new_n276_), .B(new_new_n182_), .C(new_new_n162_), .D(new_new_n160_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n278_));
  OR2        g256(.A(new_new_n275_), .B(new_new_n274_), .Y(new_new_n279_));
  OAI220     g257(.A0(new_new_n279_), .A1(i_6_), .B0(new_new_n272_), .B1(new_new_n263_), .Y(new_new_n280_));
  NO4        g258(.A(new_new_n280_), .B(new_new_n261_), .C(new_new_n199_), .D(new_new_n155_), .Y(new_new_n281_));
  NO3        g259(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n282_));
  NO3        g260(.A(i_6_), .B(new_new_n178_), .C(i_7_), .Y(new_new_n283_));
  NA2        g261(.A(new_new_n283_), .B(new_new_n182_), .Y(new_new_n284_));
  AOI210     g262(.A0(new_new_n284_), .A1(new_new_n220_), .B0(i_5_), .Y(new_new_n285_));
  NO2        g263(.A(i_2_), .B(i_3_), .Y(new_new_n286_));
  OR2        g264(.A(i_0_), .B(i_5_), .Y(new_new_n287_));
  NA2        g265(.A(new_new_n202_), .B(new_new_n287_), .Y(new_new_n288_));
  NA4        g266(.A(new_new_n288_), .B(new_new_n217_), .C(new_new_n286_), .D(i_1_), .Y(new_new_n289_));
  NA3        g267(.A(new_new_n266_), .B(new_new_n151_), .C(new_new_n105_), .Y(new_new_n290_));
  NAi21      g268(.An(i_8_), .B(i_7_), .Y(new_new_n291_));
  NA3        g269(.A(i_2_), .B(i_7_), .C(new_new_n151_), .Y(new_new_n292_));
  NA3        g270(.A(new_new_n292_), .B(new_new_n290_), .C(new_new_n289_), .Y(new_new_n293_));
  OAI210     g271(.A0(new_new_n293_), .A1(new_new_n285_), .B0(i_4_), .Y(new_new_n294_));
  NO2        g272(.A(i_12_), .B(i_10_), .Y(new_new_n295_));
  NOi21      g273(.An(i_5_), .B(i_0_), .Y(new_new_n296_));
  NO3        g274(.A(new_new_n275_), .B(new_new_n296_), .C(new_new_n119_), .Y(new_new_n297_));
  NA4        g275(.A(new_new_n77_), .B(new_new_n36_), .C(new_new_n78_), .D(i_8_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n297_), .B(new_new_n295_), .Y(new_new_n299_));
  NO2        g277(.A(i_6_), .B(i_8_), .Y(new_new_n300_));
  AN2        g278(.A(i_0_), .B(new_new_n300_), .Y(new_new_n301_));
  NO2        g279(.A(i_1_), .B(i_7_), .Y(new_new_n302_));
  NA3        g280(.A(new_new_n300_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n303_));
  NA3        g281(.A(new_new_n303_), .B(new_new_n299_), .C(new_new_n294_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n95_), .B(new_new_n115_), .Y(new_new_n305_));
  NA2        g283(.A(new_new_n305_), .B(i_3_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n85_), .B(new_new_n178_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n178_), .B(i_9_), .Y(new_new_n308_));
  AOI210     g286(.A0(new_new_n956_), .A1(new_new_n306_), .B0(new_new_n150_), .Y(new_new_n309_));
  AOI210     g287(.A0(new_new_n304_), .A1(new_new_n282_), .B0(new_new_n309_), .Y(new_new_n310_));
  NOi32      g288(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n311_));
  INV        g289(.A(new_new_n311_), .Y(new_new_n312_));
  NAi21      g290(.An(i_1_), .B(i_5_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n313_), .B(i_0_), .Y(new_new_n314_));
  NA2        g292(.A(new_new_n314_), .B(new_new_n25_), .Y(new_new_n315_));
  OAI210     g293(.A0(new_new_n315_), .A1(new_new_n147_), .B0(new_new_n225_), .Y(new_new_n316_));
  NAi41      g294(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n317_));
  OAI220     g295(.A0(new_new_n317_), .A1(new_new_n313_), .B0(new_new_n204_), .B1(new_new_n147_), .Y(new_new_n318_));
  AOI210     g296(.A0(new_new_n317_), .A1(new_new_n147_), .B0(new_new_n145_), .Y(new_new_n319_));
  NOi32      g297(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n320_), .B(new_new_n46_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n321_), .B(i_0_), .Y(new_new_n322_));
  OR3        g300(.A(new_new_n322_), .B(new_new_n319_), .C(new_new_n318_), .Y(new_new_n323_));
  NO2        g301(.A(i_1_), .B(new_new_n93_), .Y(new_new_n324_));
  NAi21      g302(.An(i_3_), .B(i_4_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n325_), .B(i_9_), .Y(new_new_n326_));
  AN2        g304(.A(i_6_), .B(i_7_), .Y(new_new_n327_));
  OAI210     g305(.A0(new_new_n327_), .A1(new_new_n324_), .B0(new_new_n326_), .Y(new_new_n328_));
  NA2        g306(.A(i_2_), .B(i_7_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n325_), .B(i_10_), .Y(new_new_n330_));
  NA3        g308(.A(new_new_n330_), .B(new_new_n329_), .C(new_new_n223_), .Y(new_new_n331_));
  AOI210     g309(.A0(new_new_n331_), .A1(new_new_n328_), .B0(new_new_n170_), .Y(new_new_n332_));
  AOI210     g310(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n333_));
  OAI210     g311(.A0(new_new_n333_), .A1(new_new_n173_), .B0(new_new_n330_), .Y(new_new_n334_));
  AOI220     g312(.A0(new_new_n330_), .A1(new_new_n302_), .B0(new_new_n219_), .B1(new_new_n173_), .Y(new_new_n335_));
  AOI210     g313(.A0(new_new_n335_), .A1(new_new_n334_), .B0(i_5_), .Y(new_new_n336_));
  NO4        g314(.A(new_new_n336_), .B(new_new_n332_), .C(new_new_n323_), .D(new_new_n316_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n337_), .B(new_new_n312_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n339_));
  AN2        g317(.A(i_12_), .B(i_5_), .Y(new_new_n340_));
  NO2        g318(.A(i_4_), .B(new_new_n26_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n342_));
  NO2        g320(.A(i_11_), .B(i_6_), .Y(new_new_n343_));
  NA3        g321(.A(new_new_n343_), .B(i_2_), .C(new_new_n208_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n344_), .B(new_new_n342_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n222_), .B(i_5_), .Y(new_new_n346_));
  NO2        g324(.A(i_5_), .B(i_10_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n133_), .B(new_new_n45_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n222_), .Y(new_new_n349_));
  OAI210     g327(.A0(new_new_n349_), .A1(new_new_n345_), .B0(new_new_n339_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n139_), .B(new_new_n78_), .Y(new_new_n352_));
  OAI210     g330(.A0(new_new_n352_), .A1(new_new_n345_), .B0(new_new_n351_), .Y(new_new_n353_));
  NO2        g331(.A(i_11_), .B(i_12_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n347_), .B(new_new_n218_), .Y(new_new_n355_));
  OAI220     g333(.A0(new_new_n36_), .A1(new_new_n204_), .B0(new_new_n355_), .B1(new_new_n298_), .Y(new_new_n356_));
  NAi21      g334(.An(i_13_), .B(i_0_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(new_new_n220_), .Y(new_new_n358_));
  NA2        g336(.A(new_new_n356_), .B(new_new_n358_), .Y(new_new_n359_));
  NA3        g337(.A(new_new_n359_), .B(new_new_n353_), .C(new_new_n350_), .Y(new_new_n360_));
  NO2        g338(.A(i_0_), .B(i_11_), .Y(new_new_n361_));
  AN2        g339(.A(i_1_), .B(i_6_), .Y(new_new_n362_));
  NOi21      g340(.An(i_2_), .B(i_12_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n131_), .B(i_9_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n364_), .B(i_4_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n363_), .B(new_new_n365_), .Y(new_new_n366_));
  NAi21      g344(.An(i_9_), .B(i_4_), .Y(new_new_n367_));
  OR2        g345(.A(i_13_), .B(i_10_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n158_), .B(new_new_n114_), .Y(new_new_n369_));
  BUFFER     g347(.A(new_new_n200_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n371_));
  NA2        g349(.A(new_new_n262_), .B(new_new_n371_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n256_), .B(new_new_n195_), .Y(new_new_n373_));
  OAI220     g351(.A0(new_new_n373_), .A1(new_new_n370_), .B0(new_new_n372_), .B1(new_new_n95_), .Y(new_new_n374_));
  INV        g352(.A(new_new_n374_), .Y(new_new_n375_));
  AOI210     g353(.A0(new_new_n375_), .A1(new_new_n366_), .B0(new_new_n26_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n290_), .B(new_new_n289_), .Y(new_new_n377_));
  AOI220     g355(.A0(new_new_n269_), .A1(i_2_), .B0(new_new_n266_), .B1(i_7_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(i_5_), .Y(new_new_n379_));
  AOI220     g357(.A0(i_3_), .A1(i_1_), .B0(i_3_), .B1(new_new_n195_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n380_), .B(new_new_n264_), .Y(new_new_n381_));
  NO3        g359(.A(new_new_n381_), .B(new_new_n379_), .C(new_new_n377_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n180_), .B(new_new_n88_), .Y(new_new_n383_));
  NA3        g361(.A(i_2_), .B(new_new_n151_), .C(new_new_n78_), .Y(new_new_n384_));
  AOI210     g362(.A0(new_new_n384_), .A1(new_new_n383_), .B0(new_new_n291_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n178_), .B(i_10_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n63_), .B(i_2_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n269_), .B(i_2_), .Y(new_new_n388_));
  OAI220     g366(.A0(new_new_n388_), .A1(new_new_n168_), .B0(new_new_n387_), .B1(new_new_n386_), .Y(new_new_n389_));
  NA3        g367(.A(new_new_n302_), .B(new_new_n301_), .C(i_5_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n283_), .B(new_new_n288_), .Y(new_new_n391_));
  OAI210     g369(.A0(new_new_n391_), .A1(new_new_n174_), .B0(new_new_n390_), .Y(new_new_n392_));
  NO3        g370(.A(new_new_n392_), .B(new_new_n389_), .C(new_new_n385_), .Y(new_new_n393_));
  AOI210     g371(.A0(new_new_n393_), .A1(new_new_n382_), .B0(new_new_n251_), .Y(new_new_n394_));
  NO4        g372(.A(new_new_n394_), .B(new_new_n376_), .C(new_new_n360_), .D(new_new_n338_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n68_), .B(i_13_), .Y(new_new_n396_));
  NA3        g374(.A(new_new_n396_), .B(i_1_), .C(i_2_), .Y(new_new_n397_));
  NO2        g375(.A(i_10_), .B(i_9_), .Y(new_new_n398_));
  NAi21      g376(.An(i_12_), .B(i_8_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(i_3_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n400_), .B(new_new_n398_), .Y(new_new_n401_));
  OAI220     g379(.A0(i_4_), .A1(new_new_n189_), .B0(new_new_n401_), .B1(new_new_n397_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n278_), .B(i_0_), .Y(new_new_n403_));
  NO3        g381(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n246_), .B(new_new_n89_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n405_), .B(new_new_n404_), .Y(new_new_n406_));
  NA2        g384(.A(i_8_), .B(i_9_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n262_), .B(new_new_n190_), .Y(new_new_n408_));
  OAI220     g386(.A0(new_new_n408_), .A1(new_new_n407_), .B0(new_new_n406_), .B1(new_new_n403_), .Y(new_new_n409_));
  NO3        g387(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n410_));
  NA3        g388(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n411_));
  NA4        g389(.A(new_new_n134_), .B(new_new_n108_), .C(new_new_n75_), .D(new_new_n23_), .Y(new_new_n412_));
  NO2        g390(.A(new_new_n412_), .B(new_new_n411_), .Y(new_new_n413_));
  NO3        g391(.A(new_new_n413_), .B(new_new_n409_), .C(new_new_n402_), .Y(new_new_n414_));
  OR2        g392(.A(new_new_n192_), .B(new_new_n215_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n88_), .B(i_13_), .Y(new_new_n416_));
  NA2        g394(.A(i_3_), .B(new_new_n339_), .Y(new_new_n417_));
  NO2        g395(.A(i_2_), .B(i_13_), .Y(new_new_n418_));
  NA3        g396(.A(new_new_n418_), .B(new_new_n149_), .C(new_new_n91_), .Y(new_new_n419_));
  OAI220     g397(.A0(new_new_n419_), .A1(new_new_n218_), .B0(new_new_n417_), .B1(new_new_n416_), .Y(new_new_n420_));
  NO3        g398(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n421_));
  NO2        g399(.A(i_6_), .B(i_7_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n422_), .B(new_new_n421_), .Y(new_new_n423_));
  OR2        g401(.A(i_11_), .B(i_8_), .Y(new_new_n424_));
  NOi21      g402(.An(i_2_), .B(i_7_), .Y(new_new_n425_));
  NAi31      g403(.An(new_new_n424_), .B(new_new_n425_), .C(i_0_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n368_), .B(new_new_n426_), .Y(new_new_n427_));
  NO2        g405(.A(i_6_), .B(i_10_), .Y(new_new_n428_));
  NA4        g406(.A(new_new_n428_), .B(new_new_n282_), .C(i_8_), .D(new_new_n218_), .Y(new_new_n429_));
  NO2        g407(.A(new_new_n429_), .B(new_new_n143_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n224_), .B(new_new_n157_), .C(new_new_n121_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n145_), .B(i_3_), .Y(new_new_n433_));
  NAi31      g411(.An(new_new_n432_), .B(new_new_n433_), .C(new_new_n209_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n434_), .B(new_new_n431_), .Y(new_new_n435_));
  NO4        g413(.A(new_new_n435_), .B(new_new_n430_), .C(new_new_n427_), .D(new_new_n420_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n410_), .B(new_new_n347_), .Y(new_new_n437_));
  NO2        g415(.A(new_new_n437_), .B(new_new_n207_), .Y(new_new_n438_));
  NAi21      g416(.An(new_new_n200_), .B(new_new_n354_), .Y(new_new_n439_));
  NO2        g417(.A(new_new_n26_), .B(i_5_), .Y(new_new_n440_));
  NA3        g418(.A(i_6_), .B(new_new_n440_), .C(new_new_n131_), .Y(new_new_n441_));
  OR3        g419(.A(new_new_n275_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n442_));
  OAI220     g420(.A0(new_new_n442_), .A1(new_new_n441_), .B0(i_1_), .B1(new_new_n439_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n27_), .B(i_10_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n282_), .B(new_new_n219_), .Y(new_new_n445_));
  OAI220     g423(.A0(new_new_n445_), .A1(new_new_n387_), .B0(new_new_n444_), .B1(new_new_n416_), .Y(new_new_n446_));
  NA4        g424(.A(new_new_n276_), .B(new_new_n206_), .C(new_new_n68_), .D(new_new_n218_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n447_), .B(new_new_n423_), .Y(new_new_n448_));
  NO4        g426(.A(new_new_n448_), .B(new_new_n446_), .C(new_new_n443_), .D(new_new_n438_), .Y(new_new_n449_));
  NA4        g427(.A(new_new_n449_), .B(new_new_n436_), .C(new_new_n415_), .D(new_new_n414_), .Y(new_new_n450_));
  NA3        g428(.A(new_new_n276_), .B(new_new_n162_), .C(new_new_n160_), .Y(new_new_n451_));
  OAI210     g429(.A0(new_new_n274_), .A1(new_new_n166_), .B0(new_new_n451_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n217_), .B(new_new_n452_), .Y(new_new_n453_));
  AN2        g431(.A(new_new_n57_), .B(new_new_n404_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n282_), .B(i_0_), .Y(new_new_n455_));
  OAI210     g433(.A0(new_new_n455_), .A1(new_new_n215_), .B0(new_new_n277_), .Y(new_new_n456_));
  AOI220     g434(.A0(new_new_n456_), .A1(i_7_), .B0(new_new_n454_), .B1(new_new_n278_), .Y(new_new_n457_));
  NA4        g435(.A(new_new_n396_), .B(i_1_), .C(new_new_n187_), .D(i_2_), .Y(new_new_n458_));
  INV        g436(.A(new_new_n458_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n340_), .B(new_new_n208_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n311_), .B(new_new_n68_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n327_), .B(new_new_n320_), .Y(new_new_n462_));
  AO210      g440(.A0(new_new_n461_), .A1(new_new_n460_), .B0(new_new_n462_), .Y(new_new_n463_));
  INV        g441(.A(new_new_n463_), .Y(new_new_n464_));
  AOI210     g442(.A0(new_new_n459_), .A1(new_new_n188_), .B0(new_new_n464_), .Y(new_new_n465_));
  NO2        g443(.A(i_7_), .B(new_new_n183_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n168_), .B(new_new_n78_), .Y(new_new_n467_));
  AOI220     g445(.A0(new_new_n467_), .A1(new_new_n466_), .B0(new_new_n949_), .B1(new_new_n369_), .Y(new_new_n468_));
  NA4        g446(.A(new_new_n468_), .B(new_new_n465_), .C(new_new_n457_), .D(new_new_n453_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n346_), .B(i_1_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n342_), .B(new_new_n470_), .Y(new_new_n471_));
  NO2        g449(.A(i_12_), .B(new_new_n178_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n472_), .B(new_new_n208_), .Y(new_new_n473_));
  NO2        g451(.A(i_10_), .B(new_new_n473_), .Y(new_new_n474_));
  NOi31      g452(.An(new_new_n283_), .B(new_new_n368_), .C(new_new_n38_), .Y(new_new_n475_));
  OAI210     g453(.A0(new_new_n475_), .A1(new_new_n474_), .B0(new_new_n471_), .Y(new_new_n476_));
  NO2        g454(.A(i_8_), .B(i_7_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n44_), .B(i_10_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n478_), .B(i_6_), .Y(new_new_n479_));
  NA3        g457(.A(new_new_n479_), .B(i_2_), .C(new_new_n477_), .Y(new_new_n480_));
  OAI220     g458(.A0(new_new_n168_), .A1(new_new_n242_), .B0(new_new_n416_), .B1(new_new_n122_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n481_), .B(new_new_n245_), .Y(new_new_n482_));
  NOi31      g460(.An(new_new_n266_), .B(new_new_n274_), .C(new_new_n166_), .Y(new_new_n483_));
  NA3        g461(.A(new_new_n276_), .B(new_new_n160_), .C(new_new_n88_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n145_), .B(i_5_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n485_), .B(new_new_n286_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(new_new_n484_), .Y(new_new_n487_));
  OAI210     g465(.A0(new_new_n487_), .A1(new_new_n483_), .B0(new_new_n410_), .Y(new_new_n488_));
  NA4        g466(.A(new_new_n488_), .B(new_new_n482_), .C(new_new_n480_), .D(new_new_n476_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n262_), .B(new_new_n77_), .Y(new_new_n490_));
  NO2        g468(.A(i_11_), .B(new_new_n490_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n269_), .B(i_2_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n492_), .B(new_new_n159_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n206_), .B(i_0_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n398_), .B(new_new_n205_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n494_), .B(new_new_n495_), .Y(new_new_n496_));
  NA2        g474(.A(i_0_), .B(new_new_n48_), .Y(new_new_n497_));
  NA3        g475(.A(new_new_n472_), .B(new_new_n254_), .C(new_new_n497_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n498_), .Y(new_new_n499_));
  NO4        g477(.A(new_new_n499_), .B(new_new_n496_), .C(new_new_n493_), .D(new_new_n491_), .Y(new_new_n500_));
  NO4        g478(.A(new_new_n230_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n501_));
  NO3        g479(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n216_), .B(new_new_n36_), .Y(new_new_n503_));
  AN2        g481(.A(new_new_n503_), .B(new_new_n502_), .Y(new_new_n504_));
  OA210      g482(.A0(new_new_n504_), .A1(new_new_n501_), .B0(new_new_n311_), .Y(new_new_n505_));
  NO2        g483(.A(new_new_n368_), .B(i_1_), .Y(new_new_n506_));
  AN3        g484(.A(new_new_n506_), .B(new_new_n365_), .C(i_2_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n378_), .B(new_new_n163_), .Y(new_new_n508_));
  NO3        g486(.A(new_new_n508_), .B(new_new_n507_), .C(new_new_n505_), .Y(new_new_n509_));
  NOi21      g487(.An(i_10_), .B(i_6_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n78_), .B(new_new_n25_), .Y(new_new_n511_));
  AOI220     g489(.A0(new_new_n262_), .A1(new_new_n511_), .B0(new_new_n254_), .B1(new_new_n510_), .Y(new_new_n512_));
  NO2        g490(.A(new_new_n512_), .B(new_new_n403_), .Y(new_new_n513_));
  NO2        g491(.A(new_new_n107_), .B(new_new_n23_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n283_), .B(i_0_), .Y(new_new_n515_));
  AOI220     g493(.A0(new_new_n515_), .A1(new_new_n388_), .B0(new_new_n158_), .B1(new_new_n167_), .Y(new_new_n516_));
  NOi21      g494(.An(new_new_n135_), .B(new_new_n298_), .Y(new_new_n517_));
  NO3        g495(.A(new_new_n517_), .B(new_new_n516_), .C(new_new_n513_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n461_), .B(new_new_n335_), .Y(new_new_n519_));
  INV        g497(.A(new_new_n286_), .Y(new_new_n520_));
  NO2        g498(.A(i_12_), .B(new_new_n78_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n521_), .B(new_new_n254_), .C(new_new_n497_), .Y(new_new_n522_));
  NA3        g500(.A(new_new_n343_), .B(new_new_n262_), .C(new_new_n202_), .Y(new_new_n523_));
  AOI210     g501(.A0(new_new_n523_), .A1(new_new_n522_), .B0(new_new_n520_), .Y(new_new_n524_));
  NO3        g502(.A(i_4_), .B(i_8_), .C(new_new_n274_), .Y(new_new_n525_));
  OR2        g503(.A(i_5_), .B(new_new_n362_), .Y(new_new_n526_));
  AOI210     g504(.A0(i_6_), .A1(new_new_n526_), .B0(new_new_n439_), .Y(new_new_n527_));
  NO4        g505(.A(new_new_n527_), .B(new_new_n525_), .C(new_new_n524_), .D(new_new_n519_), .Y(new_new_n528_));
  NA4        g506(.A(new_new_n528_), .B(new_new_n518_), .C(new_new_n509_), .D(new_new_n500_), .Y(new_new_n529_));
  NO4        g507(.A(new_new_n529_), .B(new_new_n489_), .C(new_new_n469_), .D(new_new_n450_), .Y(new_new_n530_));
  NA4        g508(.A(new_new_n530_), .B(new_new_n395_), .C(new_new_n310_), .D(new_new_n281_), .Y(mai7));
  NO2        g509(.A(new_new_n100_), .B(new_new_n82_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n341_), .B(new_new_n532_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n428_), .B(new_new_n77_), .Y(new_new_n534_));
  NA2        g512(.A(i_11_), .B(new_new_n178_), .Y(new_new_n535_));
  OAI210     g513(.A0(new_new_n951_), .A1(new_new_n534_), .B0(new_new_n533_), .Y(new_new_n536_));
  NA3        g514(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n218_), .B(i_4_), .Y(new_new_n538_));
  NA2        g516(.A(new_new_n538_), .B(i_8_), .Y(new_new_n539_));
  AOI210     g517(.A0(new_new_n539_), .A1(new_new_n97_), .B0(new_new_n537_), .Y(new_new_n540_));
  OAI210     g518(.A0(new_new_n81_), .A1(new_new_n187_), .B0(new_new_n188_), .Y(new_new_n541_));
  NO2        g519(.A(i_7_), .B(new_new_n37_), .Y(new_new_n542_));
  NA2        g520(.A(i_4_), .B(i_8_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n541_), .B(i_13_), .Y(new_new_n544_));
  NO3        g522(.A(new_new_n544_), .B(new_new_n540_), .C(new_new_n536_), .Y(new_new_n545_));
  AOI210     g523(.A0(new_new_n119_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n546_));
  AOI210     g524(.A0(new_new_n546_), .A1(new_new_n218_), .B0(new_new_n149_), .Y(new_new_n547_));
  OR2        g525(.A(i_6_), .B(i_10_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n548_), .B(new_new_n23_), .Y(new_new_n549_));
  OR3        g527(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n550_));
  NO3        g528(.A(new_new_n550_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n184_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n551_), .B(new_new_n549_), .Y(new_new_n553_));
  OA220      g531(.A0(new_new_n553_), .A1(new_new_n520_), .B0(new_new_n547_), .B1(new_new_n247_), .Y(new_new_n554_));
  AOI210     g532(.A0(new_new_n554_), .A1(new_new_n545_), .B0(new_new_n62_), .Y(new_new_n555_));
  NOi21      g533(.An(i_11_), .B(i_7_), .Y(new_new_n556_));
  AO210      g534(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n557_), .B(new_new_n556_), .Y(new_new_n558_));
  NA2        g536(.A(new_new_n558_), .B(new_new_n191_), .Y(new_new_n559_));
  NA3        g537(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n560_));
  NAi31      g538(.An(new_new_n560_), .B(i_12_), .C(i_11_), .Y(new_new_n561_));
  AOI210     g539(.A0(new_new_n561_), .A1(new_new_n559_), .B0(new_new_n62_), .Y(new_new_n562_));
  NA2        g540(.A(new_new_n80_), .B(new_new_n62_), .Y(new_new_n563_));
  AO210      g541(.A0(new_new_n563_), .A1(new_new_n335_), .B0(new_new_n40_), .Y(new_new_n564_));
  NO3        g542(.A(new_new_n236_), .B(new_new_n193_), .C(new_new_n535_), .Y(new_new_n565_));
  OAI210     g543(.A0(new_new_n565_), .A1(new_new_n209_), .B0(new_new_n62_), .Y(new_new_n566_));
  NA2        g544(.A(new_new_n363_), .B(new_new_n31_), .Y(new_new_n567_));
  OR2        g545(.A(new_new_n193_), .B(new_new_n100_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n568_), .B(new_new_n567_), .Y(new_new_n569_));
  NO2        g547(.A(new_new_n62_), .B(i_9_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n570_), .B(i_4_), .Y(new_new_n571_));
  NA2        g549(.A(new_new_n571_), .B(new_new_n569_), .Y(new_new_n572_));
  NO2        g550(.A(i_1_), .B(i_12_), .Y(new_new_n573_));
  NA3        g551(.A(new_new_n572_), .B(new_new_n566_), .C(new_new_n564_), .Y(new_new_n574_));
  OAI210     g552(.A0(new_new_n574_), .A1(new_new_n562_), .B0(i_6_), .Y(new_new_n575_));
  OAI210     g553(.A0(new_new_n560_), .A1(new_new_n100_), .B0(new_new_n411_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n576_), .B(new_new_n521_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n218_), .B(new_new_n78_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n578_), .B(i_11_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n577_), .B(new_new_n406_), .Y(new_new_n580_));
  NO4        g558(.A(i_12_), .B(new_new_n119_), .C(i_13_), .D(new_new_n78_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n581_), .B(new_new_n570_), .Y(new_new_n582_));
  NO3        g560(.A(new_new_n548_), .B(new_new_n216_), .C(new_new_n23_), .Y(new_new_n583_));
  AOI210     g561(.A0(i_1_), .A1(new_new_n237_), .B0(new_new_n583_), .Y(new_new_n584_));
  OAI210     g562(.A0(new_new_n584_), .A1(new_new_n44_), .B0(new_new_n582_), .Y(new_new_n585_));
  NA3        g563(.A(new_new_n477_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n586_));
  INV        g564(.A(i_2_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n127_), .B(i_9_), .Y(new_new_n588_));
  NA3        g566(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n46_), .B(i_1_), .Y(new_new_n590_));
  NA3        g568(.A(new_new_n590_), .B(new_new_n246_), .C(new_new_n44_), .Y(new_new_n591_));
  OAI220     g569(.A0(new_new_n591_), .A1(new_new_n589_), .B0(new_new_n588_), .B1(new_new_n587_), .Y(new_new_n592_));
  NA3        g570(.A(new_new_n570_), .B(new_new_n286_), .C(i_6_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n593_), .B(new_new_n23_), .Y(new_new_n594_));
  NAi21      g572(.An(new_new_n586_), .B(new_new_n84_), .Y(new_new_n595_));
  INV        g573(.A(new_new_n595_), .Y(new_new_n596_));
  OR3        g574(.A(new_new_n596_), .B(new_new_n594_), .C(new_new_n592_), .Y(new_new_n597_));
  NO3        g575(.A(new_new_n597_), .B(new_new_n585_), .C(new_new_n580_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n218_), .B(new_new_n93_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n599_), .B(new_new_n556_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n600_), .B(i_1_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n601_), .B(new_new_n550_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n367_), .B(new_new_n78_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n602_), .B(new_new_n46_), .Y(new_new_n604_));
  NA2        g582(.A(i_3_), .B(new_new_n178_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n605_), .B(new_new_n107_), .Y(new_new_n606_));
  AN2        g584(.A(new_new_n606_), .B(new_new_n479_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n216_), .B(new_new_n44_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n78_), .B(i_9_), .Y(new_new_n609_));
  NA2        g587(.A(i_1_), .B(i_3_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n407_), .B(new_new_n85_), .Y(new_new_n611_));
  AOI210     g589(.A0(new_new_n608_), .A1(new_new_n510_), .B0(new_new_n611_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n610_), .Y(new_new_n613_));
  NO2        g591(.A(new_new_n613_), .B(new_new_n607_), .Y(new_new_n614_));
  NA4        g592(.A(new_new_n614_), .B(new_new_n604_), .C(new_new_n598_), .D(new_new_n575_), .Y(new_new_n615_));
  NO3        g593(.A(new_new_n424_), .B(i_3_), .C(i_7_), .Y(new_new_n616_));
  OA210      g594(.A0(new_new_n616_), .A1(new_new_n224_), .B0(new_new_n78_), .Y(new_new_n617_));
  NA2        g595(.A(new_new_n327_), .B(new_new_n326_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n428_), .B(i_4_), .C(new_new_n46_), .Y(new_new_n619_));
  NO3        g597(.A(new_new_n425_), .B(new_new_n543_), .C(new_new_n78_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n25_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n149_), .B(new_new_n77_), .C(new_new_n78_), .Y(new_new_n622_));
  NA4        g600(.A(new_new_n622_), .B(new_new_n621_), .C(new_new_n619_), .D(new_new_n618_), .Y(new_new_n623_));
  OAI210     g601(.A0(new_new_n623_), .A1(new_new_n617_), .B0(i_1_), .Y(new_new_n624_));
  AOI210     g602(.A0(new_new_n246_), .A1(new_new_n89_), .B0(i_1_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n325_), .B(i_2_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n626_), .B(new_new_n625_), .Y(new_new_n627_));
  OAI210     g605(.A0(new_new_n593_), .A1(new_new_n399_), .B0(new_new_n627_), .Y(new_new_n628_));
  INV        g606(.A(new_new_n628_), .Y(new_new_n629_));
  AOI210     g607(.A0(new_new_n629_), .A1(new_new_n624_), .B0(i_13_), .Y(new_new_n630_));
  NA3        g608(.A(i_11_), .B(new_new_n98_), .C(new_new_n127_), .Y(new_new_n631_));
  NA2        g609(.A(new_new_n418_), .B(new_new_n149_), .Y(new_new_n632_));
  OAI210     g610(.A0(new_new_n632_), .A1(new_new_n44_), .B0(new_new_n631_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n425_), .B(new_new_n24_), .Y(new_new_n634_));
  AOI220     g612(.A0(new_new_n634_), .A1(new_new_n603_), .B0(new_new_n224_), .B1(new_new_n120_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n635_), .B(new_new_n40_), .Y(new_new_n636_));
  AOI210     g614(.A0(new_new_n633_), .A1(new_new_n300_), .B0(new_new_n636_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n343_), .B(new_new_n590_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n222_), .Y(new_new_n639_));
  AOI210     g617(.A0(new_new_n399_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n640_));
  NOi31      g618(.An(new_new_n640_), .B(new_new_n534_), .C(new_new_n44_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n118_), .B(i_13_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n589_), .B(new_new_n107_), .Y(new_new_n643_));
  INV        g621(.A(new_new_n643_), .Y(new_new_n644_));
  OAI220     g622(.A0(new_new_n644_), .A1(new_new_n66_), .B0(new_new_n642_), .B1(new_new_n625_), .Y(new_new_n645_));
  NO3        g623(.A(new_new_n66_), .B(new_new_n32_), .C(new_new_n93_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n26_), .B(new_new_n178_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n647_), .B(i_7_), .Y(new_new_n648_));
  NO3        g626(.A(new_new_n425_), .B(new_new_n218_), .C(new_new_n78_), .Y(new_new_n649_));
  AOI210     g627(.A0(new_new_n649_), .A1(new_new_n648_), .B0(new_new_n646_), .Y(new_new_n650_));
  AOI220     g628(.A0(new_new_n343_), .A1(new_new_n590_), .B0(new_new_n84_), .B1(new_new_n94_), .Y(new_new_n651_));
  OAI220     g629(.A0(new_new_n651_), .A1(new_new_n539_), .B0(new_new_n650_), .B1(new_new_n552_), .Y(new_new_n652_));
  NO4        g630(.A(new_new_n652_), .B(new_new_n645_), .C(new_new_n641_), .D(new_new_n639_), .Y(new_new_n653_));
  OR2        g631(.A(i_11_), .B(i_6_), .Y(new_new_n654_));
  NA3        g632(.A(new_new_n538_), .B(new_new_n647_), .C(i_7_), .Y(new_new_n655_));
  AOI210     g633(.A0(new_new_n655_), .A1(new_new_n644_), .B0(new_new_n654_), .Y(new_new_n656_));
  NA3        g634(.A(new_new_n363_), .B(new_new_n542_), .C(new_new_n89_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n579_), .B(i_13_), .Y(new_new_n658_));
  NAi21      g636(.An(i_11_), .B(i_12_), .Y(new_new_n659_));
  NOi41      g637(.An(new_new_n103_), .B(new_new_n659_), .C(i_13_), .D(new_new_n78_), .Y(new_new_n660_));
  NO3        g638(.A(new_new_n425_), .B(new_new_n521_), .C(new_new_n543_), .Y(new_new_n661_));
  AOI210     g639(.A0(new_new_n661_), .A1(new_new_n282_), .B0(new_new_n660_), .Y(new_new_n662_));
  NA3        g640(.A(new_new_n662_), .B(new_new_n658_), .C(new_new_n657_), .Y(new_new_n663_));
  OAI210     g641(.A0(new_new_n663_), .A1(new_new_n656_), .B0(new_new_n62_), .Y(new_new_n664_));
  NO2        g642(.A(i_2_), .B(i_12_), .Y(new_new_n665_));
  OAI210     g643(.A0(new_new_n546_), .A1(new_new_n324_), .B0(new_new_n665_), .Y(new_new_n666_));
  OAI210     g644(.A0(new_new_n218_), .A1(new_new_n326_), .B0(new_new_n324_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n119_), .B(i_2_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n668_), .B(new_new_n573_), .Y(new_new_n669_));
  NA3        g647(.A(new_new_n669_), .B(new_new_n667_), .C(new_new_n666_), .Y(new_new_n670_));
  NA3        g648(.A(new_new_n670_), .B(new_new_n45_), .C(new_new_n208_), .Y(new_new_n671_));
  NA4        g649(.A(new_new_n671_), .B(new_new_n664_), .C(new_new_n653_), .D(new_new_n637_), .Y(new_new_n672_));
  OR4        g650(.A(new_new_n672_), .B(new_new_n630_), .C(new_new_n615_), .D(new_new_n555_), .Y(mai5));
  AOI210     g651(.A0(new_new_n600_), .A1(new_new_n249_), .B0(new_new_n369_), .Y(new_new_n674_));
  AO210      g652(.A0(new_new_n24_), .A1(i_10_), .B0(new_new_n229_), .Y(new_new_n675_));
  NA3        g653(.A(new_new_n675_), .B(new_new_n665_), .C(new_new_n100_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n539_), .B(i_11_), .Y(new_new_n677_));
  OAI210     g655(.A0(new_new_n542_), .A1(new_new_n81_), .B0(new_new_n677_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n676_), .C(new_new_n674_), .Y(new_new_n679_));
  NO3        g657(.A(i_11_), .B(new_new_n218_), .C(i_13_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n681_));
  NA2        g659(.A(i_12_), .B(i_8_), .Y(new_new_n682_));
  OAI210     g660(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n682_), .Y(new_new_n683_));
  INV        g661(.A(new_new_n398_), .Y(new_new_n684_));
  AOI220     g662(.A0(new_new_n286_), .A1(new_new_n514_), .B0(new_new_n683_), .B1(new_new_n681_), .Y(new_new_n685_));
  INV        g663(.A(new_new_n685_), .Y(new_new_n686_));
  NO2        g664(.A(new_new_n686_), .B(new_new_n679_), .Y(new_new_n687_));
  INV        g665(.A(new_new_n157_), .Y(new_new_n688_));
  INV        g666(.A(new_new_n224_), .Y(new_new_n689_));
  OAI210     g667(.A0(new_new_n626_), .A1(new_new_n400_), .B0(new_new_n103_), .Y(new_new_n690_));
  AOI210     g668(.A0(new_new_n690_), .A1(new_new_n689_), .B0(new_new_n688_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n407_), .B(new_new_n26_), .Y(new_new_n692_));
  NO2        g670(.A(new_new_n692_), .B(new_new_n371_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n693_), .B(i_2_), .Y(new_new_n694_));
  INV        g672(.A(new_new_n694_), .Y(new_new_n695_));
  AOI210     g673(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n368_), .Y(new_new_n696_));
  AOI210     g674(.A0(new_new_n696_), .A1(new_new_n695_), .B0(new_new_n691_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n175_), .B(new_new_n116_), .Y(new_new_n698_));
  OAI210     g676(.A0(new_new_n698_), .A1(new_new_n681_), .B0(i_2_), .Y(new_new_n699_));
  INV        g677(.A(new_new_n158_), .Y(new_new_n700_));
  NO3        g678(.A(new_new_n557_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n701_));
  AOI210     g679(.A0(new_new_n700_), .A1(new_new_n81_), .B0(new_new_n701_), .Y(new_new_n702_));
  AOI210     g680(.A0(new_new_n702_), .A1(new_new_n699_), .B0(new_new_n178_), .Y(new_new_n703_));
  OA210      g681(.A0(new_new_n558_), .A1(new_new_n117_), .B0(i_13_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n184_), .B(new_new_n187_), .Y(new_new_n705_));
  NA2        g683(.A(new_new_n140_), .B(new_new_n535_), .Y(new_new_n706_));
  AOI210     g684(.A0(new_new_n706_), .A1(new_new_n705_), .B0(new_new_n329_), .Y(new_new_n707_));
  NA4        g685(.A(i_2_), .B(new_new_n276_), .C(new_new_n115_), .D(new_new_n42_), .Y(new_new_n708_));
  INV        g686(.A(new_new_n708_), .Y(new_new_n709_));
  NO4        g687(.A(new_new_n709_), .B(new_new_n707_), .C(new_new_n704_), .D(new_new_n703_), .Y(new_new_n710_));
  NA2        g688(.A(new_new_n514_), .B(new_new_n28_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n680_), .B(new_new_n255_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n712_), .B(new_new_n711_), .Y(new_new_n713_));
  NO2        g691(.A(new_new_n61_), .B(i_12_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n714_), .B(new_new_n117_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n715_), .B(new_new_n535_), .Y(new_new_n716_));
  AOI220     g694(.A0(new_new_n716_), .A1(new_new_n36_), .B0(new_new_n713_), .B1(new_new_n46_), .Y(new_new_n717_));
  NA4        g695(.A(new_new_n717_), .B(new_new_n710_), .C(new_new_n697_), .D(new_new_n687_), .Y(mai6));
  OAI210     g696(.A0(new_new_n25_), .A1(new_new_n959_), .B0(new_new_n668_), .Y(new_new_n719_));
  NA4        g697(.A(new_new_n347_), .B(i_8_), .C(new_new_n66_), .D(new_new_n93_), .Y(new_new_n720_));
  INV        g698(.A(new_new_n720_), .Y(new_new_n721_));
  NO2        g699(.A(new_new_n204_), .B(new_new_n432_), .Y(new_new_n722_));
  NO2        g700(.A(i_11_), .B(i_9_), .Y(new_new_n723_));
  NO3        g701(.A(new_new_n722_), .B(new_new_n721_), .C(new_new_n296_), .Y(new_new_n724_));
  AO210      g702(.A0(new_new_n724_), .A1(new_new_n719_), .B0(i_12_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n330_), .B(new_new_n302_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n521_), .B(new_new_n62_), .Y(new_new_n727_));
  NA2        g705(.A(new_new_n616_), .B(new_new_n66_), .Y(new_new_n728_));
  NA4        g706(.A(new_new_n563_), .B(new_new_n728_), .C(new_new_n727_), .D(new_new_n726_), .Y(new_new_n729_));
  INV        g707(.A(new_new_n181_), .Y(new_new_n730_));
  AOI220     g708(.A0(new_new_n730_), .A1(new_new_n723_), .B0(new_new_n729_), .B1(new_new_n68_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n947_), .B(new_new_n714_), .Y(new_new_n732_));
  AOI210     g710(.A0(new_new_n732_), .A1(new_new_n462_), .B0(new_new_n170_), .Y(new_new_n733_));
  NO2        g711(.A(new_new_n32_), .B(i_11_), .Y(new_new_n734_));
  NA3        g712(.A(new_new_n734_), .B(new_new_n422_), .C(new_new_n347_), .Y(new_new_n735_));
  OAI210     g713(.A0(new_new_n616_), .A1(new_new_n503_), .B0(new_new_n502_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n736_), .B(new_new_n735_), .Y(new_new_n737_));
  OR2        g715(.A(new_new_n737_), .B(new_new_n733_), .Y(new_new_n738_));
  NO2        g716(.A(i_11_), .B(i_2_), .Y(new_new_n739_));
  NA2        g717(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n740_));
  OAI210     g718(.A0(new_new_n740_), .A1(new_new_n362_), .B0(new_new_n315_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n741_), .B(new_new_n739_), .Y(new_new_n742_));
  NA3        g720(.A(new_new_n308_), .B(new_new_n234_), .C(i_7_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n400_), .B(new_new_n136_), .Y(new_new_n744_));
  AO210      g722(.A0(new_new_n437_), .A1(new_new_n684_), .B0(new_new_n36_), .Y(new_new_n745_));
  NA4        g723(.A(new_new_n745_), .B(new_new_n744_), .C(new_new_n743_), .D(new_new_n742_), .Y(new_new_n746_));
  AOI220     g724(.A0(new_new_n952_), .A1(new_new_n502_), .B0(new_new_n722_), .B1(new_new_n648_), .Y(new_new_n747_));
  NA3        g725(.A(new_new_n329_), .B(new_new_n219_), .C(new_new_n136_), .Y(new_new_n748_));
  NA3        g726(.A(new_new_n748_), .B(new_new_n747_), .C(new_new_n541_), .Y(new_new_n749_));
  AO210      g727(.A0(i_4_), .A1(new_new_n46_), .B0(new_new_n80_), .Y(new_new_n750_));
  NA3        g728(.A(new_new_n750_), .B(new_new_n428_), .C(new_new_n202_), .Y(new_new_n751_));
  AOI210     g729(.A0(new_new_n400_), .A1(new_new_n398_), .B0(new_new_n501_), .Y(new_new_n752_));
  OAI210     g730(.A0(new_new_n954_), .A1(new_new_n104_), .B0(new_new_n361_), .Y(new_new_n753_));
  NA2        g731(.A(i_0_), .B(new_new_n526_), .Y(new_new_n754_));
  NA3        g732(.A(new_new_n754_), .B(new_new_n295_), .C(i_7_), .Y(new_new_n755_));
  NA4        g733(.A(new_new_n755_), .B(new_new_n753_), .C(new_new_n752_), .D(new_new_n751_), .Y(new_new_n756_));
  NO4        g734(.A(new_new_n756_), .B(new_new_n749_), .C(new_new_n746_), .D(new_new_n738_), .Y(new_new_n757_));
  NA4        g735(.A(new_new_n757_), .B(new_new_n731_), .C(new_new_n725_), .D(new_new_n337_), .Y(mai3));
  NA2        g736(.A(i_6_), .B(i_7_), .Y(new_new_n759_));
  NO2        g737(.A(new_new_n759_), .B(i_0_), .Y(new_new_n760_));
  NO2        g738(.A(i_11_), .B(new_new_n218_), .Y(new_new_n761_));
  OAI210     g739(.A0(new_new_n760_), .A1(new_new_n266_), .B0(new_new_n761_), .Y(new_new_n762_));
  NO2        g740(.A(new_new_n762_), .B(new_new_n178_), .Y(new_new_n763_));
  AN2        g741(.A(new_new_n763_), .B(new_new_n160_), .Y(new_new_n764_));
  NA3        g742(.A(new_new_n748_), .B(new_new_n541_), .C(new_new_n328_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n765_), .B(new_new_n39_), .Y(new_new_n766_));
  NO3        g744(.A(new_new_n568_), .B(new_new_n407_), .C(new_new_n120_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n363_), .B(new_new_n45_), .Y(new_new_n768_));
  AN2        g746(.A(new_new_n405_), .B(new_new_n54_), .Y(new_new_n769_));
  NO2        g747(.A(new_new_n769_), .B(new_new_n767_), .Y(new_new_n770_));
  AOI210     g748(.A0(new_new_n770_), .A1(new_new_n766_), .B0(new_new_n48_), .Y(new_new_n771_));
  NO4        g749(.A(new_new_n333_), .B(new_new_n340_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n640_), .B(new_new_n609_), .Y(new_new_n773_));
  NA2        g751(.A(i_0_), .B(i_5_), .Y(new_new_n774_));
  OAI220     g752(.A0(new_new_n774_), .A1(new_new_n773_), .B0(new_new_n948_), .B1(new_new_n62_), .Y(new_new_n775_));
  NOi21      g753(.An(i_5_), .B(i_9_), .Y(new_new_n776_));
  NA2        g754(.A(new_new_n776_), .B(new_new_n396_), .Y(new_new_n777_));
  NO3        g755(.A(new_new_n364_), .B(new_new_n246_), .C(new_new_n68_), .Y(new_new_n778_));
  NO2        g756(.A(new_new_n161_), .B(new_new_n137_), .Y(new_new_n779_));
  AOI210     g757(.A0(new_new_n779_), .A1(new_new_n223_), .B0(new_new_n778_), .Y(new_new_n780_));
  OAI220     g758(.A0(new_new_n780_), .A1(new_new_n166_), .B0(new_new_n543_), .B1(new_new_n777_), .Y(new_new_n781_));
  NO4        g759(.A(new_new_n781_), .B(new_new_n775_), .C(new_new_n771_), .D(new_new_n764_), .Y(new_new_n782_));
  INV        g760(.A(new_new_n282_), .Y(new_new_n783_));
  NAi21      g761(.An(new_new_n150_), .B(i_5_), .Y(new_new_n784_));
  OAI220     g762(.A0(new_new_n784_), .A1(i_0_), .B0(new_new_n783_), .B1(new_new_n355_), .Y(new_new_n785_));
  INV        g763(.A(new_new_n785_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n511_), .B(i_0_), .Y(new_new_n787_));
  NO3        g765(.A(new_new_n787_), .B(new_new_n342_), .C(new_new_n81_), .Y(new_new_n788_));
  NO4        g766(.A(i_5_), .B(i_12_), .C(new_new_n368_), .D(new_new_n362_), .Y(new_new_n789_));
  AOI210     g767(.A0(new_new_n789_), .A1(i_11_), .B0(new_new_n788_), .Y(new_new_n790_));
  NA2        g768(.A(new_new_n680_), .B(new_new_n296_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n428_), .B(new_new_n57_), .Y(new_new_n792_));
  NO2        g770(.A(new_new_n792_), .B(new_new_n791_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n232_), .B(new_new_n141_), .Y(new_new_n794_));
  INV        g772(.A(new_new_n478_), .Y(new_new_n795_));
  NO4        g773(.A(new_new_n107_), .B(new_new_n57_), .C(new_new_n605_), .D(i_5_), .Y(new_new_n796_));
  AO220      g774(.A0(new_new_n796_), .A1(new_new_n795_), .B0(new_new_n794_), .B1(i_6_), .Y(new_new_n797_));
  AOI210     g775(.A0(i_0_), .A1(new_new_n90_), .B0(new_new_n170_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n506_), .B(i_4_), .Y(new_new_n799_));
  NA2        g777(.A(new_new_n173_), .B(new_new_n187_), .Y(new_new_n800_));
  OAI220     g778(.A0(new_new_n800_), .A1(new_new_n791_), .B0(new_new_n799_), .B1(new_new_n798_), .Y(new_new_n801_));
  NO3        g779(.A(new_new_n801_), .B(new_new_n797_), .C(new_new_n793_), .Y(new_new_n802_));
  NA3        g780(.A(new_new_n802_), .B(new_new_n790_), .C(new_new_n786_), .Y(new_new_n803_));
  NA2        g781(.A(i_11_), .B(i_9_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n48_), .B(i_7_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n351_), .B(new_new_n165_), .Y(new_new_n806_));
  NAi31      g784(.An(new_new_n243_), .B(new_new_n806_), .C(new_new_n148_), .Y(new_new_n807_));
  NO2        g785(.A(new_new_n161_), .B(i_0_), .Y(new_new_n808_));
  NA2        g786(.A(new_new_n422_), .B(new_new_n214_), .Y(new_new_n809_));
  OAI220     g787(.A0(i_12_), .A1(new_new_n777_), .B0(new_new_n809_), .B1(new_new_n161_), .Y(new_new_n810_));
  NO2        g788(.A(new_new_n810_), .B(new_new_n807_), .Y(new_new_n811_));
  AOI210     g789(.A0(new_new_n399_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n812_));
  NA2        g790(.A(new_new_n157_), .B(new_new_n95_), .Y(new_new_n813_));
  NOi32      g791(.An(new_new_n812_), .Bn(new_new_n173_), .C(new_new_n813_), .Y(new_new_n814_));
  NO2        g792(.A(new_new_n955_), .B(new_new_n768_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n815_), .B(new_new_n814_), .Y(new_new_n816_));
  NOi21      g794(.An(i_7_), .B(i_5_), .Y(new_new_n817_));
  NOi21      g795(.An(new_new_n817_), .B(new_new_n659_), .Y(new_new_n818_));
  NA3        g796(.A(new_new_n818_), .B(new_new_n341_), .C(i_6_), .Y(new_new_n819_));
  OA210      g797(.A0(new_new_n813_), .A1(new_new_n462_), .B0(new_new_n819_), .Y(new_new_n820_));
  NO3        g798(.A(new_new_n357_), .B(new_new_n317_), .C(new_new_n313_), .Y(new_new_n821_));
  NO2        g799(.A(new_new_n240_), .B(new_new_n287_), .Y(new_new_n822_));
  INV        g800(.A(new_new_n821_), .Y(new_new_n823_));
  NA4        g801(.A(new_new_n823_), .B(new_new_n820_), .C(new_new_n816_), .D(new_new_n811_), .Y(new_new_n824_));
  AN2        g802(.A(new_new_n300_), .B(new_new_n296_), .Y(new_new_n825_));
  AN2        g803(.A(new_new_n825_), .B(new_new_n779_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n826_), .B(i_10_), .Y(new_new_n827_));
  OA210      g805(.A0(new_new_n422_), .A1(new_new_n206_), .B0(new_new_n421_), .Y(new_new_n828_));
  NA3        g806(.A(new_new_n421_), .B(new_new_n363_), .C(new_new_n45_), .Y(new_new_n829_));
  OAI210     g807(.A0(new_new_n784_), .A1(new_new_n422_), .B0(new_new_n829_), .Y(new_new_n830_));
  INV        g808(.A(new_new_n172_), .Y(new_new_n831_));
  AOI220     g809(.A0(new_new_n831_), .A1(new_new_n422_), .B0(new_new_n830_), .B1(new_new_n68_), .Y(new_new_n832_));
  NA3        g810(.A(new_new_n740_), .B(new_new_n339_), .C(new_new_n578_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n85_), .B(new_new_n44_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n70_), .B(new_new_n682_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n835_), .B(new_new_n834_), .Y(new_new_n836_));
  AOI210     g814(.A0(new_new_n836_), .A1(new_new_n833_), .B0(new_new_n47_), .Y(new_new_n837_));
  NO3        g815(.A(i_5_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n838_));
  NO2        g816(.A(new_new_n485_), .B(new_new_n838_), .Y(new_new_n839_));
  NAi21      g817(.An(i_9_), .B(i_5_), .Y(new_new_n840_));
  NO2        g818(.A(new_new_n840_), .B(new_new_n357_), .Y(new_new_n841_));
  NO2        g819(.A(new_new_n537_), .B(new_new_n97_), .Y(new_new_n842_));
  AOI220     g820(.A0(new_new_n842_), .A1(i_0_), .B0(new_new_n841_), .B1(new_new_n558_), .Y(new_new_n843_));
  OAI220     g821(.A0(new_new_n843_), .A1(new_new_n78_), .B0(new_new_n839_), .B1(new_new_n158_), .Y(new_new_n844_));
  NO3        g822(.A(new_new_n844_), .B(new_new_n837_), .C(new_new_n464_), .Y(new_new_n845_));
  NA3        g823(.A(new_new_n845_), .B(new_new_n832_), .C(new_new_n827_), .Y(new_new_n846_));
  NO3        g824(.A(new_new_n846_), .B(new_new_n824_), .C(new_new_n803_), .Y(new_new_n847_));
  INV        g825(.A(new_new_n659_), .Y(new_new_n848_));
  NO3        g826(.A(new_new_n97_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n849_));
  AO220      g827(.A0(new_new_n849_), .A1(new_new_n44_), .B0(new_new_n848_), .B1(new_new_n160_), .Y(new_new_n850_));
  AOI210     g828(.A0(new_new_n727_), .A1(new_new_n618_), .B0(new_new_n813_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n850_), .A1(new_new_n307_), .B0(new_new_n851_), .Y(new_new_n852_));
  NA3        g830(.A(new_new_n135_), .B(new_new_n609_), .C(new_new_n68_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n736_), .B(new_new_n357_), .Y(new_new_n854_));
  NA3        g832(.A(new_new_n760_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n761_), .B(i_9_), .Y(new_new_n856_));
  AOI210     g834(.A0(new_new_n855_), .A1(new_new_n441_), .B0(new_new_n856_), .Y(new_new_n857_));
  NO2        g835(.A(new_new_n857_), .B(new_new_n854_), .Y(new_new_n858_));
  NA3        g836(.A(new_new_n858_), .B(new_new_n853_), .C(new_new_n852_), .Y(new_new_n859_));
  AOI210     g837(.A0(new_new_n274_), .A1(new_new_n150_), .B0(new_new_n957_), .Y(new_new_n860_));
  NA3        g838(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n861_));
  NA2        g839(.A(new_new_n805_), .B(new_new_n433_), .Y(new_new_n862_));
  AOI210     g840(.A0(new_new_n861_), .A1(new_new_n150_), .B0(new_new_n862_), .Y(new_new_n863_));
  NO2        g841(.A(new_new_n863_), .B(new_new_n860_), .Y(new_new_n864_));
  NO3        g842(.A(new_new_n194_), .B(new_new_n340_), .C(i_0_), .Y(new_new_n865_));
  OAI210     g843(.A0(new_new_n865_), .A1(new_new_n71_), .B0(i_13_), .Y(new_new_n866_));
  INV        g844(.A(new_new_n202_), .Y(new_new_n867_));
  OAI220     g845(.A0(new_new_n473_), .A1(new_new_n128_), .B0(i_12_), .B1(new_new_n552_), .Y(new_new_n868_));
  NA3        g846(.A(new_new_n868_), .B(i_7_), .C(new_new_n867_), .Y(new_new_n869_));
  NA3        g847(.A(new_new_n869_), .B(new_new_n866_), .C(new_new_n864_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n222_), .B(new_new_n85_), .Y(new_new_n871_));
  AOI210     g849(.A0(new_new_n871_), .A1(new_new_n848_), .B0(new_new_n101_), .Y(new_new_n872_));
  AOI220     g850(.A0(new_new_n817_), .A1(new_new_n433_), .B0(new_new_n760_), .B1(new_new_n151_), .Y(new_new_n873_));
  NA2        g851(.A(new_new_n308_), .B(new_new_n162_), .Y(new_new_n874_));
  OA220      g852(.A0(new_new_n874_), .A1(new_new_n873_), .B0(new_new_n872_), .B1(i_5_), .Y(new_new_n875_));
  AOI210     g853(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n161_), .Y(new_new_n876_));
  NA2        g854(.A(new_new_n876_), .B(new_new_n828_), .Y(new_new_n877_));
  NA2        g855(.A(new_new_n549_), .B(new_new_n170_), .Y(new_new_n878_));
  NA2        g856(.A(new_new_n878_), .B(new_new_n484_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n768_), .B(new_new_n53_), .C(new_new_n48_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n431_), .B(new_new_n419_), .Y(new_new_n881_));
  NO3        g859(.A(new_new_n881_), .B(new_new_n880_), .C(new_new_n879_), .Y(new_new_n882_));
  NA3        g860(.A(new_new_n347_), .B(new_new_n301_), .C(new_new_n205_), .Y(new_new_n883_));
  INV        g861(.A(new_new_n883_), .Y(new_new_n884_));
  NOi31      g862(.An(new_new_n346_), .B(i_11_), .C(new_new_n220_), .Y(new_new_n885_));
  NO3        g863(.A(new_new_n804_), .B(new_new_n202_), .C(new_new_n175_), .Y(new_new_n886_));
  NO3        g864(.A(new_new_n886_), .B(new_new_n885_), .C(new_new_n884_), .Y(new_new_n887_));
  NA4        g865(.A(new_new_n887_), .B(new_new_n882_), .C(new_new_n877_), .D(new_new_n875_), .Y(new_new_n888_));
  INV        g866(.A(new_new_n551_), .Y(new_new_n889_));
  NO3        g867(.A(new_new_n889_), .B(new_new_n497_), .C(i_7_), .Y(new_new_n890_));
  NO2        g868(.A(new_new_n78_), .B(i_5_), .Y(new_new_n891_));
  NA3        g869(.A(new_new_n761_), .B(new_new_n102_), .C(new_new_n115_), .Y(new_new_n892_));
  INV        g870(.A(new_new_n892_), .Y(new_new_n893_));
  AOI210     g871(.A0(new_new_n893_), .A1(new_new_n891_), .B0(new_new_n890_), .Y(new_new_n894_));
  NA3        g872(.A(new_new_n276_), .B(i_5_), .C(new_new_n178_), .Y(new_new_n895_));
  NO4        g873(.A(new_new_n220_), .B(new_new_n194_), .C(i_0_), .D(i_12_), .Y(new_new_n896_));
  AOI220     g874(.A0(new_new_n896_), .A1(new_new_n945_), .B0(new_new_n721_), .B1(new_new_n162_), .Y(new_new_n897_));
  BUFFER     g875(.A(new_new_n141_), .Y(new_new_n898_));
  NO4        g876(.A(new_new_n898_), .B(i_12_), .C(new_new_n586_), .D(new_new_n120_), .Y(new_new_n899_));
  NA2        g877(.A(new_new_n899_), .B(new_new_n202_), .Y(new_new_n900_));
  NA2        g878(.A(new_new_n817_), .B(new_new_n418_), .Y(new_new_n901_));
  OAI210     g879(.A0(i_6_), .A1(new_new_n895_), .B0(new_new_n901_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n902_), .B(new_new_n808_), .Y(new_new_n903_));
  NA4        g881(.A(new_new_n903_), .B(new_new_n900_), .C(new_new_n897_), .D(new_new_n894_), .Y(new_new_n904_));
  NO4        g882(.A(new_new_n904_), .B(new_new_n888_), .C(new_new_n870_), .D(new_new_n859_), .Y(new_new_n905_));
  OAI210     g883(.A0(new_new_n739_), .A1(new_new_n734_), .B0(new_new_n37_), .Y(new_new_n906_));
  NA3        g884(.A(new_new_n812_), .B(new_new_n324_), .C(i_5_), .Y(new_new_n907_));
  NA3        g885(.A(new_new_n907_), .B(new_new_n906_), .C(new_new_n547_), .Y(new_new_n908_));
  NA2        g886(.A(new_new_n908_), .B(new_new_n191_), .Y(new_new_n909_));
  NA2        g887(.A(new_new_n171_), .B(new_new_n173_), .Y(new_new_n910_));
  OAI210     g888(.A0(new_new_n551_), .A1(new_new_n549_), .B0(new_new_n286_), .Y(new_new_n911_));
  INV        g889(.A(new_new_n583_), .Y(new_new_n912_));
  NA3        g890(.A(new_new_n912_), .B(new_new_n911_), .C(new_new_n910_), .Y(new_new_n913_));
  NO2        g891(.A(new_new_n411_), .B(new_new_n246_), .Y(new_new_n914_));
  NO2        g892(.A(new_new_n914_), .B(new_new_n789_), .Y(new_new_n915_));
  INV        g893(.A(new_new_n915_), .Y(new_new_n916_));
  AOI210     g894(.A0(new_new_n913_), .A1(new_new_n48_), .B0(new_new_n916_), .Y(new_new_n917_));
  AOI210     g895(.A0(new_new_n917_), .A1(new_new_n909_), .B0(new_new_n68_), .Y(new_new_n918_));
  NO2        g896(.A(new_new_n504_), .B(new_new_n336_), .Y(new_new_n919_));
  NO2        g897(.A(new_new_n919_), .B(new_new_n688_), .Y(new_new_n920_));
  AOI210     g898(.A0(new_new_n876_), .A1(new_new_n805_), .B0(new_new_n818_), .Y(new_new_n921_));
  NO2        g899(.A(new_new_n921_), .B(new_new_n610_), .Y(new_new_n922_));
  INV        g900(.A(new_new_n56_), .Y(new_new_n923_));
  NA2        g901(.A(new_new_n923_), .B(new_new_n71_), .Y(new_new_n924_));
  NO2        g902(.A(new_new_n924_), .B(new_new_n218_), .Y(new_new_n925_));
  NO2        g903(.A(new_new_n925_), .B(new_new_n922_), .Y(new_new_n926_));
  OAI210     g904(.A0(new_new_n248_), .A1(new_new_n146_), .B0(new_new_n81_), .Y(new_new_n927_));
  NO2        g905(.A(new_new_n927_), .B(i_11_), .Y(new_new_n928_));
  OAI210     g906(.A0(new_new_n946_), .A1(new_new_n812_), .B0(new_new_n191_), .Y(new_new_n929_));
  NA2        g907(.A(i_0_), .B(i_5_), .Y(new_new_n930_));
  AOI210     g908(.A0(new_new_n929_), .A1(new_new_n705_), .B0(new_new_n930_), .Y(new_new_n931_));
  NO3        g909(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n932_));
  OAI210     g910(.A0(new_new_n822_), .A1(new_new_n953_), .B0(new_new_n932_), .Y(new_new_n933_));
  NO2        g911(.A(new_new_n933_), .B(new_new_n659_), .Y(new_new_n934_));
  NO4        g912(.A(new_new_n840_), .B(new_new_n424_), .C(new_new_n231_), .D(new_new_n230_), .Y(new_new_n935_));
  NO2        g913(.A(new_new_n935_), .B(new_new_n501_), .Y(new_new_n936_));
  INV        g914(.A(new_new_n318_), .Y(new_new_n937_));
  AOI210     g915(.A0(new_new_n937_), .A1(new_new_n936_), .B0(new_new_n40_), .Y(new_new_n938_));
  NO4        g916(.A(new_new_n938_), .B(new_new_n934_), .C(new_new_n931_), .D(new_new_n928_), .Y(new_new_n939_));
  OAI210     g917(.A0(new_new_n926_), .A1(i_4_), .B0(new_new_n939_), .Y(new_new_n940_));
  NO3        g918(.A(new_new_n940_), .B(new_new_n920_), .C(new_new_n918_), .Y(new_new_n941_));
  NA4        g919(.A(new_new_n941_), .B(new_new_n905_), .C(new_new_n847_), .D(new_new_n782_), .Y(mai4));
  INV        g920(.A(new_new_n222_), .Y(new_new_n945_));
  INV        g921(.A(i_12_), .Y(new_new_n946_));
  INV        g922(.A(i_9_), .Y(new_new_n947_));
  INV        g923(.A(new_new_n772_), .Y(new_new_n948_));
  INV        g924(.A(new_new_n120_), .Y(new_new_n949_));
  INV        g925(.A(i_1_), .Y(new_new_n950_));
  INV        g926(.A(new_new_n133_), .Y(new_new_n951_));
  INV        g927(.A(i_11_), .Y(new_new_n952_));
  INV        g928(.A(i_5_), .Y(new_new_n953_));
  INV        g929(.A(new_new_n548_), .Y(new_new_n954_));
  INV        g930(.A(new_new_n296_), .Y(new_new_n955_));
  INV        g931(.A(new_new_n190_), .Y(new_new_n956_));
  INV        g932(.A(new_new_n296_), .Y(new_new_n957_));
  INV        g933(.A(i_1_), .Y(new_new_n958_));
  INV        g934(.A(i_9_), .Y(new_new_n959_));
endmodule


