//Benchmark atmr_max1024_476_0.25

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  INV        o004(.A(ori_ori_n19_), .Y(ori_ori_n21_));
  NA2        o005(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n22_));
  INV        o006(.A(x5), .Y(ori_ori_n23_));
  NA2        o007(.A(x4), .B(x2), .Y(ori_ori_n24_));
  INV        o008(.A(ori_ori_n22_), .Y(ori_ori_n25_));
  NO2        o009(.A(x4), .B(x3), .Y(ori_ori_n26_));
  INV        o010(.A(ori_ori_n26_), .Y(ori_ori_n27_));
  NOi21      o011(.An(ori_ori_n21_), .B(ori_ori_n25_), .Y(ori00));
  NO2        o012(.A(x1), .B(x0), .Y(ori_ori_n29_));
  INV        o013(.A(x6), .Y(ori_ori_n30_));
  NO2        o014(.A(ori_ori_n30_), .B(ori_ori_n23_), .Y(ori_ori_n31_));
  NA2        o015(.A(x4), .B(x3), .Y(ori_ori_n32_));
  NO2        o016(.A(ori_ori_n21_), .B(ori_ori_n32_), .Y(ori_ori_n33_));
  NO2        o017(.A(x2), .B(x0), .Y(ori_ori_n34_));
  INV        o018(.A(x3), .Y(ori_ori_n35_));
  NO2        o019(.A(ori_ori_n35_), .B(ori_ori_n18_), .Y(ori_ori_n36_));
  INV        o020(.A(ori_ori_n36_), .Y(ori_ori_n37_));
  NO2        o021(.A(ori_ori_n31_), .B(x4), .Y(ori_ori_n38_));
  OAI210     o022(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n34_), .Y(ori_ori_n39_));
  INV        o023(.A(x4), .Y(ori_ori_n40_));
  NO2        o024(.A(ori_ori_n40_), .B(ori_ori_n17_), .Y(ori_ori_n41_));
  NA2        o025(.A(ori_ori_n41_), .B(x2), .Y(ori_ori_n42_));
  OAI210     o026(.A0(ori_ori_n42_), .A1(ori_ori_n20_), .B0(ori_ori_n39_), .Y(ori_ori_n43_));
  INV        o027(.A(ori_ori_n29_), .Y(ori_ori_n44_));
  INV        o028(.A(x2), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n45_), .B(ori_ori_n17_), .Y(ori_ori_n46_));
  NA2        o030(.A(ori_ori_n35_), .B(ori_ori_n18_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(ori_ori_n46_), .Y(ori_ori_n48_));
  OAI210     o032(.A0(ori_ori_n44_), .A1(ori_ori_n27_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  NO3        o033(.A(ori_ori_n49_), .B(ori_ori_n43_), .C(ori_ori_n33_), .Y(ori01));
  INV        o034(.A(x7), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n35_), .B(x1), .Y(ori_ori_n52_));
  INV        o036(.A(x6), .Y(ori_ori_n53_));
  NO2        o037(.A(ori_ori_n52_), .B(x5), .Y(ori_ori_n54_));
  OAI210     o038(.A0(ori_ori_n36_), .A1(ori_ori_n23_), .B0(ori_ori_n45_), .Y(ori_ori_n55_));
  OAI210     o039(.A0(ori_ori_n47_), .A1(ori_ori_n20_), .B0(ori_ori_n55_), .Y(ori_ori_n56_));
  INV        o040(.A(ori_ori_n56_), .Y(ori_ori_n57_));
  NA2        o041(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n58_));
  NA2        o042(.A(ori_ori_n40_), .B(x2), .Y(ori_ori_n59_));
  OAI210     o043(.A0(ori_ori_n59_), .A1(ori_ori_n47_), .B0(x0), .Y(ori_ori_n60_));
  NA2        o044(.A(x5), .B(x3), .Y(ori_ori_n61_));
  INV        o045(.A(x6), .Y(ori_ori_n62_));
  NO3        o046(.A(ori_ori_n61_), .B(ori_ori_n53_), .C(ori_ori_n45_), .Y(ori_ori_n63_));
  NAi21      o047(.An(x4), .B(x3), .Y(ori_ori_n64_));
  INV        o048(.A(ori_ori_n64_), .Y(ori_ori_n65_));
  NO2        o049(.A(x4), .B(x2), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n64_), .B(ori_ori_n18_), .Y(ori_ori_n67_));
  NO3        o051(.A(ori_ori_n67_), .B(ori_ori_n63_), .C(ori_ori_n60_), .Y(ori_ori_n68_));
  NA2        o052(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n69_));
  NO2        o053(.A(ori_ori_n69_), .B(ori_ori_n23_), .Y(ori_ori_n70_));
  INV        o054(.A(x8), .Y(ori_ori_n71_));
  NA2        o055(.A(x2), .B(x1), .Y(ori_ori_n72_));
  AOI210     o056(.A0(ori_ori_n47_), .A1(ori_ori_n23_), .B0(ori_ori_n45_), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n37_), .A1(ori_ori_n31_), .B0(ori_ori_n40_), .Y(ori_ori_n74_));
  NO2        o058(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  NA2        o059(.A(x4), .B(ori_ori_n35_), .Y(ori_ori_n76_));
  NO2        o060(.A(ori_ori_n40_), .B(ori_ori_n45_), .Y(ori_ori_n77_));
  NO2        o061(.A(ori_ori_n76_), .B(x1), .Y(ori_ori_n78_));
  NA2        o062(.A(ori_ori_n45_), .B(x1), .Y(ori_ori_n79_));
  OAI210     o063(.A0(ori_ori_n79_), .A1(ori_ori_n32_), .B0(ori_ori_n17_), .Y(ori_ori_n80_));
  NO3        o064(.A(ori_ori_n80_), .B(ori_ori_n78_), .C(ori_ori_n75_), .Y(ori_ori_n81_));
  AO210      o065(.A0(ori_ori_n68_), .A1(ori_ori_n58_), .B0(ori_ori_n81_), .Y(ori02));
  BUFFER     o066(.A(x0), .Y(ori_ori_n83_));
  INV        o067(.A(ori_ori_n83_), .Y(ori_ori_n84_));
  NO2        o068(.A(x4), .B(x1), .Y(ori_ori_n85_));
  NA2        o069(.A(ori_ori_n85_), .B(x2), .Y(ori_ori_n86_));
  NOi21      o070(.An(x0), .B(x1), .Y(ori_ori_n87_));
  NOi21      o071(.An(x0), .B(x4), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n86_), .B(ori_ori_n61_), .Y(ori_ori_n89_));
  NO2        o073(.A(x5), .B(ori_ori_n40_), .Y(ori_ori_n90_));
  NA2        o074(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n91_));
  AOI210     o075(.A0(ori_ori_n91_), .A1(ori_ori_n79_), .B0(x3), .Y(ori_ori_n92_));
  OAI210     o076(.A0(ori_ori_n92_), .A1(ori_ori_n29_), .B0(ori_ori_n90_), .Y(ori_ori_n93_));
  NAi21      o077(.An(x0), .B(x4), .Y(ori_ori_n94_));
  NO2        o078(.A(x7), .B(x0), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n66_), .B(ori_ori_n77_), .Y(ori_ori_n96_));
  NO2        o080(.A(ori_ori_n96_), .B(x3), .Y(ori_ori_n97_));
  NA2        o081(.A(ori_ori_n95_), .B(ori_ori_n97_), .Y(ori_ori_n98_));
  NA2        o082(.A(x5), .B(x0), .Y(ori_ori_n99_));
  NO2        o083(.A(ori_ori_n40_), .B(x2), .Y(ori_ori_n100_));
  NA3        o084(.A(ori_ori_n98_), .B(ori_ori_n93_), .C(ori_ori_n30_), .Y(ori_ori_n101_));
  NO2        o085(.A(ori_ori_n101_), .B(ori_ori_n89_), .Y(ori_ori_n102_));
  NO3        o086(.A(ori_ori_n61_), .B(ori_ori_n59_), .C(ori_ori_n22_), .Y(ori_ori_n103_));
  NO2        o087(.A(ori_ori_n24_), .B(ori_ori_n23_), .Y(ori_ori_n104_));
  NO2        o088(.A(ori_ori_n76_), .B(x5), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n106_));
  INV        o090(.A(x7), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n107_), .B(ori_ori_n18_), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n108_), .B(ori_ori_n106_), .Y(ori_ori_n109_));
  NO2        o093(.A(ori_ori_n23_), .B(x4), .Y(ori_ori_n110_));
  NO2        o094(.A(ori_ori_n110_), .B(ori_ori_n88_), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n111_), .B(ori_ori_n109_), .Y(ori_ori_n112_));
  NA2        o096(.A(x5), .B(x1), .Y(ori_ori_n113_));
  INV        o097(.A(ori_ori_n113_), .Y(ori_ori_n114_));
  AOI210     o098(.A0(ori_ori_n114_), .A1(ori_ori_n88_), .B0(ori_ori_n30_), .Y(ori_ori_n115_));
  BUFFER     o099(.A(x2), .Y(ori_ori_n116_));
  NO2        o100(.A(ori_ori_n116_), .B(ori_ori_n40_), .Y(ori_ori_n117_));
  NA2        o101(.A(ori_ori_n117_), .B(ori_ori_n54_), .Y(ori_ori_n118_));
  NA2        o102(.A(ori_ori_n118_), .B(ori_ori_n115_), .Y(ori_ori_n119_));
  NO3        o103(.A(ori_ori_n119_), .B(ori_ori_n112_), .C(ori_ori_n103_), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n120_), .B(ori_ori_n102_), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n99_), .B(ori_ori_n96_), .Y(ori_ori_n122_));
  NA2        o106(.A(ori_ori_n23_), .B(ori_ori_n18_), .Y(ori_ori_n123_));
  NA2        o107(.A(ori_ori_n23_), .B(ori_ori_n17_), .Y(ori_ori_n124_));
  NA3        o108(.A(ori_ori_n124_), .B(ori_ori_n123_), .C(ori_ori_n22_), .Y(ori_ori_n125_));
  AN2        o109(.A(ori_ori_n125_), .B(ori_ori_n100_), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n107_), .B(ori_ori_n23_), .Y(ori_ori_n127_));
  NA2        o111(.A(x2), .B(x0), .Y(ori_ori_n128_));
  NA2        o112(.A(x4), .B(x1), .Y(ori_ori_n129_));
  NAi21      o113(.An(ori_ori_n85_), .B(ori_ori_n129_), .Y(ori_ori_n130_));
  NOi31      o114(.An(ori_ori_n130_), .B(ori_ori_n110_), .C(ori_ori_n128_), .Y(ori_ori_n131_));
  NO3        o115(.A(ori_ori_n131_), .B(ori_ori_n126_), .C(ori_ori_n122_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n132_), .B(ori_ori_n35_), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n125_), .B(ori_ori_n59_), .Y(ori_ori_n134_));
  INV        o118(.A(ori_ori_n90_), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n79_), .B(ori_ori_n17_), .Y(ori_ori_n136_));
  NA3        o120(.A(ori_ori_n130_), .B(ori_ori_n135_), .C(ori_ori_n34_), .Y(ori_ori_n137_));
  OAI210     o121(.A0(ori_ori_n124_), .A1(ori_ori_n96_), .B0(ori_ori_n137_), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n138_), .B(ori_ori_n134_), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n139_), .B(x3), .Y(ori_ori_n140_));
  NO3        o124(.A(ori_ori_n140_), .B(ori_ori_n133_), .C(ori_ori_n121_), .Y(ori03));
  NO2        o125(.A(ori_ori_n40_), .B(x3), .Y(ori_ori_n142_));
  NA2        o126(.A(x6), .B(ori_ori_n23_), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n143_), .B(x4), .Y(ori_ori_n144_));
  NO2        o128(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n145_));
  NA2        o129(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n146_));
  NO2        o130(.A(x5), .B(x1), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n146_), .B(ori_ori_n123_), .Y(ori_ori_n148_));
  NO3        o132(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n149_));
  NO2        o133(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n150_), .B(x6), .Y(ori_ori_n151_));
  NOi21      o135(.An(ori_ori_n66_), .B(ori_ori_n151_), .Y(ori_ori_n152_));
  NA2        o136(.A(ori_ori_n150_), .B(x6), .Y(ori_ori_n153_));
  AOI210     o137(.A0(ori_ori_n153_), .A1(ori_ori_n152_), .B0(ori_ori_n107_), .Y(ori_ori_n154_));
  OR2        o138(.A(ori_ori_n154_), .B(ori_ori_n127_), .Y(ori_ori_n155_));
  NA2        o139(.A(ori_ori_n35_), .B(ori_ori_n45_), .Y(ori_ori_n156_));
  NA2        o140(.A(ori_ori_n100_), .B(ori_ori_n70_), .Y(ori_ori_n157_));
  NA2        o141(.A(x6), .B(ori_ori_n40_), .Y(ori_ori_n158_));
  OAI210     o142(.A0(ori_ori_n84_), .A1(ori_ori_n62_), .B0(x4), .Y(ori_ori_n159_));
  AOI210     o143(.A0(ori_ori_n159_), .A1(ori_ori_n158_), .B0(ori_ori_n61_), .Y(ori_ori_n160_));
  OAI210     o144(.A0(ori_ori_n54_), .A1(ori_ori_n160_), .B0(x2), .Y(ori_ori_n161_));
  NA3        o145(.A(ori_ori_n161_), .B(ori_ori_n157_), .C(ori_ori_n155_), .Y(ori_ori_n162_));
  INV        o146(.A(ori_ori_n162_), .Y(ori_ori_n163_));
  INV        o147(.A(x3), .Y(ori_ori_n164_));
  NA2        o148(.A(ori_ori_n164_), .B(ori_ori_n144_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n69_), .B(ori_ori_n23_), .Y(ori_ori_n166_));
  AOI210     o150(.A0(ori_ori_n151_), .A1(ori_ori_n110_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  AOI210     o151(.A0(ori_ori_n167_), .A1(ori_ori_n165_), .B0(x2), .Y(ori_ori_n168_));
  AOI220     o152(.A0(ori_ori_n144_), .A1(ori_ori_n136_), .B0(x2), .B1(ori_ori_n54_), .Y(ori_ori_n169_));
  NA2        o153(.A(ori_ori_n35_), .B(ori_ori_n17_), .Y(ori_ori_n170_));
  NA2        o154(.A(ori_ori_n146_), .B(x6), .Y(ori_ori_n171_));
  NO2        o155(.A(ori_ori_n146_), .B(x6), .Y(ori_ori_n172_));
  INV        o156(.A(ori_ori_n172_), .Y(ori_ori_n173_));
  NA3        o157(.A(ori_ori_n173_), .B(ori_ori_n171_), .C(ori_ori_n104_), .Y(ori_ori_n174_));
  NA3        o158(.A(ori_ori_n174_), .B(ori_ori_n169_), .C(ori_ori_n107_), .Y(ori_ori_n175_));
  BUFFER     o159(.A(x1), .Y(ori_ori_n176_));
  NA2        o160(.A(x6), .B(x2), .Y(ori_ori_n177_));
  NA2        o161(.A(x4), .B(x0), .Y(ori_ori_n178_));
  NO2        o162(.A(ori_ori_n175_), .B(ori_ori_n168_), .Y(ori_ori_n179_));
  NA2        o163(.A(ori_ori_n172_), .B(x2), .Y(ori_ori_n180_));
  OAI210     o164(.A0(x0), .A1(x6), .B0(ori_ori_n36_), .Y(ori_ori_n181_));
  AOI210     o165(.A0(ori_ori_n181_), .A1(ori_ori_n180_), .B0(ori_ori_n135_), .Y(ori_ori_n182_));
  NOi21      o166(.An(ori_ori_n177_), .B(ori_ori_n17_), .Y(ori_ori_n183_));
  NA3        o167(.A(ori_ori_n183_), .B(ori_ori_n147_), .C(ori_ori_n32_), .Y(ori_ori_n184_));
  AOI210     o168(.A0(ori_ori_n30_), .A1(ori_ori_n45_), .B0(x0), .Y(ori_ori_n185_));
  NA3        o169(.A(ori_ori_n185_), .B(ori_ori_n114_), .C(ori_ori_n27_), .Y(ori_ori_n186_));
  NA2        o170(.A(x3), .B(x2), .Y(ori_ori_n187_));
  AOI220     o171(.A0(ori_ori_n187_), .A1(ori_ori_n156_), .B0(ori_ori_n186_), .B1(ori_ori_n184_), .Y(ori_ori_n188_));
  NAi21      o172(.An(x4), .B(x0), .Y(ori_ori_n189_));
  NO3        o173(.A(ori_ori_n189_), .B(ori_ori_n36_), .C(x2), .Y(ori_ori_n190_));
  OAI210     o174(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n190_), .Y(ori_ori_n191_));
  NO2        o175(.A(ori_ori_n185_), .B(ori_ori_n183_), .Y(ori_ori_n192_));
  AOI220     o176(.A0(ori_ori_n192_), .A1(ori_ori_n65_), .B0(ori_ori_n18_), .B1(ori_ori_n26_), .Y(ori_ori_n193_));
  AOI210     o177(.A0(ori_ori_n193_), .A1(ori_ori_n191_), .B0(ori_ori_n23_), .Y(ori_ori_n194_));
  NO2        o178(.A(ori_ori_n185_), .B(ori_ori_n183_), .Y(ori_ori_n195_));
  INV        o179(.A(ori_ori_n148_), .Y(ori_ori_n196_));
  NA2        o180(.A(ori_ori_n30_), .B(ori_ori_n35_), .Y(ori_ori_n197_));
  OR2        o181(.A(ori_ori_n197_), .B(ori_ori_n178_), .Y(ori_ori_n198_));
  OAI220     o182(.A0(ori_ori_n198_), .A1(ori_ori_n113_), .B0(ori_ori_n158_), .B1(ori_ori_n196_), .Y(ori_ori_n199_));
  AO210      o183(.A0(ori_ori_n195_), .A1(ori_ori_n105_), .B0(ori_ori_n199_), .Y(ori_ori_n200_));
  NO4        o184(.A(ori_ori_n200_), .B(ori_ori_n194_), .C(ori_ori_n188_), .D(ori_ori_n182_), .Y(ori_ori_n201_));
  OAI210     o185(.A0(ori_ori_n179_), .A1(ori_ori_n163_), .B0(ori_ori_n201_), .Y(ori04));
  NO2        o186(.A(x2), .B(x1), .Y(ori_ori_n203_));
  OAI210     o187(.A0(ori_ori_n170_), .A1(ori_ori_n203_), .B0(ori_ori_n30_), .Y(ori_ori_n204_));
  INV        o188(.A(ori_ori_n189_), .Y(ori_ori_n205_));
  OAI210     o189(.A0(ori_ori_n45_), .A1(ori_ori_n205_), .B0(ori_ori_n164_), .Y(ori_ori_n206_));
  NO2        o190(.A(ori_ori_n187_), .B(ori_ori_n145_), .Y(ori_ori_n207_));
  INV        o191(.A(ori_ori_n207_), .Y(ori_ori_n208_));
  NA3        o192(.A(ori_ori_n208_), .B(x6), .C(ori_ori_n206_), .Y(ori_ori_n209_));
  NA2        o193(.A(ori_ori_n209_), .B(ori_ori_n204_), .Y(ori_ori_n210_));
  INV        o194(.A(x7), .Y(ori_ori_n211_));
  XO2        o195(.A(x4), .B(x0), .Y(ori_ori_n212_));
  NA2        o196(.A(x4), .B(ori_ori_n72_), .Y(ori_ori_n213_));
  NO2        o197(.A(ori_ori_n213_), .B(x3), .Y(ori_ori_n214_));
  INV        o198(.A(ori_ori_n72_), .Y(ori_ori_n215_));
  NA2        o199(.A(ori_ori_n88_), .B(ori_ori_n215_), .Y(ori_ori_n216_));
  NO2        o200(.A(ori_ori_n212_), .B(x2), .Y(ori_ori_n217_));
  INV        o201(.A(ori_ori_n217_), .Y(ori_ori_n218_));
  NA3        o202(.A(ori_ori_n218_), .B(ori_ori_n216_), .C(x6), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n128_), .B(ori_ori_n71_), .Y(ori_ori_n220_));
  NA2        o204(.A(ori_ori_n220_), .B(ori_ori_n52_), .Y(ori_ori_n221_));
  NO2        o205(.A(x8), .B(ori_ori_n64_), .Y(ori_ori_n222_));
  NO2        o206(.A(ori_ori_n29_), .B(x2), .Y(ori_ori_n223_));
  NA2        o207(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  NA2        o208(.A(ori_ori_n221_), .B(ori_ori_n224_), .Y(ori_ori_n225_));
  OAI220     o209(.A0(ori_ori_n225_), .A1(x6), .B0(ori_ori_n219_), .B1(ori_ori_n214_), .Y(ori_ori_n226_));
  AO220      o210(.A0(x7), .A1(ori_ori_n226_), .B0(ori_ori_n211_), .B1(ori_ori_n210_), .Y(ori_ori_n227_));
  NA2        o211(.A(ori_ori_n149_), .B(ori_ori_n41_), .Y(ori_ori_n228_));
  NA2        o212(.A(ori_ori_n228_), .B(ori_ori_n227_), .Y(ori_ori_n229_));
  NA3        o213(.A(ori_ori_n17_), .B(ori_ori_n142_), .C(ori_ori_n107_), .Y(ori_ori_n230_));
  NA3        o214(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n231_));
  NO2        o215(.A(ori_ori_n231_), .B(ori_ori_n215_), .Y(ori_ori_n232_));
  INV        o216(.A(ori_ori_n232_), .Y(ori_ori_n233_));
  AOI210     o217(.A0(ori_ori_n233_), .A1(ori_ori_n230_), .B0(ori_ori_n23_), .Y(ori_ori_n234_));
  NA2        o218(.A(ori_ori_n234_), .B(x6), .Y(ori_ori_n235_));
  INV        o219(.A(ori_ori_n94_), .Y(ori_ori_n236_));
  NO2        o220(.A(ori_ori_n236_), .B(ori_ori_n35_), .Y(ori_ori_n237_));
  AOI210     o221(.A0(ori_ori_n176_), .A1(ori_ori_n51_), .B0(ori_ori_n87_), .Y(ori_ori_n238_));
  NO2        o222(.A(ori_ori_n238_), .B(x3), .Y(ori_ori_n239_));
  NO3        o223(.A(ori_ori_n239_), .B(ori_ori_n237_), .C(x2), .Y(ori_ori_n240_));
  OAI210     o224(.A0(ori_ori_n189_), .A1(ori_ori_n35_), .B0(ori_ori_n212_), .Y(ori_ori_n241_));
  AOI220     o225(.A0(x7), .A1(ori_ori_n71_), .B0(ori_ori_n241_), .B1(ori_ori_n107_), .Y(ori_ori_n242_));
  NO2        o226(.A(ori_ori_n242_), .B(ori_ori_n45_), .Y(ori_ori_n243_));
  NO2        o227(.A(ori_ori_n243_), .B(ori_ori_n240_), .Y(ori_ori_n244_));
  AOI210     o228(.A0(ori_ori_n244_), .A1(ori_ori_n42_), .B0(ori_ori_n23_), .Y(ori_ori_n245_));
  NA2        o229(.A(ori_ori_n245_), .B(ori_ori_n30_), .Y(ori_ori_n246_));
  INV        o230(.A(ori_ori_n145_), .Y(ori_ori_n247_));
  NO4        o231(.A(ori_ori_n247_), .B(ori_ori_n61_), .C(x4), .D(ori_ori_n45_), .Y(ori_ori_n248_));
  INV        o232(.A(ori_ori_n69_), .Y(ori_ori_n249_));
  NA2        o233(.A(ori_ori_n249_), .B(ori_ori_n127_), .Y(ori_ori_n250_));
  NO2        o234(.A(ori_ori_n113_), .B(ori_ori_n35_), .Y(ori_ori_n251_));
  NA2        o235(.A(x3), .B(ori_ori_n45_), .Y(ori_ori_n252_));
  NO2        o236(.A(ori_ori_n108_), .B(ori_ori_n252_), .Y(ori_ori_n253_));
  AOI220     o237(.A0(ori_ori_n253_), .A1(x0), .B0(ori_ori_n251_), .B1(ori_ori_n95_), .Y(ori_ori_n254_));
  AOI210     o238(.A0(ori_ori_n254_), .A1(ori_ori_n250_), .B0(ori_ori_n158_), .Y(ori_ori_n255_));
  NO2        o239(.A(ori_ori_n255_), .B(ori_ori_n248_), .Y(ori_ori_n256_));
  NA3        o240(.A(ori_ori_n256_), .B(ori_ori_n246_), .C(ori_ori_n235_), .Y(ori_ori_n257_));
  AOI210     o241(.A0(ori_ori_n229_), .A1(ori_ori_n23_), .B0(ori_ori_n257_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  NO3        m047(.A(mai_mai_n36_), .B(mai_mai_n61_), .C(mai_mai_n60_), .Y(mai_mai_n64_));
  NO2        m048(.A(x7), .B(x6), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(x8), .B(x2), .Y(mai_mai_n67_));
  OA210      m051(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n69_), .Y(mai_mai_n70_));
  NAi31      m054(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n71_));
  NO2        m055(.A(mai_mai_n70_), .B(mai_mai_n68_), .Y(mai_mai_n72_));
  OAI210     m056(.A0(mai_mai_n72_), .A1(mai_mai_n64_), .B0(x4), .Y(mai_mai_n73_));
  NA2        m057(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n74_));
  OAI210     m058(.A0(mai_mai_n74_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n75_));
  NA2        m059(.A(x5), .B(x3), .Y(mai_mai_n76_));
  NO2        m060(.A(x8), .B(x6), .Y(mai_mai_n77_));
  NO4        m061(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(mai_mai_n65_), .D(mai_mai_n54_), .Y(mai_mai_n78_));
  NAi21      m062(.An(x4), .B(x3), .Y(mai_mai_n79_));
  INV        m063(.A(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n80_), .B(mai_mai_n22_), .Y(mai_mai_n81_));
  NO2        m065(.A(x4), .B(x2), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(x3), .Y(mai_mai_n83_));
  NO3        m067(.A(mai_mai_n83_), .B(mai_mai_n81_), .C(mai_mai_n18_), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n78_), .C(mai_mai_n75_), .Y(mai_mai_n85_));
  NO4        m069(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n43_), .D(x1), .Y(mai_mai_n86_));
  NA2        m070(.A(mai_mai_n62_), .B(mai_mai_n48_), .Y(mai_mai_n87_));
  INV        m071(.A(mai_mai_n87_), .Y(mai_mai_n88_));
  OAI210     m072(.A0(mai_mai_n86_), .A1(mai_mai_n66_), .B0(mai_mai_n88_), .Y(mai_mai_n89_));
  NA2        m073(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n25_), .Y(mai_mai_n91_));
  INV        m075(.A(x8), .Y(mai_mai_n92_));
  NA2        m076(.A(x2), .B(x1), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n92_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n91_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n26_), .Y(mai_mai_n96_));
  AOI210     m080(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n97_));
  OAI210     m081(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n98_));
  NO3        m082(.A(mai_mai_n98_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n99_));
  NA2        m083(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n100_));
  NO2        m084(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n101_));
  OAI210     m085(.A0(mai_mai_n101_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n102_));
  AOI210     m086(.A0(mai_mai_n100_), .A1(mai_mai_n52_), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m087(.A(x3), .B(x2), .Y(mai_mai_n104_));
  NA3        m088(.A(mai_mai_n104_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n105_));
  AOI210     m089(.A0(x8), .A1(x6), .B0(mai_mai_n105_), .Y(mai_mai_n106_));
  NA2        m090(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n107_));
  OAI210     m091(.A0(mai_mai_n107_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n108_));
  NO4        m092(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n103_), .D(mai_mai_n99_), .Y(mai_mai_n109_));
  AO220      m093(.A0(mai_mai_n109_), .A1(mai_mai_n89_), .B0(mai_mai_n85_), .B1(mai_mai_n73_), .Y(mai02));
  NO2        m094(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n111_));
  NO2        m095(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n112_));
  NA2        m096(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n113_));
  OAI210     m097(.A0(mai_mai_n87_), .A1(x0), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  AOI220     m098(.A0(mai_mai_n114_), .A1(mai_mai_n112_), .B0(mai_mai_n111_), .B1(x4), .Y(mai_mai_n115_));
  NO3        m099(.A(mai_mai_n115_), .B(x7), .C(x5), .Y(mai_mai_n116_));
  OR2        m100(.A(x8), .B(x0), .Y(mai_mai_n117_));
  INV        m101(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NAi21      m102(.An(x2), .B(x8), .Y(mai_mai_n119_));
  INV        m103(.A(mai_mai_n119_), .Y(mai_mai_n120_));
  NO2        m104(.A(x4), .B(x1), .Y(mai_mai_n121_));
  NOi21      m105(.An(x0), .B(x1), .Y(mai_mai_n122_));
  NO3        m106(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n123_));
  NOi21      m107(.An(x0), .B(x4), .Y(mai_mai_n124_));
  NO2        m108(.A(x8), .B(mai_mai_n62_), .Y(mai_mai_n125_));
  AOI220     m109(.A0(mai_mai_n125_), .A1(mai_mai_n124_), .B0(mai_mai_n123_), .B1(mai_mai_n122_), .Y(mai_mai_n126_));
  NO2        m110(.A(mai_mai_n126_), .B(mai_mai_n76_), .Y(mai_mai_n127_));
  NO2        m111(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n128_));
  NA2        m112(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n129_));
  AOI210     m113(.A0(mai_mai_n129_), .A1(mai_mai_n107_), .B0(mai_mai_n113_), .Y(mai_mai_n130_));
  OAI210     m114(.A0(mai_mai_n130_), .A1(mai_mai_n35_), .B0(mai_mai_n128_), .Y(mai_mai_n131_));
  NAi21      m115(.An(x0), .B(x4), .Y(mai_mai_n132_));
  NO2        m116(.A(mai_mai_n132_), .B(x1), .Y(mai_mai_n133_));
  NO2        m117(.A(x7), .B(x0), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n82_), .B(mai_mai_n101_), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n135_), .B(x3), .Y(mai_mai_n136_));
  OAI210     m120(.A0(mai_mai_n134_), .A1(mai_mai_n133_), .B0(mai_mai_n136_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n138_));
  NA2        m122(.A(x5), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n140_));
  NA3        m124(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n138_), .Y(mai_mai_n141_));
  NA4        m125(.A(mai_mai_n141_), .B(mai_mai_n137_), .C(mai_mai_n131_), .D(mai_mai_n36_), .Y(mai_mai_n142_));
  NO3        m126(.A(mai_mai_n142_), .B(mai_mai_n127_), .C(mai_mai_n116_), .Y(mai_mai_n143_));
  NO2        m127(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n144_));
  AOI220     m128(.A0(mai_mai_n122_), .A1(mai_mai_n144_), .B0(mai_mai_n66_), .B1(mai_mai_n17_), .Y(mai_mai_n145_));
  NO3        m129(.A(mai_mai_n145_), .B(mai_mai_n60_), .C(mai_mai_n62_), .Y(mai_mai_n146_));
  NA2        m130(.A(x7), .B(x3), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n100_), .B(x5), .Y(mai_mai_n148_));
  NO2        m132(.A(x9), .B(x7), .Y(mai_mai_n149_));
  NOi21      m133(.An(x8), .B(x0), .Y(mai_mai_n150_));
  NO2        m134(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n151_));
  INV        m135(.A(x7), .Y(mai_mai_n152_));
  AOI210     m136(.A0(mai_mai_n111_), .A1(mai_mai_n38_), .B0(mai_mai_n151_), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n154_));
  NO2        m138(.A(mai_mai_n154_), .B(mai_mai_n124_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n155_), .B(mai_mai_n153_), .Y(mai_mai_n156_));
  AOI210     m140(.A0(mai_mai_n150_), .A1(mai_mai_n148_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  OAI210     m141(.A0(mai_mai_n147_), .A1(mai_mai_n50_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  NA2        m142(.A(x5), .B(x1), .Y(mai_mai_n159_));
  INV        m143(.A(mai_mai_n159_), .Y(mai_mai_n160_));
  AOI210     m144(.A0(mai_mai_n160_), .A1(mai_mai_n124_), .B0(mai_mai_n36_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n62_), .B(mai_mai_n92_), .Y(mai_mai_n162_));
  NAi21      m146(.An(x2), .B(x7), .Y(mai_mai_n163_));
  NAi31      m147(.An(mai_mai_n76_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n164_));
  NA2        m148(.A(mai_mai_n164_), .B(mai_mai_n161_), .Y(mai_mai_n165_));
  NO3        m149(.A(mai_mai_n165_), .B(mai_mai_n158_), .C(mai_mai_n146_), .Y(mai_mai_n166_));
  NO2        m150(.A(mai_mai_n166_), .B(mai_mai_n143_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n139_), .B(mai_mai_n135_), .Y(mai_mai_n168_));
  NA2        m152(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n169_));
  NA2        m153(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n170_));
  NA3        m154(.A(mai_mai_n170_), .B(mai_mai_n169_), .C(mai_mai_n24_), .Y(mai_mai_n171_));
  AN2        m155(.A(mai_mai_n171_), .B(mai_mai_n140_), .Y(mai_mai_n172_));
  NA2        m156(.A(x8), .B(x0), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n152_), .B(mai_mai_n25_), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n122_), .B(x4), .Y(mai_mai_n175_));
  NA2        m159(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  AOI210     m160(.A0(mai_mai_n173_), .A1(mai_mai_n129_), .B0(mai_mai_n176_), .Y(mai_mai_n177_));
  NA2        m161(.A(x2), .B(x0), .Y(mai_mai_n178_));
  NA2        m162(.A(x4), .B(x1), .Y(mai_mai_n179_));
  NAi21      m163(.An(mai_mai_n121_), .B(mai_mai_n179_), .Y(mai_mai_n180_));
  NOi31      m164(.An(mai_mai_n180_), .B(mai_mai_n154_), .C(mai_mai_n178_), .Y(mai_mai_n181_));
  NO4        m165(.A(mai_mai_n181_), .B(mai_mai_n177_), .C(mai_mai_n172_), .D(mai_mai_n168_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n182_), .B(mai_mai_n43_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n171_), .B(mai_mai_n74_), .Y(mai_mai_n184_));
  INV        m168(.A(mai_mai_n128_), .Y(mai_mai_n185_));
  NO3        m169(.A(mai_mai_n410_), .B(mai_mai_n185_), .C(x7), .Y(mai_mai_n186_));
  NA3        m170(.A(mai_mai_n180_), .B(mai_mai_n185_), .C(mai_mai_n42_), .Y(mai_mai_n187_));
  OAI210     m171(.A0(mai_mai_n170_), .A1(mai_mai_n135_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  NO3        m172(.A(mai_mai_n188_), .B(mai_mai_n186_), .C(mai_mai_n184_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n189_), .B(x3), .Y(mai_mai_n190_));
  NO3        m174(.A(mai_mai_n190_), .B(mai_mai_n183_), .C(mai_mai_n167_), .Y(mai03));
  NO2        m175(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n192_));
  NO2        m176(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n194_));
  OAI210     m178(.A0(mai_mai_n194_), .A1(mai_mai_n25_), .B0(mai_mai_n63_), .Y(mai_mai_n195_));
  OAI220     m179(.A0(mai_mai_n195_), .A1(mai_mai_n17_), .B0(x6), .B1(mai_mai_n107_), .Y(mai_mai_n196_));
  NA2        m180(.A(mai_mai_n196_), .B(mai_mai_n192_), .Y(mai_mai_n197_));
  NO2        m181(.A(mai_mai_n76_), .B(x6), .Y(mai_mai_n198_));
  NA2        m182(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n199_));
  NO2        m183(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n200_));
  NA2        m184(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n201_), .B(mai_mai_n199_), .Y(mai_mai_n202_));
  NA2        m186(.A(x9), .B(mai_mai_n54_), .Y(mai_mai_n203_));
  NA2        m187(.A(mai_mai_n199_), .B(mai_mai_n79_), .Y(mai_mai_n204_));
  AOI210     m188(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n178_), .Y(mai_mai_n205_));
  AOI210     m189(.A0(mai_mai_n205_), .A1(mai_mai_n204_), .B0(mai_mai_n202_), .Y(mai_mai_n206_));
  NO3        m190(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n207_));
  NO2        m191(.A(x5), .B(x1), .Y(mai_mai_n208_));
  AOI220     m192(.A0(mai_mai_n208_), .A1(mai_mai_n17_), .B0(mai_mai_n104_), .B1(x5), .Y(mai_mai_n209_));
  NO2        m193(.A(mai_mai_n201_), .B(mai_mai_n169_), .Y(mai_mai_n210_));
  NO3        m194(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n211_));
  AOI220     m195(.A0(mai_mai_n413_), .A1(mai_mai_n48_), .B0(mai_mai_n207_), .B1(mai_mai_n128_), .Y(mai_mai_n212_));
  NA3        m196(.A(mai_mai_n212_), .B(mai_mai_n206_), .C(mai_mai_n197_), .Y(mai_mai_n213_));
  NO2        m197(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n214_));
  NA2        m198(.A(mai_mai_n214_), .B(mai_mai_n19_), .Y(mai_mai_n215_));
  NO2        m199(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n216_), .B(x6), .Y(mai_mai_n217_));
  NOi21      m201(.An(mai_mai_n82_), .B(mai_mai_n217_), .Y(mai_mai_n218_));
  NA2        m202(.A(mai_mai_n62_), .B(mai_mai_n92_), .Y(mai_mai_n219_));
  NO2        m203(.A(mai_mai_n218_), .B(mai_mai_n152_), .Y(mai_mai_n220_));
  AO210      m204(.A0(mai_mai_n220_), .A1(mai_mai_n215_), .B0(mai_mai_n174_), .Y(mai_mai_n221_));
  NA2        m205(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n222_));
  NO3        m206(.A(mai_mai_n179_), .B(mai_mai_n62_), .C(x6), .Y(mai_mai_n223_));
  AOI220     m207(.A0(mai_mai_n223_), .A1(mai_mai_n54_), .B0(mai_mai_n140_), .B1(mai_mai_n91_), .Y(mai_mai_n224_));
  NA2        m208(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n225_));
  NO2        m209(.A(mai_mai_n159_), .B(mai_mai_n43_), .Y(mai_mai_n226_));
  OAI210     m210(.A0(mai_mai_n226_), .A1(mai_mai_n210_), .B0(mai_mai_n409_), .Y(mai_mai_n227_));
  NA2        m211(.A(mai_mai_n193_), .B(mai_mai_n133_), .Y(mai_mai_n228_));
  NA2        m212(.A(mai_mai_n128_), .B(x6), .Y(mai_mai_n229_));
  OAI210     m213(.A0(mai_mai_n92_), .A1(mai_mai_n36_), .B0(mai_mai_n66_), .Y(mai_mai_n230_));
  NA4        m214(.A(mai_mai_n230_), .B(mai_mai_n229_), .C(mai_mai_n228_), .D(mai_mai_n227_), .Y(mai_mai_n231_));
  NA2        m215(.A(mai_mai_n231_), .B(x2), .Y(mai_mai_n232_));
  NA3        m216(.A(mai_mai_n232_), .B(mai_mai_n224_), .C(mai_mai_n221_), .Y(mai_mai_n233_));
  AOI210     m217(.A0(mai_mai_n213_), .A1(x8), .B0(mai_mai_n233_), .Y(mai_mai_n234_));
  NO2        m218(.A(mai_mai_n92_), .B(x3), .Y(mai_mai_n235_));
  NO3        m219(.A(mai_mai_n90_), .B(mai_mai_n77_), .C(mai_mai_n25_), .Y(mai_mai_n236_));
  NO2        m220(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n237_));
  NA2        m221(.A(mai_mai_n237_), .B(mai_mai_n66_), .Y(mai_mai_n238_));
  NA3        m222(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n239_));
  AOI210     m223(.A0(mai_mai_n239_), .A1(mai_mai_n139_), .B0(x9), .Y(mai_mai_n240_));
  NA2        m224(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n241_));
  NA2        m225(.A(mai_mai_n240_), .B(mai_mai_n121_), .Y(mai_mai_n242_));
  INV        m226(.A(x6), .Y(mai_mai_n243_));
  NO2        m227(.A(mai_mai_n201_), .B(x6), .Y(mai_mai_n244_));
  NA2        m228(.A(mai_mai_n243_), .B(mai_mai_n144_), .Y(mai_mai_n245_));
  NA4        m229(.A(mai_mai_n245_), .B(mai_mai_n242_), .C(mai_mai_n238_), .D(mai_mai_n152_), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n193_), .B(mai_mai_n216_), .Y(mai_mai_n247_));
  NO2        m231(.A(x9), .B(x6), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n139_), .B(mai_mai_n18_), .Y(mai_mai_n249_));
  NAi21      m233(.An(mai_mai_n249_), .B(mai_mai_n239_), .Y(mai_mai_n250_));
  NAi21      m234(.An(x1), .B(x4), .Y(mai_mai_n251_));
  AOI210     m235(.A0(x3), .A1(x2), .B0(mai_mai_n48_), .Y(mai_mai_n252_));
  OAI210     m236(.A0(mai_mai_n139_), .A1(x3), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  AOI220     m237(.A0(mai_mai_n253_), .A1(mai_mai_n251_), .B0(mai_mai_n250_), .B1(mai_mai_n248_), .Y(mai_mai_n254_));
  NA2        m238(.A(mai_mai_n254_), .B(mai_mai_n247_), .Y(mai_mai_n255_));
  NO3        m239(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n256_));
  INV        m240(.A(mai_mai_n256_), .Y(mai_mai_n257_));
  OAI220     m241(.A0(mai_mai_n257_), .A1(mai_mai_n43_), .B0(mai_mai_n175_), .B1(mai_mai_n46_), .Y(mai_mai_n258_));
  OAI210     m242(.A0(mai_mai_n258_), .A1(mai_mai_n193_), .B0(mai_mai_n255_), .Y(mai_mai_n259_));
  OR2        m243(.A(mai_mai_n198_), .B(mai_mai_n148_), .Y(mai_mai_n260_));
  NA2        m244(.A(x4), .B(x0), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n260_), .B(mai_mai_n42_), .Y(mai_mai_n262_));
  AOI210     m246(.A0(mai_mai_n262_), .A1(mai_mai_n259_), .B0(x8), .Y(mai_mai_n263_));
  OAI210     m247(.A0(mai_mai_n249_), .A1(mai_mai_n208_), .B0(x6), .Y(mai_mai_n264_));
  INV        m248(.A(mai_mai_n173_), .Y(mai_mai_n265_));
  OAI210     m249(.A0(mai_mai_n265_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n266_));
  AOI210     m250(.A0(mai_mai_n266_), .A1(mai_mai_n264_), .B0(mai_mai_n222_), .Y(mai_mai_n267_));
  NO4        m251(.A(mai_mai_n267_), .B(mai_mai_n263_), .C(mai_mai_n246_), .D(mai_mai_n236_), .Y(mai_mai_n268_));
  NO2        m252(.A(mai_mai_n162_), .B(x1), .Y(mai_mai_n269_));
  NO2        m253(.A(x3), .B(mai_mai_n36_), .Y(mai_mai_n270_));
  OAI210     m254(.A0(mai_mai_n270_), .A1(mai_mai_n244_), .B0(x2), .Y(mai_mai_n271_));
  OAI210     m255(.A0(mai_mai_n265_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n272_));
  AOI210     m256(.A0(mai_mai_n272_), .A1(mai_mai_n271_), .B0(mai_mai_n185_), .Y(mai_mai_n273_));
  NA3        m257(.A(x0), .B(mai_mai_n208_), .C(mai_mai_n40_), .Y(mai_mai_n274_));
  AOI210     m258(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n275_));
  NA3        m259(.A(mai_mai_n275_), .B(mai_mai_n160_), .C(mai_mai_n32_), .Y(mai_mai_n276_));
  NA2        m260(.A(x3), .B(x2), .Y(mai_mai_n277_));
  AOI220     m261(.A0(mai_mai_n277_), .A1(mai_mai_n222_), .B0(mai_mai_n276_), .B1(mai_mai_n274_), .Y(mai_mai_n278_));
  NAi21      m262(.An(x4), .B(x0), .Y(mai_mai_n279_));
  NO3        m263(.A(mai_mai_n279_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n280_));
  OAI210     m264(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  OAI220     m265(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n282_));
  AOI220     m266(.A0(mai_mai_n36_), .A1(mai_mai_n80_), .B0(mai_mai_n282_), .B1(mai_mai_n31_), .Y(mai_mai_n283_));
  AOI210     m267(.A0(mai_mai_n283_), .A1(mai_mai_n281_), .B0(mai_mai_n25_), .Y(mai_mai_n284_));
  NA3        m268(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n285_));
  INV        m269(.A(mai_mai_n210_), .Y(mai_mai_n286_));
  NA2        m270(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n287_));
  OR2        m271(.A(mai_mai_n287_), .B(mai_mai_n261_), .Y(mai_mai_n288_));
  OAI220     m272(.A0(mai_mai_n288_), .A1(mai_mai_n159_), .B0(mai_mai_n225_), .B1(mai_mai_n286_), .Y(mai_mai_n289_));
  NO4        m273(.A(mai_mai_n289_), .B(mai_mai_n284_), .C(mai_mai_n278_), .D(mai_mai_n273_), .Y(mai_mai_n290_));
  OAI210     m274(.A0(mai_mai_n268_), .A1(mai_mai_n234_), .B0(mai_mai_n290_), .Y(mai04));
  NA2        m275(.A(mai_mai_n256_), .B(mai_mai_n83_), .Y(mai_mai_n292_));
  NO2        m276(.A(mai_mai_n277_), .B(mai_mai_n200_), .Y(mai_mai_n293_));
  NA2        m277(.A(x9), .B(x0), .Y(mai_mai_n294_));
  NO2        m278(.A(mai_mai_n90_), .B(mai_mai_n294_), .Y(mai_mai_n295_));
  OAI210     m279(.A0(mai_mai_n295_), .A1(mai_mai_n293_), .B0(mai_mai_n92_), .Y(mai_mai_n296_));
  INV        m280(.A(mai_mai_n296_), .Y(mai_mai_n297_));
  NA2        m281(.A(mai_mai_n297_), .B(x6), .Y(mai_mai_n298_));
  NO3        m282(.A(x9), .B(mai_mai_n119_), .C(mai_mai_n18_), .Y(mai_mai_n299_));
  INV        m283(.A(mai_mai_n299_), .Y(mai_mai_n300_));
  OAI210     m284(.A0(mai_mai_n117_), .A1(mai_mai_n107_), .B0(mai_mai_n173_), .Y(mai_mai_n301_));
  NA3        m285(.A(mai_mai_n301_), .B(x6), .C(x3), .Y(mai_mai_n302_));
  OAI210     m286(.A0(x9), .A1(mai_mai_n285_), .B0(mai_mai_n287_), .Y(mai_mai_n303_));
  AOI210     m287(.A0(mai_mai_n150_), .A1(mai_mai_n63_), .B0(mai_mai_n303_), .Y(mai_mai_n304_));
  NA2        m288(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n305_));
  NA4        m289(.A(mai_mai_n411_), .B(mai_mai_n304_), .C(mai_mai_n302_), .D(mai_mai_n300_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n112_), .A1(x3), .B0(mai_mai_n280_), .Y(mai_mai_n307_));
  NA3        m291(.A(mai_mai_n219_), .B(mai_mai_n207_), .C(mai_mai_n82_), .Y(mai_mai_n308_));
  NA3        m292(.A(mai_mai_n308_), .B(mai_mai_n307_), .C(mai_mai_n152_), .Y(mai_mai_n309_));
  AOI210     m293(.A0(mai_mai_n306_), .A1(x4), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  NOi21      m294(.An(x4), .B(x0), .Y(mai_mai_n311_));
  AOI210     m295(.A0(x2), .A1(x8), .B0(mai_mai_n311_), .Y(mai_mai_n312_));
  AOI210     m296(.A0(mai_mai_n312_), .A1(mai_mai_n279_), .B0(x3), .Y(mai_mai_n313_));
  NO2        m297(.A(mai_mai_n92_), .B(x4), .Y(mai_mai_n314_));
  NA2        m298(.A(mai_mai_n314_), .B(mai_mai_n44_), .Y(mai_mai_n315_));
  NO2        m299(.A(mai_mai_n28_), .B(mai_mai_n24_), .Y(mai_mai_n316_));
  INV        m300(.A(mai_mai_n316_), .Y(mai_mai_n317_));
  NA4        m301(.A(mai_mai_n317_), .B(mai_mai_n315_), .C(mai_mai_n215_), .D(x6), .Y(mai_mai_n318_));
  NO2        m302(.A(mai_mai_n150_), .B(mai_mai_n107_), .Y(mai_mai_n319_));
  AOI210     m303(.A0(mai_mai_n412_), .A1(mai_mai_n61_), .B0(mai_mai_n319_), .Y(mai_mai_n320_));
  NO2        m304(.A(mai_mai_n150_), .B(mai_mai_n79_), .Y(mai_mai_n321_));
  NO2        m305(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n322_));
  NOi21      m306(.An(mai_mai_n121_), .B(mai_mai_n27_), .Y(mai_mai_n323_));
  AOI210     m307(.A0(mai_mai_n322_), .A1(mai_mai_n321_), .B0(mai_mai_n323_), .Y(mai_mai_n324_));
  OAI210     m308(.A0(mai_mai_n320_), .A1(mai_mai_n62_), .B0(mai_mai_n324_), .Y(mai_mai_n325_));
  OAI220     m309(.A0(mai_mai_n325_), .A1(x6), .B0(mai_mai_n318_), .B1(mai_mai_n313_), .Y(mai_mai_n326_));
  OAI210     m310(.A0(mai_mai_n414_), .A1(mai_mai_n92_), .B0(mai_mai_n288_), .Y(mai_mai_n327_));
  AOI210     m311(.A0(mai_mai_n327_), .A1(mai_mai_n18_), .B0(mai_mai_n152_), .Y(mai_mai_n328_));
  AO220      m312(.A0(mai_mai_n328_), .A1(mai_mai_n326_), .B0(mai_mai_n310_), .B1(mai_mai_n298_), .Y(mai_mai_n329_));
  NA2        m313(.A(mai_mai_n322_), .B(x6), .Y(mai_mai_n330_));
  AOI210     m314(.A0(x6), .A1(x1), .B0(mai_mai_n151_), .Y(mai_mai_n331_));
  NA2        m315(.A(mai_mai_n314_), .B(x0), .Y(mai_mai_n332_));
  NA2        m316(.A(mai_mai_n82_), .B(x6), .Y(mai_mai_n333_));
  OAI210     m317(.A0(mai_mai_n332_), .A1(mai_mai_n331_), .B0(mai_mai_n333_), .Y(mai_mai_n334_));
  AOI220     m318(.A0(mai_mai_n334_), .A1(mai_mai_n330_), .B0(mai_mai_n211_), .B1(mai_mai_n49_), .Y(mai_mai_n335_));
  NA3        m319(.A(mai_mai_n335_), .B(mai_mai_n329_), .C(mai_mai_n292_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(mai_mai_n194_), .A1(x8), .B0(mai_mai_n112_), .Y(mai_mai_n337_));
  NA2        m321(.A(mai_mai_n337_), .B(mai_mai_n305_), .Y(mai_mai_n338_));
  NA3        m322(.A(mai_mai_n338_), .B(mai_mai_n192_), .C(mai_mai_n152_), .Y(mai_mai_n339_));
  AO210      m323(.A0(mai_mai_n111_), .A1(x4), .B0(mai_mai_n149_), .Y(mai_mai_n340_));
  NA2        m324(.A(mai_mai_n214_), .B(x0), .Y(mai_mai_n341_));
  NO2        m325(.A(mai_mai_n341_), .B(mai_mai_n203_), .Y(mai_mai_n342_));
  AOI210     m326(.A0(mai_mai_n340_), .A1(mai_mai_n118_), .B0(mai_mai_n342_), .Y(mai_mai_n343_));
  AOI210     m327(.A0(mai_mai_n343_), .A1(mai_mai_n339_), .B0(mai_mai_n25_), .Y(mai_mai_n344_));
  NA3        m328(.A(mai_mai_n120_), .B(mai_mai_n214_), .C(x0), .Y(mai_mai_n345_));
  OAI210     m329(.A0(mai_mai_n192_), .A1(mai_mai_n67_), .B0(mai_mai_n200_), .Y(mai_mai_n346_));
  NA3        m330(.A(mai_mai_n194_), .B(mai_mai_n216_), .C(x8), .Y(mai_mai_n347_));
  AOI210     m331(.A0(mai_mai_n347_), .A1(mai_mai_n346_), .B0(mai_mai_n25_), .Y(mai_mai_n348_));
  AOI210     m332(.A0(mai_mai_n119_), .A1(mai_mai_n117_), .B0(mai_mai_n42_), .Y(mai_mai_n349_));
  NOi31      m333(.An(mai_mai_n349_), .B(x3), .C(mai_mai_n179_), .Y(mai_mai_n350_));
  OAI210     m334(.A0(mai_mai_n350_), .A1(mai_mai_n348_), .B0(mai_mai_n149_), .Y(mai_mai_n351_));
  NAi31      m335(.An(mai_mai_n50_), .B(mai_mai_n269_), .C(mai_mai_n174_), .Y(mai_mai_n352_));
  NA3        m336(.A(mai_mai_n352_), .B(mai_mai_n351_), .C(mai_mai_n345_), .Y(mai_mai_n353_));
  OAI210     m337(.A0(mai_mai_n353_), .A1(mai_mai_n344_), .B0(x6), .Y(mai_mai_n354_));
  INV        m338(.A(mai_mai_n134_), .Y(mai_mai_n355_));
  NA3        m339(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n356_));
  AOI220     m340(.A0(mai_mai_n356_), .A1(mai_mai_n355_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n357_));
  NA2        m341(.A(mai_mai_n192_), .B(mai_mai_n152_), .Y(mai_mai_n358_));
  INV        m342(.A(x1), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n358_), .A1(x8), .B0(mai_mai_n359_), .Y(mai_mai_n360_));
  NAi31      m344(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n361_));
  OAI210     m345(.A0(mai_mai_n361_), .A1(x4), .B0(mai_mai_n163_), .Y(mai_mai_n362_));
  NA3        m346(.A(mai_mai_n362_), .B(mai_mai_n147_), .C(x9), .Y(mai_mai_n363_));
  NO4        m347(.A(x8), .B(mai_mai_n279_), .C(x9), .D(x2), .Y(mai_mai_n364_));
  NOi21      m348(.An(mai_mai_n123_), .B(mai_mai_n178_), .Y(mai_mai_n365_));
  NO3        m349(.A(mai_mai_n365_), .B(mai_mai_n364_), .C(mai_mai_n18_), .Y(mai_mai_n366_));
  NO3        m350(.A(x9), .B(mai_mai_n152_), .C(x0), .Y(mai_mai_n367_));
  AOI220     m351(.A0(mai_mai_n367_), .A1(mai_mai_n235_), .B0(mai_mai_n321_), .B1(mai_mai_n152_), .Y(mai_mai_n368_));
  NA4        m352(.A(mai_mai_n368_), .B(mai_mai_n366_), .C(mai_mai_n363_), .D(mai_mai_n50_), .Y(mai_mai_n369_));
  OAI210     m353(.A0(mai_mai_n360_), .A1(mai_mai_n357_), .B0(mai_mai_n369_), .Y(mai_mai_n370_));
  NO2        m354(.A(mai_mai_n123_), .B(mai_mai_n43_), .Y(mai_mai_n371_));
  NOi31      m355(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n372_));
  AOI210     m356(.A0(mai_mai_n124_), .A1(x3), .B0(mai_mai_n311_), .Y(mai_mai_n373_));
  NA2        m357(.A(x3), .B(mai_mai_n373_), .Y(mai_mai_n374_));
  NO3        m358(.A(mai_mai_n374_), .B(mai_mai_n371_), .C(x2), .Y(mai_mai_n375_));
  INV        m359(.A(mai_mai_n375_), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n376_), .A1(mai_mai_n370_), .B0(mai_mai_n25_), .Y(mai_mai_n377_));
  NA4        m361(.A(mai_mai_n31_), .B(mai_mai_n92_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n378_));
  NO3        m362(.A(mai_mai_n67_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n379_));
  AOI220     m363(.A0(mai_mai_n379_), .A1(mai_mai_n252_), .B0(mai_mai_n415_), .B1(mai_mai_n349_), .Y(mai_mai_n380_));
  NO2        m364(.A(mai_mai_n380_), .B(mai_mai_n104_), .Y(mai_mai_n381_));
  NA2        m365(.A(mai_mai_n381_), .B(x7), .Y(mai_mai_n382_));
  NA2        m366(.A(mai_mai_n219_), .B(x7), .Y(mai_mai_n383_));
  NA3        m367(.A(mai_mai_n383_), .B(mai_mai_n151_), .C(mai_mai_n133_), .Y(mai_mai_n384_));
  NA3        m368(.A(mai_mai_n384_), .B(mai_mai_n382_), .C(mai_mai_n378_), .Y(mai_mai_n385_));
  OAI210     m369(.A0(mai_mai_n385_), .A1(mai_mai_n377_), .B0(mai_mai_n36_), .Y(mai_mai_n386_));
  NO2        m370(.A(mai_mai_n367_), .B(mai_mai_n200_), .Y(mai_mai_n387_));
  NO4        m371(.A(mai_mai_n387_), .B(mai_mai_n76_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n388_));
  NA2        m372(.A(mai_mai_n241_), .B(mai_mai_n21_), .Y(mai_mai_n389_));
  NO2        m373(.A(mai_mai_n159_), .B(mai_mai_n134_), .Y(mai_mai_n390_));
  NA2        m374(.A(mai_mai_n390_), .B(mai_mai_n389_), .Y(mai_mai_n391_));
  AOI210     m375(.A0(mai_mai_n391_), .A1(mai_mai_n164_), .B0(mai_mai_n28_), .Y(mai_mai_n392_));
  AOI220     m376(.A0(x3), .A1(mai_mai_n92_), .B0(mai_mai_n150_), .B1(mai_mai_n194_), .Y(mai_mai_n393_));
  NA3        m377(.A(mai_mai_n393_), .B(mai_mai_n361_), .C(mai_mai_n90_), .Y(mai_mai_n394_));
  NA2        m378(.A(mai_mai_n394_), .B(mai_mai_n174_), .Y(mai_mai_n395_));
  AOI210     m379(.A0(mai_mai_n163_), .A1(mai_mai_n27_), .B0(mai_mai_n71_), .Y(mai_mai_n396_));
  NO3        m380(.A(mai_mai_n372_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n397_));
  NO2        m381(.A(mai_mai_n397_), .B(mai_mai_n396_), .Y(mai_mai_n398_));
  INV        m382(.A(mai_mai_n398_), .Y(mai_mai_n399_));
  AOI220     m383(.A0(mai_mai_n399_), .A1(x0), .B0(x5), .B1(mai_mai_n134_), .Y(mai_mai_n400_));
  AOI210     m384(.A0(mai_mai_n400_), .A1(mai_mai_n395_), .B0(mai_mai_n225_), .Y(mai_mai_n401_));
  NA2        m385(.A(x9), .B(x5), .Y(mai_mai_n402_));
  NO4        m386(.A(mai_mai_n107_), .B(mai_mai_n402_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n403_));
  NO4        m387(.A(mai_mai_n403_), .B(mai_mai_n401_), .C(mai_mai_n392_), .D(mai_mai_n388_), .Y(mai_mai_n404_));
  NA3        m388(.A(mai_mai_n404_), .B(mai_mai_n386_), .C(mai_mai_n354_), .Y(mai_mai_n405_));
  AOI210     m389(.A0(mai_mai_n336_), .A1(mai_mai_n25_), .B0(mai_mai_n405_), .Y(mai05));
  INV        m390(.A(x6), .Y(mai_mai_n409_));
  INV        m391(.A(mai_mai_n35_), .Y(mai_mai_n410_));
  INV        m392(.A(mai_mai_n77_), .Y(mai_mai_n411_));
  INV        m393(.A(mai_mai_n178_), .Y(mai_mai_n412_));
  INV        m394(.A(mai_mai_n209_), .Y(mai_mai_n413_));
  INV        m395(.A(mai_mai_n42_), .Y(mai_mai_n414_));
  INV        m396(.A(x4), .Y(mai_mai_n415_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  NOi21      u016(.An(men_men_n23_), .B(men_men_n30_), .Y(men00));
  NO2        u017(.A(x1), .B(x0), .Y(men_men_n34_));
  INV        u018(.A(x6), .Y(men_men_n35_));
  NO2        u019(.A(men_men_n35_), .B(men_men_n25_), .Y(men_men_n36_));
  AN2        u020(.A(x8), .B(x7), .Y(men_men_n37_));
  NA3        u021(.A(men_men_n37_), .B(men_men_n36_), .C(men_men_n34_), .Y(men_men_n38_));
  NA2        u022(.A(x4), .B(x3), .Y(men_men_n39_));
  AOI210     u023(.A0(men_men_n38_), .A1(men_men_n23_), .B0(men_men_n39_), .Y(men_men_n40_));
  NO2        u024(.A(x2), .B(x0), .Y(men_men_n41_));
  INV        u025(.A(x3), .Y(men_men_n42_));
  NO2        u026(.A(men_men_n42_), .B(men_men_n18_), .Y(men_men_n43_));
  INV        u027(.A(men_men_n43_), .Y(men_men_n44_));
  NO2        u028(.A(men_men_n36_), .B(x4), .Y(men_men_n45_));
  OAI210     u029(.A0(men_men_n45_), .A1(men_men_n44_), .B0(men_men_n41_), .Y(men_men_n46_));
  INV        u030(.A(x4), .Y(men_men_n47_));
  NO2        u031(.A(men_men_n47_), .B(men_men_n17_), .Y(men_men_n48_));
  NA2        u032(.A(men_men_n48_), .B(x2), .Y(men_men_n49_));
  OAI210     u033(.A0(men_men_n49_), .A1(men_men_n20_), .B0(men_men_n46_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n51_));
  AOI220     u035(.A0(men_men_n51_), .A1(men_men_n34_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n52_));
  INV        u036(.A(x2), .Y(men_men_n53_));
  NO2        u037(.A(men_men_n53_), .B(men_men_n17_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n42_), .B(men_men_n18_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  OAI210     u040(.A0(men_men_n52_), .A1(men_men_n32_), .B0(men_men_n56_), .Y(men_men_n57_));
  NO3        u041(.A(men_men_n57_), .B(men_men_n50_), .C(men_men_n40_), .Y(men01));
  NA2        u042(.A(x8), .B(x7), .Y(men_men_n59_));
  NA2        u043(.A(men_men_n42_), .B(x1), .Y(men_men_n60_));
  INV        u044(.A(x9), .Y(men_men_n61_));
  NO2        u045(.A(men_men_n61_), .B(men_men_n35_), .Y(men_men_n62_));
  INV        u046(.A(men_men_n62_), .Y(men_men_n63_));
  NO3        u047(.A(men_men_n63_), .B(men_men_n60_), .C(men_men_n59_), .Y(men_men_n64_));
  NO2        u048(.A(x7), .B(x6), .Y(men_men_n65_));
  NO2        u049(.A(men_men_n60_), .B(x5), .Y(men_men_n66_));
  NO2        u050(.A(x8), .B(x2), .Y(men_men_n67_));
  INV        u051(.A(men_men_n67_), .Y(men_men_n68_));
  NO2        u052(.A(men_men_n68_), .B(x1), .Y(men_men_n69_));
  OA210      u053(.A0(men_men_n69_), .A1(men_men_n66_), .B0(men_men_n65_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n43_), .A1(men_men_n25_), .B0(men_men_n53_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n55_), .A1(men_men_n20_), .B0(men_men_n71_), .Y(men_men_n72_));
  NAi31      u056(.An(x1), .B(x9), .C(x5), .Y(men_men_n73_));
  OAI220     u057(.A0(men_men_n73_), .A1(men_men_n42_), .B0(men_men_n72_), .B1(men_men_n70_), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n64_), .B0(x4), .Y(men_men_n75_));
  NA2        u059(.A(men_men_n47_), .B(x2), .Y(men_men_n76_));
  OAI210     u060(.A0(men_men_n76_), .A1(men_men_n55_), .B0(x0), .Y(men_men_n77_));
  NA2        u061(.A(x5), .B(x3), .Y(men_men_n78_));
  NO2        u062(.A(x8), .B(x6), .Y(men_men_n79_));
  NO4        u063(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n65_), .D(men_men_n53_), .Y(men_men_n80_));
  NAi21      u064(.An(x4), .B(x3), .Y(men_men_n81_));
  INV        u065(.A(men_men_n81_), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(men_men_n22_), .Y(men_men_n83_));
  NO2        u067(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u068(.A(men_men_n84_), .B(x3), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n83_), .C(men_men_n18_), .Y(men_men_n86_));
  NO3        u070(.A(men_men_n86_), .B(men_men_n80_), .C(men_men_n77_), .Y(men_men_n87_));
  NO4        u071(.A(men_men_n21_), .B(x6), .C(men_men_n42_), .D(x1), .Y(men_men_n88_));
  NA2        u072(.A(men_men_n61_), .B(men_men_n47_), .Y(men_men_n89_));
  INV        u073(.A(men_men_n89_), .Y(men_men_n90_));
  OAI210     u074(.A0(men_men_n88_), .A1(men_men_n66_), .B0(men_men_n90_), .Y(men_men_n91_));
  NA2        u075(.A(x3), .B(men_men_n18_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n25_), .Y(men_men_n93_));
  INV        u077(.A(x8), .Y(men_men_n94_));
  NA2        u078(.A(x2), .B(x1), .Y(men_men_n95_));
  AOI210     u079(.A0(men_men_n55_), .A1(men_men_n25_), .B0(men_men_n53_), .Y(men_men_n96_));
  OAI210     u080(.A0(men_men_n44_), .A1(men_men_n36_), .B0(men_men_n47_), .Y(men_men_n97_));
  NO3        u081(.A(men_men_n97_), .B(men_men_n96_), .C(men_men_n461_), .Y(men_men_n98_));
  NA2        u082(.A(x4), .B(men_men_n42_), .Y(men_men_n99_));
  NO2        u083(.A(men_men_n47_), .B(men_men_n53_), .Y(men_men_n100_));
  OAI210     u084(.A0(men_men_n100_), .A1(men_men_n42_), .B0(men_men_n18_), .Y(men_men_n101_));
  AOI210     u085(.A0(men_men_n99_), .A1(men_men_n51_), .B0(men_men_n101_), .Y(men_men_n102_));
  NO2        u086(.A(x3), .B(x2), .Y(men_men_n103_));
  NA2        u087(.A(men_men_n53_), .B(x1), .Y(men_men_n104_));
  OAI210     u088(.A0(men_men_n104_), .A1(men_men_n39_), .B0(men_men_n17_), .Y(men_men_n105_));
  NO4        u089(.A(men_men_n105_), .B(men_men_n103_), .C(men_men_n102_), .D(men_men_n98_), .Y(men_men_n106_));
  AO220      u090(.A0(men_men_n106_), .A1(men_men_n91_), .B0(men_men_n87_), .B1(men_men_n75_), .Y(men02));
  NO2        u091(.A(x3), .B(men_men_n53_), .Y(men_men_n108_));
  NO2        u092(.A(x8), .B(men_men_n18_), .Y(men_men_n109_));
  NA2        u093(.A(men_men_n53_), .B(men_men_n17_), .Y(men_men_n110_));
  NA2        u094(.A(men_men_n42_), .B(x0), .Y(men_men_n111_));
  OAI210     u095(.A0(men_men_n89_), .A1(men_men_n110_), .B0(men_men_n111_), .Y(men_men_n112_));
  AOI220     u096(.A0(men_men_n112_), .A1(men_men_n109_), .B0(men_men_n108_), .B1(x4), .Y(men_men_n113_));
  NO3        u097(.A(men_men_n113_), .B(x7), .C(x5), .Y(men_men_n114_));
  NA2        u098(.A(x9), .B(x2), .Y(men_men_n115_));
  OR2        u099(.A(x8), .B(x0), .Y(men_men_n116_));
  INV        u100(.A(men_men_n116_), .Y(men_men_n117_));
  NAi21      u101(.An(x2), .B(x8), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  OAI220     u103(.A0(men_men_n119_), .A1(men_men_n117_), .B0(men_men_n115_), .B1(x7), .Y(men_men_n120_));
  NO2        u104(.A(x4), .B(x1), .Y(men_men_n121_));
  NA3        u105(.A(men_men_n121_), .B(men_men_n120_), .C(men_men_n59_), .Y(men_men_n122_));
  NOi21      u106(.An(x0), .B(x1), .Y(men_men_n123_));
  NO3        u107(.A(x9), .B(x8), .C(x7), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x4), .Y(men_men_n125_));
  NAi21      u109(.An(x8), .B(x7), .Y(men_men_n126_));
  NO2        u110(.A(men_men_n126_), .B(men_men_n61_), .Y(men_men_n127_));
  AOI220     u111(.A0(men_men_n127_), .A1(men_men_n125_), .B0(men_men_n124_), .B1(men_men_n123_), .Y(men_men_n128_));
  AOI210     u112(.A0(men_men_n128_), .A1(men_men_n122_), .B0(men_men_n78_), .Y(men_men_n129_));
  NO2        u113(.A(x5), .B(men_men_n47_), .Y(men_men_n130_));
  NA2        u114(.A(x2), .B(men_men_n18_), .Y(men_men_n131_));
  NA2        u115(.A(men_men_n34_), .B(men_men_n130_), .Y(men_men_n132_));
  NAi21      u116(.An(x0), .B(x4), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n133_), .B(x1), .Y(men_men_n134_));
  NO2        u118(.A(x7), .B(x0), .Y(men_men_n135_));
  NO2        u119(.A(men_men_n84_), .B(men_men_n100_), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x3), .Y(men_men_n137_));
  OAI210     u121(.A0(men_men_n135_), .A1(men_men_n134_), .B0(men_men_n137_), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n21_), .B(men_men_n42_), .Y(men_men_n139_));
  NA2        u123(.A(x5), .B(x0), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n47_), .B(x2), .Y(men_men_n141_));
  NA3        u125(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n139_), .Y(men_men_n142_));
  NA4        u126(.A(men_men_n142_), .B(men_men_n138_), .C(men_men_n132_), .D(men_men_n35_), .Y(men_men_n143_));
  NO3        u127(.A(men_men_n143_), .B(men_men_n129_), .C(men_men_n114_), .Y(men_men_n144_));
  NO3        u128(.A(men_men_n78_), .B(men_men_n76_), .C(men_men_n24_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n146_));
  NO3        u130(.A(men_men_n464_), .B(men_men_n59_), .C(men_men_n61_), .Y(men_men_n147_));
  NA2        u131(.A(x7), .B(x3), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n99_), .B(x5), .Y(men_men_n149_));
  NO2        u133(.A(x9), .B(x7), .Y(men_men_n150_));
  NOi21      u134(.An(x8), .B(x0), .Y(men_men_n151_));
  OA210      u135(.A0(men_men_n150_), .A1(x1), .B0(men_men_n151_), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n42_), .B(x2), .Y(men_men_n153_));
  INV        u137(.A(x7), .Y(men_men_n154_));
  AOI220     u138(.A0(x1), .A1(men_men_n153_), .B0(men_men_n108_), .B1(men_men_n37_), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n25_), .B(x4), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n156_), .B(men_men_n125_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n157_), .B(men_men_n155_), .Y(men_men_n158_));
  AOI210     u142(.A0(men_men_n152_), .A1(men_men_n149_), .B0(men_men_n158_), .Y(men_men_n159_));
  OAI210     u143(.A0(men_men_n148_), .A1(men_men_n49_), .B0(men_men_n159_), .Y(men_men_n160_));
  NA2        u144(.A(x5), .B(x1), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n61_), .B(men_men_n94_), .Y(men_men_n162_));
  NAi21      u146(.An(x2), .B(x7), .Y(men_men_n163_));
  NO3        u147(.A(men_men_n163_), .B(men_men_n162_), .C(men_men_n47_), .Y(men_men_n164_));
  NA2        u148(.A(men_men_n164_), .B(men_men_n66_), .Y(men_men_n165_));
  NAi31      u149(.An(men_men_n78_), .B(men_men_n37_), .C(men_men_n34_), .Y(men_men_n166_));
  NA3        u150(.A(men_men_n166_), .B(men_men_n165_), .C(x6), .Y(men_men_n167_));
  NO4        u151(.A(men_men_n167_), .B(men_men_n160_), .C(men_men_n147_), .D(men_men_n145_), .Y(men_men_n168_));
  NO2        u152(.A(men_men_n168_), .B(men_men_n144_), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n140_), .B(men_men_n136_), .Y(men_men_n170_));
  NA2        u154(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n172_));
  NA3        u156(.A(men_men_n172_), .B(men_men_n171_), .C(men_men_n24_), .Y(men_men_n173_));
  AN2        u157(.A(men_men_n173_), .B(men_men_n141_), .Y(men_men_n174_));
  NA2        u158(.A(x8), .B(x0), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n154_), .B(men_men_n25_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n123_), .B(x4), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n177_), .B(men_men_n176_), .Y(men_men_n178_));
  AOI210     u162(.A0(men_men_n175_), .A1(men_men_n131_), .B0(men_men_n178_), .Y(men_men_n179_));
  NA2        u163(.A(x2), .B(x0), .Y(men_men_n180_));
  NA2        u164(.A(x4), .B(x1), .Y(men_men_n181_));
  NO3        u165(.A(men_men_n179_), .B(men_men_n174_), .C(men_men_n170_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n182_), .B(men_men_n42_), .Y(men_men_n183_));
  NO2        u167(.A(men_men_n173_), .B(men_men_n76_), .Y(men_men_n184_));
  INV        u168(.A(men_men_n130_), .Y(men_men_n185_));
  NO2        u169(.A(men_men_n104_), .B(men_men_n17_), .Y(men_men_n186_));
  AOI210     u170(.A0(men_men_n34_), .A1(men_men_n94_), .B0(men_men_n186_), .Y(men_men_n187_));
  NO3        u171(.A(men_men_n187_), .B(men_men_n185_), .C(x7), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n172_), .B(men_men_n136_), .Y(men_men_n189_));
  NO3        u173(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n184_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(x3), .Y(men_men_n191_));
  NO3        u175(.A(men_men_n191_), .B(men_men_n183_), .C(men_men_n169_), .Y(men03));
  NO2        u176(.A(men_men_n47_), .B(x3), .Y(men_men_n193_));
  NO2        u177(.A(x6), .B(men_men_n25_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n53_), .B(x1), .Y(men_men_n195_));
  OAI220     u179(.A0(men_men_n35_), .A1(men_men_n17_), .B0(men_men_n25_), .B1(men_men_n104_), .Y(men_men_n196_));
  NA2        u180(.A(men_men_n196_), .B(men_men_n193_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n78_), .B(x6), .Y(men_men_n198_));
  NA2        u182(.A(x6), .B(men_men_n25_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n199_), .B(x4), .Y(men_men_n200_));
  NO2        u184(.A(men_men_n18_), .B(x0), .Y(men_men_n201_));
  AO220      u185(.A0(men_men_n201_), .A1(men_men_n200_), .B0(men_men_n198_), .B1(men_men_n54_), .Y(men_men_n202_));
  NA2        u186(.A(men_men_n202_), .B(men_men_n61_), .Y(men_men_n203_));
  NA2        u187(.A(x3), .B(men_men_n17_), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n204_), .B(men_men_n199_), .Y(men_men_n205_));
  NA2        u189(.A(x9), .B(men_men_n53_), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n206_), .B(x4), .Y(men_men_n207_));
  NA2        u191(.A(men_men_n199_), .B(men_men_n81_), .Y(men_men_n208_));
  AOI210     u192(.A0(men_men_n25_), .A1(x3), .B0(men_men_n180_), .Y(men_men_n209_));
  AOI220     u193(.A0(men_men_n209_), .A1(men_men_n208_), .B0(men_men_n207_), .B1(men_men_n205_), .Y(men_men_n210_));
  NO3        u194(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n211_));
  NO2        u195(.A(x5), .B(x1), .Y(men_men_n212_));
  AOI220     u196(.A0(men_men_n212_), .A1(men_men_n17_), .B0(men_men_n103_), .B1(x5), .Y(men_men_n213_));
  NO2        u197(.A(men_men_n204_), .B(men_men_n171_), .Y(men_men_n214_));
  NO3        u198(.A(x3), .B(x2), .C(x1), .Y(men_men_n215_));
  NO2        u199(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n216_));
  OAI210     u200(.A0(men_men_n213_), .A1(men_men_n63_), .B0(men_men_n216_), .Y(men_men_n217_));
  AOI220     u201(.A0(men_men_n217_), .A1(men_men_n47_), .B0(men_men_n211_), .B1(men_men_n130_), .Y(men_men_n218_));
  NA4        u202(.A(men_men_n218_), .B(men_men_n210_), .C(men_men_n203_), .D(men_men_n197_), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n47_), .B(men_men_n42_), .Y(men_men_n220_));
  NA2        u204(.A(men_men_n220_), .B(men_men_n19_), .Y(men_men_n221_));
  NO2        u205(.A(x3), .B(men_men_n17_), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n222_), .B(x6), .Y(men_men_n223_));
  NOi21      u207(.An(men_men_n84_), .B(men_men_n223_), .Y(men_men_n224_));
  NA2        u208(.A(men_men_n61_), .B(men_men_n94_), .Y(men_men_n225_));
  NA3        u209(.A(men_men_n225_), .B(men_men_n222_), .C(x6), .Y(men_men_n226_));
  AOI210     u210(.A0(men_men_n226_), .A1(men_men_n224_), .B0(men_men_n154_), .Y(men_men_n227_));
  AO210      u211(.A0(men_men_n227_), .A1(men_men_n221_), .B0(men_men_n176_), .Y(men_men_n228_));
  NA2        u212(.A(men_men_n42_), .B(men_men_n53_), .Y(men_men_n229_));
  OAI210     u213(.A0(men_men_n229_), .A1(men_men_n25_), .B0(men_men_n172_), .Y(men_men_n230_));
  NO3        u214(.A(men_men_n181_), .B(men_men_n61_), .C(x6), .Y(men_men_n231_));
  AOI220     u215(.A0(men_men_n231_), .A1(men_men_n230_), .B0(men_men_n141_), .B1(men_men_n93_), .Y(men_men_n232_));
  NA2        u216(.A(x6), .B(men_men_n47_), .Y(men_men_n233_));
  OAI210     u217(.A0(men_men_n117_), .A1(men_men_n79_), .B0(x4), .Y(men_men_n234_));
  AOI210     u218(.A0(men_men_n234_), .A1(men_men_n233_), .B0(men_men_n78_), .Y(men_men_n235_));
  NO2        u219(.A(men_men_n61_), .B(x6), .Y(men_men_n236_));
  OAI210     u220(.A0(x1), .A1(men_men_n214_), .B0(men_men_n236_), .Y(men_men_n237_));
  NA2        u221(.A(men_men_n194_), .B(men_men_n134_), .Y(men_men_n238_));
  NA3        u222(.A(men_men_n204_), .B(men_men_n130_), .C(x6), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n94_), .A1(men_men_n35_), .B0(men_men_n66_), .Y(men_men_n240_));
  NA4        u224(.A(men_men_n240_), .B(men_men_n239_), .C(men_men_n238_), .D(men_men_n237_), .Y(men_men_n241_));
  OAI210     u225(.A0(men_men_n241_), .A1(men_men_n235_), .B0(x2), .Y(men_men_n242_));
  NA3        u226(.A(men_men_n242_), .B(men_men_n232_), .C(men_men_n228_), .Y(men_men_n243_));
  AOI210     u227(.A0(men_men_n219_), .A1(x8), .B0(men_men_n243_), .Y(men_men_n244_));
  NO2        u228(.A(men_men_n94_), .B(x3), .Y(men_men_n245_));
  NA2        u229(.A(men_men_n245_), .B(men_men_n200_), .Y(men_men_n246_));
  NO3        u230(.A(men_men_n92_), .B(men_men_n79_), .C(men_men_n25_), .Y(men_men_n247_));
  AOI210     u231(.A0(men_men_n223_), .A1(men_men_n156_), .B0(men_men_n247_), .Y(men_men_n248_));
  AOI210     u232(.A0(men_men_n248_), .A1(men_men_n246_), .B0(x2), .Y(men_men_n249_));
  NO2        u233(.A(x4), .B(men_men_n53_), .Y(men_men_n250_));
  AOI220     u234(.A0(men_men_n200_), .A1(men_men_n186_), .B0(men_men_n250_), .B1(men_men_n66_), .Y(men_men_n251_));
  NA2        u235(.A(men_men_n61_), .B(x6), .Y(men_men_n252_));
  NA3        u236(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n253_));
  AOI210     u237(.A0(men_men_n253_), .A1(men_men_n140_), .B0(men_men_n252_), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n42_), .B(men_men_n17_), .Y(men_men_n255_));
  NO2        u239(.A(men_men_n255_), .B(men_men_n25_), .Y(men_men_n256_));
  OAI210     u240(.A0(men_men_n256_), .A1(men_men_n254_), .B0(men_men_n121_), .Y(men_men_n257_));
  NA2        u241(.A(men_men_n204_), .B(x6), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n204_), .B(x6), .Y(men_men_n259_));
  NAi21      u243(.An(men_men_n162_), .B(men_men_n259_), .Y(men_men_n260_));
  NA3        u244(.A(men_men_n260_), .B(men_men_n258_), .C(men_men_n146_), .Y(men_men_n261_));
  NA4        u245(.A(men_men_n261_), .B(men_men_n257_), .C(men_men_n251_), .D(men_men_n154_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n194_), .B(men_men_n222_), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n140_), .B(men_men_n18_), .Y(men_men_n264_));
  NAi21      u248(.An(men_men_n264_), .B(men_men_n253_), .Y(men_men_n265_));
  NAi21      u249(.An(x1), .B(x4), .Y(men_men_n266_));
  AOI210     u250(.A0(x3), .A1(x2), .B0(men_men_n47_), .Y(men_men_n267_));
  OAI210     u251(.A0(men_men_n140_), .A1(x3), .B0(men_men_n267_), .Y(men_men_n268_));
  AOI210     u252(.A0(men_men_n268_), .A1(men_men_n266_), .B0(men_men_n265_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n269_), .B(men_men_n263_), .Y(men_men_n270_));
  NA2        u254(.A(men_men_n61_), .B(x2), .Y(men_men_n271_));
  NO2        u255(.A(men_men_n271_), .B(men_men_n263_), .Y(men_men_n272_));
  NO3        u256(.A(x9), .B(x6), .C(x0), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n104_), .B(men_men_n25_), .Y(men_men_n274_));
  NA2        u258(.A(x6), .B(x2), .Y(men_men_n275_));
  NO2        u259(.A(men_men_n275_), .B(men_men_n171_), .Y(men_men_n276_));
  AOI210     u260(.A0(men_men_n274_), .A1(men_men_n273_), .B0(men_men_n276_), .Y(men_men_n277_));
  OAI220     u261(.A0(men_men_n277_), .A1(men_men_n42_), .B0(men_men_n177_), .B1(men_men_n45_), .Y(men_men_n278_));
  OAI210     u262(.A0(men_men_n278_), .A1(men_men_n272_), .B0(men_men_n270_), .Y(men_men_n279_));
  NA2        u263(.A(x9), .B(men_men_n42_), .Y(men_men_n280_));
  NO2        u264(.A(men_men_n280_), .B(men_men_n199_), .Y(men_men_n281_));
  OR3        u265(.A(men_men_n281_), .B(men_men_n198_), .C(men_men_n149_), .Y(men_men_n282_));
  NA2        u266(.A(x4), .B(x0), .Y(men_men_n283_));
  NO3        u267(.A(men_men_n73_), .B(men_men_n283_), .C(x6), .Y(men_men_n284_));
  AOI210     u268(.A0(men_men_n282_), .A1(men_men_n41_), .B0(men_men_n284_), .Y(men_men_n285_));
  AOI210     u269(.A0(men_men_n285_), .A1(men_men_n279_), .B0(x8), .Y(men_men_n286_));
  INV        u270(.A(men_men_n252_), .Y(men_men_n287_));
  OAI210     u271(.A0(men_men_n264_), .A1(men_men_n212_), .B0(men_men_n287_), .Y(men_men_n288_));
  INV        u272(.A(men_men_n175_), .Y(men_men_n289_));
  AOI210     u273(.A0(men_men_n465_), .A1(men_men_n288_), .B0(men_men_n229_), .Y(men_men_n290_));
  NO4        u274(.A(men_men_n290_), .B(men_men_n286_), .C(men_men_n262_), .D(men_men_n249_), .Y(men_men_n291_));
  NO2        u275(.A(men_men_n162_), .B(x1), .Y(men_men_n292_));
  NO3        u276(.A(men_men_n292_), .B(x3), .C(men_men_n35_), .Y(men_men_n293_));
  OAI210     u277(.A0(men_men_n293_), .A1(men_men_n259_), .B0(x2), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n289_), .A1(x6), .B0(men_men_n43_), .Y(men_men_n295_));
  AOI210     u279(.A0(men_men_n295_), .A1(men_men_n294_), .B0(men_men_n185_), .Y(men_men_n296_));
  NOi21      u280(.An(men_men_n275_), .B(men_men_n17_), .Y(men_men_n297_));
  AOI210     u281(.A0(men_men_n35_), .A1(men_men_n53_), .B0(x0), .Y(men_men_n298_));
  NAi21      u282(.An(x4), .B(x0), .Y(men_men_n299_));
  NO3        u283(.A(men_men_n299_), .B(men_men_n43_), .C(x2), .Y(men_men_n300_));
  OAI210     u284(.A0(x6), .A1(men_men_n18_), .B0(men_men_n300_), .Y(men_men_n301_));
  NO2        u285(.A(x9), .B(x8), .Y(men_men_n302_));
  NA3        u286(.A(men_men_n302_), .B(men_men_n35_), .C(men_men_n53_), .Y(men_men_n303_));
  OAI210     u287(.A0(men_men_n298_), .A1(men_men_n297_), .B0(men_men_n303_), .Y(men_men_n304_));
  NA2        u288(.A(men_men_n304_), .B(men_men_n82_), .Y(men_men_n305_));
  AOI210     u289(.A0(men_men_n305_), .A1(men_men_n301_), .B0(men_men_n25_), .Y(men_men_n306_));
  NA3        u290(.A(men_men_n35_), .B(x1), .C(men_men_n17_), .Y(men_men_n307_));
  OAI210     u291(.A0(men_men_n298_), .A1(men_men_n297_), .B0(men_men_n307_), .Y(men_men_n308_));
  NA2        u292(.A(men_men_n35_), .B(men_men_n42_), .Y(men_men_n309_));
  OR2        u293(.A(men_men_n309_), .B(men_men_n283_), .Y(men_men_n310_));
  AN2        u294(.A(men_men_n308_), .B(men_men_n149_), .Y(men_men_n311_));
  NO3        u295(.A(men_men_n311_), .B(men_men_n306_), .C(men_men_n296_), .Y(men_men_n312_));
  OAI210     u296(.A0(men_men_n291_), .A1(men_men_n244_), .B0(men_men_n312_), .Y(men04));
  OAI210     u297(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n314_));
  NA3        u298(.A(men_men_n314_), .B(men_men_n273_), .C(men_men_n85_), .Y(men_men_n315_));
  NO2        u299(.A(x2), .B(x1), .Y(men_men_n316_));
  OAI210     u300(.A0(men_men_n255_), .A1(men_men_n316_), .B0(men_men_n35_), .Y(men_men_n317_));
  NO2        u301(.A(men_men_n316_), .B(men_men_n299_), .Y(men_men_n318_));
  AOI210     u302(.A0(men_men_n61_), .A1(x4), .B0(men_men_n110_), .Y(men_men_n319_));
  OAI210     u303(.A0(men_men_n319_), .A1(men_men_n318_), .B0(men_men_n245_), .Y(men_men_n320_));
  NO2        u304(.A(men_men_n271_), .B(men_men_n92_), .Y(men_men_n321_));
  NO2        u305(.A(men_men_n321_), .B(men_men_n35_), .Y(men_men_n322_));
  NA2        u306(.A(x9), .B(x0), .Y(men_men_n323_));
  AOI210     u307(.A0(men_men_n92_), .A1(men_men_n76_), .B0(men_men_n323_), .Y(men_men_n324_));
  NA2        u308(.A(men_men_n324_), .B(men_men_n94_), .Y(men_men_n325_));
  NA3        u309(.A(men_men_n325_), .B(men_men_n322_), .C(men_men_n320_), .Y(men_men_n326_));
  NA2        u310(.A(men_men_n326_), .B(men_men_n317_), .Y(men_men_n327_));
  NO2        u311(.A(men_men_n206_), .B(men_men_n111_), .Y(men_men_n328_));
  NO3        u312(.A(men_men_n252_), .B(men_men_n118_), .C(men_men_n18_), .Y(men_men_n329_));
  NO2        u313(.A(men_men_n329_), .B(men_men_n328_), .Y(men_men_n330_));
  NA3        u314(.A(men_men_n462_), .B(x6), .C(x3), .Y(men_men_n331_));
  NOi21      u315(.An(men_men_n151_), .B(men_men_n131_), .Y(men_men_n332_));
  AOI210     u316(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n333_));
  OAI220     u317(.A0(men_men_n333_), .A1(men_men_n309_), .B0(men_men_n271_), .B1(men_men_n307_), .Y(men_men_n334_));
  AOI210     u318(.A0(men_men_n332_), .A1(men_men_n62_), .B0(men_men_n334_), .Y(men_men_n335_));
  NA2        u319(.A(x2), .B(men_men_n17_), .Y(men_men_n336_));
  OAI210     u320(.A0(men_men_n104_), .A1(men_men_n17_), .B0(men_men_n336_), .Y(men_men_n337_));
  AOI220     u321(.A0(men_men_n337_), .A1(men_men_n79_), .B0(men_men_n321_), .B1(men_men_n94_), .Y(men_men_n338_));
  NA4        u322(.A(men_men_n338_), .B(men_men_n335_), .C(men_men_n331_), .D(men_men_n330_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n109_), .A1(x3), .B0(men_men_n300_), .Y(men_men_n340_));
  NA3        u324(.A(men_men_n225_), .B(men_men_n211_), .C(men_men_n84_), .Y(men_men_n341_));
  NA3        u325(.A(men_men_n341_), .B(men_men_n340_), .C(men_men_n154_), .Y(men_men_n342_));
  AOI210     u326(.A0(men_men_n339_), .A1(x4), .B0(men_men_n342_), .Y(men_men_n343_));
  NA3        u327(.A(men_men_n318_), .B(men_men_n206_), .C(men_men_n94_), .Y(men_men_n344_));
  NOi21      u328(.An(x4), .B(x0), .Y(men_men_n345_));
  XO2        u329(.A(x4), .B(x0), .Y(men_men_n346_));
  OAI210     u330(.A0(men_men_n346_), .A1(men_men_n115_), .B0(men_men_n266_), .Y(men_men_n347_));
  NA2        u331(.A(men_men_n347_), .B(x8), .Y(men_men_n348_));
  AOI210     u332(.A0(men_men_n348_), .A1(men_men_n344_), .B0(x3), .Y(men_men_n349_));
  INV        u333(.A(men_men_n95_), .Y(men_men_n350_));
  NO2        u334(.A(men_men_n94_), .B(x4), .Y(men_men_n351_));
  AOI220     u335(.A0(men_men_n351_), .A1(men_men_n43_), .B0(men_men_n125_), .B1(men_men_n350_), .Y(men_men_n352_));
  NO3        u336(.A(men_men_n346_), .B(men_men_n162_), .C(x2), .Y(men_men_n353_));
  NO3        u337(.A(men_men_n225_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n354_));
  NO2        u338(.A(men_men_n354_), .B(men_men_n353_), .Y(men_men_n355_));
  NA4        u339(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n221_), .D(x6), .Y(men_men_n356_));
  NO2        u340(.A(men_men_n299_), .B(men_men_n92_), .Y(men_men_n357_));
  NO2        u341(.A(men_men_n42_), .B(x0), .Y(men_men_n358_));
  OR2        u342(.A(men_men_n351_), .B(men_men_n358_), .Y(men_men_n359_));
  NO2        u343(.A(men_men_n151_), .B(men_men_n104_), .Y(men_men_n360_));
  AOI220     u344(.A0(men_men_n360_), .A1(men_men_n359_), .B0(men_men_n357_), .B1(men_men_n60_), .Y(men_men_n361_));
  NO2        u345(.A(men_men_n151_), .B(men_men_n81_), .Y(men_men_n362_));
  NO2        u346(.A(men_men_n34_), .B(x2), .Y(men_men_n363_));
  NOi21      u347(.An(men_men_n121_), .B(men_men_n27_), .Y(men_men_n364_));
  INV        u348(.A(men_men_n364_), .Y(men_men_n365_));
  OAI210     u349(.A0(men_men_n361_), .A1(men_men_n61_), .B0(men_men_n365_), .Y(men_men_n366_));
  OAI220     u350(.A0(men_men_n366_), .A1(x6), .B0(men_men_n356_), .B1(men_men_n349_), .Y(men_men_n367_));
  OAI210     u351(.A0(men_men_n62_), .A1(men_men_n47_), .B0(men_men_n41_), .Y(men_men_n368_));
  OAI210     u352(.A0(men_men_n368_), .A1(men_men_n94_), .B0(men_men_n310_), .Y(men_men_n369_));
  AOI210     u353(.A0(men_men_n369_), .A1(men_men_n18_), .B0(men_men_n154_), .Y(men_men_n370_));
  AO220      u354(.A0(men_men_n370_), .A1(men_men_n367_), .B0(men_men_n343_), .B1(men_men_n327_), .Y(men_men_n371_));
  NA2        u355(.A(men_men_n363_), .B(x6), .Y(men_men_n372_));
  NA2        u356(.A(men_men_n351_), .B(x0), .Y(men_men_n373_));
  NA2        u357(.A(men_men_n84_), .B(x6), .Y(men_men_n374_));
  OAI210     u358(.A0(men_men_n373_), .A1(x2), .B0(men_men_n374_), .Y(men_men_n375_));
  AOI220     u359(.A0(men_men_n375_), .A1(men_men_n372_), .B0(men_men_n215_), .B1(men_men_n48_), .Y(men_men_n376_));
  NA3        u360(.A(men_men_n376_), .B(men_men_n371_), .C(men_men_n315_), .Y(men_men_n377_));
  NA3        u361(.A(men_men_n463_), .B(men_men_n193_), .C(men_men_n154_), .Y(men_men_n378_));
  OAI210     u362(.A0(men_men_n28_), .A1(x1), .B0(men_men_n229_), .Y(men_men_n379_));
  AO220      u363(.A0(men_men_n379_), .A1(men_men_n150_), .B0(men_men_n108_), .B1(x4), .Y(men_men_n380_));
  NA3        u364(.A(x7), .B(x3), .C(x0), .Y(men_men_n381_));
  NA2        u365(.A(men_men_n220_), .B(x0), .Y(men_men_n382_));
  OAI220     u366(.A0(men_men_n382_), .A1(men_men_n206_), .B0(men_men_n381_), .B1(men_men_n350_), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n380_), .A1(men_men_n117_), .B0(men_men_n383_), .Y(men_men_n384_));
  AOI210     u368(.A0(men_men_n384_), .A1(men_men_n378_), .B0(men_men_n25_), .Y(men_men_n385_));
  NA3        u369(.A(men_men_n119_), .B(men_men_n220_), .C(x0), .Y(men_men_n386_));
  OAI210     u370(.A0(men_men_n193_), .A1(men_men_n67_), .B0(men_men_n201_), .Y(men_men_n387_));
  NA3        u371(.A(men_men_n195_), .B(men_men_n222_), .C(x8), .Y(men_men_n388_));
  AOI210     u372(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n25_), .Y(men_men_n389_));
  AOI210     u373(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n41_), .Y(men_men_n390_));
  NOi31      u374(.An(men_men_n390_), .B(men_men_n358_), .C(men_men_n181_), .Y(men_men_n391_));
  OAI210     u375(.A0(men_men_n391_), .A1(men_men_n389_), .B0(men_men_n150_), .Y(men_men_n392_));
  NAi31      u376(.An(men_men_n49_), .B(men_men_n292_), .C(men_men_n176_), .Y(men_men_n393_));
  NA3        u377(.A(men_men_n393_), .B(men_men_n392_), .C(men_men_n386_), .Y(men_men_n394_));
  OAI210     u378(.A0(men_men_n394_), .A1(men_men_n385_), .B0(x6), .Y(men_men_n395_));
  OAI210     u379(.A0(men_men_n162_), .A1(men_men_n47_), .B0(men_men_n135_), .Y(men_men_n396_));
  NA3        u380(.A(men_men_n54_), .B(men_men_n37_), .C(men_men_n31_), .Y(men_men_n397_));
  AOI220     u381(.A0(men_men_n397_), .A1(men_men_n396_), .B0(men_men_n39_), .B1(men_men_n32_), .Y(men_men_n398_));
  NO2        u382(.A(men_men_n154_), .B(x0), .Y(men_men_n399_));
  AOI220     u383(.A0(men_men_n399_), .A1(men_men_n220_), .B0(men_men_n193_), .B1(men_men_n154_), .Y(men_men_n400_));
  AOI210     u384(.A0(men_men_n127_), .A1(men_men_n250_), .B0(x1), .Y(men_men_n401_));
  OAI210     u385(.A0(men_men_n400_), .A1(x8), .B0(men_men_n401_), .Y(men_men_n402_));
  OAI210     u386(.A0(x2), .A1(x4), .B0(men_men_n163_), .Y(men_men_n403_));
  NA3        u387(.A(men_men_n403_), .B(men_men_n148_), .C(x9), .Y(men_men_n404_));
  NO4        u388(.A(men_men_n126_), .B(men_men_n299_), .C(x9), .D(x2), .Y(men_men_n405_));
  NOi21      u389(.An(men_men_n124_), .B(men_men_n180_), .Y(men_men_n406_));
  NO3        u390(.A(men_men_n406_), .B(men_men_n405_), .C(men_men_n18_), .Y(men_men_n407_));
  NO3        u391(.A(x9), .B(men_men_n154_), .C(x0), .Y(men_men_n408_));
  AOI220     u392(.A0(men_men_n408_), .A1(men_men_n245_), .B0(men_men_n362_), .B1(men_men_n154_), .Y(men_men_n409_));
  NA4        u393(.A(men_men_n409_), .B(men_men_n407_), .C(men_men_n404_), .D(men_men_n49_), .Y(men_men_n410_));
  OAI210     u394(.A0(men_men_n402_), .A1(men_men_n398_), .B0(men_men_n410_), .Y(men_men_n411_));
  NOi31      u395(.An(men_men_n399_), .B(men_men_n32_), .C(x8), .Y(men_men_n412_));
  AOI210     u396(.A0(men_men_n37_), .A1(x9), .B0(men_men_n133_), .Y(men_men_n413_));
  NO3        u397(.A(men_men_n413_), .B(men_men_n124_), .C(men_men_n42_), .Y(men_men_n414_));
  NOi31      u398(.An(x1), .B(x8), .C(x7), .Y(men_men_n415_));
  AOI220     u399(.A0(men_men_n415_), .A1(men_men_n345_), .B0(men_men_n125_), .B1(x3), .Y(men_men_n416_));
  AOI210     u400(.A0(men_men_n266_), .A1(men_men_n59_), .B0(men_men_n123_), .Y(men_men_n417_));
  OAI210     u401(.A0(men_men_n417_), .A1(x3), .B0(men_men_n416_), .Y(men_men_n418_));
  NO3        u402(.A(men_men_n418_), .B(men_men_n414_), .C(x2), .Y(men_men_n419_));
  OAI220     u403(.A0(men_men_n346_), .A1(men_men_n302_), .B0(men_men_n299_), .B1(men_men_n42_), .Y(men_men_n420_));
  AOI210     u404(.A0(x9), .A1(men_men_n47_), .B0(men_men_n381_), .Y(men_men_n421_));
  AOI220     u405(.A0(men_men_n421_), .A1(men_men_n94_), .B0(men_men_n420_), .B1(men_men_n154_), .Y(men_men_n422_));
  NO2        u406(.A(men_men_n422_), .B(men_men_n53_), .Y(men_men_n423_));
  NO3        u407(.A(men_men_n423_), .B(men_men_n419_), .C(men_men_n412_), .Y(men_men_n424_));
  AOI210     u408(.A0(men_men_n424_), .A1(men_men_n411_), .B0(men_men_n25_), .Y(men_men_n425_));
  NA4        u409(.A(men_men_n31_), .B(men_men_n94_), .C(x2), .D(men_men_n17_), .Y(men_men_n426_));
  NO3        u410(.A(men_men_n61_), .B(x4), .C(x1), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n67_), .B(men_men_n18_), .C(x0), .Y(men_men_n428_));
  AOI220     u412(.A0(men_men_n428_), .A1(men_men_n267_), .B0(men_men_n427_), .B1(men_men_n390_), .Y(men_men_n429_));
  NO2        u413(.A(men_men_n429_), .B(men_men_n103_), .Y(men_men_n430_));
  NO3        u414(.A(men_men_n271_), .B(men_men_n175_), .C(men_men_n39_), .Y(men_men_n431_));
  OAI210     u415(.A0(men_men_n431_), .A1(men_men_n430_), .B0(x7), .Y(men_men_n432_));
  NA2        u416(.A(men_men_n225_), .B(x7), .Y(men_men_n433_));
  NA3        u417(.A(men_men_n433_), .B(men_men_n153_), .C(men_men_n134_), .Y(men_men_n434_));
  NA3        u418(.A(men_men_n434_), .B(men_men_n432_), .C(men_men_n426_), .Y(men_men_n435_));
  OAI210     u419(.A0(men_men_n435_), .A1(men_men_n425_), .B0(men_men_n35_), .Y(men_men_n436_));
  NO2        u420(.A(men_men_n408_), .B(men_men_n201_), .Y(men_men_n437_));
  NO4        u421(.A(men_men_n437_), .B(men_men_n78_), .C(x4), .D(men_men_n53_), .Y(men_men_n438_));
  NA2        u422(.A(men_men_n255_), .B(men_men_n21_), .Y(men_men_n439_));
  NO2        u423(.A(men_men_n161_), .B(men_men_n135_), .Y(men_men_n440_));
  NA2        u424(.A(men_men_n440_), .B(men_men_n439_), .Y(men_men_n441_));
  AOI210     u425(.A0(men_men_n441_), .A1(men_men_n166_), .B0(men_men_n28_), .Y(men_men_n442_));
  NA3        u426(.A(x0), .B(x2), .C(men_men_n92_), .Y(men_men_n443_));
  NA2        u427(.A(men_men_n443_), .B(men_men_n176_), .Y(men_men_n444_));
  OAI220     u428(.A0(men_men_n280_), .A1(men_men_n68_), .B0(men_men_n161_), .B1(men_men_n42_), .Y(men_men_n445_));
  NA2        u429(.A(x3), .B(men_men_n53_), .Y(men_men_n446_));
  AOI210     u430(.A0(men_men_n163_), .A1(men_men_n27_), .B0(men_men_n73_), .Y(men_men_n447_));
  OAI210     u431(.A0(men_men_n150_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n448_));
  NO3        u432(.A(men_men_n415_), .B(x3), .C(men_men_n53_), .Y(men_men_n449_));
  AOI210     u433(.A0(men_men_n449_), .A1(men_men_n448_), .B0(men_men_n447_), .Y(men_men_n450_));
  OAI210     u434(.A0(x1), .A1(men_men_n446_), .B0(men_men_n450_), .Y(men_men_n451_));
  AOI220     u435(.A0(men_men_n451_), .A1(x0), .B0(men_men_n445_), .B1(men_men_n135_), .Y(men_men_n452_));
  AOI210     u436(.A0(men_men_n452_), .A1(men_men_n444_), .B0(men_men_n233_), .Y(men_men_n453_));
  NA2        u437(.A(x9), .B(x5), .Y(men_men_n454_));
  NO4        u438(.A(men_men_n104_), .B(men_men_n454_), .C(men_men_n59_), .D(men_men_n32_), .Y(men_men_n455_));
  NO4        u439(.A(men_men_n455_), .B(men_men_n453_), .C(men_men_n442_), .D(men_men_n438_), .Y(men_men_n456_));
  NA3        u440(.A(men_men_n456_), .B(men_men_n436_), .C(men_men_n395_), .Y(men_men_n457_));
  AOI210     u441(.A0(men_men_n377_), .A1(men_men_n25_), .B0(men_men_n457_), .Y(men05));
  INV        u442(.A(men_men_n26_), .Y(men_men_n461_));
  INV        u443(.A(men_men_n116_), .Y(men_men_n462_));
  INV        u444(.A(men_men_n17_), .Y(men_men_n463_));
  INV        u445(.A(x2), .Y(men_men_n464_));
  INV        u446(.A(men_men_n20_), .Y(men_men_n465_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule