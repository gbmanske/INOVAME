//Benchmark atmr_alu4_1266_0.0313

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n924_, ori_ori_n925_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1007_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1058_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NO2        o034(.A(i_1_), .B(i_6_), .Y(ori_ori_n57_));
  NA2        o035(.A(i_8_), .B(i_7_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n57_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n60_));
  NAi21      o038(.An(i_2_), .B(i_7_), .Y(ori_ori_n61_));
  INV        o039(.A(i_1_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NA3        o041(.A(ori_ori_n63_), .B(ori_ori_n61_), .C(ori_ori_n31_), .Y(ori_ori_n64_));
  NA2        o042(.A(i_1_), .B(i_10_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(i_6_), .Y(ori_ori_n66_));
  NAi31      o044(.An(ori_ori_n66_), .B(ori_ori_n64_), .C(ori_ori_n60_), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n69_));
  NA2        o047(.A(i_1_), .B(i_6_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n70_), .B(ori_ori_n25_), .Y(ori_ori_n71_));
  INV        o049(.A(i_0_), .Y(ori_ori_n72_));
  NAi21      o050(.An(i_5_), .B(i_10_), .Y(ori_ori_n73_));
  NA2        o051(.A(i_5_), .B(i_9_), .Y(ori_ori_n74_));
  AOI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n73_), .B0(ori_ori_n72_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n71_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n69_), .A1(ori_ori_n68_), .B0(ori_ori_n76_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n77_), .A1(ori_ori_n67_), .B0(i_0_), .Y(ori_ori_n78_));
  NA2        o056(.A(i_12_), .B(i_5_), .Y(ori_ori_n79_));
  NO2        o057(.A(i_3_), .B(i_9_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_3_), .B(i_7_), .Y(ori_ori_n81_));
  NO3        o059(.A(ori_ori_n81_), .B(ori_ori_n80_), .C(ori_ori_n62_), .Y(ori_ori_n82_));
  INV        o060(.A(i_6_), .Y(ori_ori_n83_));
  OR4        o061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n84_), .Y(ori_ori_n85_));
  NO2        o063(.A(i_2_), .B(i_7_), .Y(ori_ori_n86_));
  NO2        o064(.A(ori_ori_n85_), .B(ori_ori_n86_), .Y(ori_ori_n87_));
  NA2        o065(.A(ori_ori_n82_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  NAi21      o066(.An(i_6_), .B(i_10_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_6_), .B(i_9_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n62_), .Y(ori_ori_n91_));
  NA2        o069(.A(i_2_), .B(i_6_), .Y(ori_ori_n92_));
  NO3        o070(.A(ori_ori_n92_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(ori_ori_n91_), .Y(ori_ori_n94_));
  AOI210     o072(.A0(ori_ori_n94_), .A1(ori_ori_n88_), .B0(ori_ori_n79_), .Y(ori_ori_n95_));
  AN3        o073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n96_));
  NAi21      o074(.An(i_6_), .B(i_11_), .Y(ori_ori_n97_));
  NO2        o075(.A(i_5_), .B(i_8_), .Y(ori_ori_n98_));
  NOi21      o076(.An(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  AOI220     o077(.A0(ori_ori_n99_), .A1(ori_ori_n61_), .B0(ori_ori_n96_), .B1(ori_ori_n32_), .Y(ori_ori_n100_));
  INV        o078(.A(i_7_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n46_), .B(ori_ori_n101_), .Y(ori_ori_n102_));
  NO2        o080(.A(i_0_), .B(i_5_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n103_), .B(ori_ori_n83_), .Y(ori_ori_n104_));
  NA2        o082(.A(i_12_), .B(i_3_), .Y(ori_ori_n105_));
  INV        o083(.A(ori_ori_n105_), .Y(ori_ori_n106_));
  NA3        o084(.A(ori_ori_n106_), .B(ori_ori_n104_), .C(ori_ori_n102_), .Y(ori_ori_n107_));
  NAi21      o085(.An(i_7_), .B(i_11_), .Y(ori_ori_n108_));
  AN2        o086(.A(i_2_), .B(i_10_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n109_), .B(i_7_), .Y(ori_ori_n110_));
  OR2        o088(.A(ori_ori_n79_), .B(ori_ori_n57_), .Y(ori_ori_n111_));
  NO2        o089(.A(i_8_), .B(ori_ori_n101_), .Y(ori_ori_n112_));
  NO3        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .C(ori_ori_n110_), .Y(ori_ori_n113_));
  NA2        o091(.A(i_12_), .B(i_7_), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n62_), .B(ori_ori_n26_), .Y(ori_ori_n115_));
  NA2        o093(.A(ori_ori_n115_), .B(i_0_), .Y(ori_ori_n116_));
  NA2        o094(.A(i_11_), .B(i_12_), .Y(ori_ori_n117_));
  OAI210     o095(.A0(ori_ori_n116_), .A1(ori_ori_n114_), .B0(ori_ori_n117_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n118_), .B(ori_ori_n113_), .Y(ori_ori_n119_));
  NA3        o097(.A(ori_ori_n119_), .B(ori_ori_n107_), .C(ori_ori_n100_), .Y(ori_ori_n120_));
  NOi21      o098(.An(i_1_), .B(i_5_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n121_), .B(i_11_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n101_), .B(ori_ori_n37_), .Y(ori_ori_n123_));
  NA2        o101(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(ori_ori_n123_), .Y(ori_ori_n125_));
  NO2        o103(.A(ori_ori_n125_), .B(ori_ori_n46_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n90_), .B(ori_ori_n89_), .Y(ori_ori_n127_));
  NAi21      o105(.An(i_3_), .B(i_8_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n61_), .Y(ori_ori_n129_));
  NOi31      o107(.An(ori_ori_n129_), .B(ori_ori_n127_), .C(ori_ori_n126_), .Y(ori_ori_n130_));
  NO2        o108(.A(i_1_), .B(ori_ori_n83_), .Y(ori_ori_n131_));
  NO2        o109(.A(i_6_), .B(i_5_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(i_3_), .Y(ori_ori_n133_));
  AO210      o111(.A0(ori_ori_n133_), .A1(ori_ori_n47_), .B0(ori_ori_n131_), .Y(ori_ori_n134_));
  OAI220     o112(.A0(ori_ori_n134_), .A1(ori_ori_n108_), .B0(ori_ori_n130_), .B1(ori_ori_n122_), .Y(ori_ori_n135_));
  NO3        o113(.A(ori_ori_n135_), .B(ori_ori_n120_), .C(ori_ori_n95_), .Y(ori_ori_n136_));
  NA3        o114(.A(ori_ori_n136_), .B(ori_ori_n78_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o115(.A(ori_ori_n62_), .B(ori_ori_n37_), .Y(ori_ori_n138_));
  INV        o116(.A(i_6_), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n139_), .B(ori_ori_n138_), .Y(ori_ori_n140_));
  NA4        o118(.A(ori_ori_n140_), .B(ori_ori_n76_), .C(ori_ori_n68_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o119(.A(i_8_), .B(i_7_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n142_), .B(i_6_), .Y(ori_ori_n143_));
  NO2        o121(.A(i_12_), .B(i_13_), .Y(ori_ori_n144_));
  NAi21      o122(.An(i_5_), .B(i_11_), .Y(ori_ori_n145_));
  NOi21      o123(.An(ori_ori_n144_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NO2        o124(.A(i_0_), .B(i_1_), .Y(ori_ori_n147_));
  NA2        o125(.A(i_2_), .B(i_3_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n148_), .B(i_4_), .Y(ori_ori_n149_));
  NA3        o127(.A(ori_ori_n149_), .B(ori_ori_n147_), .C(ori_ori_n146_), .Y(ori_ori_n150_));
  AN2        o128(.A(ori_ori_n144_), .B(ori_ori_n80_), .Y(ori_ori_n151_));
  NA2        o129(.A(i_1_), .B(i_5_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n72_), .B(ori_ori_n46_), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n153_), .B(ori_ori_n36_), .Y(ori_ori_n154_));
  OR2        o132(.A(i_0_), .B(i_1_), .Y(ori_ori_n155_));
  NO3        o133(.A(ori_ori_n155_), .B(ori_ori_n79_), .C(i_13_), .Y(ori_ori_n156_));
  NAi32      o134(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n157_));
  NAi21      o135(.An(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  NOi21      o136(.An(i_4_), .B(i_10_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n159_), .B(ori_ori_n40_), .Y(ori_ori_n160_));
  NO2        o138(.A(i_3_), .B(i_5_), .Y(ori_ori_n161_));
  NO3        o139(.A(ori_ori_n72_), .B(i_2_), .C(i_1_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n162_), .B(ori_ori_n161_), .Y(ori_ori_n163_));
  OAI210     o141(.A0(ori_ori_n163_), .A1(ori_ori_n160_), .B0(ori_ori_n158_), .Y(ori_ori_n164_));
  INV        o142(.A(ori_ori_n164_), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n165_), .B(ori_ori_n143_), .Y(ori_ori_n166_));
  NOi21      o144(.An(i_4_), .B(i_9_), .Y(ori_ori_n167_));
  NOi21      o145(.An(i_11_), .B(i_13_), .Y(ori_ori_n168_));
  NA2        o146(.A(ori_ori_n168_), .B(ori_ori_n167_), .Y(ori_ori_n169_));
  NO2        o147(.A(i_4_), .B(i_5_), .Y(ori_ori_n170_));
  NAi21      o148(.An(i_12_), .B(i_11_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n171_), .B(i_13_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n72_), .B(ori_ori_n62_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n173_), .B(ori_ori_n46_), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n36_), .B(i_5_), .Y(ori_ori_n175_));
  NAi31      o153(.An(ori_ori_n175_), .B(ori_ori_n151_), .C(i_11_), .Y(ori_ori_n176_));
  NA2        o154(.A(i_3_), .B(i_5_), .Y(ori_ori_n177_));
  OR2        o155(.A(ori_ori_n177_), .B(ori_ori_n169_), .Y(ori_ori_n178_));
  AOI210     o156(.A0(ori_ori_n178_), .A1(ori_ori_n176_), .B0(ori_ori_n174_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n180_));
  NO2        o158(.A(i_13_), .B(i_10_), .Y(ori_ori_n181_));
  NA3        o159(.A(ori_ori_n181_), .B(ori_ori_n180_), .C(ori_ori_n44_), .Y(ori_ori_n182_));
  NO2        o160(.A(i_2_), .B(i_1_), .Y(ori_ori_n183_));
  NAi21      o161(.An(i_4_), .B(i_12_), .Y(ori_ori_n184_));
  INV        o162(.A(ori_ori_n179_), .Y(ori_ori_n185_));
  INV        o163(.A(i_8_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n186_), .B(i_7_), .Y(ori_ori_n187_));
  NA2        o165(.A(ori_ori_n187_), .B(i_6_), .Y(ori_ori_n188_));
  NO3        o166(.A(i_3_), .B(ori_ori_n83_), .C(ori_ori_n48_), .Y(ori_ori_n189_));
  NO3        o167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n190_));
  NO3        o168(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n191_));
  NO2        o169(.A(i_3_), .B(i_8_), .Y(ori_ori_n192_));
  NO3        o170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n193_));
  NA3        o171(.A(ori_ori_n193_), .B(ori_ori_n192_), .C(ori_ori_n40_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n103_), .B(ori_ori_n57_), .Y(ori_ori_n195_));
  INV        o173(.A(ori_ori_n195_), .Y(ori_ori_n196_));
  NO2        o174(.A(i_13_), .B(i_9_), .Y(ori_ori_n197_));
  NAi21      o175(.An(i_12_), .B(i_3_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n199_));
  NO3        o177(.A(i_0_), .B(i_2_), .C(ori_ori_n62_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n196_), .B(ori_ori_n194_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n201_), .B(i_7_), .Y(ori_ori_n202_));
  OAI220     o180(.A0(ori_ori_n202_), .A1(i_4_), .B0(ori_ori_n188_), .B1(ori_ori_n185_), .Y(ori_ori_n203_));
  NAi21      o181(.An(i_12_), .B(i_7_), .Y(ori_ori_n204_));
  NA3        o182(.A(i_13_), .B(ori_ori_n186_), .C(i_10_), .Y(ori_ori_n205_));
  NA2        o183(.A(i_0_), .B(i_5_), .Y(ori_ori_n206_));
  NAi31      o184(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n207_));
  NO2        o185(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n208_));
  NO2        o186(.A(ori_ori_n72_), .B(ori_ori_n26_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n46_), .B(ori_ori_n62_), .Y(ori_ori_n210_));
  NA3        o188(.A(ori_ori_n210_), .B(ori_ori_n209_), .C(ori_ori_n208_), .Y(ori_ori_n211_));
  INV        o189(.A(i_13_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_12_), .B(ori_ori_n212_), .Y(ori_ori_n213_));
  NA3        o191(.A(ori_ori_n213_), .B(ori_ori_n190_), .C(ori_ori_n189_), .Y(ori_ori_n214_));
  OAI210     o192(.A0(ori_ori_n211_), .A1(ori_ori_n207_), .B0(ori_ori_n214_), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n215_), .B(ori_ori_n142_), .Y(ori_ori_n216_));
  NO2        o194(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n217_));
  OR2        o195(.A(i_8_), .B(i_7_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n53_), .B(i_1_), .Y(ori_ori_n219_));
  INV        o197(.A(i_12_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n44_), .B(ori_ori_n220_), .Y(ori_ori_n221_));
  NO3        o199(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n222_));
  NA2        o200(.A(i_2_), .B(i_1_), .Y(ori_ori_n223_));
  NO3        o201(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n224_));
  NAi21      o202(.An(i_4_), .B(i_3_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n225_), .B(ori_ori_n74_), .Y(ori_ori_n226_));
  NO2        o204(.A(i_0_), .B(i_6_), .Y(ori_ori_n227_));
  NOi41      o205(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n223_), .B(ori_ori_n177_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_11_), .B(ori_ori_n212_), .Y(ori_ori_n230_));
  NOi21      o208(.An(i_1_), .B(i_6_), .Y(ori_ori_n231_));
  NAi21      o209(.An(i_3_), .B(i_7_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n220_), .B(i_9_), .Y(ori_ori_n233_));
  NA2        o211(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n234_));
  NAi21      o212(.An(i_7_), .B(i_10_), .Y(ori_ori_n235_));
  INV        o213(.A(ori_ori_n143_), .Y(ori_ori_n236_));
  NA2        o214(.A(ori_ori_n220_), .B(i_13_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n237_), .B(ori_ori_n74_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n238_), .B(ori_ori_n236_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n218_), .B(ori_ori_n37_), .Y(ori_ori_n240_));
  NA2        o218(.A(i_12_), .B(i_6_), .Y(ori_ori_n241_));
  OR2        o219(.A(i_13_), .B(i_9_), .Y(ori_ori_n242_));
  NO3        o220(.A(ori_ori_n242_), .B(ori_ori_n241_), .C(ori_ori_n48_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n225_), .B(i_2_), .Y(ori_ori_n244_));
  NA3        o222(.A(ori_ori_n244_), .B(ori_ori_n243_), .C(ori_ori_n44_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n230_), .B(i_9_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n234_), .B(ori_ori_n63_), .Y(ori_ori_n247_));
  OAI210     o225(.A0(ori_ori_n247_), .A1(ori_ori_n246_), .B0(ori_ori_n245_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n153_), .B(ori_ori_n62_), .Y(ori_ori_n249_));
  NO3        o227(.A(i_11_), .B(ori_ori_n212_), .C(ori_ori_n25_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n232_), .B(i_8_), .Y(ori_ori_n251_));
  NO2        o229(.A(i_6_), .B(ori_ori_n48_), .Y(ori_ori_n252_));
  NA3        o230(.A(ori_ori_n252_), .B(ori_ori_n251_), .C(ori_ori_n250_), .Y(ori_ori_n253_));
  NO3        o231(.A(ori_ori_n26_), .B(ori_ori_n83_), .C(i_5_), .Y(ori_ori_n254_));
  NA3        o232(.A(ori_ori_n254_), .B(ori_ori_n240_), .C(ori_ori_n213_), .Y(ori_ori_n255_));
  AOI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n253_), .B0(ori_ori_n249_), .Y(ori_ori_n256_));
  AOI210     o234(.A0(ori_ori_n248_), .A1(ori_ori_n240_), .B0(ori_ori_n256_), .Y(ori_ori_n257_));
  NA3        o235(.A(ori_ori_n257_), .B(ori_ori_n239_), .C(ori_ori_n216_), .Y(ori_ori_n258_));
  NO3        o236(.A(i_12_), .B(ori_ori_n212_), .C(ori_ori_n37_), .Y(ori_ori_n259_));
  INV        o237(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NA2        o238(.A(i_8_), .B(ori_ori_n101_), .Y(ori_ori_n261_));
  NO3        o239(.A(i_0_), .B(ori_ori_n46_), .C(i_1_), .Y(ori_ori_n262_));
  AOI220     o240(.A0(ori_ori_n262_), .A1(ori_ori_n189_), .B0(ori_ori_n161_), .B1(ori_ori_n219_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n263_), .B(ori_ori_n261_), .Y(ori_ori_n264_));
  NO3        o242(.A(i_0_), .B(i_2_), .C(ori_ori_n62_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n223_), .B(i_0_), .Y(ori_ori_n266_));
  AOI220     o244(.A0(ori_ori_n266_), .A1(ori_ori_n187_), .B0(ori_ori_n265_), .B1(ori_ori_n142_), .Y(ori_ori_n267_));
  NA2        o245(.A(ori_ori_n252_), .B(ori_ori_n26_), .Y(ori_ori_n268_));
  NO2        o246(.A(ori_ori_n268_), .B(ori_ori_n267_), .Y(ori_ori_n269_));
  NA2        o247(.A(i_0_), .B(i_1_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n270_), .B(i_2_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n58_), .B(i_6_), .Y(ori_ori_n272_));
  NO2        o250(.A(ori_ori_n163_), .B(ori_ori_n143_), .Y(ori_ori_n273_));
  NO3        o251(.A(ori_ori_n273_), .B(ori_ori_n269_), .C(ori_ori_n264_), .Y(ori_ori_n274_));
  NO2        o252(.A(i_3_), .B(i_10_), .Y(ori_ori_n275_));
  NO2        o253(.A(i_2_), .B(ori_ori_n101_), .Y(ori_ori_n276_));
  NA2        o254(.A(i_1_), .B(ori_ori_n36_), .Y(ori_ori_n277_));
  AN2        o255(.A(i_3_), .B(i_10_), .Y(ori_ori_n278_));
  NO2        o256(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n274_), .B(ori_ori_n260_), .Y(ori_ori_n281_));
  NO4        o259(.A(ori_ori_n281_), .B(ori_ori_n258_), .C(ori_ori_n203_), .D(ori_ori_n166_), .Y(ori_ori_n282_));
  NO3        o260(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n58_), .B(ori_ori_n83_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n266_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  NO3        o263(.A(i_6_), .B(ori_ori_n186_), .C(i_7_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n286_), .B(ori_ori_n190_), .Y(ori_ori_n287_));
  AOI210     o265(.A0(ori_ori_n287_), .A1(ori_ori_n285_), .B0(i_5_), .Y(ori_ori_n288_));
  NO2        o266(.A(i_2_), .B(i_3_), .Y(ori_ori_n289_));
  OR2        o267(.A(i_0_), .B(i_5_), .Y(ori_ori_n290_));
  NA3        o268(.A(ori_ori_n266_), .B(ori_ori_n161_), .C(ori_ori_n112_), .Y(ori_ori_n291_));
  NO2        o269(.A(ori_ori_n155_), .B(ori_ori_n46_), .Y(ori_ori_n292_));
  INV        o270(.A(ori_ori_n291_), .Y(ori_ori_n293_));
  OAI210     o271(.A0(ori_ori_n293_), .A1(ori_ori_n288_), .B0(i_4_), .Y(ori_ori_n294_));
  NO2        o272(.A(i_12_), .B(i_10_), .Y(ori_ori_n295_));
  NOi21      o273(.An(i_5_), .B(i_0_), .Y(ori_ori_n296_));
  NO2        o274(.A(i_2_), .B(ori_ori_n101_), .Y(ori_ori_n297_));
  NO4        o275(.A(ori_ori_n297_), .B(ori_ori_n277_), .C(ori_ori_n296_), .D(ori_ori_n128_), .Y(ori_ori_n298_));
  NA4        o276(.A(ori_ori_n81_), .B(ori_ori_n36_), .C(ori_ori_n83_), .D(i_8_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n298_), .B(ori_ori_n295_), .Y(ori_ori_n300_));
  NO2        o278(.A(i_6_), .B(i_8_), .Y(ori_ori_n301_));
  NOi21      o279(.An(i_0_), .B(i_2_), .Y(ori_ori_n302_));
  AN2        o280(.A(ori_ori_n302_), .B(ori_ori_n301_), .Y(ori_ori_n303_));
  NO2        o281(.A(i_1_), .B(i_7_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n300_), .B(ori_ori_n294_), .Y(ori_ori_n305_));
  NOi21      o283(.An(ori_ori_n152_), .B(ori_ori_n104_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n306_), .B(ori_ori_n124_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n307_), .B(i_3_), .Y(ori_ori_n308_));
  INV        o286(.A(ori_ori_n92_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n186_), .B(i_9_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n310_), .B(ori_ori_n195_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n311_), .B(ori_ori_n46_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n312_), .B(ori_ori_n269_), .Y(ori_ori_n313_));
  AOI210     o291(.A0(ori_ori_n313_), .A1(ori_ori_n308_), .B0(ori_ori_n160_), .Y(ori_ori_n314_));
  AOI210     o292(.A0(ori_ori_n305_), .A1(ori_ori_n283_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  NOi32      o293(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n316_));
  INV        o294(.A(ori_ori_n316_), .Y(ori_ori_n317_));
  NO2        o295(.A(ori_ori_n207_), .B(ori_ori_n157_), .Y(ori_ori_n318_));
  NO2        o296(.A(ori_ori_n157_), .B(ori_ori_n155_), .Y(ori_ori_n319_));
  NOi32      o297(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n320_));
  NAi21      o298(.An(i_6_), .B(i_1_), .Y(ori_ori_n321_));
  NA3        o299(.A(ori_ori_n321_), .B(ori_ori_n320_), .C(ori_ori_n46_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n322_), .B(i_0_), .Y(ori_ori_n323_));
  OR3        o301(.A(ori_ori_n323_), .B(ori_ori_n319_), .C(ori_ori_n318_), .Y(ori_ori_n324_));
  NO2        o302(.A(i_1_), .B(ori_ori_n101_), .Y(ori_ori_n325_));
  NAi21      o303(.An(i_3_), .B(i_4_), .Y(ori_ori_n326_));
  NO2        o304(.A(ori_ori_n326_), .B(i_9_), .Y(ori_ori_n327_));
  AN2        o305(.A(i_6_), .B(i_7_), .Y(ori_ori_n328_));
  OAI210     o306(.A0(ori_ori_n328_), .A1(ori_ori_n325_), .B0(ori_ori_n327_), .Y(ori_ori_n329_));
  NA2        o307(.A(i_2_), .B(i_7_), .Y(ori_ori_n330_));
  NO2        o308(.A(ori_ori_n326_), .B(i_10_), .Y(ori_ori_n331_));
  NA3        o309(.A(ori_ori_n331_), .B(ori_ori_n330_), .C(ori_ori_n227_), .Y(ori_ori_n332_));
  AOI210     o310(.A0(ori_ori_n332_), .A1(ori_ori_n329_), .B0(ori_ori_n180_), .Y(ori_ori_n333_));
  AOI210     o311(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n334_));
  OAI210     o312(.A0(ori_ori_n334_), .A1(ori_ori_n183_), .B0(ori_ori_n331_), .Y(ori_ori_n335_));
  AOI220     o313(.A0(ori_ori_n331_), .A1(ori_ori_n304_), .B0(ori_ori_n222_), .B1(ori_ori_n183_), .Y(ori_ori_n336_));
  AOI210     o314(.A0(ori_ori_n336_), .A1(ori_ori_n335_), .B0(i_5_), .Y(ori_ori_n337_));
  NO3        o315(.A(ori_ori_n337_), .B(ori_ori_n333_), .C(ori_ori_n324_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n338_), .B(ori_ori_n317_), .Y(ori_ori_n339_));
  NO2        o317(.A(ori_ori_n58_), .B(ori_ori_n25_), .Y(ori_ori_n340_));
  AN2        o318(.A(i_12_), .B(i_5_), .Y(ori_ori_n341_));
  NO2        o319(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n342_));
  NA2        o320(.A(ori_ori_n342_), .B(ori_ori_n341_), .Y(ori_ori_n343_));
  NO2        o321(.A(i_11_), .B(i_6_), .Y(ori_ori_n344_));
  NA3        o322(.A(ori_ori_n344_), .B(ori_ori_n292_), .C(ori_ori_n212_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n345_), .B(ori_ori_n343_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n225_), .B(i_5_), .Y(ori_ori_n347_));
  NO2        o325(.A(i_5_), .B(i_10_), .Y(ori_ori_n348_));
  AOI220     o326(.A0(ori_ori_n348_), .A1(ori_ori_n244_), .B0(ori_ori_n347_), .B1(ori_ori_n190_), .Y(ori_ori_n349_));
  NA2        o327(.A(ori_ori_n144_), .B(ori_ori_n45_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n350_), .B(ori_ori_n349_), .Y(ori_ori_n351_));
  OAI210     o329(.A0(ori_ori_n351_), .A1(ori_ori_n346_), .B0(ori_ori_n340_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n353_));
  NO2        o331(.A(ori_ori_n150_), .B(ori_ori_n83_), .Y(ori_ori_n354_));
  OAI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n346_), .B0(ori_ori_n353_), .Y(ori_ori_n355_));
  NO3        o333(.A(ori_ori_n83_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n356_));
  NA3        o334(.A(ori_ori_n275_), .B(ori_ori_n74_), .C(ori_ori_n54_), .Y(ori_ori_n357_));
  NO2        o335(.A(i_11_), .B(i_12_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n358_), .B(ori_ori_n36_), .Y(ori_ori_n359_));
  NO2        o337(.A(ori_ori_n357_), .B(ori_ori_n359_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n348_), .B(ori_ori_n220_), .Y(ori_ori_n361_));
  NAi21      o339(.An(i_13_), .B(i_0_), .Y(ori_ori_n362_));
  NO2        o340(.A(ori_ori_n362_), .B(ori_ori_n223_), .Y(ori_ori_n363_));
  NA2        o341(.A(ori_ori_n360_), .B(ori_ori_n363_), .Y(ori_ori_n364_));
  NA3        o342(.A(ori_ori_n364_), .B(ori_ori_n355_), .C(ori_ori_n352_), .Y(ori_ori_n365_));
  NA2        o343(.A(ori_ori_n44_), .B(ori_ori_n212_), .Y(ori_ori_n366_));
  NO2        o344(.A(i_0_), .B(i_11_), .Y(ori_ori_n367_));
  AN2        o345(.A(i_1_), .B(i_6_), .Y(ori_ori_n368_));
  NOi21      o346(.An(i_2_), .B(i_12_), .Y(ori_ori_n369_));
  NA2        o347(.A(ori_ori_n142_), .B(i_9_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n370_), .B(i_4_), .Y(ori_ori_n371_));
  NAi21      o349(.An(i_9_), .B(i_4_), .Y(ori_ori_n372_));
  OR2        o350(.A(i_13_), .B(i_10_), .Y(ori_ori_n373_));
  NO3        o351(.A(ori_ori_n373_), .B(ori_ori_n117_), .C(ori_ori_n372_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n169_), .B(ori_ori_n123_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n101_), .B(ori_ori_n25_), .Y(ori_ori_n376_));
  NA2        o354(.A(ori_ori_n259_), .B(ori_ori_n376_), .Y(ori_ori_n377_));
  NO2        o355(.A(ori_ori_n377_), .B(ori_ori_n306_), .Y(ori_ori_n378_));
  INV        o356(.A(ori_ori_n378_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n379_), .B(ori_ori_n26_), .Y(ori_ori_n380_));
  INV        o358(.A(ori_ori_n291_), .Y(ori_ori_n381_));
  NO2        o359(.A(ori_ori_n177_), .B(ori_ori_n83_), .Y(ori_ori_n382_));
  AOI220     o360(.A0(ori_ori_n382_), .A1(ori_ori_n271_), .B0(ori_ori_n254_), .B1(ori_ori_n200_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n383_), .B(ori_ori_n261_), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n384_), .B(ori_ori_n381_), .Y(ori_ori_n385_));
  NA2        o363(.A(ori_ori_n189_), .B(ori_ori_n96_), .Y(ori_ori_n386_));
  NA3        o364(.A(ori_ori_n292_), .B(ori_ori_n161_), .C(ori_ori_n83_), .Y(ori_ori_n387_));
  AOI210     o365(.A0(ori_ori_n387_), .A1(ori_ori_n386_), .B0(i_8_), .Y(ori_ori_n388_));
  NA3        o366(.A(ori_ori_n234_), .B(ori_ori_n63_), .C(i_2_), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n272_), .B(ori_ori_n219_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n390_), .B(ori_ori_n177_), .Y(ori_ori_n391_));
  NO2        o369(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n392_));
  NA3        o370(.A(ori_ori_n304_), .B(ori_ori_n303_), .C(ori_ori_n392_), .Y(ori_ori_n393_));
  INV        o371(.A(ori_ori_n393_), .Y(ori_ori_n394_));
  NO3        o372(.A(ori_ori_n394_), .B(ori_ori_n391_), .C(ori_ori_n388_), .Y(ori_ori_n395_));
  AOI210     o373(.A0(ori_ori_n395_), .A1(ori_ori_n385_), .B0(ori_ori_n246_), .Y(ori_ori_n396_));
  NO4        o374(.A(ori_ori_n396_), .B(ori_ori_n380_), .C(ori_ori_n365_), .D(ori_ori_n339_), .Y(ori_ori_n397_));
  NO2        o375(.A(ori_ori_n72_), .B(i_13_), .Y(ori_ori_n398_));
  NO2        o376(.A(i_10_), .B(i_9_), .Y(ori_ori_n399_));
  NAi21      o377(.An(i_12_), .B(i_8_), .Y(ori_ori_n400_));
  NO2        o378(.A(ori_ori_n400_), .B(i_3_), .Y(ori_ori_n401_));
  NO2        o379(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n402_), .B(ori_ori_n104_), .Y(ori_ori_n403_));
  NO2        o381(.A(ori_ori_n403_), .B(ori_ori_n194_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n280_), .B(i_0_), .Y(ori_ori_n405_));
  NO3        o383(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n406_));
  NA2        o384(.A(ori_ori_n241_), .B(ori_ori_n97_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n407_), .B(ori_ori_n406_), .Y(ori_ori_n408_));
  NA2        o386(.A(i_8_), .B(i_9_), .Y(ori_ori_n409_));
  AOI210     o387(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n410_));
  OR2        o388(.A(ori_ori_n410_), .B(ori_ori_n409_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n259_), .B(ori_ori_n195_), .Y(ori_ori_n412_));
  OAI220     o390(.A0(ori_ori_n412_), .A1(ori_ori_n411_), .B0(ori_ori_n408_), .B1(ori_ori_n405_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n230_), .B(ori_ori_n279_), .Y(ori_ori_n414_));
  NO3        o392(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n415_));
  INV        o393(.A(ori_ori_n415_), .Y(ori_ori_n416_));
  NA3        o394(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n417_));
  NA4        o395(.A(ori_ori_n145_), .B(ori_ori_n115_), .C(ori_ori_n79_), .D(ori_ori_n23_), .Y(ori_ori_n418_));
  OAI220     o396(.A0(ori_ori_n418_), .A1(ori_ori_n417_), .B0(ori_ori_n416_), .B1(ori_ori_n414_), .Y(ori_ori_n419_));
  NO3        o397(.A(ori_ori_n419_), .B(ori_ori_n413_), .C(ori_ori_n404_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n96_), .B(i_13_), .Y(ori_ori_n421_));
  NA2        o399(.A(ori_ori_n382_), .B(ori_ori_n340_), .Y(ori_ori_n422_));
  NO2        o400(.A(i_2_), .B(i_13_), .Y(ori_ori_n423_));
  NO2        o401(.A(ori_ori_n422_), .B(ori_ori_n421_), .Y(ori_ori_n424_));
  NO3        o402(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n425_));
  NO2        o403(.A(i_6_), .B(i_7_), .Y(ori_ori_n426_));
  NO2        o404(.A(i_11_), .B(i_1_), .Y(ori_ori_n427_));
  NOi21      o405(.An(i_2_), .B(i_7_), .Y(ori_ori_n428_));
  NO2        o406(.A(i_3_), .B(ori_ori_n186_), .Y(ori_ori_n429_));
  NO2        o407(.A(i_6_), .B(i_10_), .Y(ori_ori_n430_));
  NA3        o408(.A(ori_ori_n228_), .B(ori_ori_n168_), .C(ori_ori_n132_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n432_));
  NO2        o410(.A(ori_ori_n155_), .B(i_3_), .Y(ori_ori_n433_));
  NAi31      o411(.An(ori_ori_n432_), .B(ori_ori_n433_), .C(ori_ori_n213_), .Y(ori_ori_n434_));
  NA3        o412(.A(ori_ori_n353_), .B(ori_ori_n173_), .C(ori_ori_n149_), .Y(ori_ori_n435_));
  NA3        o413(.A(ori_ori_n435_), .B(ori_ori_n434_), .C(ori_ori_n431_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n436_), .B(ori_ori_n424_), .Y(ori_ori_n437_));
  NA2        o415(.A(ori_ori_n406_), .B(ori_ori_n341_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n415_), .B(ori_ori_n348_), .Y(ori_ori_n439_));
  NO2        o417(.A(ori_ori_n439_), .B(ori_ori_n211_), .Y(ori_ori_n440_));
  NAi21      o418(.An(ori_ori_n205_), .B(ori_ori_n358_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n304_), .B(ori_ori_n206_), .Y(ori_ori_n442_));
  NO2        o420(.A(ori_ori_n442_), .B(ori_ori_n441_), .Y(ori_ori_n443_));
  NA2        o421(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n283_), .B(ori_ori_n222_), .Y(ori_ori_n445_));
  OAI220     o423(.A0(ori_ori_n445_), .A1(ori_ori_n389_), .B0(ori_ori_n444_), .B1(ori_ori_n421_), .Y(ori_ori_n446_));
  NO3        o424(.A(ori_ori_n446_), .B(ori_ori_n443_), .C(ori_ori_n440_), .Y(ori_ori_n447_));
  NA3        o425(.A(ori_ori_n447_), .B(ori_ori_n437_), .C(ori_ori_n420_), .Y(ori_ori_n448_));
  NA2        o426(.A(ori_ori_n122_), .B(ori_ori_n111_), .Y(ori_ori_n449_));
  AN2        o427(.A(ori_ori_n449_), .B(ori_ori_n406_), .Y(ori_ori_n450_));
  NA2        o428(.A(ori_ori_n450_), .B(ori_ori_n280_), .Y(ori_ori_n451_));
  NA2        o429(.A(ori_ori_n341_), .B(ori_ori_n212_), .Y(ori_ori_n452_));
  NA2        o430(.A(ori_ori_n316_), .B(ori_ori_n72_), .Y(ori_ori_n453_));
  NA2        o431(.A(ori_ori_n328_), .B(ori_ori_n320_), .Y(ori_ori_n454_));
  OR2        o432(.A(ori_ori_n452_), .B(ori_ori_n454_), .Y(ori_ori_n455_));
  NO2        o433(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n456_));
  AOI210     o434(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n374_), .Y(ori_ori_n457_));
  NA2        o435(.A(ori_ori_n457_), .B(ori_ori_n455_), .Y(ori_ori_n458_));
  INV        o436(.A(ori_ori_n458_), .Y(ori_ori_n459_));
  NA2        o437(.A(ori_ori_n234_), .B(ori_ori_n63_), .Y(ori_ori_n460_));
  OAI210     o438(.A0(i_8_), .A1(ori_ori_n460_), .B0(ori_ori_n134_), .Y(ori_ori_n461_));
  NA2        o439(.A(ori_ori_n461_), .B(ori_ori_n375_), .Y(ori_ori_n462_));
  NA3        o440(.A(ori_ori_n462_), .B(ori_ori_n459_), .C(ori_ori_n451_), .Y(ori_ori_n463_));
  NO2        o441(.A(i_12_), .B(ori_ori_n186_), .Y(ori_ori_n464_));
  NO2        o442(.A(i_8_), .B(i_7_), .Y(ori_ori_n465_));
  OAI210     o443(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(ori_ori_n466_));
  NA2        o444(.A(ori_ori_n466_), .B(ori_ori_n210_), .Y(ori_ori_n467_));
  NO2        o445(.A(ori_ori_n467_), .B(ori_ori_n225_), .Y(ori_ori_n468_));
  NA2        o446(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n469_));
  NO2        o447(.A(ori_ori_n469_), .B(i_6_), .Y(ori_ori_n470_));
  NA3        o448(.A(ori_ori_n470_), .B(ori_ori_n468_), .C(ori_ori_n465_), .Y(ori_ori_n471_));
  AOI220     o449(.A0(ori_ori_n382_), .A1(ori_ori_n292_), .B0(ori_ori_n229_), .B1(ori_ori_n227_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n472_), .B(ori_ori_n237_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n473_), .B(ori_ori_n240_), .Y(ori_ori_n474_));
  NA3        o452(.A(ori_ori_n278_), .B(ori_ori_n170_), .C(ori_ori_n96_), .Y(ori_ori_n475_));
  NO2        o453(.A(ori_ori_n208_), .B(ori_ori_n44_), .Y(ori_ori_n476_));
  NO2        o454(.A(ori_ori_n155_), .B(i_5_), .Y(ori_ori_n477_));
  NA3        o455(.A(ori_ori_n477_), .B(ori_ori_n366_), .C(ori_ori_n289_), .Y(ori_ori_n478_));
  OAI210     o456(.A0(ori_ori_n478_), .A1(ori_ori_n476_), .B0(ori_ori_n475_), .Y(ori_ori_n479_));
  NA2        o457(.A(ori_ori_n479_), .B(ori_ori_n415_), .Y(ori_ori_n480_));
  NA3        o458(.A(ori_ori_n480_), .B(ori_ori_n474_), .C(ori_ori_n471_), .Y(ori_ori_n481_));
  AOI210     o459(.A0(ori_ori_n321_), .A1(ori_ori_n46_), .B0(ori_ori_n325_), .Y(ori_ori_n482_));
  NA2        o460(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n483_));
  NA3        o461(.A(ori_ori_n464_), .B(ori_ori_n250_), .C(ori_ori_n483_), .Y(ori_ori_n484_));
  NO2        o462(.A(ori_ori_n482_), .B(ori_ori_n484_), .Y(ori_ori_n485_));
  INV        o463(.A(ori_ori_n485_), .Y(ori_ori_n486_));
  NO3        o464(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n487_));
  NO2        o465(.A(ori_ori_n218_), .B(ori_ori_n36_), .Y(ori_ori_n488_));
  NO2        o466(.A(ori_ori_n373_), .B(i_1_), .Y(ori_ori_n489_));
  NOi31      o467(.An(ori_ori_n489_), .B(ori_ori_n407_), .C(ori_ori_n72_), .Y(ori_ori_n490_));
  AN4        o468(.A(ori_ori_n490_), .B(ori_ori_n371_), .C(i_3_), .D(i_2_), .Y(ori_ori_n491_));
  INV        o469(.A(ori_ori_n491_), .Y(ori_ori_n492_));
  NOi21      o470(.An(i_10_), .B(i_6_), .Y(ori_ori_n493_));
  NO2        o471(.A(ori_ori_n83_), .B(ori_ori_n25_), .Y(ori_ori_n494_));
  AOI220     o472(.A0(ori_ori_n259_), .A1(ori_ori_n494_), .B0(ori_ori_n250_), .B1(ori_ori_n493_), .Y(ori_ori_n495_));
  NO2        o473(.A(ori_ori_n495_), .B(ori_ori_n405_), .Y(ori_ori_n496_));
  NO2        o474(.A(ori_ori_n114_), .B(ori_ori_n23_), .Y(ori_ori_n497_));
  NA2        o475(.A(ori_ori_n286_), .B(ori_ori_n162_), .Y(ori_ori_n498_));
  AOI220     o476(.A0(ori_ori_n498_), .A1(ori_ori_n390_), .B0(ori_ori_n178_), .B1(ori_ori_n176_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n190_), .B(ori_ori_n37_), .Y(ori_ori_n500_));
  NOi31      o478(.An(ori_ori_n146_), .B(ori_ori_n500_), .C(ori_ori_n299_), .Y(ori_ori_n501_));
  NO3        o479(.A(ori_ori_n501_), .B(ori_ori_n499_), .C(ori_ori_n496_), .Y(ori_ori_n502_));
  NO2        o480(.A(ori_ori_n453_), .B(ori_ori_n336_), .Y(ori_ori_n503_));
  INV        o481(.A(ori_ori_n289_), .Y(ori_ori_n504_));
  NO2        o482(.A(i_12_), .B(ori_ori_n83_), .Y(ori_ori_n505_));
  NA3        o483(.A(ori_ori_n505_), .B(ori_ori_n250_), .C(ori_ori_n483_), .Y(ori_ori_n506_));
  NA3        o484(.A(ori_ori_n344_), .B(ori_ori_n259_), .C(ori_ori_n206_), .Y(ori_ori_n507_));
  AOI210     o485(.A0(ori_ori_n507_), .A1(ori_ori_n506_), .B0(ori_ori_n504_), .Y(ori_ori_n508_));
  OR2        o486(.A(i_2_), .B(i_5_), .Y(ori_ori_n509_));
  OR2        o487(.A(ori_ori_n509_), .B(ori_ori_n368_), .Y(ori_ori_n510_));
  NA2        o488(.A(ori_ori_n330_), .B(ori_ori_n227_), .Y(ori_ori_n511_));
  AOI210     o489(.A0(ori_ori_n511_), .A1(ori_ori_n510_), .B0(ori_ori_n441_), .Y(ori_ori_n512_));
  NO3        o490(.A(ori_ori_n512_), .B(ori_ori_n508_), .C(ori_ori_n503_), .Y(ori_ori_n513_));
  NA4        o491(.A(ori_ori_n513_), .B(ori_ori_n502_), .C(ori_ori_n492_), .D(ori_ori_n486_), .Y(ori_ori_n514_));
  NO4        o492(.A(ori_ori_n514_), .B(ori_ori_n481_), .C(ori_ori_n463_), .D(ori_ori_n448_), .Y(ori_ori_n515_));
  NA4        o493(.A(ori_ori_n515_), .B(ori_ori_n397_), .C(ori_ori_n315_), .D(ori_ori_n282_), .Y(ori7));
  NO2        o494(.A(ori_ori_n92_), .B(ori_ori_n54_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n108_), .B(ori_ori_n89_), .Y(ori_ori_n518_));
  NA2        o496(.A(ori_ori_n342_), .B(ori_ori_n518_), .Y(ori_ori_n519_));
  NA2        o497(.A(ori_ori_n430_), .B(ori_ori_n81_), .Y(ori_ori_n520_));
  NA2        o498(.A(i_11_), .B(ori_ori_n186_), .Y(ori_ori_n521_));
  INV        o499(.A(ori_ori_n519_), .Y(ori_ori_n522_));
  NA3        o500(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n523_));
  NO2        o501(.A(ori_ori_n220_), .B(i_4_), .Y(ori_ori_n524_));
  NA2        o502(.A(ori_ori_n524_), .B(i_8_), .Y(ori_ori_n525_));
  NO2        o503(.A(ori_ori_n105_), .B(ori_ori_n523_), .Y(ori_ori_n526_));
  NA2        o504(.A(i_2_), .B(ori_ori_n83_), .Y(ori_ori_n527_));
  OAI210     o505(.A0(ori_ori_n86_), .A1(ori_ori_n192_), .B0(ori_ori_n193_), .Y(ori_ori_n528_));
  NO2        o506(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n529_));
  NA2        o507(.A(i_4_), .B(i_8_), .Y(ori_ori_n530_));
  AOI210     o508(.A0(ori_ori_n530_), .A1(ori_ori_n278_), .B0(ori_ori_n529_), .Y(ori_ori_n531_));
  OAI220     o509(.A0(ori_ori_n531_), .A1(ori_ori_n527_), .B0(ori_ori_n528_), .B1(i_13_), .Y(ori_ori_n532_));
  NO4        o510(.A(ori_ori_n532_), .B(ori_ori_n526_), .C(ori_ori_n522_), .D(ori_ori_n517_), .Y(ori_ori_n533_));
  AOI210     o511(.A0(ori_ori_n128_), .A1(ori_ori_n61_), .B0(i_10_), .Y(ori_ori_n534_));
  AOI210     o512(.A0(ori_ori_n534_), .A1(ori_ori_n220_), .B0(ori_ori_n159_), .Y(ori_ori_n535_));
  OR2        o513(.A(i_6_), .B(i_10_), .Y(ori_ori_n536_));
  OR3        o514(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n537_));
  INV        o515(.A(ori_ori_n191_), .Y(ori_ori_n538_));
  OR2        o516(.A(ori_ori_n535_), .B(ori_ori_n242_), .Y(ori_ori_n539_));
  AOI210     o517(.A0(ori_ori_n539_), .A1(ori_ori_n533_), .B0(ori_ori_n62_), .Y(ori_ori_n540_));
  NOi21      o518(.An(i_11_), .B(i_7_), .Y(ori_ori_n541_));
  AO210      o519(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n542_));
  NO2        o520(.A(ori_ori_n542_), .B(ori_ori_n541_), .Y(ori_ori_n543_));
  NA2        o521(.A(ori_ori_n543_), .B(ori_ori_n197_), .Y(ori_ori_n544_));
  NA3        o522(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n545_));
  NAi31      o523(.An(ori_ori_n545_), .B(ori_ori_n204_), .C(i_11_), .Y(ori_ori_n546_));
  AOI210     o524(.A0(ori_ori_n546_), .A1(ori_ori_n544_), .B0(ori_ori_n62_), .Y(ori_ori_n547_));
  NA2        o525(.A(ori_ori_n85_), .B(ori_ori_n62_), .Y(ori_ori_n548_));
  AO210      o526(.A0(ori_ori_n548_), .A1(ori_ori_n336_), .B0(ori_ori_n41_), .Y(ori_ori_n549_));
  NO3        o527(.A(ori_ori_n235_), .B(ori_ori_n198_), .C(ori_ori_n521_), .Y(ori_ori_n550_));
  OAI210     o528(.A0(ori_ori_n550_), .A1(ori_ori_n213_), .B0(ori_ori_n62_), .Y(ori_ori_n551_));
  NA2        o529(.A(ori_ori_n369_), .B(ori_ori_n31_), .Y(ori_ori_n552_));
  OR2        o530(.A(ori_ori_n198_), .B(ori_ori_n108_), .Y(ori_ori_n553_));
  NA2        o531(.A(ori_ori_n553_), .B(ori_ori_n552_), .Y(ori_ori_n554_));
  NO2        o532(.A(i_1_), .B(i_4_), .Y(ori_ori_n555_));
  NA2        o533(.A(ori_ori_n555_), .B(ori_ori_n554_), .Y(ori_ori_n556_));
  NO2        o534(.A(i_1_), .B(i_12_), .Y(ori_ori_n557_));
  NA3        o535(.A(ori_ori_n557_), .B(ori_ori_n109_), .C(ori_ori_n24_), .Y(ori_ori_n558_));
  BUFFER     o536(.A(ori_ori_n558_), .Y(ori_ori_n559_));
  NA4        o537(.A(ori_ori_n559_), .B(ori_ori_n556_), .C(ori_ori_n551_), .D(ori_ori_n549_), .Y(ori_ori_n560_));
  OAI210     o538(.A0(ori_ori_n560_), .A1(ori_ori_n547_), .B0(i_6_), .Y(ori_ori_n561_));
  NO2        o539(.A(ori_ori_n545_), .B(ori_ori_n108_), .Y(ori_ori_n562_));
  NA2        o540(.A(ori_ori_n562_), .B(ori_ori_n505_), .Y(ori_ori_n563_));
  NO2        o541(.A(ori_ori_n220_), .B(ori_ori_n83_), .Y(ori_ori_n564_));
  NO2        o542(.A(ori_ori_n564_), .B(i_11_), .Y(ori_ori_n565_));
  NA2        o543(.A(ori_ori_n563_), .B(ori_ori_n408_), .Y(ori_ori_n566_));
  NO3        o544(.A(ori_ori_n536_), .B(ori_ori_n218_), .C(ori_ori_n23_), .Y(ori_ori_n567_));
  NA3        o545(.A(ori_ori_n465_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n568_));
  INV        o546(.A(i_2_), .Y(ori_ori_n569_));
  NA2        o547(.A(ori_ori_n138_), .B(i_9_), .Y(ori_ori_n570_));
  NO2        o548(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n571_));
  NO2        o549(.A(ori_ori_n570_), .B(ori_ori_n569_), .Y(ori_ori_n572_));
  AOI210     o550(.A0(ori_ori_n427_), .A1(ori_ori_n376_), .B0(ori_ori_n224_), .Y(ori_ori_n573_));
  NO2        o551(.A(ori_ori_n573_), .B(ori_ori_n527_), .Y(ori_ori_n574_));
  NAi21      o552(.An(ori_ori_n568_), .B(ori_ori_n91_), .Y(ori_ori_n575_));
  NA2        o553(.A(ori_ori_n571_), .B(ori_ori_n241_), .Y(ori_ori_n576_));
  NO2        o554(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n577_), .B(ori_ori_n24_), .Y(ori_ori_n578_));
  OAI210     o556(.A0(ori_ori_n578_), .A1(ori_ori_n576_), .B0(ori_ori_n575_), .Y(ori_ori_n579_));
  OR3        o557(.A(ori_ori_n579_), .B(ori_ori_n574_), .C(ori_ori_n572_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n580_), .B(ori_ori_n566_), .Y(ori_ori_n581_));
  NO2        o559(.A(ori_ori_n220_), .B(ori_ori_n101_), .Y(ori_ori_n582_));
  NO2        o560(.A(ori_ori_n582_), .B(ori_ori_n541_), .Y(ori_ori_n583_));
  NA2        o561(.A(ori_ori_n583_), .B(i_1_), .Y(ori_ori_n584_));
  NO2        o562(.A(ori_ori_n584_), .B(ori_ori_n537_), .Y(ori_ori_n585_));
  NO2        o563(.A(ori_ori_n372_), .B(ori_ori_n83_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n585_), .B(ori_ori_n46_), .Y(ori_ori_n587_));
  NA2        o565(.A(i_3_), .B(ori_ori_n186_), .Y(ori_ori_n588_));
  NO2        o566(.A(ori_ori_n588_), .B(ori_ori_n114_), .Y(ori_ori_n589_));
  AN2        o567(.A(ori_ori_n589_), .B(ori_ori_n470_), .Y(ori_ori_n590_));
  NO2        o568(.A(ori_ori_n218_), .B(ori_ori_n44_), .Y(ori_ori_n591_));
  NO3        o569(.A(ori_ori_n591_), .B(ori_ori_n280_), .C(ori_ori_n221_), .Y(ori_ori_n592_));
  NO2        o570(.A(ori_ori_n117_), .B(ori_ori_n37_), .Y(ori_ori_n593_));
  NO2        o571(.A(ori_ori_n593_), .B(i_6_), .Y(ori_ori_n594_));
  NO2        o572(.A(ori_ori_n83_), .B(i_9_), .Y(ori_ori_n595_));
  NO2        o573(.A(ori_ori_n595_), .B(ori_ori_n62_), .Y(ori_ori_n596_));
  NO2        o574(.A(ori_ori_n596_), .B(ori_ori_n557_), .Y(ori_ori_n597_));
  NO4        o575(.A(ori_ori_n597_), .B(ori_ori_n594_), .C(ori_ori_n592_), .D(i_4_), .Y(ori_ori_n598_));
  NA2        o576(.A(i_1_), .B(i_3_), .Y(ori_ori_n599_));
  NO2        o577(.A(ori_ori_n409_), .B(ori_ori_n92_), .Y(ori_ori_n600_));
  AOI210     o578(.A0(ori_ori_n591_), .A1(ori_ori_n493_), .B0(ori_ori_n600_), .Y(ori_ori_n601_));
  NO2        o579(.A(ori_ori_n601_), .B(ori_ori_n599_), .Y(ori_ori_n602_));
  NO3        o580(.A(ori_ori_n602_), .B(ori_ori_n598_), .C(ori_ori_n590_), .Y(ori_ori_n603_));
  NA4        o581(.A(ori_ori_n603_), .B(ori_ori_n587_), .C(ori_ori_n581_), .D(ori_ori_n561_), .Y(ori_ori_n604_));
  NO3        o582(.A(i_11_), .B(i_3_), .C(i_7_), .Y(ori_ori_n605_));
  NOi21      o583(.An(ori_ori_n605_), .B(i_10_), .Y(ori_ori_n606_));
  OA210      o584(.A0(ori_ori_n606_), .A1(ori_ori_n228_), .B0(ori_ori_n83_), .Y(ori_ori_n607_));
  NO3        o585(.A(ori_ori_n428_), .B(ori_ori_n530_), .C(ori_ori_n83_), .Y(ori_ori_n608_));
  NA2        o586(.A(ori_ori_n608_), .B(ori_ori_n25_), .Y(ori_ori_n609_));
  INV        o587(.A(ori_ori_n609_), .Y(ori_ori_n610_));
  OAI210     o588(.A0(ori_ori_n610_), .A1(ori_ori_n607_), .B0(i_1_), .Y(ori_ori_n611_));
  AOI210     o589(.A0(ori_ori_n241_), .A1(ori_ori_n97_), .B0(i_1_), .Y(ori_ori_n612_));
  NO2        o590(.A(ori_ori_n326_), .B(i_2_), .Y(ori_ori_n613_));
  NA2        o591(.A(ori_ori_n613_), .B(ori_ori_n612_), .Y(ori_ori_n614_));
  AOI210     o592(.A0(ori_ori_n614_), .A1(ori_ori_n611_), .B0(i_13_), .Y(ori_ori_n615_));
  OR2        o593(.A(i_11_), .B(i_7_), .Y(ori_ori_n616_));
  NA3        o594(.A(ori_ori_n616_), .B(ori_ori_n106_), .C(ori_ori_n138_), .Y(ori_ori_n617_));
  AOI220     o595(.A0(ori_ori_n423_), .A1(ori_ori_n159_), .B0(ori_ori_n402_), .B1(ori_ori_n138_), .Y(ori_ori_n618_));
  OAI210     o596(.A0(ori_ori_n618_), .A1(ori_ori_n44_), .B0(ori_ori_n617_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n620_));
  NO2        o598(.A(ori_ori_n428_), .B(ori_ori_n24_), .Y(ori_ori_n621_));
  NA2        o599(.A(ori_ori_n621_), .B(ori_ori_n586_), .Y(ori_ori_n622_));
  OAI220     o600(.A0(ori_ori_n622_), .A1(ori_ori_n41_), .B0(ori_ori_n924_), .B1(ori_ori_n92_), .Y(ori_ori_n623_));
  AOI210     o601(.A0(ori_ori_n619_), .A1(ori_ori_n301_), .B0(ori_ori_n623_), .Y(ori_ori_n624_));
  NA2        o602(.A(ori_ori_n344_), .B(ori_ori_n571_), .Y(ori_ori_n625_));
  NO2        o603(.A(ori_ori_n625_), .B(ori_ori_n225_), .Y(ori_ori_n626_));
  AOI210     o604(.A0(ori_ori_n400_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n627_));
  NOi31      o605(.An(ori_ori_n627_), .B(ori_ori_n520_), .C(ori_ori_n44_), .Y(ori_ori_n628_));
  NA2        o606(.A(ori_ori_n127_), .B(i_13_), .Y(ori_ori_n629_));
  NO2        o607(.A(ori_ori_n629_), .B(ori_ori_n612_), .Y(ori_ori_n630_));
  NO3        o608(.A(ori_ori_n70_), .B(ori_ori_n32_), .C(ori_ori_n101_), .Y(ori_ori_n631_));
  NA2        o609(.A(ori_ori_n26_), .B(ori_ori_n186_), .Y(ori_ori_n632_));
  NA2        o610(.A(ori_ori_n632_), .B(i_7_), .Y(ori_ori_n633_));
  AOI220     o611(.A0(ori_ori_n344_), .A1(ori_ori_n571_), .B0(ori_ori_n91_), .B1(ori_ori_n102_), .Y(ori_ori_n634_));
  OAI220     o612(.A0(ori_ori_n634_), .A1(ori_ori_n525_), .B0(ori_ori_n925_), .B1(ori_ori_n538_), .Y(ori_ori_n635_));
  NO4        o613(.A(ori_ori_n635_), .B(ori_ori_n630_), .C(ori_ori_n628_), .D(ori_ori_n626_), .Y(ori_ori_n636_));
  OR2        o614(.A(i_11_), .B(i_6_), .Y(ori_ori_n637_));
  NA3        o615(.A(ori_ori_n524_), .B(ori_ori_n632_), .C(i_7_), .Y(ori_ori_n638_));
  NO2        o616(.A(ori_ori_n638_), .B(ori_ori_n637_), .Y(ori_ori_n639_));
  NA3        o617(.A(ori_ori_n369_), .B(ori_ori_n529_), .C(ori_ori_n97_), .Y(ori_ori_n640_));
  NA2        o618(.A(ori_ori_n565_), .B(i_13_), .Y(ori_ori_n641_));
  NA2        o619(.A(ori_ori_n102_), .B(ori_ori_n632_), .Y(ori_ori_n642_));
  NAi21      o620(.An(i_11_), .B(i_12_), .Y(ori_ori_n643_));
  NOi41      o621(.An(ori_ori_n110_), .B(ori_ori_n643_), .C(i_13_), .D(ori_ori_n83_), .Y(ori_ori_n644_));
  NO3        o622(.A(ori_ori_n428_), .B(ori_ori_n505_), .C(ori_ori_n530_), .Y(ori_ori_n645_));
  AOI220     o623(.A0(ori_ori_n645_), .A1(ori_ori_n283_), .B0(ori_ori_n644_), .B1(ori_ori_n642_), .Y(ori_ori_n646_));
  NA3        o624(.A(ori_ori_n646_), .B(ori_ori_n641_), .C(ori_ori_n640_), .Y(ori_ori_n647_));
  OAI210     o625(.A0(ori_ori_n647_), .A1(ori_ori_n639_), .B0(ori_ori_n62_), .Y(ori_ori_n648_));
  NO2        o626(.A(i_2_), .B(i_12_), .Y(ori_ori_n649_));
  NA2        o627(.A(ori_ori_n325_), .B(ori_ori_n649_), .Y(ori_ori_n650_));
  NO2        o628(.A(ori_ori_n128_), .B(i_2_), .Y(ori_ori_n651_));
  NA2        o629(.A(ori_ori_n651_), .B(ori_ori_n557_), .Y(ori_ori_n652_));
  NA2        o630(.A(ori_ori_n652_), .B(ori_ori_n650_), .Y(ori_ori_n653_));
  NA3        o631(.A(ori_ori_n653_), .B(ori_ori_n45_), .C(ori_ori_n212_), .Y(ori_ori_n654_));
  NA4        o632(.A(ori_ori_n654_), .B(ori_ori_n648_), .C(ori_ori_n636_), .D(ori_ori_n624_), .Y(ori_ori_n655_));
  OR4        o633(.A(ori_ori_n655_), .B(ori_ori_n615_), .C(ori_ori_n604_), .D(ori_ori_n540_), .Y(ori5));
  NA2        o634(.A(ori_ori_n583_), .B(ori_ori_n244_), .Y(ori_ori_n657_));
  AN2        o635(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n658_));
  NA3        o636(.A(ori_ori_n658_), .B(ori_ori_n649_), .C(ori_ori_n108_), .Y(ori_ori_n659_));
  NO2        o637(.A(ori_ori_n525_), .B(i_11_), .Y(ori_ori_n660_));
  NA2        o638(.A(ori_ori_n86_), .B(ori_ori_n660_), .Y(ori_ori_n661_));
  NA3        o639(.A(ori_ori_n661_), .B(ori_ori_n659_), .C(ori_ori_n657_), .Y(ori_ori_n662_));
  NO3        o640(.A(i_11_), .B(ori_ori_n220_), .C(i_13_), .Y(ori_ori_n663_));
  NO2        o641(.A(ori_ori_n124_), .B(ori_ori_n23_), .Y(ori_ori_n664_));
  NA2        o642(.A(i_12_), .B(i_8_), .Y(ori_ori_n665_));
  OAI210     o643(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n665_), .Y(ori_ori_n666_));
  INV        o644(.A(ori_ori_n399_), .Y(ori_ori_n667_));
  AOI220     o645(.A0(ori_ori_n289_), .A1(ori_ori_n497_), .B0(ori_ori_n666_), .B1(ori_ori_n664_), .Y(ori_ori_n668_));
  INV        o646(.A(ori_ori_n668_), .Y(ori_ori_n669_));
  NO2        o647(.A(ori_ori_n669_), .B(ori_ori_n662_), .Y(ori_ori_n670_));
  INV        o648(.A(ori_ori_n168_), .Y(ori_ori_n671_));
  INV        o649(.A(ori_ori_n228_), .Y(ori_ori_n672_));
  OAI210     o650(.A0(ori_ori_n613_), .A1(ori_ori_n401_), .B0(ori_ori_n110_), .Y(ori_ori_n673_));
  AOI210     o651(.A0(ori_ori_n673_), .A1(ori_ori_n672_), .B0(ori_ori_n671_), .Y(ori_ori_n674_));
  NO2        o652(.A(ori_ori_n409_), .B(ori_ori_n26_), .Y(ori_ori_n675_));
  NO2        o653(.A(ori_ori_n675_), .B(ori_ori_n376_), .Y(ori_ori_n676_));
  NA2        o654(.A(ori_ori_n676_), .B(i_2_), .Y(ori_ori_n677_));
  INV        o655(.A(ori_ori_n677_), .Y(ori_ori_n678_));
  AOI210     o656(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n373_), .Y(ori_ori_n679_));
  AOI210     o657(.A0(ori_ori_n679_), .A1(ori_ori_n678_), .B0(ori_ori_n674_), .Y(ori_ori_n680_));
  NO2        o658(.A(ori_ori_n184_), .B(ori_ori_n125_), .Y(ori_ori_n681_));
  OAI210     o659(.A0(ori_ori_n681_), .A1(ori_ori_n664_), .B0(i_2_), .Y(ori_ori_n682_));
  INV        o660(.A(ori_ori_n169_), .Y(ori_ori_n683_));
  NO3        o661(.A(ori_ori_n542_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n684_));
  AOI210     o662(.A0(ori_ori_n683_), .A1(ori_ori_n86_), .B0(ori_ori_n684_), .Y(ori_ori_n685_));
  AOI210     o663(.A0(ori_ori_n685_), .A1(ori_ori_n682_), .B0(ori_ori_n186_), .Y(ori_ori_n686_));
  OA210      o664(.A0(ori_ori_n543_), .A1(ori_ori_n126_), .B0(i_13_), .Y(ori_ori_n687_));
  NA2        o665(.A(ori_ori_n191_), .B(ori_ori_n192_), .Y(ori_ori_n688_));
  NA2        o666(.A(ori_ori_n151_), .B(ori_ori_n521_), .Y(ori_ori_n689_));
  AOI210     o667(.A0(ori_ori_n689_), .A1(ori_ori_n688_), .B0(ori_ori_n330_), .Y(ori_ori_n690_));
  AOI210     o668(.A0(ori_ori_n198_), .A1(ori_ori_n148_), .B0(ori_ori_n456_), .Y(ori_ori_n691_));
  NA2        o669(.A(ori_ori_n691_), .B(ori_ori_n376_), .Y(ori_ori_n692_));
  NO2        o670(.A(ori_ori_n102_), .B(ori_ori_n44_), .Y(ori_ori_n693_));
  INV        o671(.A(ori_ori_n276_), .Y(ori_ori_n694_));
  NA4        o672(.A(ori_ori_n694_), .B(ori_ori_n278_), .C(ori_ori_n124_), .D(ori_ori_n42_), .Y(ori_ori_n695_));
  OAI210     o673(.A0(ori_ori_n695_), .A1(ori_ori_n693_), .B0(ori_ori_n692_), .Y(ori_ori_n696_));
  NO4        o674(.A(ori_ori_n696_), .B(ori_ori_n690_), .C(ori_ori_n687_), .D(ori_ori_n686_), .Y(ori_ori_n697_));
  NA2        o675(.A(ori_ori_n497_), .B(ori_ori_n28_), .Y(ori_ori_n698_));
  NA2        o676(.A(ori_ori_n663_), .B(ori_ori_n251_), .Y(ori_ori_n699_));
  NA2        o677(.A(ori_ori_n699_), .B(ori_ori_n698_), .Y(ori_ori_n700_));
  NO2        o678(.A(ori_ori_n61_), .B(i_12_), .Y(ori_ori_n701_));
  NO2        o679(.A(ori_ori_n701_), .B(ori_ori_n126_), .Y(ori_ori_n702_));
  NO2        o680(.A(ori_ori_n702_), .B(ori_ori_n521_), .Y(ori_ori_n703_));
  AOI220     o681(.A0(ori_ori_n703_), .A1(ori_ori_n36_), .B0(ori_ori_n700_), .B1(ori_ori_n46_), .Y(ori_ori_n704_));
  NA4        o682(.A(ori_ori_n704_), .B(ori_ori_n697_), .C(ori_ori_n680_), .D(ori_ori_n670_), .Y(ori6));
  NO3        o683(.A(i_9_), .B(ori_ori_n279_), .C(i_1_), .Y(ori_ori_n706_));
  NA2        o684(.A(ori_ori_n706_), .B(ori_ori_n651_), .Y(ori_ori_n707_));
  NA4        o685(.A(ori_ori_n348_), .B(ori_ori_n429_), .C(ori_ori_n70_), .D(ori_ori_n101_), .Y(ori_ori_n708_));
  INV        o686(.A(ori_ori_n708_), .Y(ori_ori_n709_));
  NO2        o687(.A(ori_ori_n207_), .B(ori_ori_n432_), .Y(ori_ori_n710_));
  NO2        o688(.A(ori_ori_n709_), .B(ori_ori_n296_), .Y(ori_ori_n711_));
  AO210      o689(.A0(ori_ori_n711_), .A1(ori_ori_n707_), .B0(i_12_), .Y(ori_ori_n712_));
  NA2        o690(.A(ori_ori_n505_), .B(ori_ori_n62_), .Y(ori_ori_n713_));
  NA2        o691(.A(ori_ori_n606_), .B(ori_ori_n70_), .Y(ori_ori_n714_));
  BUFFER     o692(.A(ori_ori_n548_), .Y(ori_ori_n715_));
  NA3        o693(.A(ori_ori_n715_), .B(ori_ori_n714_), .C(ori_ori_n713_), .Y(ori_ori_n716_));
  NA2        o694(.A(ori_ori_n716_), .B(ori_ori_n72_), .Y(ori_ori_n717_));
  INV        o695(.A(ori_ori_n295_), .Y(ori_ori_n718_));
  NA2        o696(.A(ori_ori_n74_), .B(ori_ori_n131_), .Y(ori_ori_n719_));
  INV        o697(.A(ori_ori_n124_), .Y(ori_ori_n720_));
  NA2        o698(.A(ori_ori_n720_), .B(ori_ori_n46_), .Y(ori_ori_n721_));
  AOI210     o699(.A0(ori_ori_n721_), .A1(ori_ori_n719_), .B0(ori_ori_n718_), .Y(ori_ori_n722_));
  NO2        o700(.A(ori_ori_n231_), .B(i_9_), .Y(ori_ori_n723_));
  NA2        o701(.A(ori_ori_n723_), .B(ori_ori_n701_), .Y(ori_ori_n724_));
  AOI210     o702(.A0(ori_ori_n724_), .A1(ori_ori_n454_), .B0(ori_ori_n180_), .Y(ori_ori_n725_));
  NO2        o703(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n726_));
  NA3        o704(.A(ori_ori_n726_), .B(ori_ori_n426_), .C(ori_ori_n348_), .Y(ori_ori_n727_));
  NAi32      o705(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n728_));
  NO2        o706(.A(ori_ori_n637_), .B(ori_ori_n728_), .Y(ori_ori_n729_));
  OAI210     o707(.A0(ori_ori_n605_), .A1(ori_ori_n488_), .B0(ori_ori_n487_), .Y(ori_ori_n730_));
  NAi31      o708(.An(ori_ori_n729_), .B(ori_ori_n730_), .C(ori_ori_n727_), .Y(ori_ori_n731_));
  OR3        o709(.A(ori_ori_n731_), .B(ori_ori_n725_), .C(ori_ori_n722_), .Y(ori_ori_n732_));
  NO2        o710(.A(ori_ori_n616_), .B(i_2_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n734_));
  NO2        o712(.A(ori_ori_n734_), .B(ori_ori_n368_), .Y(ori_ori_n735_));
  NA2        o713(.A(ori_ori_n735_), .B(ori_ori_n733_), .Y(ori_ori_n736_));
  OR2        o714(.A(ori_ori_n543_), .B(ori_ori_n401_), .Y(ori_ori_n737_));
  NA3        o715(.A(ori_ori_n737_), .B(ori_ori_n147_), .C(ori_ori_n68_), .Y(ori_ori_n738_));
  AO210      o716(.A0(ori_ori_n439_), .A1(ori_ori_n667_), .B0(ori_ori_n36_), .Y(ori_ori_n739_));
  NA3        o717(.A(ori_ori_n739_), .B(ori_ori_n738_), .C(ori_ori_n736_), .Y(ori_ori_n740_));
  OAI210     o718(.A0(ori_ori_n564_), .A1(i_11_), .B0(ori_ori_n84_), .Y(ori_ori_n741_));
  AOI220     o719(.A0(ori_ori_n741_), .A1(ori_ori_n487_), .B0(ori_ori_n710_), .B1(ori_ori_n633_), .Y(ori_ori_n742_));
  NA3        o720(.A(ori_ori_n330_), .B(ori_ori_n222_), .C(ori_ori_n147_), .Y(ori_ori_n743_));
  NA2        o721(.A(ori_ori_n356_), .B(ori_ori_n69_), .Y(ori_ori_n744_));
  NA4        o722(.A(ori_ori_n744_), .B(ori_ori_n743_), .C(ori_ori_n742_), .D(ori_ori_n528_), .Y(ori_ori_n745_));
  AO210      o723(.A0(ori_ori_n456_), .A1(ori_ori_n46_), .B0(ori_ori_n85_), .Y(ori_ori_n746_));
  NA3        o724(.A(ori_ori_n746_), .B(ori_ori_n430_), .C(ori_ori_n206_), .Y(ori_ori_n747_));
  NA2        o725(.A(ori_ori_n401_), .B(ori_ori_n399_), .Y(ori_ori_n748_));
  NO2        o726(.A(ori_ori_n536_), .B(ori_ori_n102_), .Y(ori_ori_n749_));
  OAI210     o727(.A0(ori_ori_n749_), .A1(ori_ori_n111_), .B0(ori_ori_n367_), .Y(ori_ori_n750_));
  NA2        o728(.A(ori_ori_n227_), .B(ori_ori_n46_), .Y(ori_ori_n751_));
  INV        o729(.A(ori_ori_n510_), .Y(ori_ori_n752_));
  NA3        o730(.A(ori_ori_n752_), .B(ori_ori_n295_), .C(i_7_), .Y(ori_ori_n753_));
  NA4        o731(.A(ori_ori_n753_), .B(ori_ori_n750_), .C(ori_ori_n748_), .D(ori_ori_n747_), .Y(ori_ori_n754_));
  NO4        o732(.A(ori_ori_n754_), .B(ori_ori_n745_), .C(ori_ori_n740_), .D(ori_ori_n732_), .Y(ori_ori_n755_));
  NA4        o733(.A(ori_ori_n755_), .B(ori_ori_n717_), .C(ori_ori_n712_), .D(ori_ori_n338_), .Y(ori3));
  NA3        o734(.A(ori_ori_n743_), .B(ori_ori_n528_), .C(ori_ori_n329_), .Y(ori_ori_n757_));
  NA2        o735(.A(ori_ori_n757_), .B(ori_ori_n40_), .Y(ori_ori_n758_));
  NOi21      o736(.An(ori_ori_n96_), .B(ori_ori_n676_), .Y(ori_ori_n759_));
  NO3        o737(.A(ori_ori_n553_), .B(ori_ori_n409_), .C(ori_ori_n131_), .Y(ori_ori_n760_));
  NA2        o738(.A(ori_ori_n369_), .B(ori_ori_n45_), .Y(ori_ori_n761_));
  AN2        o739(.A(ori_ori_n407_), .B(ori_ori_n55_), .Y(ori_ori_n762_));
  NO3        o740(.A(ori_ori_n762_), .B(ori_ori_n760_), .C(ori_ori_n759_), .Y(ori_ori_n763_));
  AOI210     o741(.A0(ori_ori_n763_), .A1(ori_ori_n758_), .B0(ori_ori_n48_), .Y(ori_ori_n764_));
  NO4        o742(.A(ori_ori_n334_), .B(ori_ori_n341_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n765_));
  NA2        o743(.A(ori_ori_n180_), .B(ori_ori_n493_), .Y(ori_ori_n766_));
  NOi21      o744(.An(ori_ori_n766_), .B(ori_ori_n765_), .Y(ori_ori_n767_));
  NA2        o745(.A(ori_ori_n627_), .B(ori_ori_n595_), .Y(ori_ori_n768_));
  NA2        o746(.A(ori_ori_n302_), .B(ori_ori_n392_), .Y(ori_ori_n769_));
  OAI220     o747(.A0(ori_ori_n769_), .A1(ori_ori_n768_), .B0(ori_ori_n767_), .B1(ori_ori_n62_), .Y(ori_ori_n770_));
  NOi21      o748(.An(i_5_), .B(i_9_), .Y(ori_ori_n771_));
  NA2        o749(.A(ori_ori_n771_), .B(ori_ori_n398_), .Y(ori_ori_n772_));
  BUFFER     o750(.A(ori_ori_n241_), .Y(ori_ori_n773_));
  AOI210     o751(.A0(ori_ori_n773_), .A1(ori_ori_n427_), .B0(ori_ori_n608_), .Y(ori_ori_n774_));
  NO3        o752(.A(ori_ori_n370_), .B(ori_ori_n241_), .C(ori_ori_n72_), .Y(ori_ori_n775_));
  NO2        o753(.A(ori_ori_n171_), .B(ori_ori_n148_), .Y(ori_ori_n776_));
  AOI210     o754(.A0(ori_ori_n776_), .A1(ori_ori_n227_), .B0(ori_ori_n775_), .Y(ori_ori_n777_));
  OAI220     o755(.A0(ori_ori_n777_), .A1(ori_ori_n175_), .B0(ori_ori_n774_), .B1(ori_ori_n772_), .Y(ori_ori_n778_));
  NO3        o756(.A(ori_ori_n778_), .B(ori_ori_n770_), .C(ori_ori_n764_), .Y(ori_ori_n779_));
  NA2        o757(.A(ori_ori_n180_), .B(ori_ori_n24_), .Y(ori_ori_n780_));
  NO2        o758(.A(ori_ori_n593_), .B(ori_ori_n518_), .Y(ori_ori_n781_));
  NO2        o759(.A(ori_ori_n781_), .B(ori_ori_n780_), .Y(ori_ori_n782_));
  NA2        o760(.A(ori_ori_n283_), .B(ori_ori_n129_), .Y(ori_ori_n783_));
  NAi21      o761(.An(ori_ori_n160_), .B(ori_ori_n392_), .Y(ori_ori_n784_));
  OAI220     o762(.A0(ori_ori_n784_), .A1(ori_ori_n751_), .B0(ori_ori_n783_), .B1(ori_ori_n361_), .Y(ori_ori_n785_));
  NO2        o763(.A(ori_ori_n785_), .B(ori_ori_n782_), .Y(ori_ori_n786_));
  NA2        o764(.A(ori_ori_n494_), .B(i_0_), .Y(ori_ori_n787_));
  NO3        o765(.A(ori_ori_n787_), .B(ori_ori_n343_), .C(ori_ori_n86_), .Y(ori_ori_n788_));
  NO4        o766(.A(ori_ori_n509_), .B(ori_ori_n204_), .C(ori_ori_n373_), .D(ori_ori_n368_), .Y(ori_ori_n789_));
  AOI210     o767(.A0(ori_ori_n789_), .A1(i_11_), .B0(ori_ori_n788_), .Y(ori_ori_n790_));
  INV        o768(.A(ori_ori_n426_), .Y(ori_ori_n791_));
  AN2        o769(.A(ori_ori_n96_), .B(ori_ori_n226_), .Y(ori_ori_n792_));
  NA2        o770(.A(ori_ori_n663_), .B(ori_ori_n296_), .Y(ori_ori_n793_));
  AOI210     o771(.A0(ori_ori_n430_), .A1(ori_ori_n86_), .B0(ori_ori_n57_), .Y(ori_ori_n794_));
  OAI220     o772(.A0(ori_ori_n794_), .A1(ori_ori_n793_), .B0(ori_ori_n578_), .B1(ori_ori_n467_), .Y(ori_ori_n795_));
  NO2        o773(.A(ori_ori_n233_), .B(ori_ori_n152_), .Y(ori_ori_n796_));
  NA2        o774(.A(i_0_), .B(i_10_), .Y(ori_ori_n797_));
  INV        o775(.A(ori_ori_n469_), .Y(ori_ori_n798_));
  NO4        o776(.A(ori_ori_n114_), .B(ori_ori_n57_), .C(ori_ori_n588_), .D(i_5_), .Y(ori_ori_n799_));
  AO220      o777(.A0(ori_ori_n799_), .A1(ori_ori_n798_), .B0(ori_ori_n796_), .B1(i_6_), .Y(ori_ori_n800_));
  NA2        o778(.A(ori_ori_n183_), .B(ori_ori_n192_), .Y(ori_ori_n801_));
  NO2        o779(.A(ori_ori_n801_), .B(ori_ori_n793_), .Y(ori_ori_n802_));
  NO4        o780(.A(ori_ori_n802_), .B(ori_ori_n800_), .C(ori_ori_n795_), .D(ori_ori_n792_), .Y(ori_ori_n803_));
  NA3        o781(.A(ori_ori_n803_), .B(ori_ori_n790_), .C(ori_ori_n786_), .Y(ori_ori_n804_));
  NO2        o782(.A(ori_ori_n103_), .B(ori_ori_n37_), .Y(ori_ori_n805_));
  NA2        o783(.A(i_11_), .B(i_9_), .Y(ori_ori_n806_));
  NO3        o784(.A(i_12_), .B(ori_ori_n806_), .C(ori_ori_n527_), .Y(ori_ori_n807_));
  AN2        o785(.A(ori_ori_n807_), .B(ori_ori_n805_), .Y(ori_ori_n808_));
  NO2        o786(.A(ori_ori_n48_), .B(i_7_), .Y(ori_ori_n809_));
  NA2        o787(.A(ori_ori_n353_), .B(ori_ori_n173_), .Y(ori_ori_n810_));
  NA2        o788(.A(ori_ori_n810_), .B(ori_ori_n158_), .Y(ori_ori_n811_));
  NO2        o789(.A(ori_ori_n171_), .B(i_0_), .Y(ori_ori_n812_));
  NO2        o790(.A(ori_ori_n811_), .B(ori_ori_n808_), .Y(ori_ori_n813_));
  NA2        o791(.A(ori_ori_n577_), .B(ori_ori_n121_), .Y(ori_ori_n814_));
  NO2        o792(.A(i_6_), .B(ori_ori_n814_), .Y(ori_ori_n815_));
  AOI210     o793(.A0(ori_ori_n400_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n816_));
  NA2        o794(.A(ori_ori_n168_), .B(ori_ori_n103_), .Y(ori_ori_n817_));
  NOi32      o795(.An(ori_ori_n816_), .Bn(ori_ori_n183_), .C(ori_ori_n817_), .Y(ori_ori_n818_));
  NA2        o796(.A(ori_ori_n529_), .B(ori_ori_n296_), .Y(ori_ori_n819_));
  NO2        o797(.A(ori_ori_n819_), .B(ori_ori_n761_), .Y(ori_ori_n820_));
  NO3        o798(.A(ori_ori_n820_), .B(ori_ori_n818_), .C(ori_ori_n815_), .Y(ori_ori_n821_));
  NOi21      o799(.An(i_7_), .B(i_5_), .Y(ori_ori_n822_));
  NOi31      o800(.An(ori_ori_n822_), .B(i_0_), .C(ori_ori_n643_), .Y(ori_ori_n823_));
  NA3        o801(.A(ori_ori_n823_), .B(ori_ori_n342_), .C(i_6_), .Y(ori_ori_n824_));
  OA210      o802(.A0(ori_ori_n817_), .A1(ori_ori_n454_), .B0(ori_ori_n824_), .Y(ori_ori_n825_));
  INV        o803(.A(ori_ori_n290_), .Y(ori_ori_n826_));
  NA3        o804(.A(ori_ori_n825_), .B(ori_ori_n821_), .C(ori_ori_n813_), .Y(ori_ori_n827_));
  OA210      o805(.A0(ori_ori_n426_), .A1(ori_ori_n210_), .B0(ori_ori_n425_), .Y(ori_ori_n828_));
  NA3        o806(.A(ori_ori_n425_), .B(ori_ori_n369_), .C(ori_ori_n45_), .Y(ori_ori_n829_));
  OAI210     o807(.A0(ori_ori_n784_), .A1(ori_ori_n791_), .B0(ori_ori_n829_), .Y(ori_ori_n830_));
  NO2        o808(.A(i_3_), .B(ori_ori_n182_), .Y(ori_ori_n831_));
  AOI220     o809(.A0(ori_ori_n831_), .A1(ori_ori_n426_), .B0(ori_ori_n830_), .B1(ori_ori_n72_), .Y(ori_ori_n832_));
  NA3        o810(.A(ori_ori_n734_), .B(ori_ori_n340_), .C(ori_ori_n564_), .Y(ori_ori_n833_));
  NA2        o811(.A(ori_ori_n92_), .B(ori_ori_n44_), .Y(ori_ori_n834_));
  NO2        o812(.A(ori_ori_n74_), .B(ori_ori_n665_), .Y(ori_ori_n835_));
  AOI220     o813(.A0(ori_ori_n835_), .A1(ori_ori_n834_), .B0(ori_ori_n170_), .B1(ori_ori_n518_), .Y(ori_ori_n836_));
  AOI210     o814(.A0(ori_ori_n836_), .A1(ori_ori_n833_), .B0(ori_ori_n47_), .Y(ori_ori_n837_));
  NO2        o815(.A(ori_ori_n837_), .B(ori_ori_n458_), .Y(ori_ori_n838_));
  NA2        o816(.A(ori_ori_n838_), .B(ori_ori_n832_), .Y(ori_ori_n839_));
  NO3        o817(.A(ori_ori_n839_), .B(ori_ori_n827_), .C(ori_ori_n804_), .Y(ori_ori_n840_));
  NO2        o818(.A(i_0_), .B(ori_ori_n643_), .Y(ori_ori_n841_));
  NA2        o819(.A(ori_ori_n72_), .B(ori_ori_n44_), .Y(ori_ori_n842_));
  AN2        o820(.A(ori_ori_n841_), .B(ori_ori_n170_), .Y(ori_ori_n843_));
  NO2        o821(.A(ori_ori_n713_), .B(ori_ori_n817_), .Y(ori_ori_n844_));
  AOI210     o822(.A0(ori_ori_n843_), .A1(ori_ori_n309_), .B0(ori_ori_n844_), .Y(ori_ori_n845_));
  NO2        o823(.A(ori_ori_n730_), .B(ori_ori_n362_), .Y(ori_ori_n846_));
  NA2        o824(.A(ori_ori_n227_), .B(ori_ori_n217_), .Y(ori_ori_n847_));
  AOI210     o825(.A0(ori_ori_n847_), .A1(ori_ori_n787_), .B0(ori_ori_n152_), .Y(ori_ori_n848_));
  NO2        o826(.A(ori_ori_n848_), .B(ori_ori_n846_), .Y(ori_ori_n849_));
  NA2        o827(.A(ori_ori_n849_), .B(ori_ori_n845_), .Y(ori_ori_n850_));
  NO3        o828(.A(ori_ori_n797_), .B(ori_ori_n771_), .C(ori_ori_n184_), .Y(ori_ori_n851_));
  AOI220     o829(.A0(ori_ori_n851_), .A1(i_11_), .B0(ori_ori_n490_), .B1(ori_ori_n74_), .Y(ori_ori_n852_));
  NO3        o830(.A(ori_ori_n199_), .B(ori_ori_n341_), .C(i_0_), .Y(ori_ori_n853_));
  OAI210     o831(.A0(ori_ori_n853_), .A1(ori_ori_n75_), .B0(i_13_), .Y(ori_ori_n854_));
  NA2        o832(.A(ori_ori_n854_), .B(ori_ori_n852_), .Y(ori_ori_n855_));
  AOI210     o833(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n171_), .Y(ori_ori_n856_));
  NA2        o834(.A(ori_ori_n856_), .B(ori_ori_n828_), .Y(ori_ori_n857_));
  INV        o835(.A(ori_ori_n475_), .Y(ori_ori_n858_));
  NO3        o836(.A(ori_ori_n761_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n859_));
  NA2        o837(.A(ori_ori_n438_), .B(ori_ori_n431_), .Y(ori_ori_n860_));
  NO3        o838(.A(ori_ori_n860_), .B(ori_ori_n859_), .C(ori_ori_n858_), .Y(ori_ori_n861_));
  NA3        o839(.A(ori_ori_n348_), .B(ori_ori_n168_), .C(ori_ori_n167_), .Y(ori_ori_n862_));
  NA3        o840(.A(ori_ori_n809_), .B(ori_ori_n266_), .C(ori_ori_n217_), .Y(ori_ori_n863_));
  NA2        o841(.A(ori_ori_n863_), .B(ori_ori_n862_), .Y(ori_ori_n864_));
  NA3        o842(.A(ori_ori_n348_), .B(ori_ori_n303_), .C(ori_ori_n208_), .Y(ori_ori_n865_));
  INV        o843(.A(ori_ori_n865_), .Y(ori_ori_n866_));
  NOi31      o844(.An(ori_ori_n347_), .B(ori_ori_n842_), .C(ori_ori_n223_), .Y(ori_ori_n867_));
  NO3        o845(.A(ori_ori_n806_), .B(ori_ori_n206_), .C(ori_ori_n184_), .Y(ori_ori_n868_));
  NO4        o846(.A(ori_ori_n868_), .B(ori_ori_n867_), .C(ori_ori_n866_), .D(ori_ori_n864_), .Y(ori_ori_n869_));
  NA3        o847(.A(ori_ori_n869_), .B(ori_ori_n861_), .C(ori_ori_n857_), .Y(ori_ori_n870_));
  NA3        o848(.A(ori_ori_n278_), .B(i_5_), .C(ori_ori_n186_), .Y(ori_ori_n871_));
  NAi31      o849(.An(ori_ori_n224_), .B(ori_ori_n871_), .C(ori_ori_n225_), .Y(ori_ori_n872_));
  NO4        o850(.A(ori_ori_n223_), .B(ori_ori_n199_), .C(i_0_), .D(i_12_), .Y(ori_ori_n873_));
  AOI220     o851(.A0(ori_ori_n873_), .A1(ori_ori_n872_), .B0(ori_ori_n709_), .B1(ori_ori_n172_), .Y(ori_ori_n874_));
  AN2        o852(.A(ori_ori_n797_), .B(ori_ori_n152_), .Y(ori_ori_n875_));
  NO4        o853(.A(ori_ori_n875_), .B(i_12_), .C(ori_ori_n568_), .D(ori_ori_n131_), .Y(ori_ori_n876_));
  NA2        o854(.A(ori_ori_n876_), .B(ori_ori_n206_), .Y(ori_ori_n877_));
  NA3        o855(.A(ori_ori_n98_), .B(ori_ori_n493_), .C(i_11_), .Y(ori_ori_n878_));
  NO2        o856(.A(ori_ori_n878_), .B(ori_ori_n154_), .Y(ori_ori_n879_));
  NA2        o857(.A(ori_ori_n822_), .B(ori_ori_n423_), .Y(ori_ori_n880_));
  NA2        o858(.A(ori_ori_n63_), .B(ori_ori_n101_), .Y(ori_ori_n881_));
  OAI220     o859(.A0(ori_ori_n881_), .A1(ori_ori_n871_), .B0(ori_ori_n880_), .B1(ori_ori_n596_), .Y(ori_ori_n882_));
  AOI210     o860(.A0(ori_ori_n882_), .A1(ori_ori_n812_), .B0(ori_ori_n879_), .Y(ori_ori_n883_));
  NA3        o861(.A(ori_ori_n883_), .B(ori_ori_n877_), .C(ori_ori_n874_), .Y(ori_ori_n884_));
  NO4        o862(.A(ori_ori_n884_), .B(ori_ori_n870_), .C(ori_ori_n855_), .D(ori_ori_n850_), .Y(ori_ori_n885_));
  OAI210     o863(.A0(ori_ori_n733_), .A1(ori_ori_n726_), .B0(ori_ori_n37_), .Y(ori_ori_n886_));
  NA3        o864(.A(ori_ori_n816_), .B(ori_ori_n325_), .C(i_5_), .Y(ori_ori_n887_));
  NA3        o865(.A(ori_ori_n887_), .B(ori_ori_n886_), .C(ori_ori_n535_), .Y(ori_ori_n888_));
  NA2        o866(.A(ori_ori_n888_), .B(ori_ori_n197_), .Y(ori_ori_n889_));
  AN2        o867(.A(ori_ori_n616_), .B(ori_ori_n326_), .Y(ori_ori_n890_));
  NA2        o868(.A(ori_ori_n181_), .B(ori_ori_n183_), .Y(ori_ori_n891_));
  AO210      o869(.A0(ori_ori_n890_), .A1(ori_ori_n33_), .B0(ori_ori_n891_), .Y(ori_ori_n892_));
  NAi31      o870(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n893_));
  AOI210     o871(.A0(ori_ori_n117_), .A1(ori_ori_n69_), .B0(ori_ori_n893_), .Y(ori_ori_n894_));
  NO2        o872(.A(ori_ori_n894_), .B(ori_ori_n567_), .Y(ori_ori_n895_));
  NA2        o873(.A(ori_ori_n895_), .B(ori_ori_n892_), .Y(ori_ori_n896_));
  NO2        o874(.A(ori_ori_n417_), .B(ori_ori_n241_), .Y(ori_ori_n897_));
  NO2        o875(.A(ori_ori_n897_), .B(ori_ori_n789_), .Y(ori_ori_n898_));
  OAI210     o876(.A0(ori_ori_n878_), .A1(ori_ori_n148_), .B0(ori_ori_n898_), .Y(ori_ori_n899_));
  AOI210     o877(.A0(ori_ori_n896_), .A1(ori_ori_n48_), .B0(ori_ori_n899_), .Y(ori_ori_n900_));
  AOI210     o878(.A0(ori_ori_n900_), .A1(ori_ori_n889_), .B0(ori_ori_n72_), .Y(ori_ori_n901_));
  INV        o879(.A(ori_ori_n337_), .Y(ori_ori_n902_));
  NO2        o880(.A(ori_ori_n902_), .B(ori_ori_n671_), .Y(ori_ori_n903_));
  OAI210     o881(.A0(ori_ori_n79_), .A1(ori_ori_n54_), .B0(ori_ori_n108_), .Y(ori_ori_n904_));
  NA2        o882(.A(ori_ori_n904_), .B(ori_ori_n75_), .Y(ori_ori_n905_));
  AOI210     o883(.A0(ori_ori_n856_), .A1(ori_ori_n809_), .B0(ori_ori_n823_), .Y(ori_ori_n906_));
  AOI210     o884(.A0(ori_ori_n906_), .A1(ori_ori_n905_), .B0(ori_ori_n599_), .Y(ori_ori_n907_));
  INV        o885(.A(ori_ori_n907_), .Y(ori_ori_n908_));
  OAI210     o886(.A0(ori_ori_n243_), .A1(ori_ori_n156_), .B0(ori_ori_n86_), .Y(ori_ori_n909_));
  NO2        o887(.A(ori_ori_n909_), .B(i_11_), .Y(ori_ori_n910_));
  NA2        o888(.A(ori_ori_n530_), .B(ori_ori_n204_), .Y(ori_ori_n911_));
  OAI210     o889(.A0(ori_ori_n911_), .A1(ori_ori_n816_), .B0(ori_ori_n197_), .Y(ori_ori_n912_));
  NA2        o890(.A(ori_ori_n162_), .B(i_5_), .Y(ori_ori_n913_));
  NO2        o891(.A(ori_ori_n912_), .B(ori_ori_n913_), .Y(ori_ori_n914_));
  NO3        o892(.A(ori_ori_n58_), .B(ori_ori_n57_), .C(i_4_), .Y(ori_ori_n915_));
  OAI210     o893(.A0(ori_ori_n826_), .A1(ori_ori_n279_), .B0(ori_ori_n915_), .Y(ori_ori_n916_));
  NO2        o894(.A(ori_ori_n916_), .B(ori_ori_n643_), .Y(ori_ori_n917_));
  NO3        o895(.A(ori_ori_n917_), .B(ori_ori_n914_), .C(ori_ori_n910_), .Y(ori_ori_n918_));
  OAI210     o896(.A0(ori_ori_n908_), .A1(i_4_), .B0(ori_ori_n918_), .Y(ori_ori_n919_));
  NO3        o897(.A(ori_ori_n919_), .B(ori_ori_n903_), .C(ori_ori_n901_), .Y(ori_ori_n920_));
  NA4        o898(.A(ori_ori_n920_), .B(ori_ori_n885_), .C(ori_ori_n840_), .D(ori_ori_n779_), .Y(ori4));
  INV        o899(.A(ori_ori_n620_), .Y(ori_ori_n924_));
  INV        o900(.A(ori_ori_n631_), .Y(ori_ori_n925_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m021(.A(mai_mai_n35_), .Y(mai1));
  INV        m022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m064(.A(i_6_), .Y(mai_mai_n87_));
  OR4        m065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n88_));
  INV        m066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_2_), .B(i_7_), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  OAI210     m069(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NAi21      m070(.An(i_6_), .B(i_10_), .Y(mai_mai_n93_));
  NA2        m071(.A(i_6_), .B(i_9_), .Y(mai_mai_n94_));
  AOI210     m072(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n64_), .Y(mai_mai_n95_));
  NA2        m073(.A(i_2_), .B(i_6_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n97_), .B(mai_mai_n95_), .Y(mai_mai_n98_));
  AOI210     m076(.A0(mai_mai_n98_), .A1(mai_mai_n92_), .B0(mai_mai_n81_), .Y(mai_mai_n99_));
  AN3        m077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n100_));
  NAi21      m078(.An(i_6_), .B(i_11_), .Y(mai_mai_n101_));
  NO2        m079(.A(i_5_), .B(i_8_), .Y(mai_mai_n102_));
  NOi21      m080(.An(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  AOI220     m081(.A0(mai_mai_n103_), .A1(mai_mai_n63_), .B0(mai_mai_n100_), .B1(mai_mai_n32_), .Y(mai_mai_n104_));
  INV        m082(.A(i_7_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n47_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  NO2        m084(.A(i_0_), .B(i_5_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(mai_mai_n87_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_12_), .B(i_3_), .Y(mai_mai_n109_));
  INV        m087(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NA3        m088(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n106_), .Y(mai_mai_n111_));
  NAi21      m089(.An(i_7_), .B(i_11_), .Y(mai_mai_n112_));
  NO3        m090(.A(mai_mai_n112_), .B(mai_mai_n93_), .C(mai_mai_n54_), .Y(mai_mai_n113_));
  AN2        m091(.A(i_2_), .B(i_10_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n114_), .B(i_7_), .Y(mai_mai_n115_));
  OR2        m093(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n116_));
  NO2        m094(.A(i_8_), .B(mai_mai_n105_), .Y(mai_mai_n117_));
  NO3        m095(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(mai_mai_n115_), .Y(mai_mai_n118_));
  NA2        m096(.A(i_12_), .B(i_7_), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n120_), .B(i_0_), .Y(mai_mai_n121_));
  NA2        m099(.A(i_11_), .B(i_12_), .Y(mai_mai_n122_));
  OAI210     m100(.A0(mai_mai_n121_), .A1(mai_mai_n119_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n123_), .B(mai_mai_n118_), .Y(mai_mai_n124_));
  NAi41      m102(.An(mai_mai_n113_), .B(mai_mai_n124_), .C(mai_mai_n111_), .D(mai_mai_n104_), .Y(mai_mai_n125_));
  NOi21      m103(.An(i_1_), .B(i_5_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n126_), .B(i_11_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n105_), .B(mai_mai_n37_), .Y(mai_mai_n128_));
  NA2        m106(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n129_), .B(mai_mai_n128_), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n130_), .B(mai_mai_n47_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n132_));
  NAi21      m110(.An(i_3_), .B(i_8_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n63_), .Y(mai_mai_n134_));
  NOi31      m112(.An(mai_mai_n134_), .B(mai_mai_n132_), .C(mai_mai_n131_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n136_));
  NO2        m114(.A(i_6_), .B(i_5_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n137_), .B(i_3_), .Y(mai_mai_n138_));
  AO210      m116(.A0(mai_mai_n138_), .A1(mai_mai_n48_), .B0(mai_mai_n136_), .Y(mai_mai_n139_));
  OAI220     m117(.A0(mai_mai_n139_), .A1(mai_mai_n112_), .B0(mai_mai_n135_), .B1(mai_mai_n127_), .Y(mai_mai_n140_));
  NO3        m118(.A(mai_mai_n140_), .B(mai_mai_n125_), .C(mai_mai_n99_), .Y(mai_mai_n141_));
  NA3        m119(.A(mai_mai_n141_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m120(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n143_));
  NA2        m121(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  NA4        m123(.A(mai_mai_n145_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m124(.A(i_8_), .B(i_7_), .Y(mai_mai_n147_));
  NA2        m125(.A(mai_mai_n147_), .B(i_6_), .Y(mai_mai_n148_));
  NO2        m126(.A(i_12_), .B(i_13_), .Y(mai_mai_n149_));
  NAi21      m127(.An(i_5_), .B(i_11_), .Y(mai_mai_n150_));
  NOi21      m128(.An(mai_mai_n149_), .B(mai_mai_n150_), .Y(mai_mai_n151_));
  NO2        m129(.A(i_0_), .B(i_1_), .Y(mai_mai_n152_));
  NA2        m130(.A(i_2_), .B(i_3_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n153_), .B(i_4_), .Y(mai_mai_n154_));
  NA3        m132(.A(mai_mai_n154_), .B(mai_mai_n152_), .C(mai_mai_n151_), .Y(mai_mai_n155_));
  OR2        m133(.A(mai_mai_n155_), .B(mai_mai_n25_), .Y(mai_mai_n156_));
  AN2        m134(.A(mai_mai_n149_), .B(mai_mai_n84_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n157_), .B(mai_mai_n27_), .Y(mai_mai_n158_));
  NA2        m136(.A(i_1_), .B(i_5_), .Y(mai_mai_n159_));
  NO2        m137(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n160_), .B(mai_mai_n36_), .Y(mai_mai_n161_));
  NO3        m139(.A(mai_mai_n161_), .B(mai_mai_n159_), .C(mai_mai_n158_), .Y(mai_mai_n162_));
  OR2        m140(.A(i_0_), .B(i_1_), .Y(mai_mai_n163_));
  NAi32      m141(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_4_), .B(i_10_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n40_), .Y(mai_mai_n166_));
  NO2        m144(.A(i_3_), .B(i_5_), .Y(mai_mai_n167_));
  INV        m145(.A(mai_mai_n162_), .Y(mai_mai_n168_));
  AOI210     m146(.A0(mai_mai_n168_), .A1(mai_mai_n156_), .B0(mai_mai_n148_), .Y(mai_mai_n169_));
  NA3        m147(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n170_));
  NA2        m148(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n171_));
  NOi21      m149(.An(i_4_), .B(i_9_), .Y(mai_mai_n172_));
  NOi21      m150(.An(i_11_), .B(i_13_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  OR2        m152(.A(mai_mai_n174_), .B(mai_mai_n171_), .Y(mai_mai_n175_));
  NO2        m153(.A(i_4_), .B(i_5_), .Y(mai_mai_n176_));
  NAi21      m154(.An(i_12_), .B(i_11_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n177_), .B(i_13_), .Y(mai_mai_n178_));
  NA3        m156(.A(mai_mai_n178_), .B(mai_mai_n176_), .C(mai_mai_n84_), .Y(mai_mai_n179_));
  AOI210     m157(.A0(mai_mai_n179_), .A1(mai_mai_n175_), .B0(mai_mai_n170_), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n181_));
  NA2        m159(.A(mai_mai_n181_), .B(mai_mai_n47_), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n183_));
  NA2        m161(.A(i_3_), .B(i_5_), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n185_));
  NO2        m163(.A(i_13_), .B(i_10_), .Y(mai_mai_n186_));
  NA3        m164(.A(mai_mai_n186_), .B(mai_mai_n185_), .C(mai_mai_n45_), .Y(mai_mai_n187_));
  NO2        m165(.A(i_2_), .B(i_1_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(i_3_), .Y(mai_mai_n189_));
  NAi21      m167(.An(i_4_), .B(i_12_), .Y(mai_mai_n190_));
  NO4        m168(.A(mai_mai_n190_), .B(mai_mai_n189_), .C(mai_mai_n187_), .D(mai_mai_n25_), .Y(mai_mai_n191_));
  NO2        m169(.A(mai_mai_n191_), .B(mai_mai_n180_), .Y(mai_mai_n192_));
  INV        m170(.A(i_8_), .Y(mai_mai_n193_));
  NO3        m171(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(mai_mai_n117_), .Y(mai_mai_n195_));
  NO3        m173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n196_));
  NA3        m174(.A(mai_mai_n196_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n197_));
  NO3        m175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n198_));
  OAI210     m176(.A0(mai_mai_n100_), .A1(i_12_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  AOI210     m177(.A0(mai_mai_n199_), .A1(mai_mai_n197_), .B0(mai_mai_n195_), .Y(mai_mai_n200_));
  NO2        m178(.A(i_3_), .B(i_8_), .Y(mai_mai_n201_));
  NO3        m179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n107_), .B(mai_mai_n59_), .Y(mai_mai_n203_));
  NO2        m181(.A(i_13_), .B(i_9_), .Y(mai_mai_n204_));
  NA3        m182(.A(mai_mai_n204_), .B(i_6_), .C(mai_mai_n193_), .Y(mai_mai_n205_));
  NAi21      m183(.An(i_12_), .B(i_3_), .Y(mai_mai_n206_));
  OR2        m184(.A(mai_mai_n206_), .B(mai_mai_n205_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n208_));
  NO3        m186(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n209_));
  NA2        m187(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n210_), .B(mai_mai_n207_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n211_), .B(mai_mai_n200_), .Y(mai_mai_n212_));
  OAI220     m190(.A0(mai_mai_n212_), .A1(i_4_), .B0(i_7_), .B1(mai_mai_n192_), .Y(mai_mai_n213_));
  NAi21      m191(.An(i_12_), .B(i_7_), .Y(mai_mai_n214_));
  NA3        m192(.A(i_13_), .B(mai_mai_n193_), .C(i_10_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n216_));
  NA2        m194(.A(i_0_), .B(i_5_), .Y(mai_mai_n217_));
  OAI220     m195(.A0(mai_mai_n87_), .A1(mai_mai_n189_), .B0(mai_mai_n182_), .B1(mai_mai_n138_), .Y(mai_mai_n218_));
  NAi31      m196(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n220_));
  NO2        m198(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n222_));
  INV        m200(.A(i_13_), .Y(mai_mai_n223_));
  NO2        m201(.A(i_12_), .B(mai_mai_n223_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n218_), .B(mai_mai_n216_), .Y(mai_mai_n225_));
  NO2        m203(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n184_), .B(i_4_), .Y(mai_mai_n227_));
  NA2        m205(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  OR2        m206(.A(i_8_), .B(i_7_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n229_), .B(mai_mai_n87_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n231_));
  NA2        m209(.A(mai_mai_n231_), .B(mai_mai_n230_), .Y(mai_mai_n232_));
  INV        m210(.A(i_12_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n45_), .B(mai_mai_n233_), .Y(mai_mai_n234_));
  NO3        m212(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n235_));
  NA2        m213(.A(i_2_), .B(i_1_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n232_), .B(mai_mai_n228_), .Y(mai_mai_n237_));
  NO3        m215(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n238_));
  NAi21      m216(.An(i_4_), .B(i_3_), .Y(mai_mai_n239_));
  NO2        m217(.A(i_0_), .B(i_6_), .Y(mai_mai_n240_));
  NOi41      m218(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n241_), .B(mai_mai_n240_), .Y(mai_mai_n242_));
  NO2        m220(.A(mai_mai_n236_), .B(mai_mai_n184_), .Y(mai_mai_n243_));
  NAi21      m221(.An(mai_mai_n242_), .B(mai_mai_n243_), .Y(mai_mai_n244_));
  INV        m222(.A(mai_mai_n244_), .Y(mai_mai_n245_));
  AOI220     m223(.A0(mai_mai_n245_), .A1(mai_mai_n40_), .B0(mai_mai_n237_), .B1(mai_mai_n204_), .Y(mai_mai_n246_));
  NO2        m224(.A(i_11_), .B(mai_mai_n223_), .Y(mai_mai_n247_));
  NOi21      m225(.An(i_1_), .B(i_6_), .Y(mai_mai_n248_));
  NAi21      m226(.An(i_3_), .B(i_7_), .Y(mai_mai_n249_));
  NA2        m227(.A(mai_mai_n233_), .B(i_9_), .Y(mai_mai_n250_));
  OR4        m228(.A(mai_mai_n250_), .B(mai_mai_n249_), .C(mai_mai_n248_), .D(mai_mai_n185_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n252_));
  NO2        m230(.A(i_12_), .B(i_3_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n254_));
  NA2        m232(.A(i_3_), .B(i_9_), .Y(mai_mai_n255_));
  NAi21      m233(.An(i_7_), .B(i_10_), .Y(mai_mai_n256_));
  NO2        m234(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n257_));
  NA3        m235(.A(mai_mai_n257_), .B(mai_mai_n254_), .C(mai_mai_n65_), .Y(mai_mai_n258_));
  NA2        m236(.A(mai_mai_n258_), .B(mai_mai_n251_), .Y(mai_mai_n259_));
  NA3        m237(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n260_));
  INV        m238(.A(mai_mai_n148_), .Y(mai_mai_n261_));
  NA2        m239(.A(mai_mai_n233_), .B(i_13_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n262_), .B(mai_mai_n76_), .Y(mai_mai_n263_));
  AOI220     m241(.A0(mai_mai_n263_), .A1(mai_mai_n261_), .B0(mai_mai_n259_), .B1(mai_mai_n247_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n229_), .B(mai_mai_n37_), .Y(mai_mai_n265_));
  NA2        m243(.A(i_12_), .B(i_6_), .Y(mai_mai_n266_));
  OR2        m244(.A(i_13_), .B(i_9_), .Y(mai_mai_n267_));
  NO3        m245(.A(mai_mai_n267_), .B(mai_mai_n266_), .C(mai_mai_n49_), .Y(mai_mai_n268_));
  NO2        m246(.A(mai_mai_n239_), .B(i_2_), .Y(mai_mai_n269_));
  NA3        m247(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n45_), .Y(mai_mai_n270_));
  NA2        m248(.A(mai_mai_n247_), .B(i_9_), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n254_), .B(mai_mai_n65_), .Y(mai_mai_n272_));
  OAI210     m250(.A0(mai_mai_n272_), .A1(mai_mai_n271_), .B0(mai_mai_n270_), .Y(mai_mai_n273_));
  NO3        m251(.A(i_11_), .B(mai_mai_n223_), .C(mai_mai_n25_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n249_), .B(i_8_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n273_), .B(mai_mai_n265_), .Y(mai_mai_n276_));
  NA4        m254(.A(mai_mai_n276_), .B(mai_mai_n264_), .C(mai_mai_n246_), .D(mai_mai_n225_), .Y(mai_mai_n277_));
  NO3        m255(.A(i_12_), .B(mai_mai_n223_), .C(mai_mai_n37_), .Y(mai_mai_n278_));
  INV        m256(.A(mai_mai_n278_), .Y(mai_mai_n279_));
  NO3        m257(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n236_), .B(i_0_), .Y(mai_mai_n281_));
  NA2        m259(.A(i_0_), .B(i_1_), .Y(mai_mai_n282_));
  NO2        m260(.A(mai_mai_n282_), .B(i_2_), .Y(mai_mai_n283_));
  NO2        m261(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n284_));
  NA3        m262(.A(mai_mai_n284_), .B(mai_mai_n283_), .C(mai_mai_n167_), .Y(mai_mai_n285_));
  NO2        m263(.A(i_3_), .B(i_10_), .Y(mai_mai_n286_));
  NA3        m264(.A(mai_mai_n286_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n287_));
  NO2        m265(.A(i_2_), .B(mai_mai_n105_), .Y(mai_mai_n288_));
  NA2        m266(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n289_), .B(i_8_), .Y(mai_mai_n290_));
  NA2        m268(.A(mai_mai_n290_), .B(mai_mai_n288_), .Y(mai_mai_n291_));
  AN2        m269(.A(i_3_), .B(i_10_), .Y(mai_mai_n292_));
  NA4        m270(.A(mai_mai_n292_), .B(mai_mai_n196_), .C(mai_mai_n178_), .D(mai_mai_n176_), .Y(mai_mai_n293_));
  NO2        m271(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n295_));
  OR2        m273(.A(mai_mai_n291_), .B(mai_mai_n287_), .Y(mai_mai_n296_));
  OAI220     m274(.A0(mai_mai_n296_), .A1(i_6_), .B0(mai_mai_n285_), .B1(mai_mai_n279_), .Y(mai_mai_n297_));
  NO4        m275(.A(mai_mai_n297_), .B(mai_mai_n277_), .C(mai_mai_n213_), .D(mai_mai_n169_), .Y(mai_mai_n298_));
  NO3        m276(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n300_));
  NO3        m278(.A(i_6_), .B(mai_mai_n193_), .C(i_7_), .Y(mai_mai_n301_));
  NO2        m279(.A(i_2_), .B(i_3_), .Y(mai_mai_n302_));
  OR2        m280(.A(i_0_), .B(i_5_), .Y(mai_mai_n303_));
  NA2        m281(.A(mai_mai_n217_), .B(mai_mai_n303_), .Y(mai_mai_n304_));
  NA4        m282(.A(mai_mai_n304_), .B(mai_mai_n230_), .C(mai_mai_n302_), .D(i_1_), .Y(mai_mai_n305_));
  NAi21      m283(.An(i_8_), .B(i_7_), .Y(mai_mai_n306_));
  NO2        m284(.A(mai_mai_n306_), .B(i_6_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n163_), .B(mai_mai_n47_), .Y(mai_mai_n308_));
  NA3        m286(.A(mai_mai_n308_), .B(mai_mai_n307_), .C(mai_mai_n167_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n309_), .B(mai_mai_n305_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n310_), .B(i_4_), .Y(mai_mai_n311_));
  NO2        m289(.A(i_12_), .B(i_10_), .Y(mai_mai_n312_));
  NOi21      m290(.An(i_5_), .B(i_0_), .Y(mai_mai_n313_));
  NA4        m291(.A(mai_mai_n85_), .B(mai_mai_n36_), .C(mai_mai_n87_), .D(i_8_), .Y(mai_mai_n314_));
  NO2        m292(.A(i_6_), .B(i_8_), .Y(mai_mai_n315_));
  NOi21      m293(.An(i_0_), .B(i_2_), .Y(mai_mai_n316_));
  BUFFER     m294(.A(mai_mai_n316_), .Y(mai_mai_n317_));
  NO2        m295(.A(i_1_), .B(i_7_), .Y(mai_mai_n318_));
  AO220      m296(.A0(mai_mai_n318_), .A1(mai_mai_n317_), .B0(mai_mai_n307_), .B1(mai_mai_n231_), .Y(mai_mai_n319_));
  NA3        m297(.A(mai_mai_n319_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n320_));
  NA2        m298(.A(mai_mai_n320_), .B(mai_mai_n311_), .Y(mai_mai_n321_));
  NO3        m299(.A(mai_mai_n229_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n322_));
  NO3        m300(.A(mai_mai_n306_), .B(i_2_), .C(i_1_), .Y(mai_mai_n323_));
  OAI210     m301(.A0(mai_mai_n323_), .A1(mai_mai_n322_), .B0(i_6_), .Y(mai_mai_n324_));
  NA3        m302(.A(mai_mai_n248_), .B(mai_mai_n288_), .C(mai_mai_n193_), .Y(mai_mai_n325_));
  AOI210     m303(.A0(mai_mai_n325_), .A1(mai_mai_n324_), .B0(mai_mai_n304_), .Y(mai_mai_n326_));
  NA2        m304(.A(mai_mai_n326_), .B(i_3_), .Y(mai_mai_n327_));
  INV        m305(.A(mai_mai_n85_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n282_), .B(mai_mai_n82_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(mai_mai_n137_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n96_), .B(mai_mai_n193_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n331_), .B(mai_mai_n64_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n332_), .A1(mai_mai_n330_), .B0(mai_mai_n328_), .Y(mai_mai_n333_));
  NO2        m311(.A(mai_mai_n193_), .B(i_9_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n334_), .B(mai_mai_n203_), .Y(mai_mai_n335_));
  INV        m313(.A(mai_mai_n333_), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n327_), .B0(mai_mai_n166_), .Y(mai_mai_n337_));
  AOI210     m315(.A0(mai_mai_n321_), .A1(mai_mai_n299_), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  NOi32      m316(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n339_));
  INV        m317(.A(mai_mai_n339_), .Y(mai_mai_n340_));
  NAi21      m318(.An(i_0_), .B(i_6_), .Y(mai_mai_n341_));
  NAi21      m319(.An(i_1_), .B(i_5_), .Y(mai_mai_n342_));
  NA2        m320(.A(mai_mai_n342_), .B(mai_mai_n341_), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n343_), .B(mai_mai_n25_), .Y(mai_mai_n344_));
  OAI210     m322(.A0(mai_mai_n344_), .A1(mai_mai_n164_), .B0(mai_mai_n242_), .Y(mai_mai_n345_));
  NAi41      m323(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n346_));
  OAI220     m324(.A0(mai_mai_n346_), .A1(mai_mai_n342_), .B0(mai_mai_n219_), .B1(mai_mai_n164_), .Y(mai_mai_n347_));
  AOI210     m325(.A0(mai_mai_n346_), .A1(mai_mai_n164_), .B0(mai_mai_n163_), .Y(mai_mai_n348_));
  OR2        m326(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  NO2        m327(.A(i_1_), .B(mai_mai_n105_), .Y(mai_mai_n350_));
  NAi21      m328(.An(i_3_), .B(i_4_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n351_), .B(i_9_), .Y(mai_mai_n352_));
  AN2        m330(.A(i_6_), .B(i_7_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n350_), .B0(mai_mai_n352_), .Y(mai_mai_n354_));
  NA2        m332(.A(i_2_), .B(i_7_), .Y(mai_mai_n355_));
  NO2        m333(.A(mai_mai_n351_), .B(i_10_), .Y(mai_mai_n356_));
  NO2        m334(.A(mai_mai_n354_), .B(mai_mai_n185_), .Y(mai_mai_n357_));
  AOI210     m335(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n358_));
  OAI210     m336(.A0(mai_mai_n358_), .A1(mai_mai_n188_), .B0(mai_mai_n356_), .Y(mai_mai_n359_));
  AOI220     m337(.A0(mai_mai_n356_), .A1(mai_mai_n318_), .B0(mai_mai_n235_), .B1(mai_mai_n188_), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n360_), .A1(mai_mai_n359_), .B0(i_5_), .Y(mai_mai_n361_));
  NO4        m339(.A(mai_mai_n361_), .B(mai_mai_n357_), .C(mai_mai_n349_), .D(mai_mai_n345_), .Y(mai_mai_n362_));
  NO2        m340(.A(mai_mai_n362_), .B(mai_mai_n340_), .Y(mai_mai_n363_));
  AN2        m341(.A(i_12_), .B(i_5_), .Y(mai_mai_n364_));
  NO2        m342(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n365_), .B(mai_mai_n364_), .Y(mai_mai_n366_));
  NO2        m344(.A(i_11_), .B(i_6_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n239_), .B(i_5_), .Y(mai_mai_n368_));
  NO2        m346(.A(i_5_), .B(i_10_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n370_));
  NO3        m348(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n371_));
  NO2        m349(.A(i_3_), .B(mai_mai_n105_), .Y(mai_mai_n372_));
  NO2        m350(.A(i_11_), .B(i_12_), .Y(mai_mai_n373_));
  NA3        m351(.A(mai_mai_n117_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n374_));
  NO2        m352(.A(mai_mai_n374_), .B(mai_mai_n219_), .Y(mai_mai_n375_));
  NAi21      m353(.An(i_13_), .B(i_0_), .Y(mai_mai_n376_));
  NO2        m354(.A(mai_mai_n376_), .B(mai_mai_n236_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n375_), .B(mai_mai_n377_), .Y(mai_mai_n378_));
  INV        m356(.A(mai_mai_n378_), .Y(mai_mai_n379_));
  NA2        m357(.A(mai_mai_n45_), .B(mai_mai_n223_), .Y(mai_mai_n380_));
  NO3        m358(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n381_));
  NO2        m359(.A(i_0_), .B(i_11_), .Y(mai_mai_n382_));
  INV        m360(.A(i_5_), .Y(mai_mai_n383_));
  AN2        m361(.A(i_1_), .B(i_6_), .Y(mai_mai_n384_));
  NOi21      m362(.An(i_2_), .B(i_12_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n385_), .B(mai_mai_n384_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n386_), .B(mai_mai_n383_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n147_), .B(i_9_), .Y(mai_mai_n388_));
  NO2        m366(.A(mai_mai_n388_), .B(i_4_), .Y(mai_mai_n389_));
  NA2        m367(.A(mai_mai_n387_), .B(mai_mai_n389_), .Y(mai_mai_n390_));
  NAi21      m368(.An(i_9_), .B(i_4_), .Y(mai_mai_n391_));
  OR2        m369(.A(i_13_), .B(i_10_), .Y(mai_mai_n392_));
  NO3        m370(.A(mai_mai_n392_), .B(mai_mai_n122_), .C(mai_mai_n391_), .Y(mai_mai_n393_));
  OR2        m371(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n394_));
  NO2        m372(.A(mai_mai_n105_), .B(mai_mai_n25_), .Y(mai_mai_n395_));
  NA2        m373(.A(i_5_), .B(mai_mai_n209_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n396_), .B(mai_mai_n394_), .Y(mai_mai_n397_));
  INV        m375(.A(mai_mai_n397_), .Y(mai_mai_n398_));
  AOI210     m376(.A0(mai_mai_n398_), .A1(mai_mai_n390_), .B0(mai_mai_n26_), .Y(mai_mai_n399_));
  INV        m377(.A(mai_mai_n305_), .Y(mai_mai_n400_));
  AOI220     m378(.A0(mai_mai_n284_), .A1(mai_mai_n280_), .B0(mai_mai_n281_), .B1(mai_mai_n300_), .Y(mai_mai_n401_));
  NO2        m379(.A(mai_mai_n401_), .B(mai_mai_n171_), .Y(mai_mai_n402_));
  NO2        m380(.A(mai_mai_n402_), .B(mai_mai_n400_), .Y(mai_mai_n403_));
  NA2        m381(.A(mai_mai_n193_), .B(i_10_), .Y(mai_mai_n404_));
  NA3        m382(.A(mai_mai_n254_), .B(mai_mai_n65_), .C(i_2_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n405_), .B(mai_mai_n404_), .Y(mai_mai_n406_));
  NA2        m384(.A(mai_mai_n301_), .B(mai_mai_n304_), .Y(mai_mai_n407_));
  NO2        m385(.A(mai_mai_n407_), .B(mai_mai_n189_), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n408_), .B(mai_mai_n406_), .Y(mai_mai_n409_));
  AOI210     m387(.A0(mai_mai_n409_), .A1(mai_mai_n403_), .B0(mai_mai_n271_), .Y(mai_mai_n410_));
  NO4        m388(.A(mai_mai_n410_), .B(mai_mai_n399_), .C(mai_mai_n379_), .D(mai_mai_n363_), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n412_));
  NO2        m390(.A(i_10_), .B(i_9_), .Y(mai_mai_n413_));
  NAi21      m391(.An(i_12_), .B(i_8_), .Y(mai_mai_n414_));
  NO2        m392(.A(mai_mai_n414_), .B(i_3_), .Y(mai_mai_n415_));
  NA2        m393(.A(mai_mai_n295_), .B(i_0_), .Y(mai_mai_n416_));
  NO3        m394(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n417_));
  NA2        m395(.A(mai_mai_n266_), .B(mai_mai_n101_), .Y(mai_mai_n418_));
  NA2        m396(.A(mai_mai_n418_), .B(mai_mai_n417_), .Y(mai_mai_n419_));
  NA2        m397(.A(i_8_), .B(i_9_), .Y(mai_mai_n420_));
  AOI210     m398(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n421_));
  OR2        m399(.A(mai_mai_n421_), .B(mai_mai_n420_), .Y(mai_mai_n422_));
  NA2        m400(.A(mai_mai_n278_), .B(mai_mai_n203_), .Y(mai_mai_n423_));
  OAI220     m401(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n419_), .B1(mai_mai_n416_), .Y(mai_mai_n424_));
  NA2        m402(.A(mai_mai_n247_), .B(mai_mai_n294_), .Y(mai_mai_n425_));
  NO3        m403(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n426_));
  INV        m404(.A(mai_mai_n426_), .Y(mai_mai_n427_));
  NA3        m405(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n428_));
  NA4        m406(.A(mai_mai_n150_), .B(mai_mai_n120_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n429_));
  OAI220     m407(.A0(mai_mai_n429_), .A1(mai_mai_n428_), .B0(mai_mai_n427_), .B1(mai_mai_n425_), .Y(mai_mai_n430_));
  NO2        m408(.A(mai_mai_n430_), .B(mai_mai_n424_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n283_), .B(mai_mai_n112_), .Y(mai_mai_n432_));
  OR2        m410(.A(mai_mai_n432_), .B(mai_mai_n205_), .Y(mai_mai_n433_));
  OA210      m411(.A0(mai_mai_n335_), .A1(mai_mai_n105_), .B0(mai_mai_n285_), .Y(mai_mai_n434_));
  OA220      m412(.A0(mai_mai_n434_), .A1(mai_mai_n166_), .B0(mai_mai_n433_), .B1(mai_mai_n228_), .Y(mai_mai_n435_));
  NA2        m413(.A(mai_mai_n100_), .B(i_13_), .Y(mai_mai_n436_));
  NO2        m414(.A(i_2_), .B(i_13_), .Y(mai_mai_n437_));
  NO3        m415(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n438_));
  NO2        m416(.A(i_6_), .B(i_7_), .Y(mai_mai_n439_));
  NA2        m417(.A(mai_mai_n439_), .B(mai_mai_n438_), .Y(mai_mai_n440_));
  NO2        m418(.A(i_11_), .B(i_1_), .Y(mai_mai_n441_));
  OR2        m419(.A(i_11_), .B(i_8_), .Y(mai_mai_n442_));
  NOi21      m420(.An(i_2_), .B(i_7_), .Y(mai_mai_n443_));
  NAi31      m421(.An(mai_mai_n442_), .B(mai_mai_n443_), .C(i_0_), .Y(mai_mai_n444_));
  NO2        m422(.A(mai_mai_n392_), .B(i_6_), .Y(mai_mai_n445_));
  NA3        m423(.A(mai_mai_n445_), .B(i_1_), .C(mai_mai_n76_), .Y(mai_mai_n446_));
  NO2        m424(.A(mai_mai_n446_), .B(mai_mai_n444_), .Y(mai_mai_n447_));
  NO2        m425(.A(i_3_), .B(mai_mai_n193_), .Y(mai_mai_n448_));
  NO2        m426(.A(i_6_), .B(i_10_), .Y(mai_mai_n449_));
  NA4        m427(.A(mai_mai_n449_), .B(mai_mai_n299_), .C(mai_mai_n448_), .D(mai_mai_n233_), .Y(mai_mai_n450_));
  NO2        m428(.A(mai_mai_n450_), .B(mai_mai_n161_), .Y(mai_mai_n451_));
  NA3        m429(.A(mai_mai_n241_), .B(mai_mai_n173_), .C(mai_mai_n137_), .Y(mai_mai_n452_));
  NA2        m430(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n453_));
  NO2        m431(.A(mai_mai_n163_), .B(i_3_), .Y(mai_mai_n454_));
  NAi31      m432(.An(mai_mai_n453_), .B(mai_mai_n454_), .C(mai_mai_n224_), .Y(mai_mai_n455_));
  NA3        m433(.A(mai_mai_n370_), .B(mai_mai_n181_), .C(mai_mai_n154_), .Y(mai_mai_n456_));
  NA3        m434(.A(mai_mai_n456_), .B(mai_mai_n455_), .C(mai_mai_n452_), .Y(mai_mai_n457_));
  NO3        m435(.A(mai_mai_n457_), .B(mai_mai_n451_), .C(mai_mai_n447_), .Y(mai_mai_n458_));
  NA2        m436(.A(mai_mai_n417_), .B(mai_mai_n364_), .Y(mai_mai_n459_));
  NAi21      m437(.An(mai_mai_n215_), .B(mai_mai_n373_), .Y(mai_mai_n460_));
  NA2        m438(.A(mai_mai_n318_), .B(mai_mai_n217_), .Y(mai_mai_n461_));
  NO2        m439(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n462_));
  NO2        m440(.A(i_0_), .B(mai_mai_n87_), .Y(mai_mai_n463_));
  NA3        m441(.A(mai_mai_n463_), .B(mai_mai_n462_), .C(mai_mai_n147_), .Y(mai_mai_n464_));
  OR3        m442(.A(mai_mai_n289_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n465_));
  OAI220     m443(.A0(mai_mai_n465_), .A1(mai_mai_n464_), .B0(mai_mai_n461_), .B1(mai_mai_n460_), .Y(mai_mai_n466_));
  NA2        m444(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n467_));
  NA2        m445(.A(mai_mai_n299_), .B(mai_mai_n235_), .Y(mai_mai_n468_));
  OAI220     m446(.A0(mai_mai_n468_), .A1(mai_mai_n405_), .B0(mai_mai_n467_), .B1(mai_mai_n436_), .Y(mai_mai_n469_));
  NA4        m447(.A(mai_mai_n292_), .B(mai_mai_n222_), .C(mai_mai_n74_), .D(mai_mai_n233_), .Y(mai_mai_n470_));
  NO2        m448(.A(mai_mai_n470_), .B(mai_mai_n440_), .Y(mai_mai_n471_));
  NO3        m449(.A(mai_mai_n471_), .B(mai_mai_n469_), .C(mai_mai_n466_), .Y(mai_mai_n472_));
  NA4        m450(.A(mai_mai_n472_), .B(mai_mai_n458_), .C(mai_mai_n435_), .D(mai_mai_n431_), .Y(mai_mai_n473_));
  NA3        m451(.A(mai_mai_n292_), .B(mai_mai_n178_), .C(mai_mai_n176_), .Y(mai_mai_n474_));
  OAI210     m452(.A0(mai_mai_n287_), .A1(mai_mai_n183_), .B0(mai_mai_n474_), .Y(mai_mai_n475_));
  AN2        m453(.A(mai_mai_n280_), .B(mai_mai_n230_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n476_), .B(mai_mai_n475_), .Y(mai_mai_n477_));
  NA2        m455(.A(mai_mai_n127_), .B(mai_mai_n116_), .Y(mai_mai_n478_));
  AN2        m456(.A(mai_mai_n478_), .B(mai_mai_n417_), .Y(mai_mai_n479_));
  NA2        m457(.A(mai_mai_n299_), .B(i_0_), .Y(mai_mai_n480_));
  OAI210     m458(.A0(mai_mai_n480_), .A1(mai_mai_n228_), .B0(mai_mai_n293_), .Y(mai_mai_n481_));
  AOI220     m459(.A0(mai_mai_n481_), .A1(mai_mai_n307_), .B0(mai_mai_n479_), .B1(mai_mai_n295_), .Y(mai_mai_n482_));
  NA2        m460(.A(mai_mai_n339_), .B(mai_mai_n74_), .Y(mai_mai_n483_));
  NO2        m461(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n484_));
  NAi41      m462(.An(mai_mai_n483_), .B(mai_mai_n449_), .C(mai_mai_n484_), .D(mai_mai_n47_), .Y(mai_mai_n485_));
  AOI210     m463(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n393_), .Y(mai_mai_n486_));
  NA2        m464(.A(mai_mai_n486_), .B(mai_mai_n485_), .Y(mai_mai_n487_));
  INV        m465(.A(mai_mai_n487_), .Y(mai_mai_n488_));
  NO2        m466(.A(i_7_), .B(mai_mai_n197_), .Y(mai_mai_n489_));
  OR2        m467(.A(mai_mai_n184_), .B(i_4_), .Y(mai_mai_n490_));
  NO2        m468(.A(mai_mai_n490_), .B(mai_mai_n87_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n491_), .B(mai_mai_n489_), .Y(mai_mai_n492_));
  NA4        m470(.A(mai_mai_n492_), .B(mai_mai_n488_), .C(mai_mai_n482_), .D(mai_mai_n477_), .Y(mai_mai_n493_));
  NA2        m471(.A(mai_mai_n368_), .B(mai_mai_n283_), .Y(mai_mai_n494_));
  OAI210     m472(.A0(mai_mai_n366_), .A1(mai_mai_n170_), .B0(mai_mai_n494_), .Y(mai_mai_n495_));
  NO2        m473(.A(i_12_), .B(mai_mai_n193_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n496_), .B(mai_mai_n223_), .Y(mai_mai_n497_));
  NO3        m475(.A(mai_mai_n1007_), .B(mai_mai_n497_), .C(mai_mai_n432_), .Y(mai_mai_n498_));
  NOi31      m476(.An(mai_mai_n301_), .B(mai_mai_n392_), .C(mai_mai_n38_), .Y(mai_mai_n499_));
  OAI210     m477(.A0(mai_mai_n499_), .A1(mai_mai_n498_), .B0(mai_mai_n495_), .Y(mai_mai_n500_));
  AOI220     m478(.A0(mai_mai_n308_), .A1(mai_mai_n40_), .B0(mai_mai_n231_), .B1(mai_mai_n204_), .Y(mai_mai_n501_));
  NO2        m479(.A(mai_mai_n501_), .B(mai_mai_n490_), .Y(mai_mai_n502_));
  NA2        m480(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n503_));
  NO2        m481(.A(mai_mai_n503_), .B(i_6_), .Y(mai_mai_n504_));
  NA2        m482(.A(mai_mai_n504_), .B(mai_mai_n502_), .Y(mai_mai_n505_));
  NA2        m483(.A(mai_mai_n243_), .B(mai_mai_n240_), .Y(mai_mai_n506_));
  OAI220     m484(.A0(mai_mai_n506_), .A1(mai_mai_n262_), .B0(mai_mai_n436_), .B1(mai_mai_n138_), .Y(mai_mai_n507_));
  NA2        m485(.A(mai_mai_n507_), .B(mai_mai_n265_), .Y(mai_mai_n508_));
  NOi31      m486(.An(mai_mai_n281_), .B(mai_mai_n287_), .C(mai_mai_n183_), .Y(mai_mai_n509_));
  NA3        m487(.A(mai_mai_n292_), .B(mai_mai_n176_), .C(mai_mai_n100_), .Y(mai_mai_n510_));
  NO2        m488(.A(mai_mai_n220_), .B(mai_mai_n45_), .Y(mai_mai_n511_));
  NO2        m489(.A(mai_mai_n163_), .B(i_5_), .Y(mai_mai_n512_));
  NA3        m490(.A(mai_mai_n512_), .B(mai_mai_n380_), .C(mai_mai_n302_), .Y(mai_mai_n513_));
  OAI210     m491(.A0(mai_mai_n513_), .A1(mai_mai_n511_), .B0(mai_mai_n510_), .Y(mai_mai_n514_));
  OAI210     m492(.A0(mai_mai_n514_), .A1(mai_mai_n509_), .B0(mai_mai_n426_), .Y(mai_mai_n515_));
  NA4        m493(.A(mai_mai_n515_), .B(mai_mai_n508_), .C(mai_mai_n505_), .D(mai_mai_n500_), .Y(mai_mai_n516_));
  NA3        m494(.A(mai_mai_n217_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n517_));
  NA2        m495(.A(mai_mai_n278_), .B(mai_mai_n85_), .Y(mai_mai_n518_));
  AOI210     m496(.A0(mai_mai_n517_), .A1(mai_mai_n330_), .B0(mai_mai_n518_), .Y(mai_mai_n519_));
  NA2        m497(.A(mai_mai_n284_), .B(mai_mai_n280_), .Y(mai_mai_n520_));
  NO2        m498(.A(mai_mai_n520_), .B(mai_mai_n175_), .Y(mai_mai_n521_));
  NA2        m499(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n522_));
  NA2        m500(.A(mai_mai_n413_), .B(mai_mai_n220_), .Y(mai_mai_n523_));
  NO2        m501(.A(mai_mai_n522_), .B(mai_mai_n523_), .Y(mai_mai_n524_));
  AOI210     m502(.A0(i_6_), .A1(mai_mai_n47_), .B0(mai_mai_n350_), .Y(mai_mai_n525_));
  NA2        m503(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n526_));
  NA3        m504(.A(mai_mai_n496_), .B(mai_mai_n274_), .C(mai_mai_n526_), .Y(mai_mai_n527_));
  NO2        m505(.A(mai_mai_n525_), .B(mai_mai_n527_), .Y(mai_mai_n528_));
  NO4        m506(.A(mai_mai_n528_), .B(mai_mai_n524_), .C(mai_mai_n521_), .D(mai_mai_n519_), .Y(mai_mai_n529_));
  NO4        m507(.A(mai_mai_n248_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n530_));
  NO3        m508(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n229_), .B(mai_mai_n36_), .Y(mai_mai_n532_));
  AN2        m510(.A(mai_mai_n532_), .B(mai_mai_n531_), .Y(mai_mai_n533_));
  OA210      m511(.A0(mai_mai_n533_), .A1(mai_mai_n530_), .B0(mai_mai_n339_), .Y(mai_mai_n534_));
  NO2        m512(.A(mai_mai_n392_), .B(i_1_), .Y(mai_mai_n535_));
  NOi31      m513(.An(mai_mai_n535_), .B(mai_mai_n418_), .C(mai_mai_n74_), .Y(mai_mai_n536_));
  AN4        m514(.A(mai_mai_n536_), .B(mai_mai_n389_), .C(mai_mai_n462_), .D(i_2_), .Y(mai_mai_n537_));
  NO2        m515(.A(mai_mai_n401_), .B(mai_mai_n179_), .Y(mai_mai_n538_));
  NO3        m516(.A(mai_mai_n538_), .B(mai_mai_n537_), .C(mai_mai_n534_), .Y(mai_mai_n539_));
  NOi21      m517(.An(i_10_), .B(i_6_), .Y(mai_mai_n540_));
  NO2        m518(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n541_));
  AOI220     m519(.A0(mai_mai_n278_), .A1(mai_mai_n541_), .B0(mai_mai_n274_), .B1(mai_mai_n540_), .Y(mai_mai_n542_));
  NO2        m520(.A(mai_mai_n542_), .B(mai_mai_n416_), .Y(mai_mai_n543_));
  NO2        m521(.A(mai_mai_n119_), .B(mai_mai_n23_), .Y(mai_mai_n544_));
  NO2        m522(.A(mai_mai_n196_), .B(mai_mai_n37_), .Y(mai_mai_n545_));
  NOi31      m523(.An(mai_mai_n151_), .B(mai_mai_n545_), .C(mai_mai_n314_), .Y(mai_mai_n546_));
  NO2        m524(.A(mai_mai_n546_), .B(mai_mai_n543_), .Y(mai_mai_n547_));
  NO2        m525(.A(mai_mai_n483_), .B(mai_mai_n360_), .Y(mai_mai_n548_));
  INV        m526(.A(mai_mai_n302_), .Y(mai_mai_n549_));
  NO2        m527(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n550_));
  NA2        m528(.A(mai_mai_n176_), .B(i_0_), .Y(mai_mai_n551_));
  NO3        m529(.A(mai_mai_n551_), .B(mai_mai_n324_), .C(mai_mai_n287_), .Y(mai_mai_n552_));
  OR2        m530(.A(i_2_), .B(i_5_), .Y(mai_mai_n553_));
  OR2        m531(.A(mai_mai_n553_), .B(mai_mai_n384_), .Y(mai_mai_n554_));
  NO2        m532(.A(mai_mai_n554_), .B(mai_mai_n460_), .Y(mai_mai_n555_));
  NO3        m533(.A(mai_mai_n555_), .B(mai_mai_n552_), .C(mai_mai_n548_), .Y(mai_mai_n556_));
  NA4        m534(.A(mai_mai_n556_), .B(mai_mai_n547_), .C(mai_mai_n539_), .D(mai_mai_n529_), .Y(mai_mai_n557_));
  NO4        m535(.A(mai_mai_n557_), .B(mai_mai_n516_), .C(mai_mai_n493_), .D(mai_mai_n473_), .Y(mai_mai_n558_));
  NA4        m536(.A(mai_mai_n558_), .B(mai_mai_n411_), .C(mai_mai_n338_), .D(mai_mai_n298_), .Y(mai7));
  NO2        m537(.A(mai_mai_n96_), .B(mai_mai_n55_), .Y(mai_mai_n560_));
  NO2        m538(.A(mai_mai_n112_), .B(mai_mai_n93_), .Y(mai_mai_n561_));
  NA2        m539(.A(mai_mai_n365_), .B(mai_mai_n561_), .Y(mai_mai_n562_));
  NA2        m540(.A(mai_mai_n449_), .B(mai_mai_n85_), .Y(mai_mai_n563_));
  NA2        m541(.A(i_11_), .B(mai_mai_n193_), .Y(mai_mai_n564_));
  INV        m542(.A(mai_mai_n562_), .Y(mai_mai_n565_));
  NA3        m543(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n566_));
  NO2        m544(.A(mai_mai_n233_), .B(i_4_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n567_), .B(i_8_), .Y(mai_mai_n568_));
  NO2        m546(.A(mai_mai_n109_), .B(mai_mai_n566_), .Y(mai_mai_n569_));
  NA2        m547(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n570_));
  OAI210     m548(.A0(mai_mai_n90_), .A1(mai_mai_n201_), .B0(mai_mai_n202_), .Y(mai_mai_n571_));
  NO2        m549(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n572_));
  NA2        m550(.A(i_4_), .B(i_8_), .Y(mai_mai_n573_));
  AOI210     m551(.A0(mai_mai_n573_), .A1(mai_mai_n292_), .B0(mai_mai_n572_), .Y(mai_mai_n574_));
  OAI220     m552(.A0(mai_mai_n574_), .A1(mai_mai_n570_), .B0(mai_mai_n571_), .B1(i_13_), .Y(mai_mai_n575_));
  NO4        m553(.A(mai_mai_n575_), .B(mai_mai_n569_), .C(mai_mai_n565_), .D(mai_mai_n560_), .Y(mai_mai_n576_));
  AOI210     m554(.A0(mai_mai_n133_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n577_));
  AOI210     m555(.A0(mai_mai_n577_), .A1(mai_mai_n233_), .B0(mai_mai_n165_), .Y(mai_mai_n578_));
  OR2        m556(.A(i_6_), .B(i_10_), .Y(mai_mai_n579_));
  NO2        m557(.A(mai_mai_n579_), .B(mai_mai_n23_), .Y(mai_mai_n580_));
  OR3        m558(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n581_));
  NO3        m559(.A(mai_mai_n581_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n582_));
  INV        m560(.A(mai_mai_n198_), .Y(mai_mai_n583_));
  NO2        m561(.A(mai_mai_n582_), .B(mai_mai_n580_), .Y(mai_mai_n584_));
  OA220      m562(.A0(mai_mai_n584_), .A1(mai_mai_n549_), .B0(mai_mai_n578_), .B1(mai_mai_n267_), .Y(mai_mai_n585_));
  AOI210     m563(.A0(mai_mai_n585_), .A1(mai_mai_n576_), .B0(mai_mai_n64_), .Y(mai_mai_n586_));
  NOi21      m564(.An(i_11_), .B(i_7_), .Y(mai_mai_n587_));
  AO210      m565(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n588_));
  NO2        m566(.A(mai_mai_n588_), .B(mai_mai_n587_), .Y(mai_mai_n589_));
  NA2        m567(.A(mai_mai_n589_), .B(mai_mai_n204_), .Y(mai_mai_n590_));
  NO2        m568(.A(mai_mai_n590_), .B(mai_mai_n64_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n89_), .B(mai_mai_n64_), .Y(mai_mai_n592_));
  AO210      m570(.A0(mai_mai_n592_), .A1(mai_mai_n360_), .B0(mai_mai_n41_), .Y(mai_mai_n593_));
  NO3        m571(.A(mai_mai_n256_), .B(mai_mai_n206_), .C(mai_mai_n564_), .Y(mai_mai_n594_));
  OAI210     m572(.A0(mai_mai_n594_), .A1(mai_mai_n224_), .B0(mai_mai_n64_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n385_), .B(mai_mai_n31_), .Y(mai_mai_n596_));
  OR2        m574(.A(mai_mai_n206_), .B(mai_mai_n112_), .Y(mai_mai_n597_));
  NA2        m575(.A(mai_mai_n597_), .B(mai_mai_n596_), .Y(mai_mai_n598_));
  NO2        m576(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n599_));
  NO2        m577(.A(mai_mai_n599_), .B(i_4_), .Y(mai_mai_n600_));
  NA2        m578(.A(mai_mai_n600_), .B(mai_mai_n598_), .Y(mai_mai_n601_));
  NO2        m579(.A(i_1_), .B(i_12_), .Y(mai_mai_n602_));
  NA3        m580(.A(mai_mai_n602_), .B(mai_mai_n114_), .C(mai_mai_n24_), .Y(mai_mai_n603_));
  BUFFER     m581(.A(mai_mai_n603_), .Y(mai_mai_n604_));
  NA4        m582(.A(mai_mai_n604_), .B(mai_mai_n601_), .C(mai_mai_n595_), .D(mai_mai_n593_), .Y(mai_mai_n605_));
  OAI210     m583(.A0(mai_mai_n605_), .A1(mai_mai_n591_), .B0(i_6_), .Y(mai_mai_n606_));
  NO2        m584(.A(i_6_), .B(i_11_), .Y(mai_mai_n607_));
  INV        m585(.A(mai_mai_n419_), .Y(mai_mai_n608_));
  NO4        m586(.A(mai_mai_n214_), .B(mai_mai_n133_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n609_));
  NA2        m587(.A(mai_mai_n609_), .B(mai_mai_n599_), .Y(mai_mai_n610_));
  NA2        m588(.A(mai_mai_n233_), .B(i_6_), .Y(mai_mai_n611_));
  NO3        m589(.A(mai_mai_n579_), .B(mai_mai_n229_), .C(mai_mai_n23_), .Y(mai_mai_n612_));
  AOI210     m590(.A0(i_1_), .A1(mai_mai_n257_), .B0(mai_mai_n612_), .Y(mai_mai_n613_));
  OAI210     m591(.A0(mai_mai_n613_), .A1(mai_mai_n45_), .B0(mai_mai_n610_), .Y(mai_mai_n614_));
  INV        m592(.A(i_2_), .Y(mai_mai_n615_));
  NA2        m593(.A(mai_mai_n143_), .B(i_9_), .Y(mai_mai_n616_));
  NA3        m594(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n617_));
  NO2        m595(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n618_));
  NA3        m596(.A(mai_mai_n618_), .B(mai_mai_n266_), .C(mai_mai_n45_), .Y(mai_mai_n619_));
  OAI220     m597(.A0(mai_mai_n619_), .A1(mai_mai_n617_), .B0(mai_mai_n616_), .B1(mai_mai_n615_), .Y(mai_mai_n620_));
  NA3        m598(.A(mai_mai_n599_), .B(mai_mai_n302_), .C(i_6_), .Y(mai_mai_n621_));
  NO2        m599(.A(mai_mai_n621_), .B(mai_mai_n23_), .Y(mai_mai_n622_));
  AOI210     m600(.A0(mai_mai_n441_), .A1(mai_mai_n395_), .B0(mai_mai_n238_), .Y(mai_mai_n623_));
  NO2        m601(.A(mai_mai_n623_), .B(mai_mai_n570_), .Y(mai_mai_n624_));
  NO2        m602(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n625_));
  OR3        m603(.A(mai_mai_n624_), .B(mai_mai_n622_), .C(mai_mai_n620_), .Y(mai_mai_n626_));
  NO3        m604(.A(mai_mai_n626_), .B(mai_mai_n614_), .C(mai_mai_n608_), .Y(mai_mai_n627_));
  NO2        m605(.A(mai_mai_n233_), .B(mai_mai_n105_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n628_), .B(mai_mai_n587_), .Y(mai_mai_n629_));
  NA2        m607(.A(mai_mai_n629_), .B(i_1_), .Y(mai_mai_n630_));
  NO2        m608(.A(mai_mai_n630_), .B(mai_mai_n581_), .Y(mai_mai_n631_));
  NO2        m609(.A(mai_mai_n391_), .B(mai_mai_n87_), .Y(mai_mai_n632_));
  NA2        m610(.A(mai_mai_n631_), .B(mai_mai_n47_), .Y(mai_mai_n633_));
  NA2        m611(.A(i_3_), .B(mai_mai_n193_), .Y(mai_mai_n634_));
  NO2        m612(.A(mai_mai_n634_), .B(mai_mai_n119_), .Y(mai_mai_n635_));
  AN2        m613(.A(mai_mai_n635_), .B(mai_mai_n504_), .Y(mai_mai_n636_));
  NO2        m614(.A(mai_mai_n229_), .B(mai_mai_n45_), .Y(mai_mai_n637_));
  NO3        m615(.A(mai_mai_n637_), .B(mai_mai_n295_), .C(mai_mai_n234_), .Y(mai_mai_n638_));
  NO2        m616(.A(mai_mai_n122_), .B(mai_mai_n37_), .Y(mai_mai_n639_));
  NO2        m617(.A(mai_mai_n639_), .B(i_6_), .Y(mai_mai_n640_));
  NO2        m618(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n641_));
  NO2        m619(.A(mai_mai_n641_), .B(mai_mai_n64_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n642_), .B(mai_mai_n602_), .Y(mai_mai_n643_));
  NO4        m621(.A(mai_mai_n643_), .B(mai_mai_n640_), .C(mai_mai_n638_), .D(i_4_), .Y(mai_mai_n644_));
  NA2        m622(.A(i_1_), .B(i_3_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n420_), .B(mai_mai_n96_), .Y(mai_mai_n646_));
  AOI210     m624(.A0(mai_mai_n637_), .A1(mai_mai_n540_), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  NO2        m625(.A(mai_mai_n647_), .B(mai_mai_n645_), .Y(mai_mai_n648_));
  NO3        m626(.A(mai_mai_n648_), .B(mai_mai_n644_), .C(mai_mai_n636_), .Y(mai_mai_n649_));
  NA4        m627(.A(mai_mai_n649_), .B(mai_mai_n633_), .C(mai_mai_n627_), .D(mai_mai_n606_), .Y(mai_mai_n650_));
  NO3        m628(.A(mai_mai_n442_), .B(i_3_), .C(i_7_), .Y(mai_mai_n651_));
  NOi21      m629(.An(mai_mai_n651_), .B(i_10_), .Y(mai_mai_n652_));
  OA210      m630(.A0(mai_mai_n652_), .A1(mai_mai_n241_), .B0(mai_mai_n87_), .Y(mai_mai_n653_));
  NA2        m631(.A(mai_mai_n353_), .B(mai_mai_n352_), .Y(mai_mai_n654_));
  NA3        m632(.A(mai_mai_n449_), .B(mai_mai_n484_), .C(mai_mai_n47_), .Y(mai_mai_n655_));
  NA3        m633(.A(mai_mai_n165_), .B(mai_mai_n85_), .C(mai_mai_n87_), .Y(mai_mai_n656_));
  NA3        m634(.A(mai_mai_n656_), .B(mai_mai_n655_), .C(mai_mai_n654_), .Y(mai_mai_n657_));
  OAI210     m635(.A0(mai_mai_n657_), .A1(mai_mai_n653_), .B0(i_1_), .Y(mai_mai_n658_));
  AOI210     m636(.A0(mai_mai_n266_), .A1(mai_mai_n101_), .B0(i_1_), .Y(mai_mai_n659_));
  NO2        m637(.A(mai_mai_n351_), .B(i_2_), .Y(mai_mai_n660_));
  NA2        m638(.A(mai_mai_n660_), .B(mai_mai_n659_), .Y(mai_mai_n661_));
  OAI210     m639(.A0(mai_mai_n621_), .A1(mai_mai_n414_), .B0(mai_mai_n661_), .Y(mai_mai_n662_));
  INV        m640(.A(mai_mai_n662_), .Y(mai_mai_n663_));
  AOI210     m641(.A0(mai_mai_n663_), .A1(mai_mai_n658_), .B0(i_13_), .Y(mai_mai_n664_));
  NO2        m642(.A(mai_mai_n55_), .B(i_12_), .Y(mai_mai_n665_));
  INV        m643(.A(mai_mai_n665_), .Y(mai_mai_n666_));
  NO2        m644(.A(mai_mai_n443_), .B(mai_mai_n24_), .Y(mai_mai_n667_));
  AOI220     m645(.A0(mai_mai_n667_), .A1(mai_mai_n632_), .B0(mai_mai_n241_), .B1(mai_mai_n136_), .Y(mai_mai_n668_));
  OAI220     m646(.A0(mai_mai_n668_), .A1(mai_mai_n41_), .B0(mai_mai_n666_), .B1(mai_mai_n96_), .Y(mai_mai_n669_));
  INV        m647(.A(mai_mai_n669_), .Y(mai_mai_n670_));
  INV        m648(.A(mai_mai_n119_), .Y(mai_mai_n671_));
  AOI220     m649(.A0(mai_mai_n671_), .A1(mai_mai_n73_), .B0(mai_mai_n367_), .B1(mai_mai_n618_), .Y(mai_mai_n672_));
  NO2        m650(.A(mai_mai_n672_), .B(mai_mai_n239_), .Y(mai_mai_n673_));
  AOI210     m651(.A0(mai_mai_n414_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n674_));
  NOi31      m652(.An(mai_mai_n674_), .B(mai_mai_n563_), .C(mai_mai_n45_), .Y(mai_mai_n675_));
  NA2        m653(.A(mai_mai_n132_), .B(i_13_), .Y(mai_mai_n676_));
  NO2        m654(.A(mai_mai_n617_), .B(mai_mai_n119_), .Y(mai_mai_n677_));
  INV        m655(.A(mai_mai_n677_), .Y(mai_mai_n678_));
  OAI220     m656(.A0(mai_mai_n678_), .A1(mai_mai_n72_), .B0(mai_mai_n676_), .B1(mai_mai_n659_), .Y(mai_mai_n679_));
  NO3        m657(.A(mai_mai_n72_), .B(mai_mai_n32_), .C(mai_mai_n105_), .Y(mai_mai_n680_));
  NA2        m658(.A(mai_mai_n26_), .B(mai_mai_n193_), .Y(mai_mai_n681_));
  NA2        m659(.A(mai_mai_n681_), .B(i_7_), .Y(mai_mai_n682_));
  NO3        m660(.A(mai_mai_n443_), .B(mai_mai_n233_), .C(mai_mai_n87_), .Y(mai_mai_n683_));
  AOI210     m661(.A0(mai_mai_n683_), .A1(mai_mai_n682_), .B0(mai_mai_n680_), .Y(mai_mai_n684_));
  AOI220     m662(.A0(mai_mai_n367_), .A1(mai_mai_n618_), .B0(mai_mai_n95_), .B1(mai_mai_n106_), .Y(mai_mai_n685_));
  OAI220     m663(.A0(mai_mai_n685_), .A1(mai_mai_n568_), .B0(mai_mai_n684_), .B1(mai_mai_n583_), .Y(mai_mai_n686_));
  NO4        m664(.A(mai_mai_n686_), .B(mai_mai_n679_), .C(mai_mai_n675_), .D(mai_mai_n673_), .Y(mai_mai_n687_));
  OR2        m665(.A(i_11_), .B(i_6_), .Y(mai_mai_n688_));
  NA3        m666(.A(mai_mai_n567_), .B(mai_mai_n681_), .C(i_7_), .Y(mai_mai_n689_));
  AOI210     m667(.A0(mai_mai_n689_), .A1(mai_mai_n678_), .B0(mai_mai_n688_), .Y(mai_mai_n690_));
  NA3        m668(.A(mai_mai_n385_), .B(mai_mai_n572_), .C(mai_mai_n101_), .Y(mai_mai_n691_));
  NA2        m669(.A(mai_mai_n607_), .B(i_13_), .Y(mai_mai_n692_));
  NA2        m670(.A(mai_mai_n106_), .B(mai_mai_n681_), .Y(mai_mai_n693_));
  NAi21      m671(.An(i_11_), .B(i_12_), .Y(mai_mai_n694_));
  NOi41      m672(.An(mai_mai_n115_), .B(mai_mai_n694_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n695_));
  NA2        m673(.A(mai_mai_n695_), .B(mai_mai_n693_), .Y(mai_mai_n696_));
  NA3        m674(.A(mai_mai_n696_), .B(mai_mai_n692_), .C(mai_mai_n691_), .Y(mai_mai_n697_));
  OAI210     m675(.A0(mai_mai_n697_), .A1(mai_mai_n690_), .B0(mai_mai_n64_), .Y(mai_mai_n698_));
  NO2        m676(.A(i_2_), .B(i_12_), .Y(mai_mai_n699_));
  NA2        m677(.A(mai_mai_n350_), .B(mai_mai_n699_), .Y(mai_mai_n700_));
  NA2        m678(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n701_));
  NO3        m679(.A(mai_mai_n701_), .B(mai_mai_n365_), .C(mai_mai_n567_), .Y(mai_mai_n702_));
  OAI210     m680(.A0(mai_mai_n702_), .A1(mai_mai_n352_), .B0(mai_mai_n350_), .Y(mai_mai_n703_));
  NO2        m681(.A(mai_mai_n133_), .B(i_2_), .Y(mai_mai_n704_));
  NA2        m682(.A(mai_mai_n703_), .B(mai_mai_n700_), .Y(mai_mai_n705_));
  NA3        m683(.A(mai_mai_n705_), .B(mai_mai_n46_), .C(mai_mai_n223_), .Y(mai_mai_n706_));
  NA4        m684(.A(mai_mai_n706_), .B(mai_mai_n698_), .C(mai_mai_n687_), .D(mai_mai_n670_), .Y(mai_mai_n707_));
  OR4        m685(.A(mai_mai_n707_), .B(mai_mai_n664_), .C(mai_mai_n650_), .D(mai_mai_n586_), .Y(mai5));
  NA2        m686(.A(mai_mai_n629_), .B(mai_mai_n269_), .Y(mai_mai_n709_));
  AN2        m687(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n710_));
  NA3        m688(.A(mai_mai_n710_), .B(mai_mai_n699_), .C(mai_mai_n112_), .Y(mai_mai_n711_));
  NO2        m689(.A(mai_mai_n568_), .B(i_11_), .Y(mai_mai_n712_));
  NA2        m690(.A(mai_mai_n90_), .B(mai_mai_n712_), .Y(mai_mai_n713_));
  NA3        m691(.A(mai_mai_n713_), .B(mai_mai_n711_), .C(mai_mai_n709_), .Y(mai_mai_n714_));
  NO3        m692(.A(i_11_), .B(mai_mai_n233_), .C(i_13_), .Y(mai_mai_n715_));
  NO2        m693(.A(mai_mai_n129_), .B(mai_mai_n23_), .Y(mai_mai_n716_));
  NA2        m694(.A(i_12_), .B(i_8_), .Y(mai_mai_n717_));
  OAI210     m695(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  INV        m696(.A(mai_mai_n413_), .Y(mai_mai_n719_));
  AOI220     m697(.A0(mai_mai_n302_), .A1(mai_mai_n544_), .B0(mai_mai_n718_), .B1(mai_mai_n716_), .Y(mai_mai_n720_));
  INV        m698(.A(mai_mai_n720_), .Y(mai_mai_n721_));
  NO2        m699(.A(mai_mai_n721_), .B(mai_mai_n714_), .Y(mai_mai_n722_));
  INV        m700(.A(mai_mai_n173_), .Y(mai_mai_n723_));
  INV        m701(.A(mai_mai_n241_), .Y(mai_mai_n724_));
  OAI210     m702(.A0(mai_mai_n660_), .A1(mai_mai_n415_), .B0(mai_mai_n115_), .Y(mai_mai_n725_));
  AOI210     m703(.A0(mai_mai_n725_), .A1(mai_mai_n724_), .B0(mai_mai_n723_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n420_), .B(mai_mai_n26_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n727_), .B(mai_mai_n395_), .Y(mai_mai_n728_));
  NA2        m706(.A(mai_mai_n728_), .B(i_2_), .Y(mai_mai_n729_));
  INV        m707(.A(mai_mai_n729_), .Y(mai_mai_n730_));
  AOI210     m708(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n392_), .Y(mai_mai_n731_));
  AOI210     m709(.A0(mai_mai_n731_), .A1(mai_mai_n730_), .B0(mai_mai_n726_), .Y(mai_mai_n732_));
  NO2        m710(.A(mai_mai_n190_), .B(mai_mai_n130_), .Y(mai_mai_n733_));
  OAI210     m711(.A0(mai_mai_n733_), .A1(mai_mai_n716_), .B0(i_2_), .Y(mai_mai_n734_));
  INV        m712(.A(mai_mai_n174_), .Y(mai_mai_n735_));
  NO3        m713(.A(mai_mai_n588_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n736_));
  AOI210     m714(.A0(mai_mai_n735_), .A1(mai_mai_n90_), .B0(mai_mai_n736_), .Y(mai_mai_n737_));
  AOI210     m715(.A0(mai_mai_n737_), .A1(mai_mai_n734_), .B0(mai_mai_n193_), .Y(mai_mai_n738_));
  OA210      m716(.A0(mai_mai_n589_), .A1(mai_mai_n131_), .B0(i_13_), .Y(mai_mai_n739_));
  NA2        m717(.A(mai_mai_n198_), .B(mai_mai_n201_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n157_), .B(mai_mai_n564_), .Y(mai_mai_n741_));
  AOI210     m719(.A0(mai_mai_n741_), .A1(mai_mai_n740_), .B0(mai_mai_n355_), .Y(mai_mai_n742_));
  AOI210     m720(.A0(mai_mai_n206_), .A1(mai_mai_n153_), .B0(mai_mai_n484_), .Y(mai_mai_n743_));
  NA2        m721(.A(mai_mai_n743_), .B(mai_mai_n395_), .Y(mai_mai_n744_));
  NO2        m722(.A(mai_mai_n106_), .B(mai_mai_n45_), .Y(mai_mai_n745_));
  INV        m723(.A(mai_mai_n288_), .Y(mai_mai_n746_));
  NA4        m724(.A(mai_mai_n746_), .B(mai_mai_n292_), .C(mai_mai_n129_), .D(mai_mai_n43_), .Y(mai_mai_n747_));
  OAI210     m725(.A0(mai_mai_n747_), .A1(mai_mai_n745_), .B0(mai_mai_n744_), .Y(mai_mai_n748_));
  NO4        m726(.A(mai_mai_n748_), .B(mai_mai_n742_), .C(mai_mai_n739_), .D(mai_mai_n738_), .Y(mai_mai_n749_));
  NA2        m727(.A(mai_mai_n544_), .B(mai_mai_n28_), .Y(mai_mai_n750_));
  NA2        m728(.A(mai_mai_n715_), .B(mai_mai_n275_), .Y(mai_mai_n751_));
  NA2        m729(.A(mai_mai_n751_), .B(mai_mai_n750_), .Y(mai_mai_n752_));
  NO2        m730(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n753_));
  NO2        m731(.A(mai_mai_n753_), .B(mai_mai_n131_), .Y(mai_mai_n754_));
  NO2        m732(.A(mai_mai_n754_), .B(mai_mai_n564_), .Y(mai_mai_n755_));
  AOI220     m733(.A0(mai_mai_n755_), .A1(mai_mai_n36_), .B0(mai_mai_n752_), .B1(mai_mai_n47_), .Y(mai_mai_n756_));
  NA4        m734(.A(mai_mai_n756_), .B(mai_mai_n749_), .C(mai_mai_n732_), .D(mai_mai_n722_), .Y(mai6));
  NO2        m735(.A(mai_mai_n185_), .B(mai_mai_n144_), .Y(mai_mai_n758_));
  NA2        m736(.A(mai_mai_n758_), .B(mai_mai_n704_), .Y(mai_mai_n759_));
  NA4        m737(.A(mai_mai_n369_), .B(mai_mai_n448_), .C(mai_mai_n72_), .D(mai_mai_n105_), .Y(mai_mai_n760_));
  INV        m738(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  NO2        m739(.A(mai_mai_n219_), .B(mai_mai_n453_), .Y(mai_mai_n762_));
  NO2        m740(.A(i_11_), .B(i_9_), .Y(mai_mai_n763_));
  NO2        m741(.A(mai_mai_n761_), .B(mai_mai_n313_), .Y(mai_mai_n764_));
  AO210      m742(.A0(mai_mai_n764_), .A1(mai_mai_n759_), .B0(i_12_), .Y(mai_mai_n765_));
  NA2        m743(.A(mai_mai_n356_), .B(mai_mai_n318_), .Y(mai_mai_n766_));
  NA2        m744(.A(mai_mai_n550_), .B(mai_mai_n64_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n652_), .B(mai_mai_n72_), .Y(mai_mai_n768_));
  BUFFER     m746(.A(mai_mai_n592_), .Y(mai_mai_n769_));
  NA4        m747(.A(mai_mai_n769_), .B(mai_mai_n768_), .C(mai_mai_n767_), .D(mai_mai_n766_), .Y(mai_mai_n770_));
  INV        m748(.A(mai_mai_n195_), .Y(mai_mai_n771_));
  AOI220     m749(.A0(mai_mai_n771_), .A1(mai_mai_n763_), .B0(mai_mai_n770_), .B1(mai_mai_n74_), .Y(mai_mai_n772_));
  INV        m750(.A(mai_mai_n312_), .Y(mai_mai_n773_));
  NA2        m751(.A(mai_mai_n76_), .B(mai_mai_n136_), .Y(mai_mai_n774_));
  INV        m752(.A(mai_mai_n129_), .Y(mai_mai_n775_));
  NA2        m753(.A(mai_mai_n775_), .B(mai_mai_n47_), .Y(mai_mai_n776_));
  AOI210     m754(.A0(mai_mai_n776_), .A1(mai_mai_n774_), .B0(mai_mai_n773_), .Y(mai_mai_n777_));
  NO2        m755(.A(mai_mai_n248_), .B(i_9_), .Y(mai_mai_n778_));
  NA2        m756(.A(mai_mai_n778_), .B(mai_mai_n753_), .Y(mai_mai_n779_));
  NO2        m757(.A(mai_mai_n779_), .B(mai_mai_n185_), .Y(mai_mai_n780_));
  NO2        m758(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n781_));
  NA3        m759(.A(mai_mai_n781_), .B(mai_mai_n439_), .C(mai_mai_n369_), .Y(mai_mai_n782_));
  NAi32      m760(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n783_));
  NO2        m761(.A(mai_mai_n688_), .B(mai_mai_n783_), .Y(mai_mai_n784_));
  OAI210     m762(.A0(mai_mai_n651_), .A1(mai_mai_n532_), .B0(mai_mai_n531_), .Y(mai_mai_n785_));
  NAi31      m763(.An(mai_mai_n784_), .B(mai_mai_n785_), .C(mai_mai_n782_), .Y(mai_mai_n786_));
  OR3        m764(.A(mai_mai_n786_), .B(mai_mai_n780_), .C(mai_mai_n777_), .Y(mai_mai_n787_));
  AO220      m765(.A0(mai_mai_n343_), .A1(mai_mai_n334_), .B0(mai_mai_n371_), .B1(mai_mai_n564_), .Y(mai_mai_n788_));
  NA3        m766(.A(mai_mai_n788_), .B(mai_mai_n253_), .C(i_7_), .Y(mai_mai_n789_));
  BUFFER     m767(.A(mai_mai_n589_), .Y(mai_mai_n790_));
  NA3        m768(.A(mai_mai_n790_), .B(mai_mai_n152_), .C(mai_mai_n70_), .Y(mai_mai_n791_));
  OR2        m769(.A(mai_mai_n719_), .B(mai_mai_n36_), .Y(mai_mai_n792_));
  NA3        m770(.A(mai_mai_n792_), .B(mai_mai_n791_), .C(mai_mai_n789_), .Y(mai_mai_n793_));
  OAI210     m771(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n88_), .Y(mai_mai_n794_));
  AOI220     m772(.A0(mai_mai_n794_), .A1(mai_mai_n531_), .B0(mai_mai_n762_), .B1(mai_mai_n682_), .Y(mai_mai_n795_));
  NA2        m773(.A(mai_mai_n371_), .B(mai_mai_n71_), .Y(mai_mai_n796_));
  NA3        m774(.A(mai_mai_n796_), .B(mai_mai_n795_), .C(mai_mai_n571_), .Y(mai_mai_n797_));
  AO210      m775(.A0(mai_mai_n484_), .A1(mai_mai_n47_), .B0(mai_mai_n89_), .Y(mai_mai_n798_));
  NA3        m776(.A(mai_mai_n798_), .B(mai_mai_n449_), .C(mai_mai_n217_), .Y(mai_mai_n799_));
  AOI210     m777(.A0(mai_mai_n415_), .A1(mai_mai_n413_), .B0(mai_mai_n530_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n579_), .B(mai_mai_n106_), .Y(mai_mai_n801_));
  OAI210     m779(.A0(mai_mai_n801_), .A1(mai_mai_n116_), .B0(mai_mai_n382_), .Y(mai_mai_n802_));
  INV        m780(.A(mai_mai_n554_), .Y(mai_mai_n803_));
  NA3        m781(.A(mai_mai_n803_), .B(mai_mai_n312_), .C(i_7_), .Y(mai_mai_n804_));
  NA4        m782(.A(mai_mai_n804_), .B(mai_mai_n802_), .C(mai_mai_n800_), .D(mai_mai_n799_), .Y(mai_mai_n805_));
  NO4        m783(.A(mai_mai_n805_), .B(mai_mai_n797_), .C(mai_mai_n793_), .D(mai_mai_n787_), .Y(mai_mai_n806_));
  NA4        m784(.A(mai_mai_n806_), .B(mai_mai_n772_), .C(mai_mai_n765_), .D(mai_mai_n362_), .Y(mai3));
  NA2        m785(.A(i_12_), .B(i_10_), .Y(mai_mai_n808_));
  NA2        m786(.A(i_6_), .B(i_7_), .Y(mai_mai_n809_));
  NO2        m787(.A(mai_mai_n809_), .B(i_0_), .Y(mai_mai_n810_));
  NO2        m788(.A(i_11_), .B(mai_mai_n233_), .Y(mai_mai_n811_));
  OAI210     m789(.A0(mai_mai_n810_), .A1(mai_mai_n281_), .B0(mai_mai_n811_), .Y(mai_mai_n812_));
  NO2        m790(.A(mai_mai_n812_), .B(mai_mai_n193_), .Y(mai_mai_n813_));
  NO3        m791(.A(mai_mai_n416_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n814_));
  OA210      m792(.A0(mai_mai_n814_), .A1(mai_mai_n813_), .B0(mai_mai_n176_), .Y(mai_mai_n815_));
  NOi21      m793(.An(mai_mai_n100_), .B(mai_mai_n728_), .Y(mai_mai_n816_));
  NO3        m794(.A(mai_mai_n597_), .B(mai_mai_n420_), .C(mai_mai_n136_), .Y(mai_mai_n817_));
  AN2        m795(.A(mai_mai_n418_), .B(mai_mai_n56_), .Y(mai_mai_n818_));
  NO3        m796(.A(mai_mai_n818_), .B(mai_mai_n817_), .C(mai_mai_n816_), .Y(mai_mai_n819_));
  NO2        m797(.A(mai_mai_n819_), .B(mai_mai_n49_), .Y(mai_mai_n820_));
  NO4        m798(.A(mai_mai_n358_), .B(mai_mai_n364_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n821_));
  NA2        m799(.A(mai_mai_n185_), .B(mai_mai_n540_), .Y(mai_mai_n822_));
  NOi21      m800(.An(mai_mai_n822_), .B(mai_mai_n821_), .Y(mai_mai_n823_));
  NO2        m801(.A(mai_mai_n823_), .B(mai_mai_n64_), .Y(mai_mai_n824_));
  NOi21      m802(.An(i_5_), .B(i_9_), .Y(mai_mai_n825_));
  NA2        m803(.A(mai_mai_n825_), .B(mai_mai_n412_), .Y(mai_mai_n826_));
  BUFFER     m804(.A(mai_mai_n266_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n827_), .B(mai_mai_n441_), .Y(mai_mai_n828_));
  NO3        m806(.A(mai_mai_n388_), .B(mai_mai_n266_), .C(mai_mai_n74_), .Y(mai_mai_n829_));
  NO2        m807(.A(mai_mai_n177_), .B(mai_mai_n153_), .Y(mai_mai_n830_));
  AOI210     m808(.A0(mai_mai_n830_), .A1(mai_mai_n240_), .B0(mai_mai_n829_), .Y(mai_mai_n831_));
  OAI220     m809(.A0(mai_mai_n831_), .A1(mai_mai_n183_), .B0(mai_mai_n828_), .B1(mai_mai_n826_), .Y(mai_mai_n832_));
  NO4        m810(.A(mai_mai_n832_), .B(mai_mai_n824_), .C(mai_mai_n820_), .D(mai_mai_n815_), .Y(mai_mai_n833_));
  NA2        m811(.A(mai_mai_n185_), .B(mai_mai_n24_), .Y(mai_mai_n834_));
  NO2        m812(.A(mai_mai_n639_), .B(mai_mai_n561_), .Y(mai_mai_n835_));
  NO2        m813(.A(mai_mai_n835_), .B(mai_mai_n834_), .Y(mai_mai_n836_));
  INV        m814(.A(mai_mai_n836_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n369_), .B(mai_mai_n282_), .Y(mai_mai_n838_));
  NA2        m816(.A(mai_mai_n838_), .B(mai_mai_n677_), .Y(mai_mai_n839_));
  NA2        m817(.A(mai_mai_n541_), .B(i_0_), .Y(mai_mai_n840_));
  NO3        m818(.A(mai_mai_n840_), .B(mai_mai_n366_), .C(mai_mai_n90_), .Y(mai_mai_n841_));
  NO4        m819(.A(mai_mai_n553_), .B(mai_mai_n214_), .C(mai_mai_n392_), .D(mai_mai_n384_), .Y(mai_mai_n842_));
  AOI210     m820(.A0(mai_mai_n842_), .A1(i_11_), .B0(mai_mai_n841_), .Y(mai_mai_n843_));
  NA2        m821(.A(mai_mai_n715_), .B(mai_mai_n313_), .Y(mai_mai_n844_));
  AOI210     m822(.A0(mai_mai_n449_), .A1(mai_mai_n90_), .B0(mai_mai_n59_), .Y(mai_mai_n845_));
  NO2        m823(.A(mai_mai_n845_), .B(mai_mai_n844_), .Y(mai_mai_n846_));
  NO2        m824(.A(mai_mai_n250_), .B(mai_mai_n159_), .Y(mai_mai_n847_));
  NA2        m825(.A(i_0_), .B(i_10_), .Y(mai_mai_n848_));
  INV        m826(.A(mai_mai_n503_), .Y(mai_mai_n849_));
  NO4        m827(.A(mai_mai_n119_), .B(mai_mai_n59_), .C(mai_mai_n634_), .D(i_5_), .Y(mai_mai_n850_));
  AO220      m828(.A0(mai_mai_n850_), .A1(mai_mai_n849_), .B0(mai_mai_n847_), .B1(i_6_), .Y(mai_mai_n851_));
  AOI220     m829(.A0(mai_mai_n316_), .A1(mai_mai_n102_), .B0(mai_mai_n185_), .B1(mai_mai_n85_), .Y(mai_mai_n852_));
  NA2        m830(.A(mai_mai_n535_), .B(i_4_), .Y(mai_mai_n853_));
  NA2        m831(.A(mai_mai_n188_), .B(mai_mai_n201_), .Y(mai_mai_n854_));
  OAI220     m832(.A0(mai_mai_n854_), .A1(mai_mai_n844_), .B0(mai_mai_n853_), .B1(mai_mai_n852_), .Y(mai_mai_n855_));
  NO3        m833(.A(mai_mai_n855_), .B(mai_mai_n851_), .C(mai_mai_n846_), .Y(mai_mai_n856_));
  NA4        m834(.A(mai_mai_n856_), .B(mai_mai_n843_), .C(mai_mai_n839_), .D(mai_mai_n837_), .Y(mai_mai_n857_));
  NO2        m835(.A(mai_mai_n107_), .B(mai_mai_n37_), .Y(mai_mai_n858_));
  NA2        m836(.A(i_11_), .B(i_9_), .Y(mai_mai_n859_));
  NO3        m837(.A(i_12_), .B(mai_mai_n859_), .C(mai_mai_n570_), .Y(mai_mai_n860_));
  AN2        m838(.A(mai_mai_n860_), .B(mai_mai_n858_), .Y(mai_mai_n861_));
  NO2        m839(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n862_));
  NA2        m840(.A(mai_mai_n370_), .B(mai_mai_n181_), .Y(mai_mai_n863_));
  INV        m841(.A(mai_mai_n863_), .Y(mai_mai_n864_));
  NO2        m842(.A(mai_mai_n859_), .B(mai_mai_n74_), .Y(mai_mai_n865_));
  NO2        m843(.A(mai_mai_n177_), .B(i_0_), .Y(mai_mai_n866_));
  INV        m844(.A(mai_mai_n866_), .Y(mai_mai_n867_));
  NA2        m845(.A(mai_mai_n439_), .B(mai_mai_n227_), .Y(mai_mai_n868_));
  AOI210     m846(.A0(mai_mai_n353_), .A1(mai_mai_n42_), .B0(mai_mai_n381_), .Y(mai_mai_n869_));
  OAI220     m847(.A0(mai_mai_n869_), .A1(mai_mai_n826_), .B0(mai_mai_n868_), .B1(mai_mai_n867_), .Y(mai_mai_n870_));
  NO3        m848(.A(mai_mai_n870_), .B(mai_mai_n864_), .C(mai_mai_n861_), .Y(mai_mai_n871_));
  NA2        m849(.A(mai_mai_n625_), .B(mai_mai_n126_), .Y(mai_mai_n872_));
  NO2        m850(.A(i_6_), .B(mai_mai_n872_), .Y(mai_mai_n873_));
  NA2        m851(.A(mai_mai_n173_), .B(mai_mai_n107_), .Y(mai_mai_n874_));
  INV        m852(.A(mai_mai_n873_), .Y(mai_mai_n875_));
  NOi21      m853(.An(i_7_), .B(i_5_), .Y(mai_mai_n876_));
  NOi31      m854(.An(mai_mai_n876_), .B(i_0_), .C(mai_mai_n694_), .Y(mai_mai_n877_));
  NA3        m855(.A(mai_mai_n877_), .B(mai_mai_n365_), .C(i_6_), .Y(mai_mai_n878_));
  BUFFER     m856(.A(mai_mai_n878_), .Y(mai_mai_n879_));
  NO3        m857(.A(mai_mai_n376_), .B(mai_mai_n346_), .C(mai_mai_n342_), .Y(mai_mai_n880_));
  NO2        m858(.A(mai_mai_n260_), .B(mai_mai_n303_), .Y(mai_mai_n881_));
  NO2        m859(.A(mai_mai_n694_), .B(mai_mai_n255_), .Y(mai_mai_n882_));
  AOI210     m860(.A0(mai_mai_n882_), .A1(mai_mai_n881_), .B0(mai_mai_n880_), .Y(mai_mai_n883_));
  NA4        m861(.A(mai_mai_n883_), .B(mai_mai_n879_), .C(mai_mai_n875_), .D(mai_mai_n871_), .Y(mai_mai_n884_));
  NO2        m862(.A(mai_mai_n834_), .B(mai_mai_n236_), .Y(mai_mai_n885_));
  AN2        m863(.A(mai_mai_n315_), .B(mai_mai_n313_), .Y(mai_mai_n886_));
  AN2        m864(.A(mai_mai_n886_), .B(mai_mai_n830_), .Y(mai_mai_n887_));
  OAI210     m865(.A0(mai_mai_n887_), .A1(mai_mai_n885_), .B0(i_10_), .Y(mai_mai_n888_));
  NO2        m866(.A(mai_mai_n808_), .B(mai_mai_n302_), .Y(mai_mai_n889_));
  OA210      m867(.A0(mai_mai_n439_), .A1(mai_mai_n222_), .B0(mai_mai_n438_), .Y(mai_mai_n890_));
  NA2        m868(.A(mai_mai_n889_), .B(mai_mai_n865_), .Y(mai_mai_n891_));
  NA2        m869(.A(mai_mai_n865_), .B(mai_mai_n292_), .Y(mai_mai_n892_));
  OAI210     m870(.A0(i_2_), .A1(mai_mai_n187_), .B0(mai_mai_n892_), .Y(mai_mai_n893_));
  NA2        m871(.A(mai_mai_n893_), .B(mai_mai_n439_), .Y(mai_mai_n894_));
  NA2        m872(.A(mai_mai_n96_), .B(mai_mai_n45_), .Y(mai_mai_n895_));
  NO2        m873(.A(mai_mai_n76_), .B(mai_mai_n717_), .Y(mai_mai_n896_));
  AOI220     m874(.A0(mai_mai_n896_), .A1(mai_mai_n895_), .B0(mai_mai_n176_), .B1(mai_mai_n561_), .Y(mai_mai_n897_));
  NO2        m875(.A(mai_mai_n897_), .B(mai_mai_n48_), .Y(mai_mai_n898_));
  NO3        m876(.A(mai_mai_n553_), .B(mai_mai_n341_), .C(mai_mai_n24_), .Y(mai_mai_n899_));
  AOI210     m877(.A0(mai_mai_n667_), .A1(mai_mai_n512_), .B0(mai_mai_n899_), .Y(mai_mai_n900_));
  NAi21      m878(.An(i_9_), .B(i_5_), .Y(mai_mai_n901_));
  NO2        m879(.A(mai_mai_n901_), .B(mai_mai_n376_), .Y(mai_mai_n902_));
  NO2        m880(.A(mai_mai_n566_), .B(mai_mai_n109_), .Y(mai_mai_n903_));
  AOI220     m881(.A0(mai_mai_n903_), .A1(i_0_), .B0(mai_mai_n902_), .B1(mai_mai_n589_), .Y(mai_mai_n904_));
  OAI220     m882(.A0(mai_mai_n904_), .A1(mai_mai_n87_), .B0(mai_mai_n900_), .B1(mai_mai_n174_), .Y(mai_mai_n905_));
  NO3        m883(.A(mai_mai_n905_), .B(mai_mai_n898_), .C(mai_mai_n487_), .Y(mai_mai_n906_));
  NA4        m884(.A(mai_mai_n906_), .B(mai_mai_n894_), .C(mai_mai_n891_), .D(mai_mai_n888_), .Y(mai_mai_n907_));
  NO3        m885(.A(mai_mai_n907_), .B(mai_mai_n884_), .C(mai_mai_n857_), .Y(mai_mai_n908_));
  NO2        m886(.A(i_0_), .B(mai_mai_n694_), .Y(mai_mai_n909_));
  NA2        m887(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n910_));
  INV        m888(.A(mai_mai_n910_), .Y(mai_mai_n911_));
  NO3        m889(.A(mai_mai_n109_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n912_));
  AO220      m890(.A0(mai_mai_n912_), .A1(mai_mai_n911_), .B0(mai_mai_n909_), .B1(mai_mai_n176_), .Y(mai_mai_n913_));
  AOI210     m891(.A0(mai_mai_n767_), .A1(mai_mai_n654_), .B0(mai_mai_n874_), .Y(mai_mai_n914_));
  AOI210     m892(.A0(mai_mai_n913_), .A1(mai_mai_n331_), .B0(mai_mai_n914_), .Y(mai_mai_n915_));
  NA2        m893(.A(mai_mai_n704_), .B(mai_mai_n151_), .Y(mai_mai_n916_));
  INV        m894(.A(mai_mai_n916_), .Y(mai_mai_n917_));
  NA3        m895(.A(mai_mai_n917_), .B(mai_mai_n641_), .C(mai_mai_n74_), .Y(mai_mai_n918_));
  NO2        m896(.A(mai_mai_n785_), .B(mai_mai_n376_), .Y(mai_mai_n919_));
  NA3        m897(.A(mai_mai_n810_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n920_));
  NA2        m898(.A(mai_mai_n811_), .B(i_9_), .Y(mai_mai_n921_));
  AOI210     m899(.A0(mai_mai_n920_), .A1(mai_mai_n464_), .B0(mai_mai_n921_), .Y(mai_mai_n922_));
  OAI210     m900(.A0(mai_mai_n240_), .A1(i_9_), .B0(mai_mai_n226_), .Y(mai_mai_n923_));
  AOI210     m901(.A0(mai_mai_n923_), .A1(mai_mai_n840_), .B0(mai_mai_n159_), .Y(mai_mai_n924_));
  NO3        m902(.A(mai_mai_n924_), .B(mai_mai_n922_), .C(mai_mai_n919_), .Y(mai_mai_n925_));
  NA3        m903(.A(mai_mai_n925_), .B(mai_mai_n918_), .C(mai_mai_n915_), .Y(mai_mai_n926_));
  NA2        m904(.A(mai_mai_n886_), .B(mai_mai_n355_), .Y(mai_mai_n927_));
  AOI210     m905(.A0(mai_mai_n287_), .A1(mai_mai_n166_), .B0(mai_mai_n927_), .Y(mai_mai_n928_));
  NA3        m906(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n929_));
  NA2        m907(.A(mai_mai_n862_), .B(mai_mai_n454_), .Y(mai_mai_n930_));
  AOI210     m908(.A0(mai_mai_n929_), .A1(mai_mai_n166_), .B0(mai_mai_n930_), .Y(mai_mai_n931_));
  NO2        m909(.A(mai_mai_n931_), .B(mai_mai_n928_), .Y(mai_mai_n932_));
  NO3        m910(.A(mai_mai_n848_), .B(mai_mai_n825_), .C(mai_mai_n190_), .Y(mai_mai_n933_));
  AOI220     m911(.A0(mai_mai_n933_), .A1(i_11_), .B0(mai_mai_n536_), .B1(mai_mai_n76_), .Y(mai_mai_n934_));
  NO3        m912(.A(mai_mai_n208_), .B(mai_mai_n364_), .C(i_0_), .Y(mai_mai_n935_));
  OAI210     m913(.A0(mai_mai_n935_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n936_));
  INV        m914(.A(mai_mai_n217_), .Y(mai_mai_n937_));
  OAI220     m915(.A0(mai_mai_n497_), .A1(mai_mai_n144_), .B0(mai_mai_n611_), .B1(mai_mai_n583_), .Y(mai_mai_n938_));
  NA3        m916(.A(mai_mai_n938_), .B(mai_mai_n372_), .C(mai_mai_n937_), .Y(mai_mai_n939_));
  NA4        m917(.A(mai_mai_n939_), .B(mai_mai_n936_), .C(mai_mai_n934_), .D(mai_mai_n932_), .Y(mai_mai_n940_));
  NO2        m918(.A(mai_mai_n239_), .B(mai_mai_n96_), .Y(mai_mai_n941_));
  AOI210     m919(.A0(mai_mai_n941_), .A1(mai_mai_n909_), .B0(mai_mai_n113_), .Y(mai_mai_n942_));
  AOI220     m920(.A0(mai_mai_n876_), .A1(mai_mai_n454_), .B0(mai_mai_n810_), .B1(mai_mai_n167_), .Y(mai_mai_n943_));
  NA2        m921(.A(mai_mai_n334_), .B(mai_mai_n178_), .Y(mai_mai_n944_));
  OA220      m922(.A0(mai_mai_n944_), .A1(mai_mai_n943_), .B0(mai_mai_n942_), .B1(i_5_), .Y(mai_mai_n945_));
  AOI210     m923(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n177_), .Y(mai_mai_n946_));
  NA2        m924(.A(mai_mai_n946_), .B(mai_mai_n890_), .Y(mai_mai_n947_));
  NA3        m925(.A(mai_mai_n580_), .B(mai_mai_n185_), .C(mai_mai_n85_), .Y(mai_mai_n948_));
  NA2        m926(.A(mai_mai_n948_), .B(mai_mai_n510_), .Y(mai_mai_n949_));
  NA2        m927(.A(mai_mai_n459_), .B(mai_mai_n452_), .Y(mai_mai_n950_));
  NO2        m928(.A(mai_mai_n950_), .B(mai_mai_n949_), .Y(mai_mai_n951_));
  NA3        m929(.A(mai_mai_n369_), .B(mai_mai_n173_), .C(mai_mai_n172_), .Y(mai_mai_n952_));
  NA3        m930(.A(mai_mai_n862_), .B(mai_mai_n281_), .C(mai_mai_n226_), .Y(mai_mai_n953_));
  NA2        m931(.A(mai_mai_n953_), .B(mai_mai_n952_), .Y(mai_mai_n954_));
  NO3        m932(.A(mai_mai_n859_), .B(mai_mai_n217_), .C(mai_mai_n190_), .Y(mai_mai_n955_));
  NO2        m933(.A(mai_mai_n955_), .B(mai_mai_n954_), .Y(mai_mai_n956_));
  NA4        m934(.A(mai_mai_n956_), .B(mai_mai_n951_), .C(mai_mai_n947_), .D(mai_mai_n945_), .Y(mai_mai_n957_));
  INV        m935(.A(mai_mai_n582_), .Y(mai_mai_n958_));
  NO3        m936(.A(mai_mai_n958_), .B(mai_mai_n526_), .C(mai_mai_n328_), .Y(mai_mai_n959_));
  NO2        m937(.A(mai_mai_n87_), .B(i_5_), .Y(mai_mai_n960_));
  NA3        m938(.A(mai_mai_n811_), .B(mai_mai_n114_), .C(mai_mai_n129_), .Y(mai_mai_n961_));
  INV        m939(.A(mai_mai_n961_), .Y(mai_mai_n962_));
  AOI210     m940(.A0(mai_mai_n962_), .A1(mai_mai_n960_), .B0(mai_mai_n959_), .Y(mai_mai_n963_));
  NA2        m941(.A(mai_mai_n292_), .B(i_5_), .Y(mai_mai_n964_));
  NAi31      m942(.An(mai_mai_n238_), .B(mai_mai_n964_), .C(mai_mai_n239_), .Y(mai_mai_n965_));
  NO4        m943(.A(mai_mai_n236_), .B(mai_mai_n208_), .C(i_0_), .D(i_12_), .Y(mai_mai_n966_));
  AOI220     m944(.A0(mai_mai_n966_), .A1(mai_mai_n965_), .B0(mai_mai_n761_), .B1(mai_mai_n178_), .Y(mai_mai_n967_));
  NA2        m945(.A(mai_mai_n876_), .B(mai_mai_n437_), .Y(mai_mai_n968_));
  NA2        m946(.A(mai_mai_n65_), .B(mai_mai_n105_), .Y(mai_mai_n969_));
  OAI220     m947(.A0(mai_mai_n969_), .A1(mai_mai_n964_), .B0(mai_mai_n968_), .B1(mai_mai_n642_), .Y(mai_mai_n970_));
  NA2        m948(.A(mai_mai_n970_), .B(mai_mai_n866_), .Y(mai_mai_n971_));
  NA3        m949(.A(mai_mai_n971_), .B(mai_mai_n967_), .C(mai_mai_n963_), .Y(mai_mai_n972_));
  NO4        m950(.A(mai_mai_n972_), .B(mai_mai_n957_), .C(mai_mai_n940_), .D(mai_mai_n926_), .Y(mai_mai_n973_));
  INV        m951(.A(mai_mai_n578_), .Y(mai_mai_n974_));
  NA2        m952(.A(mai_mai_n974_), .B(mai_mai_n204_), .Y(mai_mai_n975_));
  OAI210     m953(.A0(mai_mai_n582_), .A1(mai_mai_n580_), .B0(mai_mai_n302_), .Y(mai_mai_n976_));
  INV        m954(.A(mai_mai_n976_), .Y(mai_mai_n977_));
  NO4        m955(.A(mai_mai_n229_), .B(mai_mai_n150_), .C(mai_mai_n645_), .D(mai_mai_n37_), .Y(mai_mai_n978_));
  AOI210     m956(.A0(mai_mai_n977_), .A1(mai_mai_n49_), .B0(mai_mai_n978_), .Y(mai_mai_n979_));
  AOI210     m957(.A0(mai_mai_n979_), .A1(mai_mai_n975_), .B0(mai_mai_n74_), .Y(mai_mai_n980_));
  NO2        m958(.A(mai_mai_n533_), .B(mai_mai_n361_), .Y(mai_mai_n981_));
  NO2        m959(.A(mai_mai_n981_), .B(mai_mai_n723_), .Y(mai_mai_n982_));
  AOI210     m960(.A0(mai_mai_n946_), .A1(mai_mai_n862_), .B0(mai_mai_n877_), .Y(mai_mai_n983_));
  NO2        m961(.A(mai_mai_n983_), .B(mai_mai_n645_), .Y(mai_mai_n984_));
  NA2        m962(.A(mai_mai_n260_), .B(mai_mai_n58_), .Y(mai_mai_n985_));
  AOI220     m963(.A0(mai_mai_n985_), .A1(mai_mai_n77_), .B0(mai_mai_n329_), .B1(mai_mai_n252_), .Y(mai_mai_n986_));
  NO2        m964(.A(mai_mai_n986_), .B(mai_mai_n233_), .Y(mai_mai_n987_));
  NA3        m965(.A(mai_mai_n100_), .B(mai_mai_n294_), .C(mai_mai_n31_), .Y(mai_mai_n988_));
  INV        m966(.A(mai_mai_n988_), .Y(mai_mai_n989_));
  NO3        m967(.A(mai_mai_n989_), .B(mai_mai_n987_), .C(mai_mai_n984_), .Y(mai_mai_n990_));
  NA2        m968(.A(mai_mai_n268_), .B(mai_mai_n90_), .Y(mai_mai_n991_));
  NA3        m969(.A(mai_mai_n727_), .B(mai_mai_n281_), .C(mai_mai_n81_), .Y(mai_mai_n992_));
  AOI210     m970(.A0(mai_mai_n992_), .A1(mai_mai_n991_), .B0(i_11_), .Y(mai_mai_n993_));
  NO3        m971(.A(mai_mai_n60_), .B(mai_mai_n59_), .C(i_4_), .Y(mai_mai_n994_));
  OAI210     m972(.A0(mai_mai_n881_), .A1(mai_mai_n294_), .B0(mai_mai_n994_), .Y(mai_mai_n995_));
  NO2        m973(.A(mai_mai_n995_), .B(mai_mai_n694_), .Y(mai_mai_n996_));
  NO4        m974(.A(mai_mai_n901_), .B(mai_mai_n442_), .C(mai_mai_n249_), .D(mai_mai_n248_), .Y(mai_mai_n997_));
  NO2        m975(.A(mai_mai_n997_), .B(mai_mai_n530_), .Y(mai_mai_n998_));
  INV        m976(.A(mai_mai_n347_), .Y(mai_mai_n999_));
  AOI210     m977(.A0(mai_mai_n999_), .A1(mai_mai_n998_), .B0(mai_mai_n41_), .Y(mai_mai_n1000_));
  NO3        m978(.A(mai_mai_n1000_), .B(mai_mai_n996_), .C(mai_mai_n993_), .Y(mai_mai_n1001_));
  OAI210     m979(.A0(mai_mai_n990_), .A1(i_4_), .B0(mai_mai_n1001_), .Y(mai_mai_n1002_));
  NO3        m980(.A(mai_mai_n1002_), .B(mai_mai_n982_), .C(mai_mai_n980_), .Y(mai_mai_n1003_));
  NA4        m981(.A(mai_mai_n1003_), .B(mai_mai_n973_), .C(mai_mai_n908_), .D(mai_mai_n833_), .Y(mai4));
  INV        m982(.A(mai_mai_n449_), .Y(mai_mai_n1007_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n51_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  NO2        u0062(.A(men_men_n83_), .B(men_men_n63_), .Y(men_men_n85_));
  INV        u0063(.A(i_6_), .Y(men_men_n86_));
  NO2        u0064(.A(i_2_), .B(i_7_), .Y(men_men_n87_));
  INV        u0065(.A(men_men_n87_), .Y(men_men_n88_));
  OAI210     u0066(.A0(men_men_n85_), .A1(men_men_n82_), .B0(men_men_n88_), .Y(men_men_n89_));
  NAi21      u0067(.An(i_6_), .B(i_10_), .Y(men_men_n90_));
  NA2        u0068(.A(i_6_), .B(i_9_), .Y(men_men_n91_));
  AOI210     u0069(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n63_), .Y(men_men_n92_));
  NA2        u0070(.A(i_2_), .B(i_6_), .Y(men_men_n93_));
  INV        u0071(.A(men_men_n92_), .Y(men_men_n94_));
  AOI210     u0072(.A0(men_men_n94_), .A1(men_men_n89_), .B0(men_men_n80_), .Y(men_men_n95_));
  AN3        u0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n96_));
  NAi21      u0074(.An(i_6_), .B(i_11_), .Y(men_men_n97_));
  NO2        u0075(.A(i_5_), .B(i_8_), .Y(men_men_n98_));
  NOi21      u0076(.An(men_men_n98_), .B(men_men_n97_), .Y(men_men_n99_));
  AOI220     u0077(.A0(men_men_n99_), .A1(men_men_n62_), .B0(men_men_n96_), .B1(men_men_n32_), .Y(men_men_n100_));
  INV        u0078(.A(i_7_), .Y(men_men_n101_));
  NA2        u0079(.A(men_men_n47_), .B(men_men_n101_), .Y(men_men_n102_));
  NO2        u0080(.A(i_0_), .B(i_5_), .Y(men_men_n103_));
  NO2        u0081(.A(men_men_n103_), .B(men_men_n86_), .Y(men_men_n104_));
  NA2        u0082(.A(i_12_), .B(i_3_), .Y(men_men_n105_));
  INV        u0083(.A(men_men_n105_), .Y(men_men_n106_));
  NA3        u0084(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n102_), .Y(men_men_n107_));
  NAi21      u0085(.An(i_7_), .B(i_11_), .Y(men_men_n108_));
  NO3        u0086(.A(men_men_n108_), .B(men_men_n90_), .C(men_men_n54_), .Y(men_men_n109_));
  AN2        u0087(.A(i_2_), .B(i_10_), .Y(men_men_n110_));
  NO2        u0088(.A(men_men_n110_), .B(i_7_), .Y(men_men_n111_));
  OR2        u0089(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n112_));
  NO2        u0090(.A(i_8_), .B(men_men_n101_), .Y(men_men_n113_));
  NO3        u0091(.A(men_men_n113_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n114_));
  NA2        u0092(.A(i_12_), .B(i_7_), .Y(men_men_n115_));
  NO2        u0093(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n116_));
  NA2        u0094(.A(i_11_), .B(i_12_), .Y(men_men_n117_));
  INV        u0095(.A(men_men_n117_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n118_), .B(men_men_n114_), .Y(men_men_n119_));
  NAi41      u0097(.An(men_men_n109_), .B(men_men_n119_), .C(men_men_n107_), .D(men_men_n100_), .Y(men_men_n120_));
  NOi21      u0098(.An(i_1_), .B(i_5_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n121_), .B(i_11_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n123_));
  NA2        u0101(.A(i_7_), .B(men_men_n25_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NO2        u0103(.A(men_men_n125_), .B(men_men_n47_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n127_));
  NAi21      u0105(.An(i_3_), .B(i_8_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(men_men_n62_), .Y(men_men_n129_));
  NOi31      u0107(.An(men_men_n129_), .B(men_men_n127_), .C(men_men_n126_), .Y(men_men_n130_));
  NO2        u0108(.A(i_1_), .B(men_men_n86_), .Y(men_men_n131_));
  NO2        u0109(.A(i_6_), .B(i_5_), .Y(men_men_n132_));
  NA2        u0110(.A(men_men_n132_), .B(i_3_), .Y(men_men_n133_));
  AO210      u0111(.A0(men_men_n133_), .A1(men_men_n48_), .B0(men_men_n131_), .Y(men_men_n134_));
  OAI220     u0112(.A0(men_men_n134_), .A1(men_men_n108_), .B0(men_men_n130_), .B1(men_men_n122_), .Y(men_men_n135_));
  NO3        u0113(.A(men_men_n135_), .B(men_men_n120_), .C(men_men_n95_), .Y(men_men_n136_));
  NA3        u0114(.A(men_men_n136_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0115(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n138_));
  NA2        u0116(.A(i_6_), .B(men_men_n25_), .Y(men_men_n139_));
  NA2        u0117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NA4        u0118(.A(men_men_n140_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0119(.A(i_8_), .B(i_7_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(i_6_), .Y(men_men_n143_));
  NO2        u0121(.A(i_12_), .B(i_13_), .Y(men_men_n144_));
  NAi21      u0122(.An(i_5_), .B(i_11_), .Y(men_men_n145_));
  NOi21      u0123(.An(men_men_n144_), .B(men_men_n145_), .Y(men_men_n146_));
  NO2        u0124(.A(i_0_), .B(i_1_), .Y(men_men_n147_));
  NA2        u0125(.A(i_2_), .B(i_3_), .Y(men_men_n148_));
  NO2        u0126(.A(men_men_n148_), .B(i_4_), .Y(men_men_n149_));
  NA3        u0127(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n150_));
  AN2        u0128(.A(men_men_n144_), .B(men_men_n83_), .Y(men_men_n151_));
  NO2        u0129(.A(men_men_n151_), .B(men_men_n27_), .Y(men_men_n152_));
  NA2        u0130(.A(i_1_), .B(i_5_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n73_), .B(men_men_n47_), .Y(men_men_n154_));
  NA2        u0132(.A(men_men_n154_), .B(men_men_n36_), .Y(men_men_n155_));
  NO3        u0133(.A(men_men_n155_), .B(men_men_n153_), .C(men_men_n152_), .Y(men_men_n156_));
  OR2        u0134(.A(i_0_), .B(i_1_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n158_));
  NAi32      u0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n159_));
  NAi21      u0137(.An(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  NOi21      u0138(.An(i_4_), .B(i_10_), .Y(men_men_n161_));
  NA2        u0139(.A(men_men_n161_), .B(men_men_n40_), .Y(men_men_n162_));
  NO2        u0140(.A(i_3_), .B(i_5_), .Y(men_men_n163_));
  NO3        u0141(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n164_));
  NA2        u0142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OAI210     u0143(.A0(men_men_n165_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n166_));
  NO2        u0144(.A(men_men_n166_), .B(men_men_n156_), .Y(men_men_n167_));
  AOI210     u0145(.A0(men_men_n167_), .A1(men_men_n150_), .B0(men_men_n143_), .Y(men_men_n168_));
  NA3        u0146(.A(men_men_n73_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n169_));
  NA2        u0147(.A(i_3_), .B(men_men_n49_), .Y(men_men_n170_));
  NOi21      u0148(.An(i_4_), .B(i_9_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_11_), .B(i_13_), .Y(men_men_n172_));
  NA2        u0150(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  OR2        u0151(.A(men_men_n173_), .B(men_men_n170_), .Y(men_men_n174_));
  NO2        u0152(.A(i_4_), .B(i_5_), .Y(men_men_n175_));
  NAi21      u0153(.An(i_12_), .B(i_11_), .Y(men_men_n176_));
  NO2        u0154(.A(men_men_n176_), .B(i_13_), .Y(men_men_n177_));
  NA3        u0155(.A(men_men_n177_), .B(men_men_n175_), .C(men_men_n83_), .Y(men_men_n178_));
  AOI210     u0156(.A0(men_men_n178_), .A1(men_men_n174_), .B0(men_men_n169_), .Y(men_men_n179_));
  NO2        u0157(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n180_));
  NA2        u0158(.A(men_men_n180_), .B(men_men_n47_), .Y(men_men_n181_));
  NAi31      u0159(.An(i_4_), .B(men_men_n151_), .C(i_11_), .Y(men_men_n182_));
  NA2        u0160(.A(i_3_), .B(i_5_), .Y(men_men_n183_));
  OR2        u0161(.A(men_men_n183_), .B(men_men_n173_), .Y(men_men_n184_));
  AOI210     u0162(.A0(men_men_n184_), .A1(men_men_n182_), .B0(men_men_n181_), .Y(men_men_n185_));
  NO2        u0163(.A(men_men_n73_), .B(i_5_), .Y(men_men_n186_));
  NO2        u0164(.A(i_13_), .B(i_10_), .Y(men_men_n187_));
  NA3        u0165(.A(men_men_n187_), .B(men_men_n186_), .C(men_men_n45_), .Y(men_men_n188_));
  NO2        u0166(.A(i_2_), .B(i_1_), .Y(men_men_n189_));
  NA2        u0167(.A(men_men_n189_), .B(i_3_), .Y(men_men_n190_));
  NAi21      u0168(.An(i_4_), .B(i_12_), .Y(men_men_n191_));
  NO4        u0169(.A(men_men_n191_), .B(men_men_n190_), .C(men_men_n188_), .D(men_men_n25_), .Y(men_men_n192_));
  NO3        u0170(.A(men_men_n192_), .B(men_men_n185_), .C(men_men_n179_), .Y(men_men_n193_));
  INV        u0171(.A(i_8_), .Y(men_men_n194_));
  NO2        u0172(.A(men_men_n194_), .B(i_7_), .Y(men_men_n195_));
  NA2        u0173(.A(men_men_n195_), .B(i_6_), .Y(men_men_n196_));
  NO3        u0174(.A(i_3_), .B(men_men_n86_), .C(men_men_n49_), .Y(men_men_n197_));
  NA2        u0175(.A(men_men_n197_), .B(men_men_n113_), .Y(men_men_n198_));
  NO3        u0176(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n199_));
  NA3        u0177(.A(men_men_n199_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n200_));
  NO3        u0178(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n201_));
  OAI210     u0179(.A0(men_men_n96_), .A1(i_12_), .B0(men_men_n201_), .Y(men_men_n202_));
  AOI210     u0180(.A0(men_men_n202_), .A1(men_men_n200_), .B0(men_men_n198_), .Y(men_men_n203_));
  NO2        u0181(.A(i_3_), .B(i_8_), .Y(men_men_n204_));
  NO3        u0182(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n205_));
  NA3        u0183(.A(men_men_n205_), .B(men_men_n204_), .C(men_men_n40_), .Y(men_men_n206_));
  NO2        u0184(.A(men_men_n103_), .B(men_men_n58_), .Y(men_men_n207_));
  INV        u0185(.A(men_men_n207_), .Y(men_men_n208_));
  NO2        u0186(.A(i_13_), .B(i_9_), .Y(men_men_n209_));
  NA3        u0187(.A(men_men_n209_), .B(i_6_), .C(men_men_n194_), .Y(men_men_n210_));
  NAi21      u0188(.An(i_12_), .B(i_3_), .Y(men_men_n211_));
  NO2        u0189(.A(men_men_n45_), .B(i_5_), .Y(men_men_n212_));
  NO3        u0190(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n213_));
  NA3        u0191(.A(men_men_n213_), .B(men_men_n212_), .C(i_10_), .Y(men_men_n214_));
  OAI220     u0192(.A0(men_men_n214_), .A1(men_men_n210_), .B0(men_men_n208_), .B1(men_men_n206_), .Y(men_men_n215_));
  AOI210     u0193(.A0(men_men_n215_), .A1(i_7_), .B0(men_men_n203_), .Y(men_men_n216_));
  OAI220     u0194(.A0(men_men_n216_), .A1(i_4_), .B0(men_men_n196_), .B1(men_men_n193_), .Y(men_men_n217_));
  NAi21      u0195(.An(i_12_), .B(i_7_), .Y(men_men_n218_));
  NA3        u0196(.A(i_13_), .B(men_men_n194_), .C(i_10_), .Y(men_men_n219_));
  NO2        u0197(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n220_));
  NA2        u0198(.A(i_0_), .B(i_5_), .Y(men_men_n221_));
  NA2        u0199(.A(men_men_n221_), .B(men_men_n104_), .Y(men_men_n222_));
  OAI220     u0200(.A0(men_men_n222_), .A1(men_men_n190_), .B0(men_men_n181_), .B1(men_men_n133_), .Y(men_men_n223_));
  NAi31      u0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n224_));
  NO2        u0202(.A(men_men_n36_), .B(i_13_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n226_));
  NO2        u0204(.A(men_men_n47_), .B(men_men_n63_), .Y(men_men_n227_));
  NA3        u0205(.A(men_men_n227_), .B(men_men_n226_), .C(men_men_n225_), .Y(men_men_n228_));
  INV        u0206(.A(i_13_), .Y(men_men_n229_));
  NO2        u0207(.A(i_12_), .B(men_men_n229_), .Y(men_men_n230_));
  NA3        u0208(.A(men_men_n230_), .B(men_men_n199_), .C(men_men_n197_), .Y(men_men_n231_));
  OAI210     u0209(.A0(men_men_n228_), .A1(men_men_n224_), .B0(men_men_n231_), .Y(men_men_n232_));
  AOI220     u0210(.A0(men_men_n232_), .A1(men_men_n142_), .B0(men_men_n223_), .B1(men_men_n220_), .Y(men_men_n233_));
  NO2        u0211(.A(i_12_), .B(men_men_n37_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n183_), .B(i_4_), .Y(men_men_n235_));
  NA2        u0213(.A(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  OR2        u0214(.A(i_8_), .B(i_7_), .Y(men_men_n237_));
  NO2        u0215(.A(men_men_n237_), .B(men_men_n86_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n54_), .B(i_1_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  INV        u0218(.A(i_12_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n45_), .B(men_men_n241_), .Y(men_men_n242_));
  NO3        u0220(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n243_));
  NA2        u0221(.A(i_2_), .B(i_1_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n240_), .B(men_men_n236_), .Y(men_men_n245_));
  NO3        u0223(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n246_));
  NAi21      u0224(.An(i_4_), .B(i_3_), .Y(men_men_n247_));
  NO2        u0225(.A(i_0_), .B(i_6_), .Y(men_men_n248_));
  NOi41      u0226(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n249_));
  NA2        u0227(.A(men_men_n249_), .B(men_men_n248_), .Y(men_men_n250_));
  NO2        u0228(.A(men_men_n244_), .B(men_men_n183_), .Y(men_men_n251_));
  NAi21      u0229(.An(men_men_n250_), .B(men_men_n251_), .Y(men_men_n252_));
  INV        u0230(.A(men_men_n252_), .Y(men_men_n253_));
  AOI210     u0231(.A0(men_men_n253_), .A1(men_men_n40_), .B0(men_men_n245_), .Y(men_men_n254_));
  NO2        u0232(.A(i_11_), .B(men_men_n229_), .Y(men_men_n255_));
  NOi21      u0233(.An(i_1_), .B(i_6_), .Y(men_men_n256_));
  NAi21      u0234(.An(i_3_), .B(i_7_), .Y(men_men_n257_));
  NA2        u0235(.A(men_men_n241_), .B(i_9_), .Y(men_men_n258_));
  OR4        u0236(.A(men_men_n258_), .B(men_men_n257_), .C(men_men_n256_), .D(men_men_n186_), .Y(men_men_n259_));
  NO2        u0237(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n260_));
  NO2        u0238(.A(i_12_), .B(i_3_), .Y(men_men_n261_));
  NA2        u0239(.A(men_men_n73_), .B(i_5_), .Y(men_men_n262_));
  NA2        u0240(.A(i_3_), .B(i_9_), .Y(men_men_n263_));
  NAi21      u0241(.An(i_7_), .B(i_10_), .Y(men_men_n264_));
  NO2        u0242(.A(men_men_n264_), .B(men_men_n263_), .Y(men_men_n265_));
  NA3        u0243(.A(men_men_n265_), .B(men_men_n262_), .C(men_men_n64_), .Y(men_men_n266_));
  NA2        u0244(.A(men_men_n266_), .B(men_men_n259_), .Y(men_men_n267_));
  NA3        u0245(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n268_));
  INV        u0246(.A(men_men_n143_), .Y(men_men_n269_));
  NA2        u0247(.A(men_men_n241_), .B(i_13_), .Y(men_men_n270_));
  NO2        u0248(.A(men_men_n270_), .B(men_men_n75_), .Y(men_men_n271_));
  AOI220     u0249(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n267_), .B1(men_men_n255_), .Y(men_men_n272_));
  NO2        u0250(.A(men_men_n237_), .B(men_men_n37_), .Y(men_men_n273_));
  NA2        u0251(.A(i_12_), .B(i_6_), .Y(men_men_n274_));
  OR2        u0252(.A(i_13_), .B(i_9_), .Y(men_men_n275_));
  NO2        u0253(.A(men_men_n247_), .B(i_2_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n255_), .B(i_9_), .Y(men_men_n277_));
  NA2        u0255(.A(men_men_n154_), .B(men_men_n63_), .Y(men_men_n278_));
  NO3        u0256(.A(i_11_), .B(men_men_n229_), .C(men_men_n25_), .Y(men_men_n279_));
  NO2        u0257(.A(men_men_n257_), .B(i_8_), .Y(men_men_n280_));
  NO2        u0258(.A(i_6_), .B(men_men_n49_), .Y(men_men_n281_));
  NA3        u0259(.A(men_men_n281_), .B(men_men_n280_), .C(men_men_n279_), .Y(men_men_n282_));
  NO3        u0260(.A(men_men_n26_), .B(men_men_n86_), .C(i_5_), .Y(men_men_n283_));
  NA3        u0261(.A(men_men_n283_), .B(men_men_n273_), .C(men_men_n230_), .Y(men_men_n284_));
  AOI210     u0262(.A0(men_men_n284_), .A1(men_men_n282_), .B0(men_men_n278_), .Y(men_men_n285_));
  INV        u0263(.A(men_men_n285_), .Y(men_men_n286_));
  NA4        u0264(.A(men_men_n286_), .B(men_men_n272_), .C(men_men_n254_), .D(men_men_n233_), .Y(men_men_n287_));
  NO3        u0265(.A(i_12_), .B(men_men_n229_), .C(men_men_n37_), .Y(men_men_n288_));
  INV        u0266(.A(men_men_n288_), .Y(men_men_n289_));
  NA2        u0267(.A(i_8_), .B(men_men_n101_), .Y(men_men_n290_));
  NOi21      u0268(.An(men_men_n163_), .B(men_men_n86_), .Y(men_men_n291_));
  NO3        u0269(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n292_));
  AOI220     u0270(.A0(men_men_n292_), .A1(men_men_n197_), .B0(men_men_n291_), .B1(men_men_n239_), .Y(men_men_n293_));
  NO2        u0271(.A(men_men_n293_), .B(men_men_n290_), .Y(men_men_n294_));
  NO3        u0272(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n244_), .B(i_0_), .Y(men_men_n296_));
  AOI220     u0274(.A0(men_men_n296_), .A1(men_men_n195_), .B0(men_men_n295_), .B1(men_men_n142_), .Y(men_men_n297_));
  NA2        u0275(.A(men_men_n281_), .B(men_men_n26_), .Y(men_men_n298_));
  NO2        u0276(.A(men_men_n298_), .B(men_men_n297_), .Y(men_men_n299_));
  NA2        u0277(.A(i_0_), .B(i_1_), .Y(men_men_n300_));
  NO2        u0278(.A(men_men_n300_), .B(i_2_), .Y(men_men_n301_));
  NO2        u0279(.A(men_men_n59_), .B(i_6_), .Y(men_men_n302_));
  NA3        u0280(.A(men_men_n302_), .B(men_men_n301_), .C(men_men_n163_), .Y(men_men_n303_));
  OAI210     u0281(.A0(men_men_n165_), .A1(men_men_n143_), .B0(men_men_n303_), .Y(men_men_n304_));
  NO3        u0282(.A(men_men_n304_), .B(men_men_n299_), .C(men_men_n294_), .Y(men_men_n305_));
  NO2        u0283(.A(i_3_), .B(i_10_), .Y(men_men_n306_));
  NA3        u0284(.A(men_men_n306_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n307_));
  NO2        u0285(.A(i_2_), .B(men_men_n101_), .Y(men_men_n308_));
  NA2        u0286(.A(i_1_), .B(men_men_n36_), .Y(men_men_n309_));
  NO2        u0287(.A(men_men_n309_), .B(i_8_), .Y(men_men_n310_));
  NOi21      u0288(.An(men_men_n221_), .B(men_men_n103_), .Y(men_men_n311_));
  NA3        u0289(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n308_), .Y(men_men_n312_));
  AN2        u0290(.A(i_3_), .B(i_10_), .Y(men_men_n313_));
  NA4        u0291(.A(men_men_n313_), .B(men_men_n199_), .C(men_men_n177_), .D(men_men_n175_), .Y(men_men_n314_));
  NO2        u0292(.A(i_5_), .B(men_men_n37_), .Y(men_men_n315_));
  NO2        u0293(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n316_));
  OR2        u0294(.A(men_men_n312_), .B(men_men_n307_), .Y(men_men_n317_));
  OAI220     u0295(.A0(men_men_n317_), .A1(i_6_), .B0(men_men_n305_), .B1(men_men_n289_), .Y(men_men_n318_));
  NO4        u0296(.A(men_men_n318_), .B(men_men_n287_), .C(men_men_n217_), .D(men_men_n168_), .Y(men_men_n319_));
  NO3        u0297(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n320_));
  NO2        u0298(.A(men_men_n59_), .B(men_men_n86_), .Y(men_men_n321_));
  NA2        u0299(.A(men_men_n296_), .B(men_men_n321_), .Y(men_men_n322_));
  NO3        u0300(.A(i_6_), .B(men_men_n194_), .C(i_7_), .Y(men_men_n323_));
  NA2        u0301(.A(men_men_n323_), .B(men_men_n199_), .Y(men_men_n324_));
  AOI210     u0302(.A0(men_men_n324_), .A1(men_men_n322_), .B0(men_men_n170_), .Y(men_men_n325_));
  NO2        u0303(.A(i_2_), .B(i_3_), .Y(men_men_n326_));
  OR2        u0304(.A(i_0_), .B(i_5_), .Y(men_men_n327_));
  NA2        u0305(.A(men_men_n221_), .B(men_men_n327_), .Y(men_men_n328_));
  NA4        u0306(.A(men_men_n328_), .B(men_men_n238_), .C(men_men_n326_), .D(i_1_), .Y(men_men_n329_));
  NA3        u0307(.A(men_men_n296_), .B(men_men_n291_), .C(men_men_n113_), .Y(men_men_n330_));
  NAi21      u0308(.An(i_8_), .B(i_7_), .Y(men_men_n331_));
  NO2        u0309(.A(men_men_n331_), .B(i_6_), .Y(men_men_n332_));
  NO2        u0310(.A(men_men_n157_), .B(men_men_n47_), .Y(men_men_n333_));
  NA3        u0311(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n163_), .Y(men_men_n334_));
  NA3        u0312(.A(men_men_n334_), .B(men_men_n330_), .C(men_men_n329_), .Y(men_men_n335_));
  OAI210     u0313(.A0(men_men_n335_), .A1(men_men_n325_), .B0(i_4_), .Y(men_men_n336_));
  NO2        u0314(.A(i_12_), .B(i_10_), .Y(men_men_n337_));
  NOi21      u0315(.An(i_5_), .B(i_0_), .Y(men_men_n338_));
  NO3        u0316(.A(men_men_n309_), .B(men_men_n338_), .C(men_men_n128_), .Y(men_men_n339_));
  NA2        u0317(.A(men_men_n339_), .B(men_men_n337_), .Y(men_men_n340_));
  NO2        u0318(.A(i_6_), .B(i_8_), .Y(men_men_n341_));
  NOi21      u0319(.An(i_0_), .B(i_2_), .Y(men_men_n342_));
  AN2        u0320(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  NO2        u0321(.A(i_1_), .B(i_7_), .Y(men_men_n344_));
  AO220      u0322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n332_), .B1(men_men_n239_), .Y(men_men_n345_));
  NA2        u0323(.A(men_men_n345_), .B(men_men_n42_), .Y(men_men_n346_));
  NA3        u0324(.A(men_men_n346_), .B(men_men_n340_), .C(men_men_n336_), .Y(men_men_n347_));
  NO3        u0325(.A(men_men_n237_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n348_));
  NO3        u0326(.A(men_men_n331_), .B(i_2_), .C(i_1_), .Y(men_men_n349_));
  OAI210     u0327(.A0(men_men_n349_), .A1(men_men_n348_), .B0(i_6_), .Y(men_men_n350_));
  NA3        u0328(.A(men_men_n256_), .B(men_men_n308_), .C(men_men_n194_), .Y(men_men_n351_));
  AOI210     u0329(.A0(men_men_n351_), .A1(men_men_n350_), .B0(men_men_n328_), .Y(men_men_n352_));
  NOi21      u0330(.An(men_men_n153_), .B(men_men_n104_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n353_), .B(men_men_n124_), .Y(men_men_n354_));
  OAI210     u0332(.A0(men_men_n354_), .A1(men_men_n352_), .B0(i_3_), .Y(men_men_n355_));
  INV        u0333(.A(men_men_n84_), .Y(men_men_n356_));
  NO2        u0334(.A(men_men_n300_), .B(men_men_n81_), .Y(men_men_n357_));
  NA2        u0335(.A(men_men_n357_), .B(men_men_n132_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n93_), .B(men_men_n194_), .Y(men_men_n359_));
  NA3        u0337(.A(men_men_n311_), .B(men_men_n359_), .C(men_men_n63_), .Y(men_men_n360_));
  AOI210     u0338(.A0(men_men_n360_), .A1(men_men_n358_), .B0(men_men_n356_), .Y(men_men_n361_));
  NO2        u0339(.A(men_men_n194_), .B(i_9_), .Y(men_men_n362_));
  NA2        u0340(.A(men_men_n362_), .B(men_men_n207_), .Y(men_men_n363_));
  NO2        u0341(.A(men_men_n363_), .B(men_men_n47_), .Y(men_men_n364_));
  NO3        u0342(.A(men_men_n364_), .B(men_men_n361_), .C(men_men_n299_), .Y(men_men_n365_));
  AOI210     u0343(.A0(men_men_n365_), .A1(men_men_n355_), .B0(men_men_n162_), .Y(men_men_n366_));
  AOI210     u0344(.A0(men_men_n347_), .A1(men_men_n320_), .B0(men_men_n366_), .Y(men_men_n367_));
  NOi32      u0345(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n368_));
  INV        u0346(.A(men_men_n368_), .Y(men_men_n369_));
  NAi21      u0347(.An(i_0_), .B(i_6_), .Y(men_men_n370_));
  NAi21      u0348(.An(i_1_), .B(i_5_), .Y(men_men_n371_));
  NA2        u0349(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  NA2        u0350(.A(men_men_n372_), .B(men_men_n25_), .Y(men_men_n373_));
  OAI210     u0351(.A0(men_men_n373_), .A1(men_men_n159_), .B0(men_men_n250_), .Y(men_men_n374_));
  NAi41      u0352(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n375_));
  OAI220     u0353(.A0(men_men_n375_), .A1(men_men_n371_), .B0(men_men_n224_), .B1(men_men_n159_), .Y(men_men_n376_));
  AOI210     u0354(.A0(men_men_n375_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n377_));
  NOi32      u0355(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n378_));
  NAi21      u0356(.An(i_6_), .B(i_1_), .Y(men_men_n379_));
  NA3        u0357(.A(men_men_n379_), .B(men_men_n378_), .C(men_men_n47_), .Y(men_men_n380_));
  NO2        u0358(.A(men_men_n380_), .B(i_0_), .Y(men_men_n381_));
  OR3        u0359(.A(men_men_n381_), .B(men_men_n377_), .C(men_men_n376_), .Y(men_men_n382_));
  NO2        u0360(.A(i_1_), .B(men_men_n101_), .Y(men_men_n383_));
  NAi21      u0361(.An(i_3_), .B(i_4_), .Y(men_men_n384_));
  NO2        u0362(.A(men_men_n384_), .B(i_9_), .Y(men_men_n385_));
  AN2        u0363(.A(i_6_), .B(i_7_), .Y(men_men_n386_));
  OAI210     u0364(.A0(men_men_n386_), .A1(men_men_n383_), .B0(men_men_n385_), .Y(men_men_n387_));
  NA2        u0365(.A(i_2_), .B(i_7_), .Y(men_men_n388_));
  NO2        u0366(.A(men_men_n384_), .B(i_10_), .Y(men_men_n389_));
  NA3        u0367(.A(men_men_n389_), .B(men_men_n388_), .C(men_men_n248_), .Y(men_men_n390_));
  AOI210     u0368(.A0(men_men_n390_), .A1(men_men_n387_), .B0(men_men_n186_), .Y(men_men_n391_));
  AOI210     u0369(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n392_));
  OAI210     u0370(.A0(men_men_n392_), .A1(men_men_n189_), .B0(men_men_n389_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n393_), .B(i_5_), .Y(men_men_n394_));
  NO4        u0372(.A(men_men_n394_), .B(men_men_n391_), .C(men_men_n382_), .D(men_men_n374_), .Y(men_men_n395_));
  NO2        u0373(.A(men_men_n395_), .B(men_men_n369_), .Y(men_men_n396_));
  NO2        u0374(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n397_));
  AN2        u0375(.A(i_12_), .B(i_5_), .Y(men_men_n398_));
  NA2        u0376(.A(i_3_), .B(men_men_n398_), .Y(men_men_n399_));
  NO2        u0377(.A(i_11_), .B(i_6_), .Y(men_men_n400_));
  NA3        u0378(.A(men_men_n400_), .B(men_men_n333_), .C(men_men_n229_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n401_), .B(men_men_n399_), .Y(men_men_n402_));
  NO2        u0380(.A(men_men_n247_), .B(i_5_), .Y(men_men_n403_));
  NO2        u0381(.A(i_5_), .B(i_10_), .Y(men_men_n404_));
  AOI220     u0382(.A0(men_men_n404_), .A1(men_men_n276_), .B0(men_men_n403_), .B1(men_men_n199_), .Y(men_men_n405_));
  NA2        u0383(.A(men_men_n144_), .B(men_men_n46_), .Y(men_men_n406_));
  NO2        u0384(.A(men_men_n406_), .B(men_men_n405_), .Y(men_men_n407_));
  OAI210     u0385(.A0(men_men_n407_), .A1(men_men_n402_), .B0(men_men_n397_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n150_), .B(men_men_n86_), .Y(men_men_n410_));
  OAI210     u0388(.A0(men_men_n410_), .A1(men_men_n402_), .B0(men_men_n409_), .Y(men_men_n411_));
  NO3        u0389(.A(men_men_n86_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n412_));
  NO2        u0390(.A(i_3_), .B(men_men_n101_), .Y(men_men_n413_));
  NA2        u0391(.A(men_men_n306_), .B(men_men_n91_), .Y(men_men_n414_));
  NO2        u0392(.A(i_11_), .B(i_12_), .Y(men_men_n415_));
  NA2        u0393(.A(men_men_n415_), .B(men_men_n36_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n414_), .B(men_men_n416_), .Y(men_men_n417_));
  NA2        u0395(.A(men_men_n404_), .B(men_men_n241_), .Y(men_men_n418_));
  NA3        u0396(.A(men_men_n113_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n419_), .B(men_men_n224_), .Y(men_men_n420_));
  NAi21      u0398(.An(i_13_), .B(i_0_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n421_), .B(men_men_n244_), .Y(men_men_n422_));
  OAI210     u0400(.A0(men_men_n420_), .A1(men_men_n417_), .B0(men_men_n422_), .Y(men_men_n423_));
  NA3        u0401(.A(men_men_n423_), .B(men_men_n411_), .C(men_men_n408_), .Y(men_men_n424_));
  NO3        u0402(.A(i_1_), .B(i_12_), .C(men_men_n86_), .Y(men_men_n425_));
  NO2        u0403(.A(i_0_), .B(i_11_), .Y(men_men_n426_));
  INV        u0404(.A(i_5_), .Y(men_men_n427_));
  AN2        u0405(.A(i_1_), .B(i_6_), .Y(men_men_n428_));
  NOi21      u0406(.An(i_2_), .B(i_12_), .Y(men_men_n429_));
  NA2        u0407(.A(men_men_n429_), .B(men_men_n428_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n430_), .B(men_men_n427_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n142_), .B(i_9_), .Y(men_men_n432_));
  NO2        u0410(.A(men_men_n432_), .B(i_4_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n431_), .B(men_men_n433_), .Y(men_men_n434_));
  NAi21      u0412(.An(i_9_), .B(i_4_), .Y(men_men_n435_));
  OR2        u0413(.A(i_13_), .B(i_10_), .Y(men_men_n436_));
  NO3        u0414(.A(men_men_n436_), .B(men_men_n117_), .C(men_men_n435_), .Y(men_men_n437_));
  NO2        u0415(.A(men_men_n173_), .B(men_men_n123_), .Y(men_men_n438_));
  OR2        u0416(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n439_));
  NO2        u0417(.A(men_men_n101_), .B(men_men_n25_), .Y(men_men_n440_));
  NA2        u0418(.A(men_men_n288_), .B(men_men_n440_), .Y(men_men_n441_));
  NA2        u0419(.A(men_men_n281_), .B(men_men_n213_), .Y(men_men_n442_));
  OAI220     u0420(.A0(men_men_n442_), .A1(men_men_n439_), .B0(men_men_n441_), .B1(men_men_n353_), .Y(men_men_n443_));
  INV        u0421(.A(men_men_n443_), .Y(men_men_n444_));
  AOI210     u0422(.A0(men_men_n444_), .A1(men_men_n434_), .B0(men_men_n26_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n330_), .B(men_men_n329_), .Y(men_men_n446_));
  AOI220     u0424(.A0(men_men_n302_), .A1(men_men_n292_), .B0(men_men_n296_), .B1(men_men_n321_), .Y(men_men_n447_));
  NO2        u0425(.A(men_men_n447_), .B(men_men_n170_), .Y(men_men_n448_));
  NO2        u0426(.A(men_men_n183_), .B(men_men_n86_), .Y(men_men_n449_));
  AOI220     u0427(.A0(men_men_n449_), .A1(men_men_n301_), .B0(men_men_n283_), .B1(men_men_n213_), .Y(men_men_n450_));
  NO2        u0428(.A(men_men_n450_), .B(men_men_n290_), .Y(men_men_n451_));
  NO3        u0429(.A(men_men_n451_), .B(men_men_n448_), .C(men_men_n446_), .Y(men_men_n452_));
  NA2        u0430(.A(men_men_n197_), .B(men_men_n96_), .Y(men_men_n453_));
  NA3        u0431(.A(men_men_n333_), .B(men_men_n163_), .C(men_men_n86_), .Y(men_men_n454_));
  AOI210     u0432(.A0(men_men_n454_), .A1(men_men_n453_), .B0(men_men_n331_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n194_), .B(i_10_), .Y(men_men_n456_));
  NA3        u0434(.A(men_men_n262_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n302_), .B(men_men_n239_), .Y(men_men_n458_));
  OAI220     u0436(.A0(men_men_n458_), .A1(men_men_n183_), .B0(men_men_n457_), .B1(men_men_n456_), .Y(men_men_n459_));
  NO2        u0437(.A(i_3_), .B(men_men_n49_), .Y(men_men_n460_));
  NA3        u0438(.A(men_men_n344_), .B(men_men_n343_), .C(men_men_n460_), .Y(men_men_n461_));
  NA2        u0439(.A(men_men_n323_), .B(men_men_n328_), .Y(men_men_n462_));
  OAI210     u0440(.A0(men_men_n462_), .A1(men_men_n190_), .B0(men_men_n461_), .Y(men_men_n463_));
  NO3        u0441(.A(men_men_n463_), .B(men_men_n459_), .C(men_men_n455_), .Y(men_men_n464_));
  AOI210     u0442(.A0(men_men_n464_), .A1(men_men_n452_), .B0(men_men_n277_), .Y(men_men_n465_));
  NO4        u0443(.A(men_men_n465_), .B(men_men_n445_), .C(men_men_n424_), .D(men_men_n396_), .Y(men_men_n466_));
  NO2        u0444(.A(men_men_n63_), .B(i_4_), .Y(men_men_n467_));
  NO2        u0445(.A(men_men_n73_), .B(i_13_), .Y(men_men_n468_));
  NO2        u0446(.A(i_10_), .B(i_9_), .Y(men_men_n469_));
  NAi21      u0447(.An(i_12_), .B(i_8_), .Y(men_men_n470_));
  NO2        u0448(.A(men_men_n470_), .B(i_3_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n47_), .B(i_4_), .Y(men_men_n472_));
  NA2        u0450(.A(men_men_n472_), .B(men_men_n104_), .Y(men_men_n473_));
  NO2        u0451(.A(men_men_n473_), .B(men_men_n206_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n316_), .B(i_0_), .Y(men_men_n475_));
  NO3        u0453(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n274_), .B(men_men_n97_), .Y(men_men_n477_));
  NA2        u0455(.A(men_men_n477_), .B(men_men_n476_), .Y(men_men_n478_));
  NA2        u0456(.A(i_8_), .B(i_9_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n255_), .B(men_men_n315_), .Y(men_men_n480_));
  NO3        u0458(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n481_));
  INV        u0459(.A(men_men_n481_), .Y(men_men_n482_));
  NA3        u0460(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n483_));
  NA4        u0461(.A(men_men_n145_), .B(men_men_n116_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n484_));
  OAI220     u0462(.A0(men_men_n484_), .A1(men_men_n483_), .B0(men_men_n482_), .B1(men_men_n480_), .Y(men_men_n485_));
  NO2        u0463(.A(men_men_n485_), .B(men_men_n474_), .Y(men_men_n486_));
  INV        u0464(.A(men_men_n301_), .Y(men_men_n487_));
  OR2        u0465(.A(men_men_n487_), .B(men_men_n210_), .Y(men_men_n488_));
  OA210      u0466(.A0(men_men_n363_), .A1(men_men_n101_), .B0(men_men_n303_), .Y(men_men_n489_));
  OA220      u0467(.A0(men_men_n489_), .A1(men_men_n162_), .B0(men_men_n488_), .B1(men_men_n236_), .Y(men_men_n490_));
  NA2        u0468(.A(men_men_n96_), .B(i_13_), .Y(men_men_n491_));
  NA2        u0469(.A(men_men_n449_), .B(men_men_n397_), .Y(men_men_n492_));
  NO2        u0470(.A(i_2_), .B(i_13_), .Y(men_men_n493_));
  NA3        u0471(.A(men_men_n493_), .B(men_men_n161_), .C(men_men_n99_), .Y(men_men_n494_));
  OAI220     u0472(.A0(men_men_n494_), .A1(men_men_n241_), .B0(men_men_n492_), .B1(men_men_n491_), .Y(men_men_n495_));
  NO3        u0473(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n496_));
  NO2        u0474(.A(i_6_), .B(i_7_), .Y(men_men_n497_));
  NA2        u0475(.A(men_men_n497_), .B(men_men_n496_), .Y(men_men_n498_));
  NO2        u0476(.A(i_11_), .B(i_1_), .Y(men_men_n499_));
  NO2        u0477(.A(men_men_n73_), .B(i_3_), .Y(men_men_n500_));
  OR2        u0478(.A(i_11_), .B(i_8_), .Y(men_men_n501_));
  NOi21      u0479(.An(i_2_), .B(i_7_), .Y(men_men_n502_));
  NAi31      u0480(.An(men_men_n501_), .B(men_men_n502_), .C(men_men_n500_), .Y(men_men_n503_));
  NO2        u0481(.A(men_men_n436_), .B(i_6_), .Y(men_men_n504_));
  NA2        u0482(.A(men_men_n504_), .B(men_men_n467_), .Y(men_men_n505_));
  NO2        u0483(.A(men_men_n505_), .B(men_men_n503_), .Y(men_men_n506_));
  NO2        u0484(.A(i_3_), .B(men_men_n194_), .Y(men_men_n507_));
  NO2        u0485(.A(i_6_), .B(i_10_), .Y(men_men_n508_));
  NA4        u0486(.A(men_men_n508_), .B(men_men_n320_), .C(men_men_n507_), .D(men_men_n241_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n509_), .B(men_men_n155_), .Y(men_men_n510_));
  NA3        u0488(.A(men_men_n249_), .B(men_men_n172_), .C(men_men_n132_), .Y(men_men_n511_));
  NA2        u0489(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n512_));
  NO2        u0490(.A(men_men_n157_), .B(i_3_), .Y(men_men_n513_));
  NAi31      u0491(.An(men_men_n512_), .B(men_men_n513_), .C(men_men_n230_), .Y(men_men_n514_));
  NA3        u0492(.A(men_men_n409_), .B(men_men_n180_), .C(men_men_n149_), .Y(men_men_n515_));
  NA3        u0493(.A(men_men_n515_), .B(men_men_n514_), .C(men_men_n511_), .Y(men_men_n516_));
  NO4        u0494(.A(men_men_n516_), .B(men_men_n510_), .C(men_men_n506_), .D(men_men_n495_), .Y(men_men_n517_));
  NA2        u0495(.A(men_men_n476_), .B(men_men_n398_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n481_), .B(men_men_n404_), .Y(men_men_n519_));
  NO2        u0497(.A(men_men_n519_), .B(men_men_n228_), .Y(men_men_n520_));
  NAi21      u0498(.An(men_men_n219_), .B(men_men_n415_), .Y(men_men_n521_));
  NO2        u0499(.A(men_men_n26_), .B(i_5_), .Y(men_men_n522_));
  NO2        u0500(.A(i_0_), .B(men_men_n86_), .Y(men_men_n523_));
  NA3        u0501(.A(men_men_n523_), .B(men_men_n522_), .C(men_men_n142_), .Y(men_men_n524_));
  OR3        u0502(.A(men_men_n309_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n525_));
  NO2        u0503(.A(men_men_n525_), .B(men_men_n524_), .Y(men_men_n526_));
  NA2        u0504(.A(men_men_n27_), .B(i_10_), .Y(men_men_n527_));
  NO2        u0505(.A(men_men_n527_), .B(men_men_n491_), .Y(men_men_n528_));
  NA4        u0506(.A(men_men_n313_), .B(men_men_n227_), .C(men_men_n73_), .D(men_men_n241_), .Y(men_men_n529_));
  NO2        u0507(.A(men_men_n529_), .B(men_men_n498_), .Y(men_men_n530_));
  NO4        u0508(.A(men_men_n530_), .B(men_men_n528_), .C(men_men_n526_), .D(men_men_n520_), .Y(men_men_n531_));
  NA4        u0509(.A(men_men_n531_), .B(men_men_n517_), .C(men_men_n490_), .D(men_men_n486_), .Y(men_men_n532_));
  NA3        u0510(.A(men_men_n313_), .B(men_men_n177_), .C(men_men_n175_), .Y(men_men_n533_));
  OAI210     u0511(.A0(men_men_n307_), .A1(i_4_), .B0(men_men_n533_), .Y(men_men_n534_));
  AN2        u0512(.A(men_men_n292_), .B(men_men_n238_), .Y(men_men_n535_));
  NA2        u0513(.A(men_men_n535_), .B(men_men_n534_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n320_), .B(men_men_n164_), .Y(men_men_n537_));
  OAI210     u0515(.A0(men_men_n537_), .A1(men_men_n236_), .B0(men_men_n314_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n538_), .B(men_men_n332_), .Y(men_men_n539_));
  NA2        u0517(.A(men_men_n398_), .B(men_men_n229_), .Y(men_men_n540_));
  NA2        u0518(.A(men_men_n386_), .B(men_men_n378_), .Y(men_men_n541_));
  OR2        u0519(.A(men_men_n540_), .B(men_men_n541_), .Y(men_men_n542_));
  NO2        u0520(.A(men_men_n36_), .B(i_8_), .Y(men_men_n543_));
  AOI210     u0521(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n437_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n544_), .B(men_men_n542_), .Y(men_men_n545_));
  INV        u0523(.A(men_men_n545_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n262_), .B(men_men_n64_), .Y(men_men_n547_));
  OAI210     u0525(.A0(i_8_), .A1(men_men_n547_), .B0(men_men_n134_), .Y(men_men_n548_));
  AOI210     u0526(.A0(men_men_n195_), .A1(i_9_), .B0(men_men_n273_), .Y(men_men_n549_));
  NO2        u0527(.A(men_men_n549_), .B(men_men_n200_), .Y(men_men_n550_));
  NO2        u0528(.A(men_men_n183_), .B(men_men_n86_), .Y(men_men_n551_));
  AOI220     u0529(.A0(men_men_n551_), .A1(men_men_n550_), .B0(men_men_n548_), .B1(men_men_n438_), .Y(men_men_n552_));
  NA4        u0530(.A(men_men_n552_), .B(men_men_n546_), .C(men_men_n539_), .D(men_men_n536_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n403_), .B(men_men_n301_), .Y(men_men_n554_));
  OAI210     u0532(.A0(men_men_n399_), .A1(men_men_n169_), .B0(men_men_n554_), .Y(men_men_n555_));
  NO2        u0533(.A(i_12_), .B(men_men_n194_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n556_), .B(men_men_n229_), .Y(men_men_n557_));
  NA2        u0535(.A(men_men_n508_), .B(men_men_n27_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n558_), .B(men_men_n557_), .Y(men_men_n559_));
  NOi31      u0537(.An(men_men_n323_), .B(men_men_n436_), .C(men_men_n38_), .Y(men_men_n560_));
  OAI210     u0538(.A0(men_men_n560_), .A1(men_men_n559_), .B0(men_men_n555_), .Y(men_men_n561_));
  NO2        u0539(.A(i_8_), .B(i_7_), .Y(men_men_n562_));
  OAI210     u0540(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n563_), .B(men_men_n227_), .Y(men_men_n564_));
  AOI220     u0542(.A0(men_men_n333_), .A1(men_men_n40_), .B0(men_men_n239_), .B1(men_men_n209_), .Y(men_men_n565_));
  OAI220     u0543(.A0(men_men_n565_), .A1(men_men_n183_), .B0(men_men_n564_), .B1(men_men_n247_), .Y(men_men_n566_));
  NA2        u0544(.A(men_men_n45_), .B(i_10_), .Y(men_men_n567_));
  NO2        u0545(.A(men_men_n567_), .B(i_6_), .Y(men_men_n568_));
  NA3        u0546(.A(men_men_n568_), .B(men_men_n566_), .C(men_men_n562_), .Y(men_men_n569_));
  NA2        u0547(.A(men_men_n449_), .B(men_men_n333_), .Y(men_men_n570_));
  OAI220     u0548(.A0(men_men_n570_), .A1(men_men_n270_), .B0(men_men_n491_), .B1(men_men_n133_), .Y(men_men_n571_));
  NA2        u0549(.A(men_men_n571_), .B(men_men_n273_), .Y(men_men_n572_));
  NOi31      u0550(.An(men_men_n296_), .B(men_men_n307_), .C(i_4_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n157_), .B(i_5_), .Y(men_men_n574_));
  NA2        u0552(.A(men_men_n573_), .B(men_men_n481_), .Y(men_men_n575_));
  NA4        u0553(.A(men_men_n575_), .B(men_men_n572_), .C(men_men_n569_), .D(men_men_n561_), .Y(men_men_n576_));
  NA3        u0554(.A(men_men_n221_), .B(men_men_n71_), .C(men_men_n45_), .Y(men_men_n577_));
  NA2        u0555(.A(men_men_n288_), .B(men_men_n84_), .Y(men_men_n578_));
  AOI210     u0556(.A0(men_men_n577_), .A1(men_men_n358_), .B0(men_men_n578_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n302_), .B(men_men_n292_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n580_), .B(men_men_n174_), .Y(men_men_n581_));
  NA2        u0559(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n582_));
  NA2        u0560(.A(men_men_n469_), .B(men_men_n225_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n582_), .B(men_men_n583_), .Y(men_men_n584_));
  AOI210     u0562(.A0(men_men_n379_), .A1(men_men_n47_), .B0(men_men_n383_), .Y(men_men_n585_));
  NA2        u0563(.A(i_0_), .B(men_men_n49_), .Y(men_men_n586_));
  NA3        u0564(.A(men_men_n556_), .B(men_men_n279_), .C(men_men_n586_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n585_), .B(men_men_n587_), .Y(men_men_n588_));
  NO4        u0566(.A(men_men_n588_), .B(men_men_n584_), .C(men_men_n581_), .D(men_men_n579_), .Y(men_men_n589_));
  NO4        u0567(.A(men_men_n256_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n590_));
  NO3        u0568(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n591_));
  NO2        u0569(.A(men_men_n237_), .B(men_men_n36_), .Y(men_men_n592_));
  AN2        u0570(.A(men_men_n592_), .B(men_men_n591_), .Y(men_men_n593_));
  OA210      u0571(.A0(men_men_n593_), .A1(men_men_n590_), .B0(men_men_n368_), .Y(men_men_n594_));
  NO2        u0572(.A(men_men_n436_), .B(i_1_), .Y(men_men_n595_));
  NOi31      u0573(.An(men_men_n595_), .B(men_men_n477_), .C(men_men_n73_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n447_), .B(men_men_n178_), .Y(men_men_n597_));
  NO2        u0575(.A(men_men_n597_), .B(men_men_n594_), .Y(men_men_n598_));
  NOi21      u0576(.An(i_10_), .B(i_6_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n600_));
  NO2        u0578(.A(men_men_n115_), .B(men_men_n23_), .Y(men_men_n601_));
  NA2        u0579(.A(men_men_n323_), .B(men_men_n164_), .Y(men_men_n602_));
  AOI220     u0580(.A0(men_men_n602_), .A1(men_men_n458_), .B0(men_men_n184_), .B1(men_men_n182_), .Y(men_men_n603_));
  INV        u0581(.A(men_men_n603_), .Y(men_men_n604_));
  INV        u0582(.A(men_men_n326_), .Y(men_men_n605_));
  NO2        u0583(.A(i_12_), .B(men_men_n86_), .Y(men_men_n606_));
  NA3        u0584(.A(men_men_n606_), .B(men_men_n279_), .C(men_men_n586_), .Y(men_men_n607_));
  NA3        u0585(.A(men_men_n400_), .B(men_men_n288_), .C(men_men_n221_), .Y(men_men_n608_));
  AOI210     u0586(.A0(men_men_n608_), .A1(men_men_n607_), .B0(men_men_n605_), .Y(men_men_n609_));
  NO3        u0587(.A(i_4_), .B(men_men_n350_), .C(men_men_n307_), .Y(men_men_n610_));
  OR2        u0588(.A(i_2_), .B(i_5_), .Y(men_men_n611_));
  OR2        u0589(.A(men_men_n611_), .B(men_men_n428_), .Y(men_men_n612_));
  AOI210     u0590(.A0(men_men_n388_), .A1(men_men_n248_), .B0(men_men_n199_), .Y(men_men_n613_));
  AOI210     u0591(.A0(men_men_n613_), .A1(men_men_n612_), .B0(men_men_n521_), .Y(men_men_n614_));
  NO3        u0592(.A(men_men_n614_), .B(men_men_n610_), .C(men_men_n609_), .Y(men_men_n615_));
  NA4        u0593(.A(men_men_n615_), .B(men_men_n604_), .C(men_men_n598_), .D(men_men_n589_), .Y(men_men_n616_));
  NO4        u0594(.A(men_men_n616_), .B(men_men_n576_), .C(men_men_n553_), .D(men_men_n532_), .Y(men_men_n617_));
  NA4        u0595(.A(men_men_n617_), .B(men_men_n466_), .C(men_men_n367_), .D(men_men_n319_), .Y(men7));
  NO2        u0596(.A(men_men_n93_), .B(men_men_n55_), .Y(men_men_n619_));
  NA2        u0597(.A(men_men_n508_), .B(men_men_n84_), .Y(men_men_n620_));
  NA2        u0598(.A(i_11_), .B(men_men_n194_), .Y(men_men_n621_));
  NA2        u0599(.A(men_men_n144_), .B(men_men_n621_), .Y(men_men_n622_));
  NO2        u0600(.A(men_men_n622_), .B(men_men_n620_), .Y(men_men_n623_));
  NA3        u0601(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n624_));
  NO2        u0602(.A(men_men_n241_), .B(i_4_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n625_), .B(i_8_), .Y(men_men_n626_));
  NO2        u0604(.A(men_men_n105_), .B(men_men_n624_), .Y(men_men_n627_));
  NA2        u0605(.A(i_2_), .B(men_men_n86_), .Y(men_men_n628_));
  OAI210     u0606(.A0(men_men_n87_), .A1(men_men_n204_), .B0(men_men_n205_), .Y(men_men_n629_));
  NO2        u0607(.A(i_7_), .B(men_men_n37_), .Y(men_men_n630_));
  NA2        u0608(.A(i_4_), .B(i_8_), .Y(men_men_n631_));
  AOI210     u0609(.A0(men_men_n631_), .A1(men_men_n313_), .B0(men_men_n630_), .Y(men_men_n632_));
  OAI220     u0610(.A0(men_men_n632_), .A1(men_men_n628_), .B0(men_men_n629_), .B1(i_13_), .Y(men_men_n633_));
  NO4        u0611(.A(men_men_n633_), .B(men_men_n627_), .C(men_men_n623_), .D(men_men_n619_), .Y(men_men_n634_));
  AOI210     u0612(.A0(men_men_n128_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n635_));
  AOI210     u0613(.A0(men_men_n635_), .A1(men_men_n241_), .B0(men_men_n161_), .Y(men_men_n636_));
  OR2        u0614(.A(i_6_), .B(i_10_), .Y(men_men_n637_));
  NO2        u0615(.A(men_men_n637_), .B(men_men_n23_), .Y(men_men_n638_));
  OR3        u0616(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n639_));
  NO3        u0617(.A(men_men_n639_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n640_));
  INV        u0618(.A(men_men_n201_), .Y(men_men_n641_));
  NO2        u0619(.A(men_men_n640_), .B(men_men_n638_), .Y(men_men_n642_));
  OA220      u0620(.A0(men_men_n642_), .A1(men_men_n605_), .B0(men_men_n636_), .B1(men_men_n275_), .Y(men_men_n643_));
  AOI210     u0621(.A0(men_men_n643_), .A1(men_men_n634_), .B0(men_men_n63_), .Y(men_men_n644_));
  NOi21      u0622(.An(i_11_), .B(i_7_), .Y(men_men_n645_));
  AO210      u0623(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n646_), .B(men_men_n645_), .Y(men_men_n647_));
  NA2        u0625(.A(men_men_n647_), .B(men_men_n209_), .Y(men_men_n648_));
  NA3        u0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n649_));
  NAi31      u0627(.An(men_men_n649_), .B(men_men_n218_), .C(i_11_), .Y(men_men_n650_));
  AOI210     u0628(.A0(men_men_n650_), .A1(men_men_n648_), .B0(men_men_n63_), .Y(men_men_n651_));
  NA2        u0629(.A(men_men_n230_), .B(men_men_n63_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n63_), .B(i_9_), .Y(men_men_n653_));
  NO2        u0631(.A(i_1_), .B(i_12_), .Y(men_men_n654_));
  INV        u0632(.A(men_men_n652_), .Y(men_men_n655_));
  OAI210     u0633(.A0(men_men_n655_), .A1(men_men_n651_), .B0(i_6_), .Y(men_men_n656_));
  NO2        u0634(.A(men_men_n649_), .B(men_men_n108_), .Y(men_men_n657_));
  NA2        u0635(.A(men_men_n657_), .B(men_men_n606_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n241_), .B(men_men_n86_), .Y(men_men_n659_));
  NO2        u0637(.A(men_men_n659_), .B(i_11_), .Y(men_men_n660_));
  NA2        u0638(.A(men_men_n658_), .B(men_men_n478_), .Y(men_men_n661_));
  NO4        u0639(.A(men_men_n218_), .B(men_men_n128_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(men_men_n653_), .Y(men_men_n663_));
  NA2        u0641(.A(men_men_n241_), .B(i_6_), .Y(men_men_n664_));
  NO3        u0642(.A(men_men_n637_), .B(men_men_n237_), .C(men_men_n23_), .Y(men_men_n665_));
  AOI210     u0643(.A0(i_1_), .A1(men_men_n265_), .B0(men_men_n665_), .Y(men_men_n666_));
  OAI210     u0644(.A0(men_men_n666_), .A1(men_men_n45_), .B0(men_men_n663_), .Y(men_men_n667_));
  NA3        u0645(.A(men_men_n562_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n668_));
  NA2        u0646(.A(men_men_n138_), .B(i_9_), .Y(men_men_n669_));
  NA3        u0647(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n670_));
  NO2        u0648(.A(men_men_n47_), .B(i_1_), .Y(men_men_n671_));
  NA3        u0649(.A(men_men_n671_), .B(men_men_n274_), .C(men_men_n45_), .Y(men_men_n672_));
  OAI220     u0650(.A0(men_men_n672_), .A1(men_men_n670_), .B0(men_men_n669_), .B1(men_men_n1058_), .Y(men_men_n673_));
  NA3        u0651(.A(men_men_n653_), .B(men_men_n326_), .C(i_6_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(men_men_n23_), .Y(men_men_n675_));
  AOI210     u0653(.A0(men_men_n499_), .A1(men_men_n440_), .B0(men_men_n246_), .Y(men_men_n676_));
  NO2        u0654(.A(men_men_n676_), .B(men_men_n628_), .Y(men_men_n677_));
  NAi21      u0655(.An(men_men_n668_), .B(men_men_n92_), .Y(men_men_n678_));
  NA2        u0656(.A(men_men_n671_), .B(men_men_n274_), .Y(men_men_n679_));
  NO2        u0657(.A(i_11_), .B(men_men_n37_), .Y(men_men_n680_));
  NA2        u0658(.A(men_men_n680_), .B(men_men_n24_), .Y(men_men_n681_));
  OAI210     u0659(.A0(men_men_n681_), .A1(men_men_n679_), .B0(men_men_n678_), .Y(men_men_n682_));
  OR4        u0660(.A(men_men_n682_), .B(men_men_n677_), .C(men_men_n675_), .D(men_men_n673_), .Y(men_men_n683_));
  NO3        u0661(.A(men_men_n683_), .B(men_men_n667_), .C(men_men_n661_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n241_), .B(men_men_n101_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n685_), .B(men_men_n645_), .Y(men_men_n686_));
  NA2        u0664(.A(men_men_n686_), .B(i_1_), .Y(men_men_n687_));
  NO2        u0665(.A(men_men_n687_), .B(men_men_n639_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n435_), .B(men_men_n86_), .Y(men_men_n689_));
  NA2        u0667(.A(men_men_n688_), .B(men_men_n47_), .Y(men_men_n690_));
  NO2        u0668(.A(men_men_n237_), .B(men_men_n45_), .Y(men_men_n691_));
  NO3        u0669(.A(men_men_n691_), .B(men_men_n316_), .C(men_men_n242_), .Y(men_men_n692_));
  NO2        u0670(.A(men_men_n117_), .B(men_men_n37_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n693_), .B(i_6_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n86_), .B(i_9_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n695_), .B(men_men_n63_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n696_), .B(men_men_n654_), .Y(men_men_n697_));
  NO4        u0675(.A(men_men_n697_), .B(men_men_n694_), .C(men_men_n692_), .D(i_4_), .Y(men_men_n698_));
  NA2        u0676(.A(i_1_), .B(i_3_), .Y(men_men_n699_));
  INV        u0677(.A(men_men_n698_), .Y(men_men_n700_));
  NA4        u0678(.A(men_men_n700_), .B(men_men_n690_), .C(men_men_n684_), .D(men_men_n656_), .Y(men_men_n701_));
  NA2        u0679(.A(men_men_n386_), .B(men_men_n385_), .Y(men_men_n702_));
  NA3        u0680(.A(men_men_n508_), .B(men_men_n543_), .C(men_men_n47_), .Y(men_men_n703_));
  NO3        u0681(.A(men_men_n502_), .B(men_men_n631_), .C(men_men_n86_), .Y(men_men_n704_));
  NA2        u0682(.A(men_men_n704_), .B(men_men_n25_), .Y(men_men_n705_));
  NA3        u0683(.A(men_men_n161_), .B(men_men_n84_), .C(men_men_n86_), .Y(men_men_n706_));
  NA4        u0684(.A(men_men_n706_), .B(men_men_n705_), .C(men_men_n703_), .D(men_men_n702_), .Y(men_men_n707_));
  NA2        u0685(.A(men_men_n707_), .B(i_1_), .Y(men_men_n708_));
  AOI210     u0686(.A0(men_men_n274_), .A1(men_men_n97_), .B0(i_1_), .Y(men_men_n709_));
  NO2        u0687(.A(men_men_n384_), .B(i_2_), .Y(men_men_n710_));
  NA2        u0688(.A(men_men_n710_), .B(men_men_n709_), .Y(men_men_n711_));
  OAI210     u0689(.A0(men_men_n674_), .A1(men_men_n470_), .B0(men_men_n711_), .Y(men_men_n712_));
  INV        u0690(.A(men_men_n712_), .Y(men_men_n713_));
  AOI210     u0691(.A0(men_men_n713_), .A1(men_men_n708_), .B0(i_13_), .Y(men_men_n714_));
  OR2        u0692(.A(i_11_), .B(i_7_), .Y(men_men_n715_));
  NA3        u0693(.A(men_men_n715_), .B(men_men_n106_), .C(men_men_n138_), .Y(men_men_n716_));
  AOI220     u0694(.A0(men_men_n493_), .A1(men_men_n161_), .B0(men_men_n472_), .B1(men_men_n138_), .Y(men_men_n717_));
  OAI210     u0695(.A0(men_men_n717_), .A1(men_men_n45_), .B0(men_men_n716_), .Y(men_men_n718_));
  NO2        u0696(.A(men_men_n55_), .B(i_12_), .Y(men_men_n719_));
  INV        u0697(.A(men_men_n719_), .Y(men_men_n720_));
  NO2        u0698(.A(men_men_n502_), .B(men_men_n24_), .Y(men_men_n721_));
  AOI220     u0699(.A0(men_men_n721_), .A1(men_men_n689_), .B0(men_men_n249_), .B1(men_men_n131_), .Y(men_men_n722_));
  OAI220     u0700(.A0(men_men_n722_), .A1(men_men_n41_), .B0(men_men_n720_), .B1(men_men_n93_), .Y(men_men_n723_));
  AOI210     u0701(.A0(men_men_n718_), .A1(men_men_n341_), .B0(men_men_n723_), .Y(men_men_n724_));
  INV        u0702(.A(men_men_n115_), .Y(men_men_n725_));
  AOI220     u0703(.A0(men_men_n725_), .A1(men_men_n72_), .B0(men_men_n400_), .B1(men_men_n671_), .Y(men_men_n726_));
  NO2        u0704(.A(men_men_n726_), .B(men_men_n247_), .Y(men_men_n727_));
  AOI210     u0705(.A0(men_men_n470_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n728_));
  NA2        u0706(.A(men_men_n127_), .B(i_13_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n670_), .B(men_men_n115_), .Y(men_men_n730_));
  INV        u0708(.A(men_men_n730_), .Y(men_men_n731_));
  OAI220     u0709(.A0(men_men_n731_), .A1(men_men_n71_), .B0(men_men_n729_), .B1(men_men_n709_), .Y(men_men_n732_));
  NA2        u0710(.A(men_men_n26_), .B(men_men_n194_), .Y(men_men_n733_));
  NA2        u0711(.A(men_men_n733_), .B(i_7_), .Y(men_men_n734_));
  NO3        u0712(.A(men_men_n502_), .B(men_men_n241_), .C(men_men_n86_), .Y(men_men_n735_));
  NA2        u0713(.A(men_men_n735_), .B(men_men_n734_), .Y(men_men_n736_));
  AOI220     u0714(.A0(men_men_n400_), .A1(men_men_n671_), .B0(men_men_n92_), .B1(men_men_n102_), .Y(men_men_n737_));
  OAI220     u0715(.A0(men_men_n737_), .A1(men_men_n626_), .B0(men_men_n736_), .B1(men_men_n641_), .Y(men_men_n738_));
  NO3        u0716(.A(men_men_n738_), .B(men_men_n732_), .C(men_men_n727_), .Y(men_men_n739_));
  OR2        u0717(.A(i_11_), .B(i_6_), .Y(men_men_n740_));
  NA3        u0718(.A(men_men_n625_), .B(men_men_n733_), .C(i_7_), .Y(men_men_n741_));
  AOI210     u0719(.A0(men_men_n741_), .A1(men_men_n731_), .B0(men_men_n740_), .Y(men_men_n742_));
  NA3        u0720(.A(men_men_n429_), .B(men_men_n630_), .C(men_men_n97_), .Y(men_men_n743_));
  NA2        u0721(.A(men_men_n660_), .B(i_13_), .Y(men_men_n744_));
  NAi21      u0722(.An(i_11_), .B(i_12_), .Y(men_men_n745_));
  NOi41      u0723(.An(men_men_n111_), .B(men_men_n745_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n746_));
  NO3        u0724(.A(men_men_n502_), .B(men_men_n606_), .C(men_men_n631_), .Y(men_men_n747_));
  AOI220     u0725(.A0(men_men_n747_), .A1(men_men_n320_), .B0(men_men_n746_), .B1(men_men_n47_), .Y(men_men_n748_));
  NA3        u0726(.A(men_men_n748_), .B(men_men_n744_), .C(men_men_n743_), .Y(men_men_n749_));
  OAI210     u0727(.A0(men_men_n749_), .A1(men_men_n742_), .B0(men_men_n63_), .Y(men_men_n750_));
  NO2        u0728(.A(i_2_), .B(i_12_), .Y(men_men_n751_));
  NA2        u0729(.A(men_men_n383_), .B(men_men_n751_), .Y(men_men_n752_));
  NA2        u0730(.A(i_8_), .B(men_men_n25_), .Y(men_men_n753_));
  NO3        u0731(.A(men_men_n753_), .B(i_3_), .C(men_men_n625_), .Y(men_men_n754_));
  OAI210     u0732(.A0(men_men_n754_), .A1(men_men_n385_), .B0(men_men_n383_), .Y(men_men_n755_));
  NO2        u0733(.A(men_men_n128_), .B(i_2_), .Y(men_men_n756_));
  NA2        u0734(.A(men_men_n756_), .B(men_men_n654_), .Y(men_men_n757_));
  NA3        u0735(.A(men_men_n757_), .B(men_men_n755_), .C(men_men_n752_), .Y(men_men_n758_));
  NA3        u0736(.A(men_men_n758_), .B(men_men_n46_), .C(men_men_n229_), .Y(men_men_n759_));
  NA4        u0737(.A(men_men_n759_), .B(men_men_n750_), .C(men_men_n739_), .D(men_men_n724_), .Y(men_men_n760_));
  OR4        u0738(.A(men_men_n760_), .B(men_men_n714_), .C(men_men_n701_), .D(men_men_n644_), .Y(men5));
  NA2        u0739(.A(men_men_n686_), .B(men_men_n276_), .Y(men_men_n762_));
  AN2        u0740(.A(men_men_n24_), .B(i_10_), .Y(men_men_n763_));
  NA3        u0741(.A(men_men_n763_), .B(men_men_n751_), .C(men_men_n108_), .Y(men_men_n764_));
  NO2        u0742(.A(men_men_n626_), .B(i_11_), .Y(men_men_n765_));
  NA2        u0743(.A(men_men_n87_), .B(men_men_n765_), .Y(men_men_n766_));
  NA3        u0744(.A(men_men_n766_), .B(men_men_n764_), .C(men_men_n762_), .Y(men_men_n767_));
  NO3        u0745(.A(i_11_), .B(men_men_n241_), .C(i_13_), .Y(men_men_n768_));
  NO2        u0746(.A(men_men_n124_), .B(men_men_n23_), .Y(men_men_n769_));
  NA2        u0747(.A(i_12_), .B(i_8_), .Y(men_men_n770_));
  OAI210     u0748(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n770_), .Y(men_men_n771_));
  INV        u0749(.A(men_men_n469_), .Y(men_men_n772_));
  AOI220     u0750(.A0(men_men_n326_), .A1(men_men_n601_), .B0(men_men_n771_), .B1(men_men_n769_), .Y(men_men_n773_));
  INV        u0751(.A(men_men_n773_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n774_), .B(men_men_n767_), .Y(men_men_n775_));
  INV        u0753(.A(men_men_n172_), .Y(men_men_n776_));
  INV        u0754(.A(men_men_n249_), .Y(men_men_n777_));
  OAI210     u0755(.A0(men_men_n710_), .A1(men_men_n471_), .B0(men_men_n111_), .Y(men_men_n778_));
  AOI210     u0756(.A0(men_men_n778_), .A1(men_men_n777_), .B0(men_men_n776_), .Y(men_men_n779_));
  NO2        u0757(.A(men_men_n479_), .B(men_men_n26_), .Y(men_men_n780_));
  NO2        u0758(.A(men_men_n780_), .B(men_men_n440_), .Y(men_men_n781_));
  NA2        u0759(.A(men_men_n781_), .B(i_2_), .Y(men_men_n782_));
  INV        u0760(.A(men_men_n782_), .Y(men_men_n783_));
  AOI210     u0761(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n436_), .Y(men_men_n784_));
  AOI210     u0762(.A0(men_men_n784_), .A1(men_men_n783_), .B0(men_men_n779_), .Y(men_men_n785_));
  NO2        u0763(.A(men_men_n191_), .B(men_men_n125_), .Y(men_men_n786_));
  OAI210     u0764(.A0(men_men_n786_), .A1(men_men_n769_), .B0(i_2_), .Y(men_men_n787_));
  INV        u0765(.A(men_men_n173_), .Y(men_men_n788_));
  NO3        u0766(.A(men_men_n646_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n789_));
  AOI210     u0767(.A0(men_men_n788_), .A1(men_men_n87_), .B0(men_men_n789_), .Y(men_men_n790_));
  AOI210     u0768(.A0(men_men_n790_), .A1(men_men_n787_), .B0(men_men_n194_), .Y(men_men_n791_));
  OA210      u0769(.A0(men_men_n647_), .A1(men_men_n126_), .B0(i_13_), .Y(men_men_n792_));
  NA2        u0770(.A(men_men_n201_), .B(men_men_n204_), .Y(men_men_n793_));
  NA2        u0771(.A(men_men_n151_), .B(men_men_n621_), .Y(men_men_n794_));
  AOI210     u0772(.A0(men_men_n794_), .A1(men_men_n793_), .B0(men_men_n388_), .Y(men_men_n795_));
  AOI210     u0773(.A0(men_men_n211_), .A1(men_men_n148_), .B0(men_men_n543_), .Y(men_men_n796_));
  NA2        u0774(.A(men_men_n796_), .B(men_men_n440_), .Y(men_men_n797_));
  NO2        u0775(.A(men_men_n102_), .B(men_men_n45_), .Y(men_men_n798_));
  INV        u0776(.A(men_men_n308_), .Y(men_men_n799_));
  NA4        u0777(.A(men_men_n799_), .B(men_men_n313_), .C(men_men_n124_), .D(men_men_n43_), .Y(men_men_n800_));
  OAI210     u0778(.A0(men_men_n800_), .A1(men_men_n798_), .B0(men_men_n797_), .Y(men_men_n801_));
  NO4        u0779(.A(men_men_n801_), .B(men_men_n795_), .C(men_men_n792_), .D(men_men_n791_), .Y(men_men_n802_));
  NA2        u0780(.A(men_men_n601_), .B(men_men_n28_), .Y(men_men_n803_));
  NA2        u0781(.A(men_men_n768_), .B(men_men_n280_), .Y(men_men_n804_));
  NA2        u0782(.A(men_men_n804_), .B(men_men_n803_), .Y(men_men_n805_));
  NO2        u0783(.A(men_men_n62_), .B(i_12_), .Y(men_men_n806_));
  NO2        u0784(.A(men_men_n806_), .B(men_men_n126_), .Y(men_men_n807_));
  NO2        u0785(.A(men_men_n807_), .B(men_men_n621_), .Y(men_men_n808_));
  AOI220     u0786(.A0(men_men_n808_), .A1(men_men_n36_), .B0(men_men_n805_), .B1(men_men_n47_), .Y(men_men_n809_));
  NA4        u0787(.A(men_men_n809_), .B(men_men_n802_), .C(men_men_n785_), .D(men_men_n775_), .Y(men6));
  NO3        u0788(.A(men_men_n260_), .B(men_men_n315_), .C(i_1_), .Y(men_men_n811_));
  NO2        u0789(.A(men_men_n186_), .B(men_men_n139_), .Y(men_men_n812_));
  OAI210     u0790(.A0(men_men_n812_), .A1(men_men_n811_), .B0(men_men_n756_), .Y(men_men_n813_));
  NO2        u0791(.A(men_men_n224_), .B(men_men_n512_), .Y(men_men_n814_));
  NO2        u0792(.A(i_11_), .B(i_9_), .Y(men_men_n815_));
  INV        u0793(.A(men_men_n338_), .Y(men_men_n816_));
  AO210      u0794(.A0(men_men_n816_), .A1(men_men_n813_), .B0(i_12_), .Y(men_men_n817_));
  NA2        u0795(.A(men_men_n389_), .B(men_men_n344_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n606_), .B(men_men_n63_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n819_), .B(men_men_n818_), .Y(men_men_n820_));
  INV        u0798(.A(men_men_n198_), .Y(men_men_n821_));
  AOI220     u0799(.A0(men_men_n821_), .A1(men_men_n815_), .B0(men_men_n820_), .B1(men_men_n73_), .Y(men_men_n822_));
  INV        u0800(.A(men_men_n337_), .Y(men_men_n823_));
  NA2        u0801(.A(men_men_n75_), .B(men_men_n131_), .Y(men_men_n824_));
  INV        u0802(.A(men_men_n124_), .Y(men_men_n825_));
  NA2        u0803(.A(men_men_n825_), .B(men_men_n47_), .Y(men_men_n826_));
  AOI210     u0804(.A0(men_men_n826_), .A1(men_men_n824_), .B0(men_men_n823_), .Y(men_men_n827_));
  NO2        u0805(.A(men_men_n256_), .B(i_9_), .Y(men_men_n828_));
  NA2        u0806(.A(men_men_n828_), .B(men_men_n806_), .Y(men_men_n829_));
  AOI210     u0807(.A0(men_men_n829_), .A1(men_men_n541_), .B0(men_men_n186_), .Y(men_men_n830_));
  NO2        u0808(.A(men_men_n32_), .B(i_11_), .Y(men_men_n831_));
  NAi32      u0809(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n740_), .B(men_men_n832_), .Y(men_men_n833_));
  OR3        u0811(.A(men_men_n833_), .B(men_men_n830_), .C(men_men_n827_), .Y(men_men_n834_));
  NO2        u0812(.A(men_men_n715_), .B(i_2_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n836_));
  NO2        u0814(.A(men_men_n836_), .B(men_men_n428_), .Y(men_men_n837_));
  NA2        u0815(.A(men_men_n837_), .B(men_men_n835_), .Y(men_men_n838_));
  AO220      u0816(.A0(men_men_n372_), .A1(men_men_n362_), .B0(men_men_n412_), .B1(men_men_n621_), .Y(men_men_n839_));
  NA3        u0817(.A(men_men_n839_), .B(men_men_n261_), .C(i_7_), .Y(men_men_n840_));
  OR2        u0818(.A(men_men_n647_), .B(men_men_n471_), .Y(men_men_n841_));
  NA3        u0819(.A(men_men_n841_), .B(men_men_n147_), .C(men_men_n69_), .Y(men_men_n842_));
  AO210      u0820(.A0(men_men_n519_), .A1(men_men_n772_), .B0(men_men_n36_), .Y(men_men_n843_));
  NA4        u0821(.A(men_men_n843_), .B(men_men_n842_), .C(men_men_n840_), .D(men_men_n838_), .Y(men_men_n844_));
  NO2        u0822(.A(men_men_n659_), .B(i_11_), .Y(men_men_n845_));
  AOI220     u0823(.A0(men_men_n845_), .A1(men_men_n591_), .B0(men_men_n814_), .B1(men_men_n734_), .Y(men_men_n846_));
  NA3        u0824(.A(men_men_n388_), .B(men_men_n243_), .C(men_men_n147_), .Y(men_men_n847_));
  NA2        u0825(.A(men_men_n412_), .B(men_men_n70_), .Y(men_men_n848_));
  NA4        u0826(.A(men_men_n848_), .B(men_men_n847_), .C(men_men_n846_), .D(men_men_n629_), .Y(men_men_n849_));
  AOI210     u0827(.A0(men_men_n471_), .A1(men_men_n469_), .B0(men_men_n590_), .Y(men_men_n850_));
  NA2        u0828(.A(men_men_n112_), .B(men_men_n426_), .Y(men_men_n851_));
  NA2        u0829(.A(men_men_n248_), .B(men_men_n47_), .Y(men_men_n852_));
  INV        u0830(.A(men_men_n612_), .Y(men_men_n853_));
  NA3        u0831(.A(men_men_n853_), .B(men_men_n337_), .C(i_7_), .Y(men_men_n854_));
  NA3        u0832(.A(men_men_n854_), .B(men_men_n851_), .C(men_men_n850_), .Y(men_men_n855_));
  NO4        u0833(.A(men_men_n855_), .B(men_men_n849_), .C(men_men_n844_), .D(men_men_n834_), .Y(men_men_n856_));
  NA4        u0834(.A(men_men_n856_), .B(men_men_n822_), .C(men_men_n817_), .D(men_men_n395_), .Y(men3));
  NA2        u0835(.A(i_12_), .B(i_10_), .Y(men_men_n858_));
  NA2        u0836(.A(i_6_), .B(i_7_), .Y(men_men_n859_));
  NO2        u0837(.A(men_men_n859_), .B(i_0_), .Y(men_men_n860_));
  NO2        u0838(.A(i_11_), .B(men_men_n241_), .Y(men_men_n861_));
  OAI210     u0839(.A0(men_men_n860_), .A1(men_men_n296_), .B0(men_men_n861_), .Y(men_men_n862_));
  NO2        u0840(.A(men_men_n862_), .B(men_men_n194_), .Y(men_men_n863_));
  NO3        u0841(.A(men_men_n475_), .B(men_men_n90_), .C(men_men_n45_), .Y(men_men_n864_));
  OA210      u0842(.A0(men_men_n864_), .A1(men_men_n863_), .B0(men_men_n175_), .Y(men_men_n865_));
  NA3        u0843(.A(men_men_n847_), .B(men_men_n629_), .C(men_men_n387_), .Y(men_men_n866_));
  NA2        u0844(.A(men_men_n866_), .B(men_men_n40_), .Y(men_men_n867_));
  NOi21      u0845(.An(men_men_n96_), .B(men_men_n781_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n429_), .B(men_men_n46_), .Y(men_men_n869_));
  INV        u0847(.A(men_men_n868_), .Y(men_men_n870_));
  AOI210     u0848(.A0(men_men_n870_), .A1(men_men_n867_), .B0(men_men_n49_), .Y(men_men_n871_));
  NO4        u0849(.A(men_men_n392_), .B(men_men_n398_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n872_));
  NA2        u0850(.A(men_men_n186_), .B(men_men_n599_), .Y(men_men_n873_));
  NOi21      u0851(.An(men_men_n873_), .B(men_men_n872_), .Y(men_men_n874_));
  NA2        u0852(.A(men_men_n728_), .B(men_men_n695_), .Y(men_men_n875_));
  NA2        u0853(.A(men_men_n342_), .B(men_men_n460_), .Y(men_men_n876_));
  OAI220     u0854(.A0(men_men_n876_), .A1(men_men_n875_), .B0(men_men_n874_), .B1(men_men_n63_), .Y(men_men_n877_));
  NOi21      u0855(.An(i_5_), .B(i_9_), .Y(men_men_n878_));
  NA2        u0856(.A(men_men_n878_), .B(men_men_n468_), .Y(men_men_n879_));
  BUFFER     u0857(.A(men_men_n274_), .Y(men_men_n880_));
  AOI210     u0858(.A0(men_men_n880_), .A1(men_men_n499_), .B0(men_men_n704_), .Y(men_men_n881_));
  NO2        u0859(.A(men_men_n176_), .B(men_men_n148_), .Y(men_men_n882_));
  NO2        u0860(.A(men_men_n881_), .B(men_men_n879_), .Y(men_men_n883_));
  NO4        u0861(.A(men_men_n883_), .B(men_men_n877_), .C(men_men_n871_), .D(men_men_n865_), .Y(men_men_n884_));
  NA2        u0862(.A(men_men_n186_), .B(men_men_n24_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n320_), .B(men_men_n129_), .Y(men_men_n886_));
  NAi21      u0864(.An(men_men_n162_), .B(men_men_n460_), .Y(men_men_n887_));
  OAI220     u0865(.A0(men_men_n887_), .A1(men_men_n852_), .B0(men_men_n886_), .B1(men_men_n418_), .Y(men_men_n888_));
  INV        u0866(.A(men_men_n888_), .Y(men_men_n889_));
  NO2        u0867(.A(men_men_n404_), .B(men_men_n300_), .Y(men_men_n890_));
  NA2        u0868(.A(men_men_n890_), .B(men_men_n730_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n600_), .B(i_0_), .Y(men_men_n892_));
  NO4        u0870(.A(men_men_n611_), .B(men_men_n218_), .C(men_men_n436_), .D(men_men_n428_), .Y(men_men_n893_));
  INV        u0871(.A(men_men_n497_), .Y(men_men_n894_));
  NA2        u0872(.A(men_men_n768_), .B(men_men_n338_), .Y(men_men_n895_));
  INV        u0873(.A(men_men_n58_), .Y(men_men_n896_));
  OAI220     u0874(.A0(men_men_n896_), .A1(men_men_n895_), .B0(men_men_n681_), .B1(men_men_n564_), .Y(men_men_n897_));
  NO2        u0875(.A(men_men_n258_), .B(men_men_n153_), .Y(men_men_n898_));
  NA2        u0876(.A(i_0_), .B(i_10_), .Y(men_men_n899_));
  AN2        u0877(.A(men_men_n898_), .B(i_6_), .Y(men_men_n900_));
  AOI220     u0878(.A0(men_men_n342_), .A1(men_men_n98_), .B0(men_men_n186_), .B1(men_men_n84_), .Y(men_men_n901_));
  NA2        u0879(.A(men_men_n595_), .B(i_4_), .Y(men_men_n902_));
  NO2        u0880(.A(men_men_n902_), .B(men_men_n901_), .Y(men_men_n903_));
  NO3        u0881(.A(men_men_n903_), .B(men_men_n900_), .C(men_men_n897_), .Y(men_men_n904_));
  NA3        u0882(.A(men_men_n904_), .B(men_men_n891_), .C(men_men_n889_), .Y(men_men_n905_));
  NA2        u0883(.A(i_11_), .B(i_9_), .Y(men_men_n906_));
  NA2        u0884(.A(men_men_n409_), .B(men_men_n180_), .Y(men_men_n907_));
  NA2        u0885(.A(men_men_n907_), .B(men_men_n160_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n906_), .B(men_men_n73_), .Y(men_men_n909_));
  NO2        u0887(.A(men_men_n176_), .B(i_0_), .Y(men_men_n910_));
  INV        u0888(.A(men_men_n910_), .Y(men_men_n911_));
  NA2        u0889(.A(men_men_n497_), .B(men_men_n235_), .Y(men_men_n912_));
  AOI210     u0890(.A0(men_men_n386_), .A1(men_men_n42_), .B0(men_men_n425_), .Y(men_men_n913_));
  OAI220     u0891(.A0(men_men_n913_), .A1(men_men_n879_), .B0(men_men_n912_), .B1(men_men_n911_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n914_), .B(men_men_n908_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n680_), .B(men_men_n121_), .Y(men_men_n916_));
  NO2        u0894(.A(i_6_), .B(men_men_n916_), .Y(men_men_n917_));
  AOI210     u0895(.A0(men_men_n470_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n172_), .B(men_men_n103_), .Y(men_men_n919_));
  NOi32      u0897(.An(men_men_n918_), .Bn(men_men_n189_), .C(men_men_n919_), .Y(men_men_n920_));
  NA2        u0898(.A(men_men_n630_), .B(men_men_n338_), .Y(men_men_n921_));
  NO2        u0899(.A(men_men_n921_), .B(men_men_n869_), .Y(men_men_n922_));
  NO3        u0900(.A(men_men_n922_), .B(men_men_n920_), .C(men_men_n917_), .Y(men_men_n923_));
  NOi21      u0901(.An(i_7_), .B(i_5_), .Y(men_men_n924_));
  OR2        u0902(.A(men_men_n919_), .B(men_men_n541_), .Y(men_men_n925_));
  NO3        u0903(.A(men_men_n421_), .B(men_men_n375_), .C(men_men_n371_), .Y(men_men_n926_));
  NO2        u0904(.A(men_men_n268_), .B(men_men_n327_), .Y(men_men_n927_));
  NO2        u0905(.A(men_men_n745_), .B(men_men_n263_), .Y(men_men_n928_));
  AOI210     u0906(.A0(men_men_n928_), .A1(men_men_n927_), .B0(men_men_n926_), .Y(men_men_n929_));
  NA4        u0907(.A(men_men_n929_), .B(men_men_n925_), .C(men_men_n923_), .D(men_men_n915_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n885_), .B(men_men_n244_), .Y(men_men_n931_));
  AN2        u0909(.A(men_men_n341_), .B(men_men_n338_), .Y(men_men_n932_));
  AN2        u0910(.A(men_men_n932_), .B(men_men_n882_), .Y(men_men_n933_));
  OAI210     u0911(.A0(men_men_n933_), .A1(men_men_n931_), .B0(i_10_), .Y(men_men_n934_));
  NO2        u0912(.A(men_men_n858_), .B(men_men_n326_), .Y(men_men_n935_));
  NA2        u0913(.A(men_men_n935_), .B(men_men_n909_), .Y(men_men_n936_));
  NA3        u0914(.A(men_men_n496_), .B(men_men_n429_), .C(men_men_n46_), .Y(men_men_n937_));
  OAI210     u0915(.A0(men_men_n887_), .A1(men_men_n894_), .B0(men_men_n937_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n261_), .B(men_men_n47_), .Y(men_men_n939_));
  NA2        u0917(.A(men_men_n909_), .B(men_men_n313_), .Y(men_men_n940_));
  OAI210     u0918(.A0(men_men_n939_), .A1(men_men_n188_), .B0(men_men_n940_), .Y(men_men_n941_));
  AOI220     u0919(.A0(men_men_n941_), .A1(men_men_n497_), .B0(men_men_n938_), .B1(men_men_n73_), .Y(men_men_n942_));
  NA3        u0920(.A(men_men_n836_), .B(men_men_n397_), .C(men_men_n659_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n943_), .B(men_men_n48_), .Y(men_men_n944_));
  NO3        u0922(.A(men_men_n611_), .B(men_men_n370_), .C(men_men_n24_), .Y(men_men_n945_));
  AOI210     u0923(.A0(men_men_n721_), .A1(men_men_n574_), .B0(men_men_n945_), .Y(men_men_n946_));
  NAi21      u0924(.An(i_9_), .B(i_5_), .Y(men_men_n947_));
  NO2        u0925(.A(men_men_n947_), .B(men_men_n421_), .Y(men_men_n948_));
  NO2        u0926(.A(men_men_n624_), .B(men_men_n105_), .Y(men_men_n949_));
  AOI220     u0927(.A0(men_men_n949_), .A1(i_0_), .B0(men_men_n948_), .B1(men_men_n647_), .Y(men_men_n950_));
  OAI220     u0928(.A0(men_men_n950_), .A1(men_men_n86_), .B0(men_men_n946_), .B1(men_men_n173_), .Y(men_men_n951_));
  NO3        u0929(.A(men_men_n951_), .B(men_men_n944_), .C(men_men_n545_), .Y(men_men_n952_));
  NA4        u0930(.A(men_men_n952_), .B(men_men_n942_), .C(men_men_n936_), .D(men_men_n934_), .Y(men_men_n953_));
  NO3        u0931(.A(men_men_n953_), .B(men_men_n930_), .C(men_men_n905_), .Y(men_men_n954_));
  NA2        u0932(.A(men_men_n73_), .B(men_men_n45_), .Y(men_men_n955_));
  NA2        u0933(.A(men_men_n899_), .B(men_men_n955_), .Y(men_men_n956_));
  NO3        u0934(.A(men_men_n105_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n957_));
  AN2        u0935(.A(men_men_n957_), .B(men_men_n956_), .Y(men_men_n958_));
  AOI210     u0936(.A0(men_men_n819_), .A1(men_men_n702_), .B0(men_men_n919_), .Y(men_men_n959_));
  AOI210     u0937(.A0(men_men_n958_), .A1(men_men_n359_), .B0(men_men_n959_), .Y(men_men_n960_));
  NA2        u0938(.A(men_men_n756_), .B(men_men_n146_), .Y(men_men_n961_));
  INV        u0939(.A(men_men_n961_), .Y(men_men_n962_));
  NA3        u0940(.A(men_men_n962_), .B(men_men_n695_), .C(men_men_n73_), .Y(men_men_n963_));
  NA3        u0941(.A(men_men_n860_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n964_));
  NA2        u0942(.A(men_men_n861_), .B(i_9_), .Y(men_men_n965_));
  AOI210     u0943(.A0(men_men_n964_), .A1(men_men_n524_), .B0(men_men_n965_), .Y(men_men_n966_));
  OAI210     u0944(.A0(men_men_n248_), .A1(i_9_), .B0(men_men_n234_), .Y(men_men_n967_));
  AOI210     u0945(.A0(men_men_n967_), .A1(men_men_n892_), .B0(men_men_n153_), .Y(men_men_n968_));
  NO2        u0946(.A(men_men_n968_), .B(men_men_n966_), .Y(men_men_n969_));
  NA3        u0947(.A(men_men_n969_), .B(men_men_n963_), .C(men_men_n960_), .Y(men_men_n970_));
  NA2        u0948(.A(men_men_n932_), .B(men_men_n388_), .Y(men_men_n971_));
  AOI210     u0949(.A0(men_men_n307_), .A1(men_men_n162_), .B0(men_men_n971_), .Y(men_men_n972_));
  NA3        u0950(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n973_));
  NA2        u0951(.A(i_5_), .B(men_men_n513_), .Y(men_men_n974_));
  AOI210     u0952(.A0(men_men_n973_), .A1(men_men_n162_), .B0(men_men_n974_), .Y(men_men_n975_));
  NO2        u0953(.A(men_men_n975_), .B(men_men_n972_), .Y(men_men_n976_));
  NO3        u0954(.A(men_men_n899_), .B(men_men_n878_), .C(men_men_n191_), .Y(men_men_n977_));
  AOI220     u0955(.A0(men_men_n977_), .A1(i_11_), .B0(men_men_n596_), .B1(men_men_n75_), .Y(men_men_n978_));
  NO3        u0956(.A(men_men_n212_), .B(men_men_n398_), .C(i_0_), .Y(men_men_n979_));
  OAI210     u0957(.A0(men_men_n979_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n980_));
  INV        u0958(.A(men_men_n221_), .Y(men_men_n981_));
  OAI220     u0959(.A0(men_men_n557_), .A1(men_men_n139_), .B0(men_men_n664_), .B1(men_men_n641_), .Y(men_men_n982_));
  NA3        u0960(.A(men_men_n982_), .B(men_men_n413_), .C(men_men_n981_), .Y(men_men_n983_));
  NA4        u0961(.A(men_men_n983_), .B(men_men_n980_), .C(men_men_n978_), .D(men_men_n976_), .Y(men_men_n984_));
  INV        u0962(.A(men_men_n109_), .Y(men_men_n985_));
  AOI220     u0963(.A0(men_men_n924_), .A1(men_men_n513_), .B0(men_men_n860_), .B1(men_men_n163_), .Y(men_men_n986_));
  NA2        u0964(.A(men_men_n362_), .B(men_men_n177_), .Y(men_men_n987_));
  OA220      u0965(.A0(men_men_n987_), .A1(men_men_n986_), .B0(men_men_n985_), .B1(i_5_), .Y(men_men_n988_));
  NA3        u0966(.A(men_men_n638_), .B(men_men_n186_), .C(men_men_n84_), .Y(men_men_n989_));
  INV        u0967(.A(men_men_n989_), .Y(men_men_n990_));
  NO3        u0968(.A(men_men_n869_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n991_));
  NA2        u0969(.A(men_men_n518_), .B(men_men_n494_), .Y(men_men_n992_));
  NO3        u0970(.A(men_men_n992_), .B(men_men_n991_), .C(men_men_n990_), .Y(men_men_n993_));
  NA3        u0971(.A(men_men_n404_), .B(men_men_n343_), .C(men_men_n225_), .Y(men_men_n994_));
  INV        u0972(.A(men_men_n994_), .Y(men_men_n995_));
  NOi31      u0973(.An(men_men_n403_), .B(men_men_n955_), .C(men_men_n244_), .Y(men_men_n996_));
  NO3        u0974(.A(men_men_n906_), .B(men_men_n221_), .C(men_men_n191_), .Y(men_men_n997_));
  NO3        u0975(.A(men_men_n997_), .B(men_men_n996_), .C(men_men_n995_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n998_), .B(men_men_n993_), .C(men_men_n988_), .Y(men_men_n999_));
  INV        u0977(.A(men_men_n640_), .Y(men_men_n1000_));
  NO3        u0978(.A(men_men_n1000_), .B(men_men_n586_), .C(men_men_n356_), .Y(men_men_n1001_));
  NO2        u0979(.A(men_men_n86_), .B(i_5_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n861_), .B(men_men_n110_), .C(men_men_n124_), .Y(men_men_n1003_));
  INV        u0981(.A(men_men_n1003_), .Y(men_men_n1004_));
  AOI210     u0982(.A0(men_men_n1004_), .A1(men_men_n1002_), .B0(men_men_n1001_), .Y(men_men_n1005_));
  AN2        u0983(.A(men_men_n899_), .B(men_men_n153_), .Y(men_men_n1006_));
  NO4        u0984(.A(men_men_n1006_), .B(i_12_), .C(men_men_n668_), .D(men_men_n131_), .Y(men_men_n1007_));
  NA2        u0985(.A(men_men_n1007_), .B(men_men_n221_), .Y(men_men_n1008_));
  NA3        u0986(.A(men_men_n98_), .B(men_men_n599_), .C(i_11_), .Y(men_men_n1009_));
  NO2        u0987(.A(men_men_n1009_), .B(men_men_n155_), .Y(men_men_n1010_));
  INV        u0988(.A(men_men_n1010_), .Y(men_men_n1011_));
  NA3        u0989(.A(men_men_n1011_), .B(men_men_n1008_), .C(men_men_n1005_), .Y(men_men_n1012_));
  NO4        u0990(.A(men_men_n1012_), .B(men_men_n999_), .C(men_men_n984_), .D(men_men_n970_), .Y(men_men_n1013_));
  OAI210     u0991(.A0(men_men_n835_), .A1(men_men_n831_), .B0(men_men_n37_), .Y(men_men_n1014_));
  NA3        u0992(.A(men_men_n918_), .B(men_men_n383_), .C(i_5_), .Y(men_men_n1015_));
  NA3        u0993(.A(men_men_n1015_), .B(men_men_n1014_), .C(men_men_n636_), .Y(men_men_n1016_));
  NA2        u0994(.A(men_men_n1016_), .B(men_men_n209_), .Y(men_men_n1017_));
  NA2        u0995(.A(men_men_n187_), .B(men_men_n189_), .Y(men_men_n1018_));
  AO210      u0996(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n1018_), .Y(men_men_n1019_));
  OAI210     u0997(.A0(men_men_n640_), .A1(men_men_n638_), .B0(men_men_n326_), .Y(men_men_n1020_));
  NAi31      u0998(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1021_));
  NO2        u0999(.A(men_men_n70_), .B(men_men_n1021_), .Y(men_men_n1022_));
  NO2        u1000(.A(men_men_n1022_), .B(men_men_n665_), .Y(men_men_n1023_));
  NA3        u1001(.A(men_men_n1023_), .B(men_men_n1020_), .C(men_men_n1019_), .Y(men_men_n1024_));
  NO2        u1002(.A(men_men_n483_), .B(men_men_n274_), .Y(men_men_n1025_));
  NO4        u1003(.A(men_men_n237_), .B(men_men_n145_), .C(men_men_n699_), .D(men_men_n37_), .Y(men_men_n1026_));
  NO3        u1004(.A(men_men_n1026_), .B(men_men_n1025_), .C(men_men_n893_), .Y(men_men_n1027_));
  OAI210     u1005(.A0(men_men_n1009_), .A1(men_men_n148_), .B0(men_men_n1027_), .Y(men_men_n1028_));
  AOI210     u1006(.A0(men_men_n1024_), .A1(men_men_n49_), .B0(men_men_n1028_), .Y(men_men_n1029_));
  AOI210     u1007(.A0(men_men_n1029_), .A1(men_men_n1017_), .B0(men_men_n73_), .Y(men_men_n1030_));
  NO2        u1008(.A(men_men_n593_), .B(men_men_n394_), .Y(men_men_n1031_));
  NO2        u1009(.A(men_men_n1031_), .B(men_men_n776_), .Y(men_men_n1032_));
  INV        u1010(.A(men_men_n76_), .Y(men_men_n1033_));
  NO2        u1011(.A(men_men_n1033_), .B(men_men_n699_), .Y(men_men_n1034_));
  NA2        u1012(.A(men_men_n268_), .B(men_men_n57_), .Y(men_men_n1035_));
  AOI220     u1013(.A0(men_men_n1035_), .A1(men_men_n76_), .B0(men_men_n357_), .B1(men_men_n260_), .Y(men_men_n1036_));
  NO2        u1014(.A(men_men_n1036_), .B(men_men_n241_), .Y(men_men_n1037_));
  NA3        u1015(.A(men_men_n96_), .B(men_men_n315_), .C(men_men_n31_), .Y(men_men_n1038_));
  INV        u1016(.A(men_men_n1038_), .Y(men_men_n1039_));
  NO3        u1017(.A(men_men_n1039_), .B(men_men_n1037_), .C(men_men_n1034_), .Y(men_men_n1040_));
  NA2        u1018(.A(men_men_n158_), .B(men_men_n87_), .Y(men_men_n1041_));
  NA3        u1019(.A(men_men_n780_), .B(men_men_n296_), .C(men_men_n80_), .Y(men_men_n1042_));
  AOI210     u1020(.A0(men_men_n1042_), .A1(men_men_n1041_), .B0(i_11_), .Y(men_men_n1043_));
  NA2        u1021(.A(men_men_n631_), .B(men_men_n218_), .Y(men_men_n1044_));
  OAI210     u1022(.A0(men_men_n1044_), .A1(men_men_n918_), .B0(men_men_n209_), .Y(men_men_n1045_));
  NA2        u1023(.A(men_men_n164_), .B(i_5_), .Y(men_men_n1046_));
  NO2        u1024(.A(men_men_n1045_), .B(men_men_n1046_), .Y(men_men_n1047_));
  NO4        u1025(.A(men_men_n947_), .B(men_men_n501_), .C(men_men_n257_), .D(men_men_n256_), .Y(men_men_n1048_));
  NO2        u1026(.A(men_men_n1048_), .B(men_men_n590_), .Y(men_men_n1049_));
  INV        u1027(.A(men_men_n376_), .Y(men_men_n1050_));
  AOI210     u1028(.A0(men_men_n1050_), .A1(men_men_n1049_), .B0(men_men_n41_), .Y(men_men_n1051_));
  NO3        u1029(.A(men_men_n1051_), .B(men_men_n1047_), .C(men_men_n1043_), .Y(men_men_n1052_));
  OAI210     u1030(.A0(men_men_n1040_), .A1(i_4_), .B0(men_men_n1052_), .Y(men_men_n1053_));
  NO3        u1031(.A(men_men_n1053_), .B(men_men_n1032_), .C(men_men_n1030_), .Y(men_men_n1054_));
  NA4        u1032(.A(men_men_n1054_), .B(men_men_n1013_), .C(men_men_n954_), .D(men_men_n884_), .Y(men4));
  INV        u1033(.A(i_2_), .Y(men_men_n1058_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule