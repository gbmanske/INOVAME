//Benchmark atmr_max1024_476_0.0313

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  INV        o012(.A(ori_ori_n24_), .Y(ori_ori_n29_));
  NO2        o013(.A(x4), .B(x3), .Y(ori_ori_n30_));
  INV        o014(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  OA210      o015(.A0(ori_ori_n31_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n32_));
  NOi31      o016(.An(ori_ori_n23_), .B(ori_ori_n32_), .C(ori_ori_n29_), .Y(ori00));
  NO2        o017(.A(x1), .B(x0), .Y(ori_ori_n34_));
  INV        o018(.A(x6), .Y(ori_ori_n35_));
  NO2        o019(.A(ori_ori_n35_), .B(ori_ori_n25_), .Y(ori_ori_n36_));
  AN2        o020(.A(x8), .B(x7), .Y(ori_ori_n37_));
  NA3        o021(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(ori_ori_n34_), .Y(ori_ori_n38_));
  NA2        o022(.A(x4), .B(x3), .Y(ori_ori_n39_));
  AOI210     o023(.A0(ori_ori_n38_), .A1(ori_ori_n23_), .B0(ori_ori_n39_), .Y(ori_ori_n40_));
  NO2        o024(.A(x2), .B(x0), .Y(ori_ori_n41_));
  INV        o025(.A(x3), .Y(ori_ori_n42_));
  NO2        o026(.A(ori_ori_n42_), .B(ori_ori_n18_), .Y(ori_ori_n43_));
  INV        o027(.A(ori_ori_n43_), .Y(ori_ori_n44_));
  NO2        o028(.A(ori_ori_n36_), .B(x4), .Y(ori_ori_n45_));
  OAI210     o029(.A0(ori_ori_n45_), .A1(ori_ori_n44_), .B0(ori_ori_n41_), .Y(ori_ori_n46_));
  INV        o030(.A(x4), .Y(ori_ori_n47_));
  NO2        o031(.A(ori_ori_n47_), .B(ori_ori_n17_), .Y(ori_ori_n48_));
  NA2        o032(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n49_));
  OAI210     o033(.A0(ori_ori_n49_), .A1(ori_ori_n20_), .B0(ori_ori_n46_), .Y(ori_ori_n50_));
  NA2        o034(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n51_));
  AOI220     o035(.A0(ori_ori_n51_), .A1(ori_ori_n34_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n52_));
  INV        o036(.A(x2), .Y(ori_ori_n53_));
  NO2        o037(.A(ori_ori_n53_), .B(ori_ori_n17_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n42_), .B(ori_ori_n18_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n55_), .B(ori_ori_n54_), .Y(ori_ori_n56_));
  OAI210     o040(.A0(ori_ori_n52_), .A1(ori_ori_n31_), .B0(ori_ori_n56_), .Y(ori_ori_n57_));
  NO3        o041(.A(ori_ori_n57_), .B(ori_ori_n50_), .C(ori_ori_n40_), .Y(ori01));
  NA2        o042(.A(x8), .B(x7), .Y(ori_ori_n59_));
  NA2        o043(.A(ori_ori_n42_), .B(x1), .Y(ori_ori_n60_));
  INV        o044(.A(x9), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n61_), .B(ori_ori_n35_), .Y(ori_ori_n62_));
  INV        o046(.A(ori_ori_n62_), .Y(ori_ori_n63_));
  NO3        o047(.A(ori_ori_n63_), .B(ori_ori_n60_), .C(ori_ori_n59_), .Y(ori_ori_n64_));
  NO2        o048(.A(x7), .B(x6), .Y(ori_ori_n65_));
  NO2        o049(.A(ori_ori_n60_), .B(x5), .Y(ori_ori_n66_));
  NO2        o050(.A(x8), .B(x2), .Y(ori_ori_n67_));
  INV        o051(.A(ori_ori_n67_), .Y(ori_ori_n68_));
  AN2        o052(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n43_), .A1(ori_ori_n25_), .B0(ori_ori_n53_), .Y(ori_ori_n70_));
  OAI210     o054(.A0(ori_ori_n55_), .A1(ori_ori_n20_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  NO2        o055(.A(ori_ori_n71_), .B(ori_ori_n69_), .Y(ori_ori_n72_));
  OAI210     o056(.A0(ori_ori_n72_), .A1(ori_ori_n64_), .B0(x4), .Y(ori_ori_n73_));
  NA2        o057(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n74_));
  OAI210     o058(.A0(ori_ori_n74_), .A1(ori_ori_n55_), .B0(x0), .Y(ori_ori_n75_));
  NA2        o059(.A(x5), .B(x3), .Y(ori_ori_n76_));
  NO2        o060(.A(x8), .B(x6), .Y(ori_ori_n77_));
  NO4        o061(.A(ori_ori_n77_), .B(ori_ori_n76_), .C(ori_ori_n65_), .D(ori_ori_n53_), .Y(ori_ori_n78_));
  NAi21      o062(.An(x4), .B(x3), .Y(ori_ori_n79_));
  INV        o063(.A(ori_ori_n79_), .Y(ori_ori_n80_));
  NO2        o064(.A(ori_ori_n80_), .B(ori_ori_n22_), .Y(ori_ori_n81_));
  NO2        o065(.A(x4), .B(x2), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n82_), .B(x3), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n81_), .C(ori_ori_n18_), .Y(ori_ori_n84_));
  NO3        o068(.A(ori_ori_n84_), .B(ori_ori_n78_), .C(ori_ori_n75_), .Y(ori_ori_n85_));
  NA2        o069(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n86_));
  NO2        o070(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n87_));
  INV        o071(.A(x8), .Y(ori_ori_n88_));
  NA2        o072(.A(x2), .B(x1), .Y(ori_ori_n89_));
  INV        o073(.A(ori_ori_n87_), .Y(ori_ori_n90_));
  NO2        o074(.A(ori_ori_n90_), .B(ori_ori_n26_), .Y(ori_ori_n91_));
  AOI210     o075(.A0(ori_ori_n55_), .A1(ori_ori_n25_), .B0(ori_ori_n53_), .Y(ori_ori_n92_));
  OAI210     o076(.A0(ori_ori_n44_), .A1(ori_ori_n36_), .B0(ori_ori_n47_), .Y(ori_ori_n93_));
  NO3        o077(.A(ori_ori_n93_), .B(ori_ori_n92_), .C(ori_ori_n91_), .Y(ori_ori_n94_));
  NA2        o078(.A(x4), .B(ori_ori_n42_), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n47_), .B(ori_ori_n53_), .Y(ori_ori_n96_));
  OAI210     o080(.A0(ori_ori_n96_), .A1(ori_ori_n42_), .B0(ori_ori_n18_), .Y(ori_ori_n97_));
  AOI210     o081(.A0(ori_ori_n95_), .A1(ori_ori_n51_), .B0(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o082(.A(x3), .B(x2), .Y(ori_ori_n99_));
  NA3        o083(.A(ori_ori_n99_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n100_));
  AOI210     o084(.A0(x8), .A1(x6), .B0(ori_ori_n100_), .Y(ori_ori_n101_));
  NA2        o085(.A(ori_ori_n53_), .B(x1), .Y(ori_ori_n102_));
  OAI210     o086(.A0(ori_ori_n102_), .A1(ori_ori_n39_), .B0(ori_ori_n17_), .Y(ori_ori_n103_));
  NO4        o087(.A(ori_ori_n103_), .B(ori_ori_n101_), .C(ori_ori_n98_), .D(ori_ori_n94_), .Y(ori_ori_n104_));
  AO210      o088(.A0(ori_ori_n85_), .A1(ori_ori_n73_), .B0(ori_ori_n104_), .Y(ori02));
  NO2        o089(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n106_));
  NO2        o090(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n53_), .B(ori_ori_n17_), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n42_), .B(x0), .Y(ori_ori_n109_));
  INV        o093(.A(ori_ori_n109_), .Y(ori_ori_n110_));
  AOI220     o094(.A0(ori_ori_n110_), .A1(ori_ori_n107_), .B0(ori_ori_n106_), .B1(x4), .Y(ori_ori_n111_));
  NO3        o095(.A(ori_ori_n111_), .B(x7), .C(x5), .Y(ori_ori_n112_));
  OR2        o096(.A(x8), .B(x0), .Y(ori_ori_n113_));
  INV        o097(.A(ori_ori_n113_), .Y(ori_ori_n114_));
  NAi21      o098(.An(x2), .B(x8), .Y(ori_ori_n115_));
  NO2        o099(.A(x4), .B(x1), .Y(ori_ori_n116_));
  NA3        o100(.A(ori_ori_n116_), .B(x2), .C(ori_ori_n59_), .Y(ori_ori_n117_));
  NOi21      o101(.An(x0), .B(x1), .Y(ori_ori_n118_));
  NO3        o102(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n119_));
  NOi21      o103(.An(x0), .B(x4), .Y(ori_ori_n120_));
  NAi21      o104(.An(x8), .B(x7), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n121_), .B(ori_ori_n61_), .Y(ori_ori_n122_));
  NA2        o106(.A(ori_ori_n122_), .B(ori_ori_n120_), .Y(ori_ori_n123_));
  AOI210     o107(.A0(ori_ori_n123_), .A1(ori_ori_n117_), .B0(ori_ori_n76_), .Y(ori_ori_n124_));
  NO2        o108(.A(x5), .B(ori_ori_n47_), .Y(ori_ori_n125_));
  NA2        o109(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n126_));
  AOI210     o110(.A0(ori_ori_n126_), .A1(ori_ori_n102_), .B0(ori_ori_n109_), .Y(ori_ori_n127_));
  OAI210     o111(.A0(ori_ori_n127_), .A1(ori_ori_n34_), .B0(ori_ori_n125_), .Y(ori_ori_n128_));
  NAi21      o112(.An(x0), .B(x4), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n129_), .B(x1), .Y(ori_ori_n130_));
  NO2        o114(.A(x7), .B(x0), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n82_), .B(ori_ori_n96_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n132_), .B(x3), .Y(ori_ori_n133_));
  OAI210     o117(.A0(ori_ori_n131_), .A1(ori_ori_n130_), .B0(ori_ori_n133_), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n21_), .B(ori_ori_n42_), .Y(ori_ori_n135_));
  NA2        o119(.A(x5), .B(x0), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n137_));
  NA3        o121(.A(ori_ori_n137_), .B(ori_ori_n136_), .C(ori_ori_n135_), .Y(ori_ori_n138_));
  NA4        o122(.A(ori_ori_n138_), .B(ori_ori_n134_), .C(ori_ori_n128_), .D(ori_ori_n35_), .Y(ori_ori_n139_));
  NO3        o123(.A(ori_ori_n139_), .B(ori_ori_n124_), .C(ori_ori_n112_), .Y(ori_ori_n140_));
  NO3        o124(.A(ori_ori_n76_), .B(ori_ori_n74_), .C(ori_ori_n24_), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n142_));
  NA2        o126(.A(x7), .B(x3), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n95_), .B(x5), .Y(ori_ori_n144_));
  NO2        o128(.A(x9), .B(x7), .Y(ori_ori_n145_));
  NOi21      o129(.An(x8), .B(x0), .Y(ori_ori_n146_));
  OA210      o130(.A0(ori_ori_n145_), .A1(x1), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n42_), .B(x2), .Y(ori_ori_n148_));
  INV        o132(.A(x7), .Y(ori_ori_n149_));
  NA2        o133(.A(ori_ori_n149_), .B(ori_ori_n18_), .Y(ori_ori_n150_));
  AOI220     o134(.A0(ori_ori_n150_), .A1(ori_ori_n148_), .B0(ori_ori_n106_), .B1(ori_ori_n37_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n152_), .B(ori_ori_n120_), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n153_), .B(ori_ori_n151_), .Y(ori_ori_n154_));
  AOI210     o138(.A0(ori_ori_n147_), .A1(ori_ori_n144_), .B0(ori_ori_n154_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n143_), .A1(ori_ori_n49_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o140(.A(x5), .B(x1), .Y(ori_ori_n157_));
  INV        o141(.A(ori_ori_n157_), .Y(ori_ori_n158_));
  AOI210     o142(.A0(ori_ori_n158_), .A1(ori_ori_n120_), .B0(ori_ori_n35_), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n61_), .B(ori_ori_n88_), .Y(ori_ori_n160_));
  NAi21      o144(.An(x2), .B(x7), .Y(ori_ori_n161_));
  NO3        o145(.A(ori_ori_n161_), .B(ori_ori_n160_), .C(ori_ori_n47_), .Y(ori_ori_n162_));
  NA2        o146(.A(ori_ori_n162_), .B(ori_ori_n66_), .Y(ori_ori_n163_));
  NAi31      o147(.An(ori_ori_n76_), .B(ori_ori_n37_), .C(ori_ori_n34_), .Y(ori_ori_n164_));
  NA3        o148(.A(ori_ori_n164_), .B(ori_ori_n163_), .C(ori_ori_n159_), .Y(ori_ori_n165_));
  NO3        o149(.A(ori_ori_n165_), .B(ori_ori_n156_), .C(ori_ori_n141_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n166_), .B(ori_ori_n140_), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n136_), .B(ori_ori_n132_), .Y(ori_ori_n168_));
  NA2        o152(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n169_));
  NA2        o153(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n170_));
  NA3        o154(.A(ori_ori_n170_), .B(ori_ori_n169_), .C(ori_ori_n24_), .Y(ori_ori_n171_));
  AN2        o155(.A(ori_ori_n171_), .B(ori_ori_n137_), .Y(ori_ori_n172_));
  NA2        o156(.A(x8), .B(x0), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n149_), .B(ori_ori_n25_), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n118_), .B(x4), .Y(ori_ori_n175_));
  NA2        o159(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  AOI210     o160(.A0(ori_ori_n173_), .A1(ori_ori_n126_), .B0(ori_ori_n176_), .Y(ori_ori_n177_));
  NA2        o161(.A(x2), .B(x0), .Y(ori_ori_n178_));
  NA2        o162(.A(x4), .B(x1), .Y(ori_ori_n179_));
  NAi21      o163(.An(ori_ori_n116_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NOi31      o164(.An(ori_ori_n180_), .B(ori_ori_n152_), .C(ori_ori_n178_), .Y(ori_ori_n181_));
  NO4        o165(.A(ori_ori_n181_), .B(ori_ori_n177_), .C(ori_ori_n172_), .D(ori_ori_n168_), .Y(ori_ori_n182_));
  NO2        o166(.A(ori_ori_n182_), .B(ori_ori_n42_), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n171_), .B(ori_ori_n74_), .Y(ori_ori_n184_));
  INV        o168(.A(ori_ori_n125_), .Y(ori_ori_n185_));
  NO2        o169(.A(ori_ori_n102_), .B(ori_ori_n17_), .Y(ori_ori_n186_));
  AOI210     o170(.A0(ori_ori_n34_), .A1(ori_ori_n88_), .B0(ori_ori_n186_), .Y(ori_ori_n187_));
  NO3        o171(.A(ori_ori_n187_), .B(ori_ori_n185_), .C(x7), .Y(ori_ori_n188_));
  NA3        o172(.A(ori_ori_n180_), .B(ori_ori_n185_), .C(ori_ori_n41_), .Y(ori_ori_n189_));
  OAI210     o173(.A0(ori_ori_n170_), .A1(ori_ori_n132_), .B0(ori_ori_n189_), .Y(ori_ori_n190_));
  NO3        o174(.A(ori_ori_n190_), .B(ori_ori_n188_), .C(ori_ori_n184_), .Y(ori_ori_n191_));
  NO2        o175(.A(ori_ori_n191_), .B(x3), .Y(ori_ori_n192_));
  NO3        o176(.A(ori_ori_n192_), .B(ori_ori_n183_), .C(ori_ori_n167_), .Y(ori03));
  NO2        o177(.A(ori_ori_n47_), .B(x3), .Y(ori_ori_n194_));
  NO2        o178(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n53_), .B(x1), .Y(ori_ori_n196_));
  NA2        o180(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n197_));
  NO2        o181(.A(ori_ori_n197_), .B(x4), .Y(ori_ori_n198_));
  NO2        o182(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n199_));
  NA2        o183(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n200_), .B(ori_ori_n197_), .Y(ori_ori_n201_));
  NA2        o185(.A(x9), .B(ori_ori_n53_), .Y(ori_ori_n202_));
  NA2        o186(.A(ori_ori_n202_), .B(x4), .Y(ori_ori_n203_));
  NA2        o187(.A(ori_ori_n197_), .B(ori_ori_n79_), .Y(ori_ori_n204_));
  AOI210     o188(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n178_), .Y(ori_ori_n205_));
  AOI220     o189(.A0(ori_ori_n205_), .A1(ori_ori_n204_), .B0(ori_ori_n203_), .B1(ori_ori_n201_), .Y(ori_ori_n206_));
  NO3        o190(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n207_));
  NO2        o191(.A(x5), .B(x1), .Y(ori_ori_n208_));
  NO2        o192(.A(ori_ori_n200_), .B(ori_ori_n169_), .Y(ori_ori_n209_));
  NO3        o193(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n210_));
  NO2        o194(.A(ori_ori_n210_), .B(ori_ori_n209_), .Y(ori_ori_n211_));
  INV        o195(.A(ori_ori_n211_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n212_), .B(ori_ori_n47_), .Y(ori_ori_n213_));
  NA2        o197(.A(ori_ori_n213_), .B(ori_ori_n206_), .Y(ori_ori_n214_));
  NO2        o198(.A(ori_ori_n47_), .B(ori_ori_n42_), .Y(ori_ori_n215_));
  NA2        o199(.A(ori_ori_n215_), .B(ori_ori_n19_), .Y(ori_ori_n216_));
  NO2        o200(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n217_));
  NO2        o201(.A(ori_ori_n217_), .B(x6), .Y(ori_ori_n218_));
  NOi21      o202(.An(ori_ori_n82_), .B(ori_ori_n218_), .Y(ori_ori_n219_));
  NA2        o203(.A(ori_ori_n61_), .B(ori_ori_n88_), .Y(ori_ori_n220_));
  NA3        o204(.A(ori_ori_n220_), .B(ori_ori_n217_), .C(x6), .Y(ori_ori_n221_));
  AOI210     o205(.A0(ori_ori_n221_), .A1(ori_ori_n219_), .B0(ori_ori_n149_), .Y(ori_ori_n222_));
  AO210      o206(.A0(ori_ori_n222_), .A1(ori_ori_n216_), .B0(ori_ori_n174_), .Y(ori_ori_n223_));
  NA2        o207(.A(ori_ori_n42_), .B(ori_ori_n53_), .Y(ori_ori_n224_));
  OAI210     o208(.A0(ori_ori_n224_), .A1(ori_ori_n25_), .B0(ori_ori_n170_), .Y(ori_ori_n225_));
  NO2        o209(.A(ori_ori_n179_), .B(x6), .Y(ori_ori_n226_));
  AOI220     o210(.A0(ori_ori_n226_), .A1(ori_ori_n225_), .B0(ori_ori_n137_), .B1(ori_ori_n87_), .Y(ori_ori_n227_));
  NA2        o211(.A(x6), .B(ori_ori_n47_), .Y(ori_ori_n228_));
  OAI210     o212(.A0(ori_ori_n114_), .A1(ori_ori_n77_), .B0(x4), .Y(ori_ori_n229_));
  AOI210     o213(.A0(ori_ori_n229_), .A1(ori_ori_n228_), .B0(ori_ori_n76_), .Y(ori_ori_n230_));
  NO2        o214(.A(ori_ori_n61_), .B(x6), .Y(ori_ori_n231_));
  NO2        o215(.A(ori_ori_n157_), .B(ori_ori_n42_), .Y(ori_ori_n232_));
  OAI210     o216(.A0(ori_ori_n232_), .A1(ori_ori_n209_), .B0(ori_ori_n231_), .Y(ori_ori_n233_));
  NA2        o217(.A(ori_ori_n195_), .B(ori_ori_n130_), .Y(ori_ori_n234_));
  NA3        o218(.A(ori_ori_n200_), .B(ori_ori_n125_), .C(x6), .Y(ori_ori_n235_));
  OAI210     o219(.A0(ori_ori_n88_), .A1(ori_ori_n35_), .B0(ori_ori_n66_), .Y(ori_ori_n236_));
  NA4        o220(.A(ori_ori_n236_), .B(ori_ori_n235_), .C(ori_ori_n234_), .D(ori_ori_n233_), .Y(ori_ori_n237_));
  OAI210     o221(.A0(ori_ori_n237_), .A1(ori_ori_n230_), .B0(x2), .Y(ori_ori_n238_));
  NA3        o222(.A(ori_ori_n238_), .B(ori_ori_n227_), .C(ori_ori_n223_), .Y(ori_ori_n239_));
  AOI210     o223(.A0(ori_ori_n214_), .A1(x8), .B0(ori_ori_n239_), .Y(ori_ori_n240_));
  NO2        o224(.A(ori_ori_n88_), .B(x3), .Y(ori_ori_n241_));
  NA2        o225(.A(ori_ori_n241_), .B(ori_ori_n198_), .Y(ori_ori_n242_));
  NO2        o226(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n243_));
  AOI210     o227(.A0(ori_ori_n218_), .A1(ori_ori_n152_), .B0(ori_ori_n243_), .Y(ori_ori_n244_));
  AOI210     o228(.A0(ori_ori_n244_), .A1(ori_ori_n242_), .B0(x2), .Y(ori_ori_n245_));
  NO2        o229(.A(x4), .B(ori_ori_n53_), .Y(ori_ori_n246_));
  AOI220     o230(.A0(ori_ori_n198_), .A1(ori_ori_n186_), .B0(ori_ori_n246_), .B1(ori_ori_n66_), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n61_), .B(x6), .Y(ori_ori_n248_));
  NA3        o232(.A(ori_ori_n25_), .B(x3), .C(x2), .Y(ori_ori_n249_));
  AOI210     o233(.A0(ori_ori_n249_), .A1(ori_ori_n136_), .B0(ori_ori_n248_), .Y(ori_ori_n250_));
  NA2        o234(.A(ori_ori_n42_), .B(ori_ori_n17_), .Y(ori_ori_n251_));
  NO2        o235(.A(ori_ori_n251_), .B(ori_ori_n25_), .Y(ori_ori_n252_));
  OAI210     o236(.A0(ori_ori_n252_), .A1(ori_ori_n250_), .B0(ori_ori_n116_), .Y(ori_ori_n253_));
  NA2        o237(.A(ori_ori_n200_), .B(x6), .Y(ori_ori_n254_));
  NO2        o238(.A(ori_ori_n200_), .B(x6), .Y(ori_ori_n255_));
  NAi21      o239(.An(ori_ori_n160_), .B(ori_ori_n255_), .Y(ori_ori_n256_));
  NA3        o240(.A(ori_ori_n256_), .B(ori_ori_n254_), .C(ori_ori_n142_), .Y(ori_ori_n257_));
  NA4        o241(.A(ori_ori_n257_), .B(ori_ori_n253_), .C(ori_ori_n247_), .D(ori_ori_n149_), .Y(ori_ori_n258_));
  NA2        o242(.A(ori_ori_n195_), .B(ori_ori_n217_), .Y(ori_ori_n259_));
  NO2        o243(.A(x9), .B(x6), .Y(ori_ori_n260_));
  NO2        o244(.A(ori_ori_n136_), .B(ori_ori_n18_), .Y(ori_ori_n261_));
  NAi21      o245(.An(ori_ori_n261_), .B(ori_ori_n249_), .Y(ori_ori_n262_));
  NAi21      o246(.An(x1), .B(x4), .Y(ori_ori_n263_));
  AOI210     o247(.A0(x3), .A1(x2), .B0(ori_ori_n47_), .Y(ori_ori_n264_));
  OAI210     o248(.A0(ori_ori_n136_), .A1(x3), .B0(ori_ori_n264_), .Y(ori_ori_n265_));
  AOI220     o249(.A0(ori_ori_n265_), .A1(ori_ori_n263_), .B0(ori_ori_n262_), .B1(ori_ori_n260_), .Y(ori_ori_n266_));
  NA2        o250(.A(ori_ori_n266_), .B(ori_ori_n259_), .Y(ori_ori_n267_));
  NA2        o251(.A(ori_ori_n61_), .B(x2), .Y(ori_ori_n268_));
  NO2        o252(.A(ori_ori_n268_), .B(ori_ori_n259_), .Y(ori_ori_n269_));
  NA2        o253(.A(x6), .B(x2), .Y(ori_ori_n270_));
  NO2        o254(.A(ori_ori_n175_), .B(ori_ori_n45_), .Y(ori_ori_n271_));
  OAI210     o255(.A0(ori_ori_n271_), .A1(ori_ori_n269_), .B0(ori_ori_n267_), .Y(ori_ori_n272_));
  NO2        o256(.A(x3), .B(ori_ori_n197_), .Y(ori_ori_n273_));
  NA2        o257(.A(x4), .B(x0), .Y(ori_ori_n274_));
  NA2        o258(.A(ori_ori_n273_), .B(ori_ori_n41_), .Y(ori_ori_n275_));
  AOI210     o259(.A0(ori_ori_n275_), .A1(ori_ori_n272_), .B0(x8), .Y(ori_ori_n276_));
  INV        o260(.A(ori_ori_n248_), .Y(ori_ori_n277_));
  OAI210     o261(.A0(ori_ori_n261_), .A1(ori_ori_n208_), .B0(ori_ori_n277_), .Y(ori_ori_n278_));
  INV        o262(.A(ori_ori_n173_), .Y(ori_ori_n279_));
  OAI210     o263(.A0(ori_ori_n279_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n280_));
  AOI210     o264(.A0(ori_ori_n280_), .A1(ori_ori_n278_), .B0(ori_ori_n224_), .Y(ori_ori_n281_));
  NO4        o265(.A(ori_ori_n281_), .B(ori_ori_n276_), .C(ori_ori_n258_), .D(ori_ori_n245_), .Y(ori_ori_n282_));
  NO2        o266(.A(ori_ori_n160_), .B(x1), .Y(ori_ori_n283_));
  NO3        o267(.A(ori_ori_n283_), .B(x3), .C(ori_ori_n35_), .Y(ori_ori_n284_));
  OAI210     o268(.A0(ori_ori_n284_), .A1(ori_ori_n255_), .B0(x2), .Y(ori_ori_n285_));
  OAI210     o269(.A0(ori_ori_n279_), .A1(x6), .B0(ori_ori_n43_), .Y(ori_ori_n286_));
  AOI210     o270(.A0(ori_ori_n286_), .A1(ori_ori_n285_), .B0(ori_ori_n185_), .Y(ori_ori_n287_));
  NOi21      o271(.An(ori_ori_n270_), .B(ori_ori_n17_), .Y(ori_ori_n288_));
  NA3        o272(.A(ori_ori_n288_), .B(ori_ori_n208_), .C(ori_ori_n39_), .Y(ori_ori_n289_));
  AOI210     o273(.A0(ori_ori_n35_), .A1(ori_ori_n53_), .B0(x0), .Y(ori_ori_n290_));
  NA3        o274(.A(ori_ori_n290_), .B(ori_ori_n158_), .C(ori_ori_n31_), .Y(ori_ori_n291_));
  NA2        o275(.A(x3), .B(x2), .Y(ori_ori_n292_));
  AOI220     o276(.A0(ori_ori_n292_), .A1(ori_ori_n224_), .B0(ori_ori_n291_), .B1(ori_ori_n289_), .Y(ori_ori_n293_));
  NAi21      o277(.An(x4), .B(x0), .Y(ori_ori_n294_));
  NO3        o278(.A(ori_ori_n294_), .B(ori_ori_n43_), .C(x2), .Y(ori_ori_n295_));
  OAI210     o279(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n295_), .Y(ori_ori_n296_));
  OAI220     o280(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n297_));
  NO2        o281(.A(x9), .B(x8), .Y(ori_ori_n298_));
  NA3        o282(.A(ori_ori_n298_), .B(ori_ori_n35_), .C(ori_ori_n53_), .Y(ori_ori_n299_));
  OAI210     o283(.A0(ori_ori_n290_), .A1(ori_ori_n288_), .B0(ori_ori_n299_), .Y(ori_ori_n300_));
  AOI220     o284(.A0(ori_ori_n300_), .A1(ori_ori_n80_), .B0(ori_ori_n297_), .B1(ori_ori_n30_), .Y(ori_ori_n301_));
  AOI210     o285(.A0(ori_ori_n301_), .A1(ori_ori_n296_), .B0(ori_ori_n25_), .Y(ori_ori_n302_));
  NA3        o286(.A(ori_ori_n35_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n303_));
  OAI210     o287(.A0(ori_ori_n290_), .A1(ori_ori_n288_), .B0(ori_ori_n303_), .Y(ori_ori_n304_));
  INV        o288(.A(ori_ori_n209_), .Y(ori_ori_n305_));
  NA2        o289(.A(ori_ori_n35_), .B(ori_ori_n42_), .Y(ori_ori_n306_));
  OR2        o290(.A(ori_ori_n306_), .B(ori_ori_n274_), .Y(ori_ori_n307_));
  OAI220     o291(.A0(ori_ori_n307_), .A1(ori_ori_n157_), .B0(ori_ori_n228_), .B1(ori_ori_n305_), .Y(ori_ori_n308_));
  AO210      o292(.A0(ori_ori_n304_), .A1(ori_ori_n144_), .B0(ori_ori_n308_), .Y(ori_ori_n309_));
  NO4        o293(.A(ori_ori_n309_), .B(ori_ori_n302_), .C(ori_ori_n293_), .D(ori_ori_n287_), .Y(ori_ori_n310_));
  OAI210     o294(.A0(ori_ori_n282_), .A1(ori_ori_n240_), .B0(ori_ori_n310_), .Y(ori04));
  NO2        o295(.A(x2), .B(x1), .Y(ori_ori_n312_));
  OAI210     o296(.A0(ori_ori_n251_), .A1(ori_ori_n312_), .B0(ori_ori_n35_), .Y(ori_ori_n313_));
  NO2        o297(.A(ori_ori_n312_), .B(ori_ori_n294_), .Y(ori_ori_n314_));
  AOI210     o298(.A0(ori_ori_n61_), .A1(x4), .B0(ori_ori_n108_), .Y(ori_ori_n315_));
  OAI210     o299(.A0(ori_ori_n315_), .A1(ori_ori_n314_), .B0(ori_ori_n241_), .Y(ori_ori_n316_));
  NO2        o300(.A(ori_ori_n268_), .B(ori_ori_n86_), .Y(ori_ori_n317_));
  NO2        o301(.A(ori_ori_n317_), .B(ori_ori_n35_), .Y(ori_ori_n318_));
  NO2        o302(.A(ori_ori_n292_), .B(ori_ori_n199_), .Y(ori_ori_n319_));
  NA2        o303(.A(x9), .B(x0), .Y(ori_ori_n320_));
  AOI210     o304(.A0(ori_ori_n86_), .A1(ori_ori_n74_), .B0(ori_ori_n320_), .Y(ori_ori_n321_));
  OAI210     o305(.A0(ori_ori_n321_), .A1(ori_ori_n319_), .B0(ori_ori_n88_), .Y(ori_ori_n322_));
  NA3        o306(.A(ori_ori_n322_), .B(ori_ori_n318_), .C(ori_ori_n316_), .Y(ori_ori_n323_));
  NA2        o307(.A(ori_ori_n323_), .B(ori_ori_n313_), .Y(ori_ori_n324_));
  NO2        o308(.A(ori_ori_n202_), .B(ori_ori_n109_), .Y(ori_ori_n325_));
  NO3        o309(.A(ori_ori_n248_), .B(ori_ori_n115_), .C(ori_ori_n18_), .Y(ori_ori_n326_));
  NO2        o310(.A(ori_ori_n326_), .B(ori_ori_n325_), .Y(ori_ori_n327_));
  OAI210     o311(.A0(ori_ori_n113_), .A1(ori_ori_n102_), .B0(ori_ori_n173_), .Y(ori_ori_n328_));
  NA3        o312(.A(ori_ori_n328_), .B(x6), .C(x3), .Y(ori_ori_n329_));
  NOi21      o313(.An(ori_ori_n146_), .B(ori_ori_n126_), .Y(ori_ori_n330_));
  AOI210     o314(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n331_));
  OAI220     o315(.A0(ori_ori_n331_), .A1(ori_ori_n306_), .B0(ori_ori_n268_), .B1(ori_ori_n303_), .Y(ori_ori_n332_));
  AOI210     o316(.A0(ori_ori_n330_), .A1(ori_ori_n62_), .B0(ori_ori_n332_), .Y(ori_ori_n333_));
  NA2        o317(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n334_));
  OAI210     o318(.A0(ori_ori_n102_), .A1(ori_ori_n17_), .B0(ori_ori_n334_), .Y(ori_ori_n335_));
  AOI220     o319(.A0(ori_ori_n335_), .A1(ori_ori_n77_), .B0(ori_ori_n317_), .B1(ori_ori_n88_), .Y(ori_ori_n336_));
  NA4        o320(.A(ori_ori_n336_), .B(ori_ori_n333_), .C(ori_ori_n329_), .D(ori_ori_n327_), .Y(ori_ori_n337_));
  OAI210     o321(.A0(ori_ori_n107_), .A1(x3), .B0(ori_ori_n295_), .Y(ori_ori_n338_));
  NA2        o322(.A(ori_ori_n207_), .B(ori_ori_n82_), .Y(ori_ori_n339_));
  NA3        o323(.A(ori_ori_n339_), .B(ori_ori_n338_), .C(ori_ori_n149_), .Y(ori_ori_n340_));
  AOI210     o324(.A0(ori_ori_n337_), .A1(x4), .B0(ori_ori_n340_), .Y(ori_ori_n341_));
  NA3        o325(.A(ori_ori_n314_), .B(ori_ori_n202_), .C(ori_ori_n88_), .Y(ori_ori_n342_));
  NOi21      o326(.An(x4), .B(x0), .Y(ori_ori_n343_));
  XO2        o327(.A(x4), .B(x0), .Y(ori_ori_n344_));
  INV        o328(.A(ori_ori_n263_), .Y(ori_ori_n345_));
  AOI220     o329(.A0(ori_ori_n345_), .A1(x8), .B0(ori_ori_n343_), .B1(ori_ori_n89_), .Y(ori_ori_n346_));
  AOI210     o330(.A0(ori_ori_n346_), .A1(ori_ori_n342_), .B0(x3), .Y(ori_ori_n347_));
  INV        o331(.A(ori_ori_n89_), .Y(ori_ori_n348_));
  NO2        o332(.A(ori_ori_n88_), .B(x4), .Y(ori_ori_n349_));
  AOI220     o333(.A0(ori_ori_n349_), .A1(ori_ori_n43_), .B0(ori_ori_n120_), .B1(ori_ori_n348_), .Y(ori_ori_n350_));
  NO3        o334(.A(ori_ori_n344_), .B(ori_ori_n160_), .C(x2), .Y(ori_ori_n351_));
  NO3        o335(.A(ori_ori_n220_), .B(ori_ori_n28_), .C(ori_ori_n24_), .Y(ori_ori_n352_));
  NO2        o336(.A(ori_ori_n352_), .B(ori_ori_n351_), .Y(ori_ori_n353_));
  NA4        o337(.A(ori_ori_n353_), .B(ori_ori_n350_), .C(ori_ori_n216_), .D(x6), .Y(ori_ori_n354_));
  OAI220     o338(.A0(ori_ori_n294_), .A1(ori_ori_n86_), .B0(ori_ori_n178_), .B1(ori_ori_n88_), .Y(ori_ori_n355_));
  NO2        o339(.A(ori_ori_n42_), .B(x0), .Y(ori_ori_n356_));
  OR2        o340(.A(ori_ori_n349_), .B(ori_ori_n356_), .Y(ori_ori_n357_));
  NO2        o341(.A(ori_ori_n146_), .B(ori_ori_n102_), .Y(ori_ori_n358_));
  AOI220     o342(.A0(ori_ori_n358_), .A1(ori_ori_n357_), .B0(ori_ori_n355_), .B1(ori_ori_n60_), .Y(ori_ori_n359_));
  NO2        o343(.A(ori_ori_n146_), .B(ori_ori_n79_), .Y(ori_ori_n360_));
  NO2        o344(.A(ori_ori_n34_), .B(x2), .Y(ori_ori_n361_));
  NOi21      o345(.An(ori_ori_n116_), .B(ori_ori_n27_), .Y(ori_ori_n362_));
  AOI210     o346(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n362_), .Y(ori_ori_n363_));
  OAI210     o347(.A0(ori_ori_n359_), .A1(ori_ori_n61_), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  OAI220     o348(.A0(ori_ori_n364_), .A1(x6), .B0(ori_ori_n354_), .B1(ori_ori_n347_), .Y(ori_ori_n365_));
  OAI210     o349(.A0(ori_ori_n62_), .A1(ori_ori_n47_), .B0(ori_ori_n41_), .Y(ori_ori_n366_));
  OAI210     o350(.A0(ori_ori_n366_), .A1(ori_ori_n88_), .B0(ori_ori_n307_), .Y(ori_ori_n367_));
  AOI210     o351(.A0(ori_ori_n367_), .A1(ori_ori_n18_), .B0(ori_ori_n149_), .Y(ori_ori_n368_));
  AO220      o352(.A0(ori_ori_n368_), .A1(ori_ori_n365_), .B0(ori_ori_n341_), .B1(ori_ori_n324_), .Y(ori_ori_n369_));
  NA2        o353(.A(ori_ori_n361_), .B(x6), .Y(ori_ori_n370_));
  AOI210     o354(.A0(x6), .A1(x1), .B0(ori_ori_n148_), .Y(ori_ori_n371_));
  NA2        o355(.A(ori_ori_n349_), .B(x0), .Y(ori_ori_n372_));
  NA2        o356(.A(ori_ori_n82_), .B(x6), .Y(ori_ori_n373_));
  OAI210     o357(.A0(ori_ori_n372_), .A1(ori_ori_n371_), .B0(ori_ori_n373_), .Y(ori_ori_n374_));
  AOI220     o358(.A0(ori_ori_n374_), .A1(ori_ori_n370_), .B0(ori_ori_n210_), .B1(ori_ori_n48_), .Y(ori_ori_n375_));
  NA2        o359(.A(ori_ori_n375_), .B(ori_ori_n369_), .Y(ori_ori_n376_));
  AOI210     o360(.A0(ori_ori_n196_), .A1(x8), .B0(ori_ori_n107_), .Y(ori_ori_n377_));
  NA2        o361(.A(ori_ori_n377_), .B(ori_ori_n334_), .Y(ori_ori_n378_));
  NA3        o362(.A(ori_ori_n378_), .B(ori_ori_n194_), .C(ori_ori_n149_), .Y(ori_ori_n379_));
  NA3        o363(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n380_));
  NA2        o364(.A(ori_ori_n215_), .B(x0), .Y(ori_ori_n381_));
  OAI220     o365(.A0(ori_ori_n381_), .A1(ori_ori_n202_), .B0(ori_ori_n380_), .B1(ori_ori_n348_), .Y(ori_ori_n382_));
  INV        o366(.A(ori_ori_n382_), .Y(ori_ori_n383_));
  AOI210     o367(.A0(ori_ori_n383_), .A1(ori_ori_n379_), .B0(ori_ori_n25_), .Y(ori_ori_n384_));
  OAI210     o368(.A0(ori_ori_n194_), .A1(ori_ori_n67_), .B0(ori_ori_n199_), .Y(ori_ori_n385_));
  NA3        o369(.A(ori_ori_n196_), .B(ori_ori_n217_), .C(x8), .Y(ori_ori_n386_));
  AOI210     o370(.A0(ori_ori_n386_), .A1(ori_ori_n385_), .B0(ori_ori_n25_), .Y(ori_ori_n387_));
  AOI210     o371(.A0(ori_ori_n115_), .A1(ori_ori_n113_), .B0(ori_ori_n41_), .Y(ori_ori_n388_));
  NOi31      o372(.An(ori_ori_n388_), .B(ori_ori_n356_), .C(ori_ori_n179_), .Y(ori_ori_n389_));
  OAI210     o373(.A0(ori_ori_n389_), .A1(ori_ori_n387_), .B0(ori_ori_n145_), .Y(ori_ori_n390_));
  NAi31      o374(.An(ori_ori_n49_), .B(ori_ori_n283_), .C(ori_ori_n174_), .Y(ori_ori_n391_));
  NA2        o375(.A(ori_ori_n391_), .B(ori_ori_n390_), .Y(ori_ori_n392_));
  OAI210     o376(.A0(ori_ori_n392_), .A1(ori_ori_n384_), .B0(x6), .Y(ori_ori_n393_));
  OAI210     o377(.A0(ori_ori_n160_), .A1(ori_ori_n47_), .B0(ori_ori_n131_), .Y(ori_ori_n394_));
  NA3        o378(.A(ori_ori_n54_), .B(ori_ori_n37_), .C(ori_ori_n30_), .Y(ori_ori_n395_));
  AOI220     o379(.A0(ori_ori_n395_), .A1(ori_ori_n394_), .B0(ori_ori_n39_), .B1(ori_ori_n31_), .Y(ori_ori_n396_));
  NO2        o380(.A(ori_ori_n149_), .B(x0), .Y(ori_ori_n397_));
  AOI220     o381(.A0(ori_ori_n397_), .A1(ori_ori_n215_), .B0(ori_ori_n194_), .B1(ori_ori_n149_), .Y(ori_ori_n398_));
  AOI210     o382(.A0(ori_ori_n122_), .A1(ori_ori_n246_), .B0(x1), .Y(ori_ori_n399_));
  OAI210     o383(.A0(ori_ori_n398_), .A1(x8), .B0(ori_ori_n399_), .Y(ori_ori_n400_));
  NAi31      o384(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n401_));
  OAI210     o385(.A0(ori_ori_n401_), .A1(x4), .B0(ori_ori_n161_), .Y(ori_ori_n402_));
  NA3        o386(.A(ori_ori_n402_), .B(ori_ori_n143_), .C(x9), .Y(ori_ori_n403_));
  NO4        o387(.A(ori_ori_n121_), .B(ori_ori_n294_), .C(x9), .D(x2), .Y(ori_ori_n404_));
  NOi21      o388(.An(ori_ori_n119_), .B(ori_ori_n178_), .Y(ori_ori_n405_));
  NO3        o389(.A(ori_ori_n405_), .B(ori_ori_n404_), .C(ori_ori_n18_), .Y(ori_ori_n406_));
  NO3        o390(.A(x9), .B(ori_ori_n149_), .C(x0), .Y(ori_ori_n407_));
  AOI220     o391(.A0(ori_ori_n407_), .A1(ori_ori_n241_), .B0(ori_ori_n360_), .B1(ori_ori_n149_), .Y(ori_ori_n408_));
  NA4        o392(.A(ori_ori_n408_), .B(ori_ori_n406_), .C(ori_ori_n403_), .D(ori_ori_n49_), .Y(ori_ori_n409_));
  OAI210     o393(.A0(ori_ori_n400_), .A1(ori_ori_n396_), .B0(ori_ori_n409_), .Y(ori_ori_n410_));
  NOi31      o394(.An(ori_ori_n397_), .B(ori_ori_n31_), .C(x8), .Y(ori_ori_n411_));
  AOI210     o395(.A0(ori_ori_n37_), .A1(x9), .B0(ori_ori_n129_), .Y(ori_ori_n412_));
  NO3        o396(.A(ori_ori_n412_), .B(ori_ori_n119_), .C(ori_ori_n42_), .Y(ori_ori_n413_));
  NOi31      o397(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n414_));
  AOI210     o398(.A0(ori_ori_n263_), .A1(ori_ori_n59_), .B0(ori_ori_n118_), .Y(ori_ori_n415_));
  NO2        o399(.A(ori_ori_n415_), .B(x3), .Y(ori_ori_n416_));
  NO3        o400(.A(ori_ori_n416_), .B(ori_ori_n413_), .C(x2), .Y(ori_ori_n417_));
  OAI220     o401(.A0(ori_ori_n344_), .A1(ori_ori_n298_), .B0(ori_ori_n294_), .B1(ori_ori_n42_), .Y(ori_ori_n418_));
  AOI210     o402(.A0(x9), .A1(ori_ori_n47_), .B0(ori_ori_n380_), .Y(ori_ori_n419_));
  AOI220     o403(.A0(ori_ori_n419_), .A1(ori_ori_n88_), .B0(ori_ori_n418_), .B1(ori_ori_n149_), .Y(ori_ori_n420_));
  NO2        o404(.A(ori_ori_n420_), .B(ori_ori_n53_), .Y(ori_ori_n421_));
  NO3        o405(.A(ori_ori_n421_), .B(ori_ori_n417_), .C(ori_ori_n411_), .Y(ori_ori_n422_));
  AOI210     o406(.A0(ori_ori_n422_), .A1(ori_ori_n410_), .B0(ori_ori_n25_), .Y(ori_ori_n423_));
  NA4        o407(.A(ori_ori_n30_), .B(ori_ori_n88_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n424_));
  NO3        o408(.A(ori_ori_n61_), .B(x4), .C(x1), .Y(ori_ori_n425_));
  NO3        o409(.A(ori_ori_n67_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n426_));
  AOI220     o410(.A0(ori_ori_n426_), .A1(ori_ori_n264_), .B0(ori_ori_n425_), .B1(ori_ori_n388_), .Y(ori_ori_n427_));
  NO2        o411(.A(ori_ori_n427_), .B(ori_ori_n99_), .Y(ori_ori_n428_));
  NO3        o412(.A(ori_ori_n268_), .B(ori_ori_n173_), .C(ori_ori_n39_), .Y(ori_ori_n429_));
  OAI210     o413(.A0(ori_ori_n429_), .A1(ori_ori_n428_), .B0(x7), .Y(ori_ori_n430_));
  NA2        o414(.A(ori_ori_n220_), .B(x7), .Y(ori_ori_n431_));
  NA3        o415(.A(ori_ori_n431_), .B(ori_ori_n148_), .C(ori_ori_n130_), .Y(ori_ori_n432_));
  NA3        o416(.A(ori_ori_n432_), .B(ori_ori_n430_), .C(ori_ori_n424_), .Y(ori_ori_n433_));
  OAI210     o417(.A0(ori_ori_n433_), .A1(ori_ori_n423_), .B0(ori_ori_n35_), .Y(ori_ori_n434_));
  NO2        o418(.A(ori_ori_n407_), .B(ori_ori_n199_), .Y(ori_ori_n435_));
  NO4        o419(.A(ori_ori_n435_), .B(ori_ori_n76_), .C(x4), .D(ori_ori_n53_), .Y(ori_ori_n436_));
  NA2        o420(.A(ori_ori_n251_), .B(ori_ori_n21_), .Y(ori_ori_n437_));
  NO2        o421(.A(ori_ori_n157_), .B(ori_ori_n131_), .Y(ori_ori_n438_));
  NA2        o422(.A(ori_ori_n438_), .B(ori_ori_n437_), .Y(ori_ori_n439_));
  AOI210     o423(.A0(ori_ori_n439_), .A1(ori_ori_n164_), .B0(ori_ori_n28_), .Y(ori_ori_n440_));
  AOI220     o424(.A0(ori_ori_n356_), .A1(ori_ori_n88_), .B0(ori_ori_n146_), .B1(ori_ori_n196_), .Y(ori_ori_n441_));
  NA3        o425(.A(ori_ori_n441_), .B(ori_ori_n401_), .C(ori_ori_n86_), .Y(ori_ori_n442_));
  NA2        o426(.A(ori_ori_n442_), .B(ori_ori_n174_), .Y(ori_ori_n443_));
  OAI220     o427(.A0(x3), .A1(ori_ori_n68_), .B0(ori_ori_n157_), .B1(ori_ori_n42_), .Y(ori_ori_n444_));
  NA2        o428(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n445_));
  OAI210     o429(.A0(ori_ori_n145_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n446_));
  NO3        o430(.A(ori_ori_n414_), .B(x3), .C(ori_ori_n53_), .Y(ori_ori_n447_));
  NA2        o431(.A(ori_ori_n447_), .B(ori_ori_n446_), .Y(ori_ori_n448_));
  OAI210     o432(.A0(ori_ori_n150_), .A1(ori_ori_n445_), .B0(ori_ori_n448_), .Y(ori_ori_n449_));
  AOI220     o433(.A0(ori_ori_n449_), .A1(x0), .B0(ori_ori_n444_), .B1(ori_ori_n131_), .Y(ori_ori_n450_));
  AOI210     o434(.A0(ori_ori_n450_), .A1(ori_ori_n443_), .B0(ori_ori_n228_), .Y(ori_ori_n451_));
  NO3        o435(.A(ori_ori_n451_), .B(ori_ori_n440_), .C(ori_ori_n436_), .Y(ori_ori_n452_));
  NA3        o436(.A(ori_ori_n452_), .B(ori_ori_n434_), .C(ori_ori_n393_), .Y(ori_ori_n453_));
  AOI210     o437(.A0(ori_ori_n376_), .A1(ori_ori_n25_), .B0(ori_ori_n453_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  INV        m047(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  NO2        m048(.A(x7), .B(x6), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(x8), .B(x2), .Y(mai_mai_n67_));
  INV        m051(.A(mai_mai_n67_), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n68_), .B(x1), .Y(mai_mai_n69_));
  OA210      m053(.A0(mai_mai_n69_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  NAi31      m056(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n73_));
  OAI220     m057(.A0(mai_mai_n73_), .A1(mai_mai_n43_), .B0(mai_mai_n72_), .B1(mai_mai_n70_), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n74_), .B(x4), .Y(mai_mai_n75_));
  NA2        m059(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n76_));
  OAI210     m060(.A0(mai_mai_n76_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n77_));
  NA2        m061(.A(x5), .B(x3), .Y(mai_mai_n78_));
  NO2        m062(.A(x8), .B(x6), .Y(mai_mai_n79_));
  NO4        m063(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(mai_mai_n65_), .D(mai_mai_n54_), .Y(mai_mai_n80_));
  NAi21      m064(.An(x4), .B(x3), .Y(mai_mai_n81_));
  INV        m065(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(mai_mai_n22_), .Y(mai_mai_n83_));
  NO2        m067(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(x3), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n83_), .C(mai_mai_n18_), .Y(mai_mai_n86_));
  NO3        m070(.A(mai_mai_n86_), .B(mai_mai_n80_), .C(mai_mai_n77_), .Y(mai_mai_n87_));
  NO4        m071(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n43_), .D(x1), .Y(mai_mai_n88_));
  NA2        m072(.A(mai_mai_n62_), .B(mai_mai_n48_), .Y(mai_mai_n89_));
  INV        m073(.A(mai_mai_n89_), .Y(mai_mai_n90_));
  OAI210     m074(.A0(mai_mai_n88_), .A1(mai_mai_n66_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  NA2        m075(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n25_), .Y(mai_mai_n93_));
  INV        m077(.A(x8), .Y(mai_mai_n94_));
  NA2        m078(.A(x2), .B(x1), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n97_));
  NO2        m081(.A(mai_mai_n97_), .B(mai_mai_n26_), .Y(mai_mai_n98_));
  AOI210     m082(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n99_));
  OAI210     m083(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n100_));
  NO3        m084(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(mai_mai_n98_), .Y(mai_mai_n101_));
  NA2        m085(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n102_));
  NO2        m086(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n103_));
  OAI210     m087(.A0(mai_mai_n103_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n104_));
  AOI210     m088(.A0(mai_mai_n102_), .A1(mai_mai_n52_), .B0(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m089(.A(x3), .B(x2), .Y(mai_mai_n106_));
  NA3        m090(.A(mai_mai_n106_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n107_));
  AOI210     m091(.A0(x8), .A1(x6), .B0(mai_mai_n107_), .Y(mai_mai_n108_));
  NA2        m092(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n109_));
  OAI210     m093(.A0(mai_mai_n109_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n110_));
  NO4        m094(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n105_), .D(mai_mai_n101_), .Y(mai_mai_n111_));
  AO220      m095(.A0(mai_mai_n111_), .A1(mai_mai_n91_), .B0(mai_mai_n87_), .B1(mai_mai_n75_), .Y(mai02));
  NO2        m096(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n113_));
  NO2        m097(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n114_));
  NA2        m098(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n115_));
  NA2        m099(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n116_));
  OAI210     m100(.A0(mai_mai_n89_), .A1(mai_mai_n115_), .B0(mai_mai_n116_), .Y(mai_mai_n117_));
  AOI220     m101(.A0(mai_mai_n117_), .A1(mai_mai_n114_), .B0(mai_mai_n113_), .B1(x4), .Y(mai_mai_n118_));
  NO3        m102(.A(mai_mai_n118_), .B(x7), .C(x5), .Y(mai_mai_n119_));
  NA2        m103(.A(x9), .B(x2), .Y(mai_mai_n120_));
  OR2        m104(.A(x8), .B(x0), .Y(mai_mai_n121_));
  INV        m105(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  NAi21      m106(.An(x2), .B(x8), .Y(mai_mai_n123_));
  INV        m107(.A(mai_mai_n123_), .Y(mai_mai_n124_));
  OAI220     m108(.A0(mai_mai_n124_), .A1(mai_mai_n122_), .B0(mai_mai_n120_), .B1(x7), .Y(mai_mai_n125_));
  NO2        m109(.A(x4), .B(x1), .Y(mai_mai_n126_));
  NA3        m110(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n60_), .Y(mai_mai_n127_));
  NOi21      m111(.An(x0), .B(x1), .Y(mai_mai_n128_));
  NO3        m112(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n129_));
  NOi21      m113(.An(x0), .B(x4), .Y(mai_mai_n130_));
  NAi21      m114(.An(x8), .B(x7), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n131_), .B(mai_mai_n62_), .Y(mai_mai_n132_));
  AOI220     m116(.A0(mai_mai_n132_), .A1(mai_mai_n130_), .B0(mai_mai_n129_), .B1(mai_mai_n128_), .Y(mai_mai_n133_));
  AOI210     m117(.A0(mai_mai_n133_), .A1(mai_mai_n127_), .B0(mai_mai_n78_), .Y(mai_mai_n134_));
  NO2        m118(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n135_));
  NA2        m119(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n136_));
  AOI210     m120(.A0(mai_mai_n136_), .A1(mai_mai_n109_), .B0(mai_mai_n116_), .Y(mai_mai_n137_));
  OAI210     m121(.A0(mai_mai_n137_), .A1(mai_mai_n35_), .B0(mai_mai_n135_), .Y(mai_mai_n138_));
  NAi21      m122(.An(x0), .B(x4), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n139_), .B(x1), .Y(mai_mai_n140_));
  NO2        m124(.A(x7), .B(x0), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n84_), .B(mai_mai_n103_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n142_), .B(x3), .Y(mai_mai_n143_));
  OAI210     m127(.A0(mai_mai_n141_), .A1(mai_mai_n140_), .B0(mai_mai_n143_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n145_));
  NA2        m129(.A(x5), .B(x0), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n147_));
  NA3        m131(.A(mai_mai_n147_), .B(mai_mai_n146_), .C(mai_mai_n145_), .Y(mai_mai_n148_));
  NA4        m132(.A(mai_mai_n148_), .B(mai_mai_n144_), .C(mai_mai_n138_), .D(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m133(.A(mai_mai_n149_), .B(mai_mai_n134_), .C(mai_mai_n119_), .Y(mai_mai_n150_));
  NO3        m134(.A(mai_mai_n78_), .B(mai_mai_n76_), .C(mai_mai_n24_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n152_));
  AOI220     m136(.A0(mai_mai_n128_), .A1(mai_mai_n152_), .B0(mai_mai_n66_), .B1(mai_mai_n17_), .Y(mai_mai_n153_));
  NO3        m137(.A(mai_mai_n153_), .B(mai_mai_n60_), .C(mai_mai_n62_), .Y(mai_mai_n154_));
  NA2        m138(.A(x7), .B(x3), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n102_), .B(x5), .Y(mai_mai_n156_));
  NO2        m140(.A(x9), .B(x7), .Y(mai_mai_n157_));
  NOi21      m141(.An(x8), .B(x0), .Y(mai_mai_n158_));
  OA210      m142(.A0(mai_mai_n157_), .A1(x1), .B0(mai_mai_n158_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n160_));
  INV        m144(.A(x7), .Y(mai_mai_n161_));
  NA2        m145(.A(mai_mai_n161_), .B(mai_mai_n18_), .Y(mai_mai_n162_));
  AOI220     m146(.A0(mai_mai_n162_), .A1(mai_mai_n160_), .B0(mai_mai_n113_), .B1(mai_mai_n38_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n164_), .B(mai_mai_n130_), .Y(mai_mai_n165_));
  NO2        m149(.A(mai_mai_n165_), .B(mai_mai_n163_), .Y(mai_mai_n166_));
  AOI210     m150(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n166_), .Y(mai_mai_n167_));
  OAI210     m151(.A0(mai_mai_n155_), .A1(mai_mai_n50_), .B0(mai_mai_n167_), .Y(mai_mai_n168_));
  NA2        m152(.A(x5), .B(x1), .Y(mai_mai_n169_));
  INV        m153(.A(mai_mai_n169_), .Y(mai_mai_n170_));
  AOI210     m154(.A0(mai_mai_n170_), .A1(mai_mai_n130_), .B0(mai_mai_n36_), .Y(mai_mai_n171_));
  NAi21      m155(.An(x2), .B(x7), .Y(mai_mai_n172_));
  NO2        m156(.A(mai_mai_n172_), .B(mai_mai_n48_), .Y(mai_mai_n173_));
  NA2        m157(.A(mai_mai_n173_), .B(mai_mai_n66_), .Y(mai_mai_n174_));
  NAi31      m158(.An(mai_mai_n78_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n175_));
  NA3        m159(.A(mai_mai_n175_), .B(mai_mai_n174_), .C(mai_mai_n171_), .Y(mai_mai_n176_));
  NO4        m160(.A(mai_mai_n176_), .B(mai_mai_n168_), .C(mai_mai_n154_), .D(mai_mai_n151_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n177_), .B(mai_mai_n150_), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n146_), .B(mai_mai_n142_), .Y(mai_mai_n179_));
  NA2        m163(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n180_));
  NA2        m164(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n181_));
  NA3        m165(.A(mai_mai_n181_), .B(mai_mai_n180_), .C(mai_mai_n24_), .Y(mai_mai_n182_));
  AN2        m166(.A(mai_mai_n182_), .B(mai_mai_n147_), .Y(mai_mai_n183_));
  NA2        m167(.A(x8), .B(x0), .Y(mai_mai_n184_));
  NO2        m168(.A(mai_mai_n161_), .B(mai_mai_n25_), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n128_), .B(x4), .Y(mai_mai_n186_));
  NA2        m170(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  AOI210     m171(.A0(mai_mai_n184_), .A1(mai_mai_n136_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  NA2        m172(.A(x2), .B(x0), .Y(mai_mai_n189_));
  NA2        m173(.A(x4), .B(x1), .Y(mai_mai_n190_));
  NAi21      m174(.An(mai_mai_n126_), .B(mai_mai_n190_), .Y(mai_mai_n191_));
  NOi31      m175(.An(mai_mai_n191_), .B(mai_mai_n164_), .C(mai_mai_n189_), .Y(mai_mai_n192_));
  NO4        m176(.A(mai_mai_n192_), .B(mai_mai_n188_), .C(mai_mai_n183_), .D(mai_mai_n179_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n193_), .B(mai_mai_n43_), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n182_), .B(mai_mai_n76_), .Y(mai_mai_n195_));
  INV        m179(.A(mai_mai_n135_), .Y(mai_mai_n196_));
  NO2        m180(.A(mai_mai_n109_), .B(mai_mai_n17_), .Y(mai_mai_n197_));
  AOI210     m181(.A0(mai_mai_n35_), .A1(mai_mai_n94_), .B0(mai_mai_n197_), .Y(mai_mai_n198_));
  NO3        m182(.A(mai_mai_n198_), .B(mai_mai_n196_), .C(x7), .Y(mai_mai_n199_));
  NA3        m183(.A(mai_mai_n191_), .B(mai_mai_n196_), .C(mai_mai_n42_), .Y(mai_mai_n200_));
  OAI210     m184(.A0(mai_mai_n181_), .A1(mai_mai_n142_), .B0(mai_mai_n200_), .Y(mai_mai_n201_));
  NO3        m185(.A(mai_mai_n201_), .B(mai_mai_n199_), .C(mai_mai_n195_), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n202_), .B(x3), .Y(mai_mai_n203_));
  NO3        m187(.A(mai_mai_n203_), .B(mai_mai_n194_), .C(mai_mai_n178_), .Y(mai03));
  NO2        m188(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n205_));
  NO2        m189(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n206_));
  INV        m190(.A(mai_mai_n206_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n208_));
  OAI210     m192(.A0(mai_mai_n208_), .A1(mai_mai_n25_), .B0(mai_mai_n63_), .Y(mai_mai_n209_));
  OAI220     m193(.A0(mai_mai_n209_), .A1(mai_mai_n17_), .B0(mai_mai_n207_), .B1(mai_mai_n109_), .Y(mai_mai_n210_));
  NA2        m194(.A(mai_mai_n210_), .B(mai_mai_n205_), .Y(mai_mai_n211_));
  NO2        m195(.A(mai_mai_n78_), .B(x6), .Y(mai_mai_n212_));
  NA2        m196(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n213_));
  NO2        m197(.A(mai_mai_n213_), .B(x4), .Y(mai_mai_n214_));
  NO2        m198(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n215_));
  AO220      m199(.A0(mai_mai_n215_), .A1(mai_mai_n214_), .B0(mai_mai_n212_), .B1(mai_mai_n55_), .Y(mai_mai_n216_));
  NA2        m200(.A(mai_mai_n216_), .B(mai_mai_n62_), .Y(mai_mai_n217_));
  NA2        m201(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n218_));
  NO2        m202(.A(mai_mai_n218_), .B(mai_mai_n213_), .Y(mai_mai_n219_));
  NA2        m203(.A(x9), .B(mai_mai_n54_), .Y(mai_mai_n220_));
  NA2        m204(.A(mai_mai_n220_), .B(x4), .Y(mai_mai_n221_));
  NA2        m205(.A(mai_mai_n213_), .B(mai_mai_n81_), .Y(mai_mai_n222_));
  AOI210     m206(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n189_), .Y(mai_mai_n223_));
  AOI220     m207(.A0(mai_mai_n223_), .A1(mai_mai_n222_), .B0(mai_mai_n221_), .B1(mai_mai_n219_), .Y(mai_mai_n224_));
  NO3        m208(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n225_));
  NO2        m209(.A(x5), .B(x1), .Y(mai_mai_n226_));
  AOI220     m210(.A0(mai_mai_n226_), .A1(mai_mai_n17_), .B0(mai_mai_n106_), .B1(x5), .Y(mai_mai_n227_));
  NO2        m211(.A(mai_mai_n218_), .B(mai_mai_n180_), .Y(mai_mai_n228_));
  NO3        m212(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n229_));
  NO2        m213(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  OAI210     m214(.A0(mai_mai_n227_), .A1(mai_mai_n64_), .B0(mai_mai_n230_), .Y(mai_mai_n231_));
  AOI220     m215(.A0(mai_mai_n231_), .A1(mai_mai_n48_), .B0(mai_mai_n225_), .B1(mai_mai_n135_), .Y(mai_mai_n232_));
  NA4        m216(.A(mai_mai_n232_), .B(mai_mai_n224_), .C(mai_mai_n217_), .D(mai_mai_n211_), .Y(mai_mai_n233_));
  NO2        m217(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n234_));
  NA2        m218(.A(mai_mai_n234_), .B(mai_mai_n19_), .Y(mai_mai_n235_));
  NO2        m219(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n236_));
  NO2        m220(.A(mai_mai_n236_), .B(x6), .Y(mai_mai_n237_));
  NOi21      m221(.An(mai_mai_n84_), .B(mai_mai_n237_), .Y(mai_mai_n238_));
  NA2        m222(.A(mai_mai_n62_), .B(mai_mai_n94_), .Y(mai_mai_n239_));
  NA3        m223(.A(mai_mai_n239_), .B(mai_mai_n236_), .C(x6), .Y(mai_mai_n240_));
  AOI210     m224(.A0(mai_mai_n240_), .A1(mai_mai_n238_), .B0(mai_mai_n161_), .Y(mai_mai_n241_));
  AO210      m225(.A0(mai_mai_n241_), .A1(mai_mai_n235_), .B0(mai_mai_n185_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n243_));
  NA2        m227(.A(mai_mai_n147_), .B(mai_mai_n93_), .Y(mai_mai_n244_));
  NA2        m228(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n245_));
  OAI210     m229(.A0(mai_mai_n122_), .A1(mai_mai_n79_), .B0(x4), .Y(mai_mai_n246_));
  AOI210     m230(.A0(mai_mai_n246_), .A1(mai_mai_n245_), .B0(mai_mai_n78_), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n169_), .B(mai_mai_n43_), .Y(mai_mai_n249_));
  OAI210     m233(.A0(mai_mai_n249_), .A1(mai_mai_n228_), .B0(mai_mai_n248_), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n206_), .B(mai_mai_n140_), .Y(mai_mai_n251_));
  NA3        m235(.A(mai_mai_n218_), .B(mai_mai_n135_), .C(x6), .Y(mai_mai_n252_));
  OAI210     m236(.A0(mai_mai_n94_), .A1(mai_mai_n36_), .B0(mai_mai_n66_), .Y(mai_mai_n253_));
  NA4        m237(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n251_), .D(mai_mai_n250_), .Y(mai_mai_n254_));
  OAI210     m238(.A0(mai_mai_n254_), .A1(mai_mai_n247_), .B0(x2), .Y(mai_mai_n255_));
  NA3        m239(.A(mai_mai_n255_), .B(mai_mai_n244_), .C(mai_mai_n242_), .Y(mai_mai_n256_));
  AOI210     m240(.A0(mai_mai_n233_), .A1(x8), .B0(mai_mai_n256_), .Y(mai_mai_n257_));
  NO2        m241(.A(mai_mai_n94_), .B(x3), .Y(mai_mai_n258_));
  NA2        m242(.A(mai_mai_n258_), .B(mai_mai_n214_), .Y(mai_mai_n259_));
  NO3        m243(.A(mai_mai_n92_), .B(mai_mai_n79_), .C(mai_mai_n25_), .Y(mai_mai_n260_));
  AOI210     m244(.A0(mai_mai_n237_), .A1(mai_mai_n164_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  AOI210     m245(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(x2), .Y(mai_mai_n262_));
  NO2        m246(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n263_));
  AOI220     m247(.A0(mai_mai_n214_), .A1(mai_mai_n197_), .B0(mai_mai_n263_), .B1(mai_mai_n66_), .Y(mai_mai_n264_));
  NA2        m248(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n265_));
  NA2        m249(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n266_));
  NO2        m250(.A(mai_mai_n266_), .B(mai_mai_n25_), .Y(mai_mai_n267_));
  NA2        m251(.A(mai_mai_n267_), .B(mai_mai_n126_), .Y(mai_mai_n268_));
  NA2        m252(.A(mai_mai_n218_), .B(x6), .Y(mai_mai_n269_));
  NO2        m253(.A(mai_mai_n218_), .B(x6), .Y(mai_mai_n270_));
  INV        m254(.A(mai_mai_n270_), .Y(mai_mai_n271_));
  NA3        m255(.A(mai_mai_n271_), .B(mai_mai_n269_), .C(mai_mai_n152_), .Y(mai_mai_n272_));
  NA4        m256(.A(mai_mai_n272_), .B(mai_mai_n268_), .C(mai_mai_n264_), .D(mai_mai_n161_), .Y(mai_mai_n273_));
  NA2        m257(.A(mai_mai_n206_), .B(mai_mai_n236_), .Y(mai_mai_n274_));
  NO2        m258(.A(mai_mai_n146_), .B(mai_mai_n18_), .Y(mai_mai_n275_));
  NAi21      m259(.An(x1), .B(x4), .Y(mai_mai_n276_));
  AOI210     m260(.A0(x3), .A1(x2), .B0(mai_mai_n48_), .Y(mai_mai_n277_));
  OAI210     m261(.A0(mai_mai_n146_), .A1(x3), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  NA2        m262(.A(mai_mai_n278_), .B(mai_mai_n276_), .Y(mai_mai_n279_));
  NA2        m263(.A(mai_mai_n279_), .B(mai_mai_n274_), .Y(mai_mai_n280_));
  NA2        m264(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n281_));
  NO2        m265(.A(mai_mai_n281_), .B(mai_mai_n274_), .Y(mai_mai_n282_));
  NO3        m266(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n283_));
  NA2        m267(.A(mai_mai_n109_), .B(mai_mai_n25_), .Y(mai_mai_n284_));
  NA2        m268(.A(x6), .B(x2), .Y(mai_mai_n285_));
  NO2        m269(.A(mai_mai_n285_), .B(mai_mai_n180_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n284_), .A1(mai_mai_n283_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  OAI220     m271(.A0(mai_mai_n287_), .A1(mai_mai_n43_), .B0(mai_mai_n186_), .B1(mai_mai_n46_), .Y(mai_mai_n288_));
  OAI210     m272(.A0(mai_mai_n288_), .A1(mai_mai_n282_), .B0(mai_mai_n280_), .Y(mai_mai_n289_));
  NA2        m273(.A(x9), .B(mai_mai_n43_), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n290_), .B(mai_mai_n213_), .Y(mai_mai_n291_));
  OR3        m275(.A(mai_mai_n291_), .B(mai_mai_n212_), .C(mai_mai_n156_), .Y(mai_mai_n292_));
  NA2        m276(.A(x4), .B(x0), .Y(mai_mai_n293_));
  NO3        m277(.A(mai_mai_n73_), .B(mai_mai_n293_), .C(x6), .Y(mai_mai_n294_));
  AOI210     m278(.A0(mai_mai_n292_), .A1(mai_mai_n42_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  AOI210     m279(.A0(mai_mai_n295_), .A1(mai_mai_n289_), .B0(x8), .Y(mai_mai_n296_));
  INV        m280(.A(mai_mai_n265_), .Y(mai_mai_n297_));
  OAI210     m281(.A0(mai_mai_n275_), .A1(mai_mai_n226_), .B0(mai_mai_n297_), .Y(mai_mai_n298_));
  INV        m282(.A(mai_mai_n184_), .Y(mai_mai_n299_));
  OAI210     m283(.A0(mai_mai_n299_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n300_));
  AOI210     m284(.A0(mai_mai_n300_), .A1(mai_mai_n298_), .B0(mai_mai_n243_), .Y(mai_mai_n301_));
  NO4        m285(.A(mai_mai_n301_), .B(mai_mai_n296_), .C(mai_mai_n273_), .D(mai_mai_n262_), .Y(mai_mai_n302_));
  INV        m286(.A(x1), .Y(mai_mai_n303_));
  NO3        m287(.A(mai_mai_n303_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n304_));
  OAI210     m288(.A0(mai_mai_n304_), .A1(mai_mai_n270_), .B0(x2), .Y(mai_mai_n305_));
  OAI210     m289(.A0(mai_mai_n299_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n306_));
  AOI210     m290(.A0(mai_mai_n306_), .A1(mai_mai_n305_), .B0(mai_mai_n196_), .Y(mai_mai_n307_));
  NOi21      m291(.An(mai_mai_n285_), .B(mai_mai_n17_), .Y(mai_mai_n308_));
  NA3        m292(.A(mai_mai_n308_), .B(mai_mai_n226_), .C(mai_mai_n40_), .Y(mai_mai_n309_));
  AOI210     m293(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n170_), .C(mai_mai_n32_), .Y(mai_mai_n311_));
  NA2        m295(.A(x3), .B(x2), .Y(mai_mai_n312_));
  AOI220     m296(.A0(mai_mai_n312_), .A1(mai_mai_n243_), .B0(mai_mai_n311_), .B1(mai_mai_n309_), .Y(mai_mai_n313_));
  NAi21      m297(.An(x4), .B(x0), .Y(mai_mai_n314_));
  NO3        m298(.A(mai_mai_n314_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n315_));
  OAI210     m299(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n315_), .Y(mai_mai_n316_));
  OAI220     m300(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n317_));
  NO2        m301(.A(mai_mai_n310_), .B(mai_mai_n308_), .Y(mai_mai_n318_));
  AOI220     m302(.A0(mai_mai_n318_), .A1(mai_mai_n82_), .B0(mai_mai_n317_), .B1(mai_mai_n31_), .Y(mai_mai_n319_));
  AOI210     m303(.A0(mai_mai_n319_), .A1(mai_mai_n316_), .B0(mai_mai_n25_), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n321_));
  OAI210     m305(.A0(mai_mai_n310_), .A1(mai_mai_n308_), .B0(mai_mai_n321_), .Y(mai_mai_n322_));
  INV        m306(.A(mai_mai_n228_), .Y(mai_mai_n323_));
  NA2        m307(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n324_));
  OR2        m308(.A(mai_mai_n324_), .B(mai_mai_n293_), .Y(mai_mai_n325_));
  OAI220     m309(.A0(mai_mai_n325_), .A1(mai_mai_n169_), .B0(mai_mai_n245_), .B1(mai_mai_n323_), .Y(mai_mai_n326_));
  AO210      m310(.A0(mai_mai_n322_), .A1(mai_mai_n156_), .B0(mai_mai_n326_), .Y(mai_mai_n327_));
  NO4        m311(.A(mai_mai_n327_), .B(mai_mai_n320_), .C(mai_mai_n313_), .D(mai_mai_n307_), .Y(mai_mai_n328_));
  OAI210     m312(.A0(mai_mai_n302_), .A1(mai_mai_n257_), .B0(mai_mai_n328_), .Y(mai04));
  OAI210     m313(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n330_));
  NA3        m314(.A(mai_mai_n330_), .B(mai_mai_n283_), .C(mai_mai_n85_), .Y(mai_mai_n331_));
  NO2        m315(.A(x2), .B(x1), .Y(mai_mai_n332_));
  OAI210     m316(.A0(mai_mai_n266_), .A1(mai_mai_n332_), .B0(mai_mai_n36_), .Y(mai_mai_n333_));
  NO2        m317(.A(mai_mai_n332_), .B(mai_mai_n314_), .Y(mai_mai_n334_));
  AOI210     m318(.A0(mai_mai_n62_), .A1(x4), .B0(mai_mai_n115_), .Y(mai_mai_n335_));
  OAI210     m319(.A0(mai_mai_n335_), .A1(mai_mai_n334_), .B0(mai_mai_n258_), .Y(mai_mai_n336_));
  NO2        m320(.A(mai_mai_n281_), .B(mai_mai_n92_), .Y(mai_mai_n337_));
  NO2        m321(.A(mai_mai_n337_), .B(mai_mai_n36_), .Y(mai_mai_n338_));
  NO2        m322(.A(mai_mai_n312_), .B(mai_mai_n215_), .Y(mai_mai_n339_));
  NA2        m323(.A(x9), .B(x0), .Y(mai_mai_n340_));
  AOI210     m324(.A0(mai_mai_n92_), .A1(mai_mai_n76_), .B0(mai_mai_n340_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n341_), .A1(mai_mai_n339_), .B0(mai_mai_n94_), .Y(mai_mai_n342_));
  NA3        m326(.A(mai_mai_n342_), .B(mai_mai_n338_), .C(mai_mai_n336_), .Y(mai_mai_n343_));
  NA2        m327(.A(mai_mai_n343_), .B(mai_mai_n333_), .Y(mai_mai_n344_));
  NO2        m328(.A(mai_mai_n220_), .B(mai_mai_n116_), .Y(mai_mai_n345_));
  NO3        m329(.A(mai_mai_n265_), .B(mai_mai_n123_), .C(mai_mai_n18_), .Y(mai_mai_n346_));
  NO2        m330(.A(mai_mai_n346_), .B(mai_mai_n345_), .Y(mai_mai_n347_));
  OAI210     m331(.A0(mai_mai_n121_), .A1(mai_mai_n109_), .B0(mai_mai_n184_), .Y(mai_mai_n348_));
  NA3        m332(.A(mai_mai_n348_), .B(x6), .C(x3), .Y(mai_mai_n349_));
  AOI210     m333(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n350_));
  OAI220     m334(.A0(mai_mai_n350_), .A1(mai_mai_n324_), .B0(mai_mai_n281_), .B1(mai_mai_n321_), .Y(mai_mai_n351_));
  INV        m335(.A(mai_mai_n351_), .Y(mai_mai_n352_));
  NA2        m336(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n353_));
  OAI210     m337(.A0(mai_mai_n109_), .A1(mai_mai_n17_), .B0(mai_mai_n353_), .Y(mai_mai_n354_));
  NA2        m338(.A(mai_mai_n354_), .B(mai_mai_n79_), .Y(mai_mai_n355_));
  NA4        m339(.A(mai_mai_n355_), .B(mai_mai_n352_), .C(mai_mai_n349_), .D(mai_mai_n347_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n114_), .A1(x3), .B0(mai_mai_n315_), .Y(mai_mai_n357_));
  NA3        m341(.A(mai_mai_n239_), .B(mai_mai_n225_), .C(mai_mai_n84_), .Y(mai_mai_n358_));
  NA3        m342(.A(mai_mai_n358_), .B(mai_mai_n357_), .C(mai_mai_n161_), .Y(mai_mai_n359_));
  AOI210     m343(.A0(mai_mai_n356_), .A1(x4), .B0(mai_mai_n359_), .Y(mai_mai_n360_));
  NA3        m344(.A(mai_mai_n334_), .B(mai_mai_n220_), .C(mai_mai_n94_), .Y(mai_mai_n361_));
  NOi21      m345(.An(x4), .B(x0), .Y(mai_mai_n362_));
  XO2        m346(.A(x4), .B(x0), .Y(mai_mai_n363_));
  OAI210     m347(.A0(mai_mai_n363_), .A1(mai_mai_n120_), .B0(mai_mai_n276_), .Y(mai_mai_n364_));
  AOI220     m348(.A0(mai_mai_n364_), .A1(x8), .B0(mai_mai_n362_), .B1(mai_mai_n95_), .Y(mai_mai_n365_));
  AOI210     m349(.A0(mai_mai_n365_), .A1(mai_mai_n361_), .B0(x3), .Y(mai_mai_n366_));
  INV        m350(.A(mai_mai_n95_), .Y(mai_mai_n367_));
  NO2        m351(.A(mai_mai_n94_), .B(x4), .Y(mai_mai_n368_));
  AOI220     m352(.A0(mai_mai_n368_), .A1(mai_mai_n44_), .B0(mai_mai_n130_), .B1(mai_mai_n367_), .Y(mai_mai_n369_));
  NO2        m353(.A(mai_mai_n363_), .B(x2), .Y(mai_mai_n370_));
  INV        m354(.A(mai_mai_n370_), .Y(mai_mai_n371_));
  NA4        m355(.A(mai_mai_n371_), .B(mai_mai_n369_), .C(mai_mai_n235_), .D(x6), .Y(mai_mai_n372_));
  OAI220     m356(.A0(mai_mai_n314_), .A1(mai_mai_n92_), .B0(mai_mai_n189_), .B1(mai_mai_n94_), .Y(mai_mai_n373_));
  NO2        m357(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n374_));
  NA2        m358(.A(mai_mai_n373_), .B(mai_mai_n61_), .Y(mai_mai_n375_));
  NO2        m359(.A(mai_mai_n158_), .B(mai_mai_n81_), .Y(mai_mai_n376_));
  NO2        m360(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n377_));
  NOi21      m361(.An(mai_mai_n126_), .B(mai_mai_n27_), .Y(mai_mai_n378_));
  AOI210     m362(.A0(mai_mai_n377_), .A1(mai_mai_n376_), .B0(mai_mai_n378_), .Y(mai_mai_n379_));
  OAI210     m363(.A0(mai_mai_n375_), .A1(mai_mai_n62_), .B0(mai_mai_n379_), .Y(mai_mai_n380_));
  OAI220     m364(.A0(mai_mai_n380_), .A1(x6), .B0(mai_mai_n372_), .B1(mai_mai_n366_), .Y(mai_mai_n381_));
  OAI210     m365(.A0(mai_mai_n63_), .A1(mai_mai_n48_), .B0(mai_mai_n42_), .Y(mai_mai_n382_));
  OAI210     m366(.A0(mai_mai_n382_), .A1(mai_mai_n94_), .B0(mai_mai_n325_), .Y(mai_mai_n383_));
  AOI210     m367(.A0(mai_mai_n383_), .A1(mai_mai_n18_), .B0(mai_mai_n161_), .Y(mai_mai_n384_));
  AO220      m368(.A0(mai_mai_n384_), .A1(mai_mai_n381_), .B0(mai_mai_n360_), .B1(mai_mai_n344_), .Y(mai_mai_n385_));
  NA2        m369(.A(mai_mai_n377_), .B(x6), .Y(mai_mai_n386_));
  AOI210     m370(.A0(x6), .A1(x1), .B0(mai_mai_n160_), .Y(mai_mai_n387_));
  NA2        m371(.A(mai_mai_n368_), .B(x0), .Y(mai_mai_n388_));
  NA2        m372(.A(mai_mai_n84_), .B(x6), .Y(mai_mai_n389_));
  OAI210     m373(.A0(mai_mai_n388_), .A1(mai_mai_n387_), .B0(mai_mai_n389_), .Y(mai_mai_n390_));
  AOI220     m374(.A0(mai_mai_n390_), .A1(mai_mai_n386_), .B0(mai_mai_n229_), .B1(mai_mai_n49_), .Y(mai_mai_n391_));
  NA3        m375(.A(mai_mai_n391_), .B(mai_mai_n385_), .C(mai_mai_n331_), .Y(mai_mai_n392_));
  AOI210     m376(.A0(mai_mai_n208_), .A1(x8), .B0(mai_mai_n114_), .Y(mai_mai_n393_));
  NA2        m377(.A(mai_mai_n393_), .B(mai_mai_n353_), .Y(mai_mai_n394_));
  NA3        m378(.A(mai_mai_n394_), .B(mai_mai_n205_), .C(mai_mai_n161_), .Y(mai_mai_n395_));
  OAI210     m379(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n243_), .Y(mai_mai_n396_));
  AO220      m380(.A0(mai_mai_n396_), .A1(mai_mai_n157_), .B0(mai_mai_n113_), .B1(x4), .Y(mai_mai_n397_));
  NA3        m381(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n398_));
  NA2        m382(.A(mai_mai_n234_), .B(x0), .Y(mai_mai_n399_));
  OAI220     m383(.A0(mai_mai_n399_), .A1(mai_mai_n220_), .B0(mai_mai_n398_), .B1(mai_mai_n367_), .Y(mai_mai_n400_));
  AOI210     m384(.A0(mai_mai_n397_), .A1(mai_mai_n122_), .B0(mai_mai_n400_), .Y(mai_mai_n401_));
  AOI210     m385(.A0(mai_mai_n401_), .A1(mai_mai_n395_), .B0(mai_mai_n25_), .Y(mai_mai_n402_));
  NA3        m386(.A(mai_mai_n124_), .B(mai_mai_n234_), .C(x0), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n123_), .A1(mai_mai_n121_), .B0(mai_mai_n42_), .Y(mai_mai_n404_));
  NOi31      m388(.An(mai_mai_n404_), .B(mai_mai_n374_), .C(mai_mai_n190_), .Y(mai_mai_n405_));
  NA2        m389(.A(mai_mai_n405_), .B(mai_mai_n157_), .Y(mai_mai_n406_));
  NA2        m390(.A(mai_mai_n406_), .B(mai_mai_n403_), .Y(mai_mai_n407_));
  OAI210     m391(.A0(mai_mai_n407_), .A1(mai_mai_n402_), .B0(x6), .Y(mai_mai_n408_));
  NA2        m392(.A(mai_mai_n48_), .B(mai_mai_n141_), .Y(mai_mai_n409_));
  NA3        m393(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n410_));
  AOI220     m394(.A0(mai_mai_n410_), .A1(mai_mai_n409_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n411_));
  NO2        m395(.A(mai_mai_n161_), .B(x0), .Y(mai_mai_n412_));
  AOI220     m396(.A0(mai_mai_n412_), .A1(mai_mai_n234_), .B0(mai_mai_n205_), .B1(mai_mai_n161_), .Y(mai_mai_n413_));
  AOI210     m397(.A0(mai_mai_n132_), .A1(mai_mai_n263_), .B0(x1), .Y(mai_mai_n414_));
  OAI210     m398(.A0(mai_mai_n413_), .A1(x8), .B0(mai_mai_n414_), .Y(mai_mai_n415_));
  NA2        m399(.A(mai_mai_n376_), .B(mai_mai_n161_), .Y(mai_mai_n416_));
  NA3        m400(.A(mai_mai_n416_), .B(x1), .C(mai_mai_n50_), .Y(mai_mai_n417_));
  OAI210     m401(.A0(mai_mai_n415_), .A1(mai_mai_n411_), .B0(mai_mai_n417_), .Y(mai_mai_n418_));
  NOi31      m402(.An(mai_mai_n412_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n419_));
  AOI210     m403(.A0(mai_mai_n38_), .A1(x9), .B0(mai_mai_n139_), .Y(mai_mai_n420_));
  NO3        m404(.A(mai_mai_n420_), .B(mai_mai_n129_), .C(mai_mai_n43_), .Y(mai_mai_n421_));
  NOi31      m405(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n422_));
  AOI220     m406(.A0(mai_mai_n422_), .A1(mai_mai_n362_), .B0(mai_mai_n130_), .B1(x3), .Y(mai_mai_n423_));
  AOI210     m407(.A0(mai_mai_n276_), .A1(mai_mai_n60_), .B0(mai_mai_n128_), .Y(mai_mai_n424_));
  OAI210     m408(.A0(mai_mai_n424_), .A1(x3), .B0(mai_mai_n423_), .Y(mai_mai_n425_));
  NO3        m409(.A(mai_mai_n425_), .B(mai_mai_n421_), .C(x2), .Y(mai_mai_n426_));
  OAI210     m410(.A0(mai_mai_n314_), .A1(mai_mai_n43_), .B0(mai_mai_n363_), .Y(mai_mai_n427_));
  AOI210     m411(.A0(x9), .A1(mai_mai_n48_), .B0(mai_mai_n398_), .Y(mai_mai_n428_));
  AOI220     m412(.A0(mai_mai_n428_), .A1(mai_mai_n94_), .B0(mai_mai_n427_), .B1(mai_mai_n161_), .Y(mai_mai_n429_));
  NO2        m413(.A(mai_mai_n429_), .B(mai_mai_n54_), .Y(mai_mai_n430_));
  NO3        m414(.A(mai_mai_n430_), .B(mai_mai_n426_), .C(mai_mai_n419_), .Y(mai_mai_n431_));
  AOI210     m415(.A0(mai_mai_n431_), .A1(mai_mai_n418_), .B0(mai_mai_n25_), .Y(mai_mai_n432_));
  NO3        m416(.A(mai_mai_n62_), .B(x4), .C(x1), .Y(mai_mai_n433_));
  NO3        m417(.A(mai_mai_n67_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n434_));
  AOI220     m418(.A0(mai_mai_n434_), .A1(mai_mai_n277_), .B0(mai_mai_n433_), .B1(mai_mai_n404_), .Y(mai_mai_n435_));
  NO2        m419(.A(mai_mai_n435_), .B(mai_mai_n106_), .Y(mai_mai_n436_));
  NO3        m420(.A(mai_mai_n281_), .B(mai_mai_n184_), .C(mai_mai_n40_), .Y(mai_mai_n437_));
  OAI210     m421(.A0(mai_mai_n437_), .A1(mai_mai_n436_), .B0(x7), .Y(mai_mai_n438_));
  NA2        m422(.A(mai_mai_n239_), .B(x7), .Y(mai_mai_n439_));
  NA3        m423(.A(mai_mai_n439_), .B(mai_mai_n160_), .C(mai_mai_n140_), .Y(mai_mai_n440_));
  NA2        m424(.A(mai_mai_n440_), .B(mai_mai_n438_), .Y(mai_mai_n441_));
  OAI210     m425(.A0(mai_mai_n441_), .A1(mai_mai_n432_), .B0(mai_mai_n36_), .Y(mai_mai_n442_));
  INV        m426(.A(mai_mai_n215_), .Y(mai_mai_n443_));
  NO4        m427(.A(mai_mai_n443_), .B(mai_mai_n78_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n444_));
  NA2        m428(.A(mai_mai_n266_), .B(mai_mai_n21_), .Y(mai_mai_n445_));
  NO2        m429(.A(mai_mai_n169_), .B(mai_mai_n141_), .Y(mai_mai_n446_));
  NA2        m430(.A(mai_mai_n446_), .B(mai_mai_n445_), .Y(mai_mai_n447_));
  AOI210     m431(.A0(mai_mai_n447_), .A1(mai_mai_n175_), .B0(mai_mai_n28_), .Y(mai_mai_n448_));
  AOI220     m432(.A0(mai_mai_n374_), .A1(mai_mai_n94_), .B0(mai_mai_n158_), .B1(mai_mai_n208_), .Y(mai_mai_n449_));
  NA2        m433(.A(mai_mai_n449_), .B(mai_mai_n92_), .Y(mai_mai_n450_));
  NA2        m434(.A(mai_mai_n450_), .B(mai_mai_n185_), .Y(mai_mai_n451_));
  OAI220     m435(.A0(mai_mai_n290_), .A1(mai_mai_n68_), .B0(mai_mai_n169_), .B1(mai_mai_n43_), .Y(mai_mai_n452_));
  NA2        m436(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n453_));
  AOI210     m437(.A0(mai_mai_n172_), .A1(mai_mai_n27_), .B0(mai_mai_n73_), .Y(mai_mai_n454_));
  OAI210     m438(.A0(mai_mai_n157_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n455_));
  NO3        m439(.A(mai_mai_n422_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n456_));
  AOI210     m440(.A0(mai_mai_n456_), .A1(mai_mai_n455_), .B0(mai_mai_n454_), .Y(mai_mai_n457_));
  OAI210     m441(.A0(mai_mai_n162_), .A1(mai_mai_n453_), .B0(mai_mai_n457_), .Y(mai_mai_n458_));
  AOI220     m442(.A0(mai_mai_n458_), .A1(x0), .B0(mai_mai_n452_), .B1(mai_mai_n141_), .Y(mai_mai_n459_));
  AOI210     m443(.A0(mai_mai_n459_), .A1(mai_mai_n451_), .B0(mai_mai_n245_), .Y(mai_mai_n460_));
  INV        m444(.A(x5), .Y(mai_mai_n461_));
  NO4        m445(.A(mai_mai_n109_), .B(mai_mai_n461_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n462_));
  NO4        m446(.A(mai_mai_n462_), .B(mai_mai_n460_), .C(mai_mai_n448_), .D(mai_mai_n444_), .Y(mai_mai_n463_));
  NA3        m447(.A(mai_mai_n463_), .B(mai_mai_n442_), .C(mai_mai_n408_), .Y(mai_mai_n464_));
  AOI210     m448(.A0(mai_mai_n392_), .A1(mai_mai_n25_), .B0(mai_mai_n464_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  NO2        u022(.A(men_men_n23_), .B(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n37_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  AOI210     u033(.A0(men_men_n22_), .A1(men_men_n19_), .B0(men_men_n35_), .Y(men_men_n50_));
  INV        u034(.A(x2), .Y(men_men_n51_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n17_), .Y(men_men_n52_));
  NA2        u036(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  OAI210     u038(.A0(men_men_n50_), .A1(men_men_n32_), .B0(men_men_n54_), .Y(men_men_n55_));
  NO3        u039(.A(men_men_n55_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u040(.A(x8), .B(x7), .Y(men_men_n57_));
  NA2        u041(.A(men_men_n41_), .B(x1), .Y(men_men_n58_));
  INV        u042(.A(x9), .Y(men_men_n59_));
  NO2        u043(.A(men_men_n59_), .B(men_men_n36_), .Y(men_men_n60_));
  INV        u044(.A(men_men_n60_), .Y(men_men_n61_));
  NO3        u045(.A(men_men_n61_), .B(men_men_n58_), .C(men_men_n57_), .Y(men_men_n62_));
  NO2        u046(.A(x7), .B(x6), .Y(men_men_n63_));
  NO2        u047(.A(men_men_n58_), .B(x5), .Y(men_men_n64_));
  NO2        u048(.A(x8), .B(x2), .Y(men_men_n65_));
  INV        u049(.A(men_men_n65_), .Y(men_men_n66_));
  NO2        u050(.A(men_men_n66_), .B(x1), .Y(men_men_n67_));
  OA210      u051(.A0(men_men_n67_), .A1(men_men_n64_), .B0(men_men_n63_), .Y(men_men_n68_));
  OAI210     u052(.A0(men_men_n42_), .A1(men_men_n25_), .B0(men_men_n51_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n53_), .A1(men_men_n20_), .B0(men_men_n69_), .Y(men_men_n70_));
  NAi31      u054(.An(x1), .B(x9), .C(x5), .Y(men_men_n71_));
  OAI220     u055(.A0(men_men_n71_), .A1(men_men_n41_), .B0(men_men_n70_), .B1(men_men_n68_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n72_), .A1(men_men_n62_), .B0(x4), .Y(men_men_n73_));
  NA2        u057(.A(men_men_n46_), .B(x2), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n53_), .B0(x0), .Y(men_men_n75_));
  NA2        u059(.A(x5), .B(x3), .Y(men_men_n76_));
  NO2        u060(.A(x8), .B(x6), .Y(men_men_n77_));
  NO4        u061(.A(men_men_n77_), .B(men_men_n76_), .C(men_men_n63_), .D(men_men_n51_), .Y(men_men_n78_));
  NAi21      u062(.An(x4), .B(x3), .Y(men_men_n79_));
  INV        u063(.A(men_men_n79_), .Y(men_men_n80_));
  NO2        u064(.A(men_men_n80_), .B(men_men_n22_), .Y(men_men_n81_));
  NO2        u065(.A(x4), .B(x2), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(x3), .Y(men_men_n83_));
  NO3        u067(.A(men_men_n83_), .B(men_men_n81_), .C(men_men_n18_), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n78_), .C(men_men_n75_), .Y(men_men_n85_));
  NO4        u069(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n86_));
  NA2        u070(.A(men_men_n59_), .B(men_men_n46_), .Y(men_men_n87_));
  INV        u071(.A(men_men_n87_), .Y(men_men_n88_));
  OAI210     u072(.A0(men_men_n86_), .A1(men_men_n64_), .B0(men_men_n88_), .Y(men_men_n89_));
  NA2        u073(.A(x3), .B(men_men_n18_), .Y(men_men_n90_));
  NO2        u074(.A(men_men_n90_), .B(men_men_n25_), .Y(men_men_n91_));
  INV        u075(.A(x8), .Y(men_men_n92_));
  NA2        u076(.A(x2), .B(x1), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n91_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n26_), .Y(men_men_n96_));
  AOI210     u080(.A0(men_men_n53_), .A1(men_men_n25_), .B0(men_men_n51_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n43_), .A1(men_men_n37_), .B0(men_men_n46_), .Y(men_men_n98_));
  NO3        u082(.A(men_men_n98_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n99_));
  NA2        u083(.A(x4), .B(men_men_n41_), .Y(men_men_n100_));
  NO2        u084(.A(men_men_n46_), .B(men_men_n51_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n100_), .B(x1), .Y(men_men_n102_));
  NO2        u086(.A(x3), .B(x2), .Y(men_men_n103_));
  NA3        u087(.A(men_men_n103_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n104_));
  AOI210     u088(.A0(x8), .A1(x6), .B0(men_men_n104_), .Y(men_men_n105_));
  NA2        u089(.A(men_men_n51_), .B(x1), .Y(men_men_n106_));
  OAI210     u090(.A0(men_men_n106_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n107_));
  NO4        u091(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n102_), .D(men_men_n99_), .Y(men_men_n108_));
  AO220      u092(.A0(men_men_n108_), .A1(men_men_n89_), .B0(men_men_n85_), .B1(men_men_n73_), .Y(men02));
  NO2        u093(.A(x3), .B(men_men_n51_), .Y(men_men_n110_));
  NO2        u094(.A(x8), .B(men_men_n18_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n51_), .B(men_men_n17_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n41_), .B(x0), .Y(men_men_n113_));
  OAI210     u097(.A0(men_men_n87_), .A1(men_men_n112_), .B0(men_men_n113_), .Y(men_men_n114_));
  AOI220     u098(.A0(men_men_n114_), .A1(men_men_n111_), .B0(men_men_n110_), .B1(x4), .Y(men_men_n115_));
  NO3        u099(.A(men_men_n115_), .B(x7), .C(x5), .Y(men_men_n116_));
  NA2        u100(.A(x9), .B(x2), .Y(men_men_n117_));
  OR2        u101(.A(x8), .B(x0), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  NAi21      u103(.An(x2), .B(x8), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  NO2        u105(.A(men_men_n121_), .B(men_men_n119_), .Y(men_men_n122_));
  NO2        u106(.A(x4), .B(x1), .Y(men_men_n123_));
  NA3        u107(.A(men_men_n123_), .B(men_men_n122_), .C(men_men_n57_), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x1), .Y(men_men_n125_));
  NO3        u109(.A(x9), .B(x8), .C(x7), .Y(men_men_n126_));
  NOi21      u110(.An(x0), .B(x4), .Y(men_men_n127_));
  NAi21      u111(.An(x8), .B(x7), .Y(men_men_n128_));
  NO2        u112(.A(men_men_n128_), .B(men_men_n59_), .Y(men_men_n129_));
  NA2        u113(.A(men_men_n126_), .B(men_men_n125_), .Y(men_men_n130_));
  AOI210     u114(.A0(men_men_n130_), .A1(men_men_n124_), .B0(men_men_n76_), .Y(men_men_n131_));
  NO2        u115(.A(x5), .B(men_men_n46_), .Y(men_men_n132_));
  NA2        u116(.A(x2), .B(men_men_n18_), .Y(men_men_n133_));
  AOI210     u117(.A0(men_men_n133_), .A1(men_men_n106_), .B0(men_men_n113_), .Y(men_men_n134_));
  OAI210     u118(.A0(men_men_n134_), .A1(men_men_n35_), .B0(men_men_n132_), .Y(men_men_n135_));
  NAi21      u119(.An(x0), .B(x4), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x1), .Y(men_men_n137_));
  NO2        u121(.A(x7), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n82_), .B(men_men_n101_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n139_), .B(x3), .Y(men_men_n140_));
  OAI210     u124(.A0(men_men_n138_), .A1(men_men_n137_), .B0(men_men_n140_), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n142_));
  NA2        u126(.A(x5), .B(x0), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n46_), .B(x2), .Y(men_men_n144_));
  NA3        u128(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n142_), .Y(men_men_n145_));
  NA4        u129(.A(men_men_n145_), .B(men_men_n141_), .C(men_men_n135_), .D(men_men_n36_), .Y(men_men_n146_));
  NO3        u130(.A(men_men_n146_), .B(men_men_n131_), .C(men_men_n116_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n76_), .B(men_men_n74_), .C(men_men_n24_), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n149_));
  AOI220     u133(.A0(men_men_n125_), .A1(men_men_n149_), .B0(men_men_n64_), .B1(men_men_n17_), .Y(men_men_n150_));
  NO3        u134(.A(men_men_n150_), .B(men_men_n57_), .C(men_men_n59_), .Y(men_men_n151_));
  NA2        u135(.A(x7), .B(x3), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n100_), .B(x5), .Y(men_men_n153_));
  NO2        u137(.A(x9), .B(x7), .Y(men_men_n154_));
  NOi21      u138(.An(x8), .B(x0), .Y(men_men_n155_));
  OA210      u139(.A0(men_men_n154_), .A1(x1), .B0(men_men_n155_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n41_), .B(x2), .Y(men_men_n157_));
  INV        u141(.A(x7), .Y(men_men_n158_));
  NA2        u142(.A(men_men_n158_), .B(men_men_n18_), .Y(men_men_n159_));
  NA2        u143(.A(men_men_n159_), .B(men_men_n157_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n25_), .B(x4), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n161_), .B(men_men_n127_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n160_), .Y(men_men_n163_));
  AOI210     u147(.A0(men_men_n156_), .A1(men_men_n153_), .B0(men_men_n163_), .Y(men_men_n164_));
  OAI210     u148(.A0(men_men_n152_), .A1(men_men_n48_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u149(.A(x5), .B(x1), .Y(men_men_n166_));
  INV        u150(.A(men_men_n166_), .Y(men_men_n167_));
  AOI210     u151(.A0(men_men_n167_), .A1(men_men_n127_), .B0(men_men_n36_), .Y(men_men_n168_));
  NO2        u152(.A(men_men_n59_), .B(men_men_n92_), .Y(men_men_n169_));
  NAi21      u153(.An(x2), .B(x7), .Y(men_men_n170_));
  NO3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n46_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n171_), .B(men_men_n64_), .Y(men_men_n172_));
  NA2        u156(.A(men_men_n172_), .B(men_men_n168_), .Y(men_men_n173_));
  NO4        u157(.A(men_men_n173_), .B(men_men_n165_), .C(men_men_n151_), .D(men_men_n148_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n174_), .B(men_men_n147_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n143_), .B(men_men_n139_), .Y(men_men_n176_));
  NA2        u160(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n178_));
  NA3        u162(.A(men_men_n178_), .B(men_men_n177_), .C(men_men_n24_), .Y(men_men_n179_));
  AN2        u163(.A(men_men_n179_), .B(men_men_n144_), .Y(men_men_n180_));
  NA2        u164(.A(x8), .B(x0), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n158_), .B(men_men_n25_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n125_), .B(x4), .Y(men_men_n183_));
  NA2        u167(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  AOI210     u168(.A0(men_men_n181_), .A1(men_men_n133_), .B0(men_men_n184_), .Y(men_men_n185_));
  NA2        u169(.A(x2), .B(x0), .Y(men_men_n186_));
  NA2        u170(.A(x4), .B(x1), .Y(men_men_n187_));
  NAi21      u171(.An(men_men_n123_), .B(men_men_n187_), .Y(men_men_n188_));
  NOi31      u172(.An(men_men_n188_), .B(men_men_n161_), .C(men_men_n186_), .Y(men_men_n189_));
  NO4        u173(.A(men_men_n189_), .B(men_men_n185_), .C(men_men_n180_), .D(men_men_n176_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(men_men_n41_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n179_), .B(men_men_n74_), .Y(men_men_n192_));
  INV        u176(.A(men_men_n132_), .Y(men_men_n193_));
  NO2        u177(.A(men_men_n106_), .B(men_men_n17_), .Y(men_men_n194_));
  AOI210     u178(.A0(men_men_n35_), .A1(men_men_n92_), .B0(men_men_n194_), .Y(men_men_n195_));
  NO3        u179(.A(men_men_n195_), .B(men_men_n193_), .C(x7), .Y(men_men_n196_));
  NA3        u180(.A(men_men_n188_), .B(men_men_n193_), .C(men_men_n40_), .Y(men_men_n197_));
  OAI210     u181(.A0(men_men_n178_), .A1(men_men_n139_), .B0(men_men_n197_), .Y(men_men_n198_));
  NO3        u182(.A(men_men_n198_), .B(men_men_n196_), .C(men_men_n192_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n199_), .B(x3), .Y(men_men_n200_));
  NO3        u184(.A(men_men_n200_), .B(men_men_n191_), .C(men_men_n175_), .Y(men03));
  NO2        u185(.A(men_men_n46_), .B(x3), .Y(men_men_n202_));
  NO2        u186(.A(x6), .B(men_men_n25_), .Y(men_men_n203_));
  INV        u187(.A(men_men_n203_), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n51_), .B(x1), .Y(men_men_n205_));
  OAI210     u189(.A0(men_men_n205_), .A1(men_men_n25_), .B0(men_men_n60_), .Y(men_men_n206_));
  OAI220     u190(.A0(men_men_n206_), .A1(men_men_n17_), .B0(men_men_n204_), .B1(men_men_n106_), .Y(men_men_n207_));
  NA2        u191(.A(men_men_n207_), .B(men_men_n202_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n76_), .B(x6), .Y(men_men_n209_));
  NA2        u193(.A(x6), .B(men_men_n25_), .Y(men_men_n210_));
  NO2        u194(.A(men_men_n210_), .B(x4), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n18_), .B(x0), .Y(men_men_n212_));
  AO220      u196(.A0(men_men_n212_), .A1(men_men_n211_), .B0(men_men_n209_), .B1(men_men_n52_), .Y(men_men_n213_));
  INV        u197(.A(men_men_n213_), .Y(men_men_n214_));
  NA2        u198(.A(x3), .B(men_men_n17_), .Y(men_men_n215_));
  NA2        u199(.A(x9), .B(men_men_n51_), .Y(men_men_n216_));
  NO2        u200(.A(x5), .B(x1), .Y(men_men_n217_));
  AOI220     u201(.A0(men_men_n217_), .A1(men_men_n17_), .B0(men_men_n103_), .B1(x5), .Y(men_men_n218_));
  NO2        u202(.A(men_men_n215_), .B(men_men_n177_), .Y(men_men_n219_));
  NO3        u203(.A(x3), .B(x2), .C(x1), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n221_));
  OAI210     u205(.A0(men_men_n218_), .A1(men_men_n61_), .B0(men_men_n221_), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n222_), .B(men_men_n46_), .Y(men_men_n223_));
  NA3        u207(.A(men_men_n223_), .B(men_men_n214_), .C(men_men_n208_), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n225_));
  NA2        u209(.A(men_men_n225_), .B(men_men_n19_), .Y(men_men_n226_));
  NO2        u210(.A(x3), .B(men_men_n17_), .Y(men_men_n227_));
  NO2        u211(.A(men_men_n227_), .B(x6), .Y(men_men_n228_));
  NOi21      u212(.An(men_men_n82_), .B(men_men_n228_), .Y(men_men_n229_));
  NA2        u213(.A(men_men_n59_), .B(men_men_n92_), .Y(men_men_n230_));
  NA3        u214(.A(men_men_n230_), .B(men_men_n227_), .C(x6), .Y(men_men_n231_));
  AOI210     u215(.A0(men_men_n231_), .A1(men_men_n229_), .B0(men_men_n158_), .Y(men_men_n232_));
  AO210      u216(.A0(men_men_n232_), .A1(men_men_n226_), .B0(men_men_n182_), .Y(men_men_n233_));
  NA2        u217(.A(men_men_n41_), .B(men_men_n51_), .Y(men_men_n234_));
  OAI210     u218(.A0(men_men_n234_), .A1(men_men_n25_), .B0(men_men_n178_), .Y(men_men_n235_));
  NO3        u219(.A(men_men_n187_), .B(men_men_n59_), .C(x6), .Y(men_men_n236_));
  AOI220     u220(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n144_), .B1(men_men_n91_), .Y(men_men_n237_));
  NA2        u221(.A(x6), .B(men_men_n46_), .Y(men_men_n238_));
  OAI210     u222(.A0(men_men_n119_), .A1(men_men_n77_), .B0(x4), .Y(men_men_n239_));
  AOI210     u223(.A0(men_men_n239_), .A1(men_men_n238_), .B0(men_men_n76_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n203_), .B(men_men_n137_), .Y(men_men_n241_));
  NA3        u225(.A(men_men_n215_), .B(men_men_n132_), .C(x6), .Y(men_men_n242_));
  OAI210     u226(.A0(men_men_n92_), .A1(men_men_n36_), .B0(men_men_n64_), .Y(men_men_n243_));
  NA3        u227(.A(men_men_n243_), .B(men_men_n242_), .C(men_men_n241_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n240_), .B0(x2), .Y(men_men_n245_));
  NA3        u229(.A(men_men_n245_), .B(men_men_n237_), .C(men_men_n233_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n224_), .A1(x8), .B0(men_men_n246_), .Y(men_men_n247_));
  NO2        u231(.A(men_men_n92_), .B(x3), .Y(men_men_n248_));
  NA2        u232(.A(men_men_n248_), .B(men_men_n211_), .Y(men_men_n249_));
  NO3        u233(.A(men_men_n90_), .B(men_men_n77_), .C(men_men_n25_), .Y(men_men_n250_));
  AOI210     u234(.A0(men_men_n228_), .A1(men_men_n161_), .B0(men_men_n250_), .Y(men_men_n251_));
  AOI210     u235(.A0(men_men_n251_), .A1(men_men_n249_), .B0(x2), .Y(men_men_n252_));
  NO2        u236(.A(x4), .B(men_men_n51_), .Y(men_men_n253_));
  AOI220     u237(.A0(men_men_n211_), .A1(men_men_n194_), .B0(men_men_n253_), .B1(men_men_n64_), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n59_), .B(x6), .Y(men_men_n255_));
  NA3        u239(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n256_));
  AOI210     u240(.A0(men_men_n256_), .A1(men_men_n143_), .B0(men_men_n255_), .Y(men_men_n257_));
  NA2        u241(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n258_), .B(men_men_n25_), .Y(men_men_n259_));
  OAI210     u243(.A0(men_men_n259_), .A1(men_men_n257_), .B0(men_men_n123_), .Y(men_men_n260_));
  NA2        u244(.A(men_men_n215_), .B(x6), .Y(men_men_n261_));
  NO2        u245(.A(men_men_n215_), .B(x6), .Y(men_men_n262_));
  NAi21      u246(.An(men_men_n169_), .B(men_men_n262_), .Y(men_men_n263_));
  NA3        u247(.A(men_men_n263_), .B(men_men_n261_), .C(men_men_n149_), .Y(men_men_n264_));
  NA4        u248(.A(men_men_n264_), .B(men_men_n260_), .C(men_men_n254_), .D(men_men_n158_), .Y(men_men_n265_));
  NO2        u249(.A(x9), .B(x6), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n143_), .B(men_men_n18_), .Y(men_men_n267_));
  NAi21      u251(.An(men_men_n267_), .B(men_men_n256_), .Y(men_men_n268_));
  NAi21      u252(.An(x1), .B(x4), .Y(men_men_n269_));
  AOI210     u253(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n270_));
  OAI210     u254(.A0(men_men_n143_), .A1(x3), .B0(men_men_n270_), .Y(men_men_n271_));
  AOI220     u255(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n268_), .B1(men_men_n266_), .Y(men_men_n272_));
  INV        u256(.A(men_men_n272_), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n59_), .B(x2), .Y(men_men_n274_));
  NO3        u258(.A(x9), .B(x6), .C(x0), .Y(men_men_n275_));
  NA2        u259(.A(men_men_n106_), .B(men_men_n25_), .Y(men_men_n276_));
  NA2        u260(.A(x6), .B(x2), .Y(men_men_n277_));
  NO2        u261(.A(men_men_n277_), .B(men_men_n177_), .Y(men_men_n278_));
  AOI210     u262(.A0(men_men_n276_), .A1(men_men_n275_), .B0(men_men_n278_), .Y(men_men_n279_));
  OAI220     u263(.A0(men_men_n279_), .A1(men_men_n41_), .B0(men_men_n183_), .B1(men_men_n44_), .Y(men_men_n280_));
  NA2        u264(.A(men_men_n280_), .B(men_men_n273_), .Y(men_men_n281_));
  NA2        u265(.A(x9), .B(men_men_n41_), .Y(men_men_n282_));
  NO2        u266(.A(men_men_n282_), .B(men_men_n210_), .Y(men_men_n283_));
  OR3        u267(.A(men_men_n283_), .B(men_men_n209_), .C(men_men_n153_), .Y(men_men_n284_));
  NA2        u268(.A(x4), .B(x0), .Y(men_men_n285_));
  NO3        u269(.A(men_men_n71_), .B(men_men_n285_), .C(x6), .Y(men_men_n286_));
  AOI210     u270(.A0(men_men_n284_), .A1(men_men_n40_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI210     u271(.A0(men_men_n287_), .A1(men_men_n281_), .B0(x8), .Y(men_men_n288_));
  INV        u272(.A(men_men_n255_), .Y(men_men_n289_));
  NA2        u273(.A(men_men_n217_), .B(men_men_n289_), .Y(men_men_n290_));
  INV        u274(.A(men_men_n181_), .Y(men_men_n291_));
  OAI210     u275(.A0(men_men_n291_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n292_));
  AOI210     u276(.A0(men_men_n292_), .A1(men_men_n290_), .B0(men_men_n234_), .Y(men_men_n293_));
  NO4        u277(.A(men_men_n293_), .B(men_men_n288_), .C(men_men_n265_), .D(men_men_n252_), .Y(men_men_n294_));
  NO2        u278(.A(men_men_n169_), .B(x1), .Y(men_men_n295_));
  NO3        u279(.A(men_men_n295_), .B(x3), .C(men_men_n36_), .Y(men_men_n296_));
  OAI210     u280(.A0(men_men_n296_), .A1(men_men_n262_), .B0(x2), .Y(men_men_n297_));
  OAI210     u281(.A0(men_men_n291_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n298_));
  AOI210     u282(.A0(men_men_n298_), .A1(men_men_n297_), .B0(men_men_n193_), .Y(men_men_n299_));
  NOi21      u283(.An(men_men_n277_), .B(men_men_n17_), .Y(men_men_n300_));
  NA3        u284(.A(men_men_n300_), .B(men_men_n217_), .C(men_men_n38_), .Y(men_men_n301_));
  AOI210     u285(.A0(men_men_n36_), .A1(men_men_n51_), .B0(x0), .Y(men_men_n302_));
  NA3        u286(.A(men_men_n302_), .B(men_men_n167_), .C(men_men_n32_), .Y(men_men_n303_));
  NA2        u287(.A(x3), .B(x2), .Y(men_men_n304_));
  AOI220     u288(.A0(men_men_n304_), .A1(men_men_n234_), .B0(men_men_n303_), .B1(men_men_n301_), .Y(men_men_n305_));
  NAi21      u289(.An(x4), .B(x0), .Y(men_men_n306_));
  NO3        u290(.A(men_men_n306_), .B(men_men_n42_), .C(x2), .Y(men_men_n307_));
  OAI210     u291(.A0(x6), .A1(men_men_n18_), .B0(men_men_n307_), .Y(men_men_n308_));
  OAI220     u292(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n309_));
  NO2        u293(.A(x9), .B(x8), .Y(men_men_n310_));
  NA3        u294(.A(men_men_n310_), .B(men_men_n36_), .C(men_men_n51_), .Y(men_men_n311_));
  OAI210     u295(.A0(men_men_n302_), .A1(men_men_n300_), .B0(men_men_n311_), .Y(men_men_n312_));
  AOI220     u296(.A0(men_men_n312_), .A1(men_men_n80_), .B0(men_men_n309_), .B1(men_men_n31_), .Y(men_men_n313_));
  AOI210     u297(.A0(men_men_n313_), .A1(men_men_n308_), .B0(men_men_n25_), .Y(men_men_n314_));
  NA3        u298(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n315_));
  OAI210     u299(.A0(men_men_n302_), .A1(men_men_n300_), .B0(men_men_n315_), .Y(men_men_n316_));
  INV        u300(.A(men_men_n219_), .Y(men_men_n317_));
  NA2        u301(.A(men_men_n36_), .B(men_men_n41_), .Y(men_men_n318_));
  OR2        u302(.A(men_men_n318_), .B(men_men_n285_), .Y(men_men_n319_));
  OAI220     u303(.A0(men_men_n319_), .A1(men_men_n166_), .B0(men_men_n238_), .B1(men_men_n317_), .Y(men_men_n320_));
  AO210      u304(.A0(men_men_n316_), .A1(men_men_n153_), .B0(men_men_n320_), .Y(men_men_n321_));
  NO4        u305(.A(men_men_n321_), .B(men_men_n314_), .C(men_men_n305_), .D(men_men_n299_), .Y(men_men_n322_));
  OAI210     u306(.A0(men_men_n294_), .A1(men_men_n247_), .B0(men_men_n322_), .Y(men04));
  OAI210     u307(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n324_));
  NA3        u308(.A(men_men_n324_), .B(men_men_n275_), .C(men_men_n83_), .Y(men_men_n325_));
  NO2        u309(.A(x2), .B(x1), .Y(men_men_n326_));
  OAI210     u310(.A0(men_men_n258_), .A1(men_men_n326_), .B0(men_men_n36_), .Y(men_men_n327_));
  NO2        u311(.A(men_men_n326_), .B(men_men_n306_), .Y(men_men_n328_));
  AOI210     u312(.A0(men_men_n59_), .A1(x4), .B0(men_men_n112_), .Y(men_men_n329_));
  OAI210     u313(.A0(men_men_n329_), .A1(men_men_n328_), .B0(men_men_n248_), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n274_), .B(men_men_n90_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n331_), .B(men_men_n36_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n304_), .B(men_men_n212_), .Y(men_men_n333_));
  NA2        u317(.A(men_men_n333_), .B(men_men_n92_), .Y(men_men_n334_));
  NA3        u318(.A(men_men_n334_), .B(men_men_n332_), .C(men_men_n330_), .Y(men_men_n335_));
  NA2        u319(.A(men_men_n335_), .B(men_men_n327_), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n216_), .B(men_men_n113_), .Y(men_men_n337_));
  NO3        u321(.A(men_men_n255_), .B(men_men_n120_), .C(men_men_n18_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n338_), .B(men_men_n337_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n118_), .A1(men_men_n106_), .B0(men_men_n181_), .Y(men_men_n340_));
  NA3        u324(.A(men_men_n340_), .B(x6), .C(x3), .Y(men_men_n341_));
  NOi21      u325(.An(men_men_n155_), .B(men_men_n133_), .Y(men_men_n342_));
  AOI210     u326(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n343_));
  OAI220     u327(.A0(men_men_n343_), .A1(men_men_n318_), .B0(men_men_n274_), .B1(men_men_n315_), .Y(men_men_n344_));
  AOI210     u328(.A0(men_men_n342_), .A1(men_men_n60_), .B0(men_men_n344_), .Y(men_men_n345_));
  NA2        u329(.A(x2), .B(men_men_n17_), .Y(men_men_n346_));
  OAI210     u330(.A0(men_men_n106_), .A1(men_men_n17_), .B0(men_men_n346_), .Y(men_men_n347_));
  AOI220     u331(.A0(men_men_n347_), .A1(men_men_n77_), .B0(men_men_n331_), .B1(men_men_n92_), .Y(men_men_n348_));
  NA4        u332(.A(men_men_n348_), .B(men_men_n345_), .C(men_men_n341_), .D(men_men_n339_), .Y(men_men_n349_));
  OAI210     u333(.A0(men_men_n111_), .A1(x3), .B0(men_men_n307_), .Y(men_men_n350_));
  NA2        u334(.A(men_men_n350_), .B(men_men_n158_), .Y(men_men_n351_));
  AOI210     u335(.A0(men_men_n349_), .A1(x4), .B0(men_men_n351_), .Y(men_men_n352_));
  NA3        u336(.A(men_men_n328_), .B(men_men_n216_), .C(men_men_n92_), .Y(men_men_n353_));
  NOi21      u337(.An(x4), .B(x0), .Y(men_men_n354_));
  XO2        u338(.A(x4), .B(x0), .Y(men_men_n355_));
  OAI210     u339(.A0(men_men_n355_), .A1(men_men_n117_), .B0(men_men_n269_), .Y(men_men_n356_));
  AOI220     u340(.A0(men_men_n356_), .A1(x8), .B0(men_men_n354_), .B1(men_men_n93_), .Y(men_men_n357_));
  AOI210     u341(.A0(men_men_n357_), .A1(men_men_n353_), .B0(x3), .Y(men_men_n358_));
  INV        u342(.A(men_men_n93_), .Y(men_men_n359_));
  NO2        u343(.A(men_men_n92_), .B(x4), .Y(men_men_n360_));
  AOI220     u344(.A0(men_men_n360_), .A1(men_men_n42_), .B0(men_men_n127_), .B1(men_men_n359_), .Y(men_men_n361_));
  NO3        u345(.A(men_men_n355_), .B(men_men_n169_), .C(x2), .Y(men_men_n362_));
  NO3        u346(.A(men_men_n230_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n363_), .B(men_men_n362_), .Y(men_men_n364_));
  NA4        u348(.A(men_men_n364_), .B(men_men_n361_), .C(men_men_n226_), .D(x6), .Y(men_men_n365_));
  OAI220     u349(.A0(men_men_n306_), .A1(men_men_n90_), .B0(men_men_n186_), .B1(men_men_n92_), .Y(men_men_n366_));
  NO2        u350(.A(men_men_n41_), .B(x0), .Y(men_men_n367_));
  OR2        u351(.A(men_men_n360_), .B(men_men_n367_), .Y(men_men_n368_));
  NO2        u352(.A(men_men_n155_), .B(men_men_n106_), .Y(men_men_n369_));
  AOI220     u353(.A0(men_men_n369_), .A1(men_men_n368_), .B0(men_men_n366_), .B1(men_men_n58_), .Y(men_men_n370_));
  NO2        u354(.A(men_men_n155_), .B(men_men_n79_), .Y(men_men_n371_));
  NO2        u355(.A(men_men_n35_), .B(x2), .Y(men_men_n372_));
  NOi21      u356(.An(men_men_n123_), .B(men_men_n27_), .Y(men_men_n373_));
  AOI210     u357(.A0(men_men_n372_), .A1(men_men_n371_), .B0(men_men_n373_), .Y(men_men_n374_));
  OAI210     u358(.A0(men_men_n370_), .A1(men_men_n59_), .B0(men_men_n374_), .Y(men_men_n375_));
  OAI220     u359(.A0(men_men_n375_), .A1(x6), .B0(men_men_n365_), .B1(men_men_n358_), .Y(men_men_n376_));
  NA2        u360(.A(men_men_n46_), .B(men_men_n40_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n377_), .A1(men_men_n92_), .B0(men_men_n319_), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n378_), .A1(men_men_n18_), .B0(men_men_n158_), .Y(men_men_n379_));
  AO220      u363(.A0(men_men_n379_), .A1(men_men_n376_), .B0(men_men_n352_), .B1(men_men_n336_), .Y(men_men_n380_));
  NA2        u364(.A(men_men_n372_), .B(x6), .Y(men_men_n381_));
  AOI210     u365(.A0(x6), .A1(x1), .B0(men_men_n157_), .Y(men_men_n382_));
  NA2        u366(.A(men_men_n360_), .B(x0), .Y(men_men_n383_));
  NA2        u367(.A(men_men_n82_), .B(x6), .Y(men_men_n384_));
  OAI210     u368(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n384_), .Y(men_men_n385_));
  AOI220     u369(.A0(men_men_n385_), .A1(men_men_n381_), .B0(men_men_n220_), .B1(men_men_n47_), .Y(men_men_n386_));
  NA3        u370(.A(men_men_n386_), .B(men_men_n380_), .C(men_men_n325_), .Y(men_men_n387_));
  AOI210     u371(.A0(men_men_n205_), .A1(x8), .B0(men_men_n111_), .Y(men_men_n388_));
  NA2        u372(.A(men_men_n388_), .B(men_men_n346_), .Y(men_men_n389_));
  NA3        u373(.A(men_men_n389_), .B(men_men_n202_), .C(men_men_n158_), .Y(men_men_n390_));
  OAI210     u374(.A0(men_men_n28_), .A1(x1), .B0(men_men_n234_), .Y(men_men_n391_));
  AO220      u375(.A0(men_men_n391_), .A1(men_men_n154_), .B0(men_men_n110_), .B1(x4), .Y(men_men_n392_));
  NA3        u376(.A(x7), .B(x3), .C(x0), .Y(men_men_n393_));
  NA2        u377(.A(men_men_n225_), .B(x0), .Y(men_men_n394_));
  OAI220     u378(.A0(men_men_n394_), .A1(men_men_n216_), .B0(men_men_n393_), .B1(men_men_n359_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n392_), .A1(men_men_n119_), .B0(men_men_n395_), .Y(men_men_n396_));
  AOI210     u380(.A0(men_men_n396_), .A1(men_men_n390_), .B0(men_men_n25_), .Y(men_men_n397_));
  NA3        u381(.A(men_men_n121_), .B(men_men_n225_), .C(x0), .Y(men_men_n398_));
  OAI210     u382(.A0(men_men_n202_), .A1(men_men_n65_), .B0(men_men_n212_), .Y(men_men_n399_));
  NA3        u383(.A(men_men_n205_), .B(men_men_n227_), .C(x8), .Y(men_men_n400_));
  AOI210     u384(.A0(men_men_n400_), .A1(men_men_n399_), .B0(men_men_n25_), .Y(men_men_n401_));
  NA2        u385(.A(men_men_n401_), .B(men_men_n154_), .Y(men_men_n402_));
  NAi31      u386(.An(men_men_n48_), .B(men_men_n295_), .C(men_men_n182_), .Y(men_men_n403_));
  NA3        u387(.A(men_men_n403_), .B(men_men_n402_), .C(men_men_n398_), .Y(men_men_n404_));
  OAI210     u388(.A0(men_men_n404_), .A1(men_men_n397_), .B0(x6), .Y(men_men_n405_));
  OAI210     u389(.A0(men_men_n169_), .A1(men_men_n46_), .B0(men_men_n138_), .Y(men_men_n406_));
  AOI210     u390(.A0(men_men_n38_), .A1(men_men_n32_), .B0(men_men_n406_), .Y(men_men_n407_));
  NO2        u391(.A(men_men_n158_), .B(x0), .Y(men_men_n408_));
  AOI220     u392(.A0(men_men_n408_), .A1(men_men_n225_), .B0(men_men_n202_), .B1(men_men_n158_), .Y(men_men_n409_));
  AOI210     u393(.A0(men_men_n129_), .A1(men_men_n253_), .B0(x1), .Y(men_men_n410_));
  OAI210     u394(.A0(men_men_n409_), .A1(x8), .B0(men_men_n410_), .Y(men_men_n411_));
  NAi31      u395(.An(x2), .B(x8), .C(x0), .Y(men_men_n412_));
  OAI210     u396(.A0(men_men_n412_), .A1(x4), .B0(men_men_n170_), .Y(men_men_n413_));
  NA3        u397(.A(men_men_n413_), .B(men_men_n152_), .C(x9), .Y(men_men_n414_));
  NO4        u398(.A(men_men_n128_), .B(men_men_n306_), .C(x9), .D(x2), .Y(men_men_n415_));
  NOi21      u399(.An(men_men_n126_), .B(men_men_n186_), .Y(men_men_n416_));
  NO3        u400(.A(men_men_n416_), .B(men_men_n415_), .C(men_men_n18_), .Y(men_men_n417_));
  NO3        u401(.A(x9), .B(men_men_n158_), .C(x0), .Y(men_men_n418_));
  AOI220     u402(.A0(men_men_n418_), .A1(men_men_n248_), .B0(men_men_n371_), .B1(men_men_n158_), .Y(men_men_n419_));
  NA4        u403(.A(men_men_n419_), .B(men_men_n417_), .C(men_men_n414_), .D(men_men_n48_), .Y(men_men_n420_));
  OAI210     u404(.A0(men_men_n411_), .A1(men_men_n407_), .B0(men_men_n420_), .Y(men_men_n421_));
  NOi31      u405(.An(men_men_n408_), .B(men_men_n32_), .C(x8), .Y(men_men_n422_));
  INV        u406(.A(men_men_n136_), .Y(men_men_n423_));
  NO3        u407(.A(men_men_n423_), .B(men_men_n126_), .C(men_men_n41_), .Y(men_men_n424_));
  NOi31      u408(.An(x1), .B(x8), .C(x7), .Y(men_men_n425_));
  AOI220     u409(.A0(men_men_n425_), .A1(men_men_n354_), .B0(men_men_n127_), .B1(x3), .Y(men_men_n426_));
  AOI210     u410(.A0(men_men_n269_), .A1(men_men_n57_), .B0(men_men_n125_), .Y(men_men_n427_));
  OAI210     u411(.A0(men_men_n427_), .A1(x3), .B0(men_men_n426_), .Y(men_men_n428_));
  NO3        u412(.A(men_men_n428_), .B(men_men_n424_), .C(x2), .Y(men_men_n429_));
  OAI220     u413(.A0(men_men_n355_), .A1(men_men_n310_), .B0(men_men_n306_), .B1(men_men_n41_), .Y(men_men_n430_));
  INV        u414(.A(men_men_n393_), .Y(men_men_n431_));
  AOI220     u415(.A0(men_men_n431_), .A1(men_men_n92_), .B0(men_men_n430_), .B1(men_men_n158_), .Y(men_men_n432_));
  NO2        u416(.A(men_men_n432_), .B(men_men_n51_), .Y(men_men_n433_));
  NO3        u417(.A(men_men_n433_), .B(men_men_n429_), .C(men_men_n422_), .Y(men_men_n434_));
  AOI210     u418(.A0(men_men_n434_), .A1(men_men_n421_), .B0(men_men_n25_), .Y(men_men_n435_));
  NA4        u419(.A(men_men_n31_), .B(men_men_n92_), .C(x2), .D(men_men_n17_), .Y(men_men_n436_));
  NO3        u420(.A(men_men_n65_), .B(men_men_n18_), .C(x0), .Y(men_men_n437_));
  NA2        u421(.A(men_men_n437_), .B(men_men_n270_), .Y(men_men_n438_));
  NO2        u422(.A(men_men_n438_), .B(men_men_n103_), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n274_), .B(men_men_n181_), .C(men_men_n38_), .Y(men_men_n440_));
  OAI210     u424(.A0(men_men_n440_), .A1(men_men_n439_), .B0(x7), .Y(men_men_n441_));
  NA2        u425(.A(men_men_n230_), .B(x7), .Y(men_men_n442_));
  NA3        u426(.A(men_men_n442_), .B(men_men_n157_), .C(men_men_n137_), .Y(men_men_n443_));
  NA3        u427(.A(men_men_n443_), .B(men_men_n441_), .C(men_men_n436_), .Y(men_men_n444_));
  OAI210     u428(.A0(men_men_n444_), .A1(men_men_n435_), .B0(men_men_n36_), .Y(men_men_n445_));
  NO2        u429(.A(men_men_n418_), .B(men_men_n212_), .Y(men_men_n446_));
  NO4        u430(.A(men_men_n446_), .B(men_men_n76_), .C(x4), .D(men_men_n51_), .Y(men_men_n447_));
  NA2        u431(.A(men_men_n258_), .B(men_men_n21_), .Y(men_men_n448_));
  NO2        u432(.A(men_men_n166_), .B(men_men_n138_), .Y(men_men_n449_));
  NA2        u433(.A(men_men_n449_), .B(men_men_n448_), .Y(men_men_n450_));
  NO2        u434(.A(men_men_n450_), .B(men_men_n28_), .Y(men_men_n451_));
  NA2        u435(.A(men_men_n412_), .B(men_men_n90_), .Y(men_men_n452_));
  NA2        u436(.A(men_men_n452_), .B(men_men_n182_), .Y(men_men_n453_));
  OAI220     u437(.A0(men_men_n282_), .A1(men_men_n66_), .B0(men_men_n166_), .B1(men_men_n41_), .Y(men_men_n454_));
  NA2        u438(.A(x3), .B(men_men_n51_), .Y(men_men_n455_));
  AOI210     u439(.A0(men_men_n170_), .A1(men_men_n27_), .B0(men_men_n71_), .Y(men_men_n456_));
  OAI210     u440(.A0(men_men_n154_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n457_));
  NO3        u441(.A(men_men_n425_), .B(x3), .C(men_men_n51_), .Y(men_men_n458_));
  AOI210     u442(.A0(men_men_n458_), .A1(men_men_n457_), .B0(men_men_n456_), .Y(men_men_n459_));
  OAI210     u443(.A0(men_men_n159_), .A1(men_men_n455_), .B0(men_men_n459_), .Y(men_men_n460_));
  AOI220     u444(.A0(men_men_n460_), .A1(x0), .B0(men_men_n454_), .B1(men_men_n138_), .Y(men_men_n461_));
  AOI210     u445(.A0(men_men_n461_), .A1(men_men_n453_), .B0(men_men_n238_), .Y(men_men_n462_));
  NA2        u446(.A(x9), .B(x5), .Y(men_men_n463_));
  NO4        u447(.A(men_men_n106_), .B(men_men_n463_), .C(men_men_n57_), .D(men_men_n32_), .Y(men_men_n464_));
  NO4        u448(.A(men_men_n464_), .B(men_men_n462_), .C(men_men_n451_), .D(men_men_n447_), .Y(men_men_n465_));
  NA3        u449(.A(men_men_n465_), .B(men_men_n445_), .C(men_men_n405_), .Y(men_men_n466_));
  AOI210     u450(.A0(men_men_n387_), .A1(men_men_n25_), .B0(men_men_n466_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule