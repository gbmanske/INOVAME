//Benchmark atmr_prom1_2672_0.0313

module atmr_prom1(x0, x1, x2, x3, x4, x5, x6, x7, x8, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39;
 wire ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1401_, ori_ori_n1402_, ori_ori_n1403_, ori_ori_n1404_, ori_ori_n1406_, ori_ori_n1407_, ori_ori_n1408_, ori_ori_n1409_, ori_ori_n1410_, ori_ori_n1411_, ori_ori_n1412_, ori_ori_n1413_, ori_ori_n1414_, ori_ori_n1415_, ori_ori_n1416_, ori_ori_n1417_, ori_ori_n1418_, ori_ori_n1419_, ori_ori_n1420_, ori_ori_n1421_, ori_ori_n1422_, ori_ori_n1423_, ori_ori_n1424_, ori_ori_n1425_, ori_ori_n1426_, ori_ori_n1427_, ori_ori_n1428_, ori_ori_n1429_, ori_ori_n1430_, ori_ori_n1431_, ori_ori_n1432_, ori_ori_n1433_, ori_ori_n1434_, ori_ori_n1435_, ori_ori_n1436_, ori_ori_n1437_, ori_ori_n1438_, ori_ori_n1439_, ori_ori_n1440_, ori_ori_n1441_, ori_ori_n1442_, ori_ori_n1443_, ori_ori_n1444_, ori_ori_n1445_, ori_ori_n1446_, ori_ori_n1447_, ori_ori_n1448_, ori_ori_n1449_, ori_ori_n1450_, ori_ori_n1451_, ori_ori_n1452_, ori_ori_n1453_, ori_ori_n1454_, ori_ori_n1455_, ori_ori_n1456_, ori_ori_n1457_, ori_ori_n1458_, ori_ori_n1459_, ori_ori_n1460_, ori_ori_n1461_, ori_ori_n1462_, ori_ori_n1463_, ori_ori_n1464_, ori_ori_n1465_, ori_ori_n1466_, ori_ori_n1467_, ori_ori_n1468_, ori_ori_n1469_, ori_ori_n1470_, ori_ori_n1471_, ori_ori_n1472_, ori_ori_n1473_, ori_ori_n1474_, ori_ori_n1475_, ori_ori_n1476_, ori_ori_n1477_, ori_ori_n1478_, ori_ori_n1479_, ori_ori_n1480_, ori_ori_n1481_, ori_ori_n1482_, ori_ori_n1483_, ori_ori_n1484_, ori_ori_n1485_, ori_ori_n1486_, ori_ori_n1487_, ori_ori_n1488_, ori_ori_n1489_, ori_ori_n1490_, ori_ori_n1491_, ori_ori_n1492_, ori_ori_n1493_, ori_ori_n1494_, ori_ori_n1496_, ori_ori_n1497_, ori_ori_n1498_, ori_ori_n1499_, ori_ori_n1500_, ori_ori_n1501_, ori_ori_n1502_, ori_ori_n1503_, ori_ori_n1504_, ori_ori_n1505_, ori_ori_n1506_, ori_ori_n1507_, ori_ori_n1508_, ori_ori_n1509_, ori_ori_n1510_, ori_ori_n1511_, ori_ori_n1512_, ori_ori_n1513_, ori_ori_n1514_, ori_ori_n1515_, ori_ori_n1516_, ori_ori_n1517_, ori_ori_n1518_, ori_ori_n1519_, ori_ori_n1520_, ori_ori_n1521_, ori_ori_n1522_, ori_ori_n1523_, ori_ori_n1525_, ori_ori_n1526_, ori_ori_n1527_, ori_ori_n1528_, ori_ori_n1529_, ori_ori_n1530_, ori_ori_n1531_, ori_ori_n1532_, ori_ori_n1533_, ori_ori_n1534_, ori_ori_n1535_, ori_ori_n1536_, ori_ori_n1537_, ori_ori_n1538_, ori_ori_n1539_, ori_ori_n1540_, ori_ori_n1541_, ori_ori_n1542_, ori_ori_n1543_, ori_ori_n1544_, ori_ori_n1545_, ori_ori_n1546_, ori_ori_n1547_, ori_ori_n1548_, ori_ori_n1549_, ori_ori_n1550_, ori_ori_n1551_, ori_ori_n1552_, ori_ori_n1553_, ori_ori_n1554_, ori_ori_n1555_, ori_ori_n1556_, ori_ori_n1557_, ori_ori_n1558_, ori_ori_n1559_, ori_ori_n1560_, ori_ori_n1561_, ori_ori_n1562_, ori_ori_n1563_, ori_ori_n1564_, ori_ori_n1565_, ori_ori_n1566_, ori_ori_n1567_, ori_ori_n1568_, ori_ori_n1569_, ori_ori_n1570_, ori_ori_n1571_, ori_ori_n1572_, ori_ori_n1573_, ori_ori_n1574_, ori_ori_n1575_, ori_ori_n1576_, ori_ori_n1577_, ori_ori_n1578_, ori_ori_n1579_, ori_ori_n1580_, ori_ori_n1581_, ori_ori_n1582_, ori_ori_n1583_, ori_ori_n1584_, ori_ori_n1585_, ori_ori_n1586_, ori_ori_n1587_, ori_ori_n1588_, ori_ori_n1589_, ori_ori_n1590_, ori_ori_n1592_, ori_ori_n1593_, ori_ori_n1594_, ori_ori_n1595_, ori_ori_n1596_, ori_ori_n1597_, ori_ori_n1598_, ori_ori_n1599_, ori_ori_n1600_, ori_ori_n1601_, ori_ori_n1602_, ori_ori_n1603_, ori_ori_n1604_, ori_ori_n1605_, ori_ori_n1606_, ori_ori_n1607_, ori_ori_n1608_, ori_ori_n1609_, ori_ori_n1610_, ori_ori_n1611_, ori_ori_n1612_, ori_ori_n1613_, ori_ori_n1614_, ori_ori_n1615_, ori_ori_n1616_, ori_ori_n1617_, ori_ori_n1618_, ori_ori_n1619_, ori_ori_n1620_, ori_ori_n1621_, ori_ori_n1622_, ori_ori_n1623_, ori_ori_n1624_, ori_ori_n1625_, ori_ori_n1626_, ori_ori_n1627_, ori_ori_n1628_, ori_ori_n1629_, ori_ori_n1630_, ori_ori_n1631_, ori_ori_n1632_, ori_ori_n1633_, ori_ori_n1634_, ori_ori_n1635_, ori_ori_n1636_, ori_ori_n1637_, ori_ori_n1638_, ori_ori_n1639_, ori_ori_n1640_, ori_ori_n1641_, ori_ori_n1642_, ori_ori_n1643_, ori_ori_n1644_, ori_ori_n1645_, ori_ori_n1646_, ori_ori_n1647_, ori_ori_n1648_, ori_ori_n1650_, ori_ori_n1651_, ori_ori_n1652_, ori_ori_n1653_, ori_ori_n1654_, ori_ori_n1655_, ori_ori_n1656_, ori_ori_n1657_, ori_ori_n1658_, ori_ori_n1659_, ori_ori_n1660_, ori_ori_n1661_, ori_ori_n1662_, ori_ori_n1663_, ori_ori_n1664_, ori_ori_n1665_, ori_ori_n1666_, ori_ori_n1667_, ori_ori_n1668_, ori_ori_n1669_, ori_ori_n1670_, ori_ori_n1671_, ori_ori_n1672_, ori_ori_n1673_, ori_ori_n1674_, ori_ori_n1676_, ori_ori_n1677_, ori_ori_n1678_, ori_ori_n1679_, ori_ori_n1680_, ori_ori_n1681_, ori_ori_n1682_, ori_ori_n1683_, ori_ori_n1684_, ori_ori_n1685_, ori_ori_n1686_, ori_ori_n1687_, ori_ori_n1688_, ori_ori_n1689_, ori_ori_n1690_, ori_ori_n1691_, ori_ori_n1692_, ori_ori_n1693_, ori_ori_n1694_, ori_ori_n1695_, ori_ori_n1696_, ori_ori_n1697_, ori_ori_n1698_, ori_ori_n1699_, ori_ori_n1700_, ori_ori_n1701_, ori_ori_n1702_, ori_ori_n1703_, ori_ori_n1704_, ori_ori_n1705_, ori_ori_n1706_, ori_ori_n1707_, ori_ori_n1708_, ori_ori_n1709_, ori_ori_n1710_, ori_ori_n1711_, ori_ori_n1712_, ori_ori_n1713_, ori_ori_n1714_, ori_ori_n1715_, ori_ori_n1716_, ori_ori_n1717_, ori_ori_n1718_, ori_ori_n1719_, ori_ori_n1720_, ori_ori_n1721_, ori_ori_n1722_, ori_ori_n1723_, ori_ori_n1724_, ori_ori_n1725_, ori_ori_n1726_, ori_ori_n1727_, ori_ori_n1728_, ori_ori_n1729_, ori_ori_n1730_, ori_ori_n1731_, ori_ori_n1732_, ori_ori_n1733_, ori_ori_n1734_, ori_ori_n1735_, ori_ori_n1736_, ori_ori_n1737_, ori_ori_n1738_, ori_ori_n1739_, ori_ori_n1740_, ori_ori_n1741_, ori_ori_n1742_, ori_ori_n1743_, ori_ori_n1744_, ori_ori_n1745_, ori_ori_n1746_, ori_ori_n1747_, ori_ori_n1748_, ori_ori_n1749_, ori_ori_n1750_, ori_ori_n1751_, ori_ori_n1752_, ori_ori_n1753_, ori_ori_n1754_, ori_ori_n1755_, ori_ori_n1756_, ori_ori_n1757_, ori_ori_n1758_, ori_ori_n1759_, ori_ori_n1760_, ori_ori_n1761_, ori_ori_n1763_, ori_ori_n1764_, ori_ori_n1765_, ori_ori_n1766_, ori_ori_n1767_, ori_ori_n1768_, ori_ori_n1769_, ori_ori_n1770_, ori_ori_n1771_, ori_ori_n1772_, ori_ori_n1773_, ori_ori_n1774_, ori_ori_n1775_, ori_ori_n1776_, ori_ori_n1777_, ori_ori_n1778_, ori_ori_n1779_, ori_ori_n1780_, ori_ori_n1781_, ori_ori_n1782_, ori_ori_n1783_, ori_ori_n1784_, ori_ori_n1785_, ori_ori_n1786_, ori_ori_n1787_, ori_ori_n1788_, ori_ori_n1789_, ori_ori_n1790_, ori_ori_n1791_, ori_ori_n1792_, ori_ori_n1793_, ori_ori_n1794_, ori_ori_n1795_, ori_ori_n1796_, ori_ori_n1797_, ori_ori_n1798_, ori_ori_n1799_, ori_ori_n1800_, ori_ori_n1801_, ori_ori_n1802_, ori_ori_n1803_, ori_ori_n1804_, ori_ori_n1805_, ori_ori_n1806_, ori_ori_n1807_, ori_ori_n1808_, ori_ori_n1809_, ori_ori_n1810_, ori_ori_n1811_, ori_ori_n1812_, ori_ori_n1813_, ori_ori_n1814_, ori_ori_n1815_, ori_ori_n1816_, ori_ori_n1818_, ori_ori_n1819_, ori_ori_n1820_, ori_ori_n1821_, ori_ori_n1822_, ori_ori_n1823_, ori_ori_n1824_, ori_ori_n1825_, ori_ori_n1826_, ori_ori_n1827_, ori_ori_n1828_, ori_ori_n1829_, ori_ori_n1830_, ori_ori_n1831_, ori_ori_n1832_, ori_ori_n1833_, ori_ori_n1834_, ori_ori_n1835_, ori_ori_n1836_, ori_ori_n1838_, ori_ori_n1839_, ori_ori_n1840_, ori_ori_n1841_, ori_ori_n1842_, ori_ori_n1843_, ori_ori_n1844_, ori_ori_n1845_, ori_ori_n1846_, ori_ori_n1847_, ori_ori_n1848_, ori_ori_n1849_, ori_ori_n1850_, ori_ori_n1852_, ori_ori_n1853_, ori_ori_n1854_, ori_ori_n1855_, ori_ori_n1856_, ori_ori_n1857_, ori_ori_n1858_, ori_ori_n1859_, ori_ori_n1860_, ori_ori_n1861_, ori_ori_n1862_, ori_ori_n1863_, ori_ori_n1864_, ori_ori_n1865_, ori_ori_n1866_, ori_ori_n1868_, ori_ori_n1869_, ori_ori_n1870_, ori_ori_n1871_, ori_ori_n1872_, ori_ori_n1873_, ori_ori_n1874_, ori_ori_n1875_, ori_ori_n1876_, ori_ori_n1877_, ori_ori_n1878_, ori_ori_n1879_, ori_ori_n1880_, ori_ori_n1881_, ori_ori_n1882_, ori_ori_n1883_, ori_ori_n1884_, ori_ori_n1885_, ori_ori_n1886_, ori_ori_n1887_, ori_ori_n1888_, ori_ori_n1889_, ori_ori_n1890_, ori_ori_n1891_, ori_ori_n1892_, ori_ori_n1893_, ori_ori_n1894_, ori_ori_n1895_, ori_ori_n1896_, ori_ori_n1897_, ori_ori_n1898_, ori_ori_n1899_, ori_ori_n1900_, ori_ori_n1901_, ori_ori_n1902_, ori_ori_n1903_, ori_ori_n1904_, ori_ori_n1905_, ori_ori_n1906_, ori_ori_n1907_, ori_ori_n1908_, ori_ori_n1909_, ori_ori_n1910_, ori_ori_n1911_, ori_ori_n1912_, ori_ori_n1913_, ori_ori_n1914_, ori_ori_n1916_, ori_ori_n1917_, ori_ori_n1918_, ori_ori_n1919_, ori_ori_n1920_, ori_ori_n1921_, ori_ori_n1922_, ori_ori_n1923_, ori_ori_n1924_, ori_ori_n1925_, ori_ori_n1926_, ori_ori_n1927_, ori_ori_n1928_, ori_ori_n1929_, ori_ori_n1931_, ori_ori_n1932_, ori_ori_n1933_, ori_ori_n1934_, ori_ori_n1935_, ori_ori_n1936_, ori_ori_n1937_, ori_ori_n1938_, ori_ori_n1939_, ori_ori_n1940_, ori_ori_n1941_, ori_ori_n1942_, ori_ori_n1943_, ori_ori_n1944_, ori_ori_n1945_, ori_ori_n1946_, ori_ori_n1947_, ori_ori_n1948_, ori_ori_n1949_, ori_ori_n1950_, ori_ori_n1951_, ori_ori_n1952_, ori_ori_n1953_, ori_ori_n1954_, ori_ori_n1955_, ori_ori_n1956_, ori_ori_n1957_, ori_ori_n1958_, ori_ori_n1959_, ori_ori_n1960_, ori_ori_n1961_, ori_ori_n1962_, ori_ori_n1963_, ori_ori_n1964_, ori_ori_n1965_, ori_ori_n1966_, ori_ori_n1967_, ori_ori_n1968_, ori_ori_n1969_, ori_ori_n1970_, ori_ori_n1971_, ori_ori_n1972_, ori_ori_n1973_, ori_ori_n1974_, ori_ori_n1975_, ori_ori_n1976_, ori_ori_n1977_, ori_ori_n1978_, ori_ori_n1980_, ori_ori_n1981_, ori_ori_n1982_, ori_ori_n1983_, ori_ori_n1984_, ori_ori_n1985_, ori_ori_n1986_, ori_ori_n1987_, ori_ori_n1988_, ori_ori_n1989_, ori_ori_n1990_, ori_ori_n1991_, ori_ori_n1992_, ori_ori_n1993_, ori_ori_n1994_, ori_ori_n1995_, ori_ori_n1996_, ori_ori_n1997_, ori_ori_n1998_, ori_ori_n1999_, ori_ori_n2000_, ori_ori_n2001_, ori_ori_n2002_, ori_ori_n2003_, ori_ori_n2004_, ori_ori_n2005_, ori_ori_n2006_, ori_ori_n2007_, ori_ori_n2008_, ori_ori_n2009_, ori_ori_n2010_, ori_ori_n2011_, ori_ori_n2012_, ori_ori_n2013_, ori_ori_n2014_, ori_ori_n2015_, ori_ori_n2016_, ori_ori_n2017_, ori_ori_n2018_, ori_ori_n2019_, ori_ori_n2020_, ori_ori_n2021_, ori_ori_n2022_, ori_ori_n2023_, ori_ori_n2024_, ori_ori_n2025_, ori_ori_n2026_, ori_ori_n2027_, ori_ori_n2028_, ori_ori_n2029_, ori_ori_n2030_, ori_ori_n2031_, ori_ori_n2032_, ori_ori_n2033_, ori_ori_n2034_, ori_ori_n2035_, ori_ori_n2036_, ori_ori_n2037_, ori_ori_n2038_, ori_ori_n2039_, ori_ori_n2040_, ori_ori_n2041_, ori_ori_n2042_, ori_ori_n2043_, ori_ori_n2044_, ori_ori_n2045_, ori_ori_n2047_, ori_ori_n2048_, ori_ori_n2049_, ori_ori_n2050_, ori_ori_n2051_, ori_ori_n2052_, ori_ori_n2053_, ori_ori_n2054_, ori_ori_n2055_, ori_ori_n2056_, ori_ori_n2057_, ori_ori_n2058_, ori_ori_n2059_, ori_ori_n2060_, ori_ori_n2061_, ori_ori_n2062_, ori_ori_n2063_, ori_ori_n2064_, ori_ori_n2065_, ori_ori_n2066_, ori_ori_n2067_, ori_ori_n2068_, ori_ori_n2069_, ori_ori_n2070_, ori_ori_n2071_, ori_ori_n2072_, ori_ori_n2073_, ori_ori_n2074_, ori_ori_n2075_, ori_ori_n2076_, ori_ori_n2077_, ori_ori_n2078_, ori_ori_n2079_, ori_ori_n2080_, ori_ori_n2081_, ori_ori_n2082_, ori_ori_n2083_, ori_ori_n2084_, ori_ori_n2085_, ori_ori_n2086_, ori_ori_n2087_, ori_ori_n2088_, ori_ori_n2089_, ori_ori_n2090_, ori_ori_n2091_, ori_ori_n2092_, ori_ori_n2093_, ori_ori_n2094_, ori_ori_n2095_, ori_ori_n2096_, ori_ori_n2097_, ori_ori_n2098_, ori_ori_n2099_, ori_ori_n2100_, ori_ori_n2101_, ori_ori_n2102_, ori_ori_n2103_, ori_ori_n2104_, ori_ori_n2105_, ori_ori_n2106_, ori_ori_n2107_, ori_ori_n2108_, ori_ori_n2109_, ori_ori_n2110_, ori_ori_n2111_, ori_ori_n2112_, ori_ori_n2113_, ori_ori_n2114_, ori_ori_n2115_, ori_ori_n2116_, ori_ori_n2117_, ori_ori_n2118_, ori_ori_n2119_, ori_ori_n2120_, ori_ori_n2121_, ori_ori_n2122_, ori_ori_n2124_, ori_ori_n2125_, ori_ori_n2126_, ori_ori_n2127_, ori_ori_n2128_, ori_ori_n2129_, ori_ori_n2130_, ori_ori_n2131_, ori_ori_n2132_, ori_ori_n2133_, ori_ori_n2134_, ori_ori_n2135_, ori_ori_n2136_, ori_ori_n2137_, ori_ori_n2138_, ori_ori_n2139_, ori_ori_n2140_, ori_ori_n2141_, ori_ori_n2142_, ori_ori_n2143_, ori_ori_n2144_, ori_ori_n2145_, ori_ori_n2146_, ori_ori_n2147_, ori_ori_n2148_, ori_ori_n2149_, ori_ori_n2150_, ori_ori_n2151_, ori_ori_n2152_, ori_ori_n2153_, ori_ori_n2154_, ori_ori_n2155_, ori_ori_n2156_, ori_ori_n2157_, ori_ori_n2158_, ori_ori_n2159_, ori_ori_n2160_, ori_ori_n2161_, ori_ori_n2162_, ori_ori_n2163_, ori_ori_n2164_, ori_ori_n2165_, ori_ori_n2166_, ori_ori_n2167_, ori_ori_n2168_, ori_ori_n2169_, ori_ori_n2170_, ori_ori_n2171_, ori_ori_n2172_, ori_ori_n2173_, ori_ori_n2174_, ori_ori_n2175_, ori_ori_n2176_, ori_ori_n2177_, ori_ori_n2178_, ori_ori_n2179_, ori_ori_n2180_, ori_ori_n2181_, ori_ori_n2182_, ori_ori_n2183_, ori_ori_n2184_, ori_ori_n2185_, ori_ori_n2186_, ori_ori_n2187_, ori_ori_n2188_, ori_ori_n2189_, ori_ori_n2190_, ori_ori_n2191_, ori_ori_n2192_, ori_ori_n2193_, ori_ori_n2194_, ori_ori_n2195_, ori_ori_n2196_, ori_ori_n2197_, ori_ori_n2198_, ori_ori_n2200_, ori_ori_n2201_, ori_ori_n2202_, ori_ori_n2203_, ori_ori_n2204_, ori_ori_n2205_, ori_ori_n2206_, ori_ori_n2207_, ori_ori_n2208_, ori_ori_n2209_, ori_ori_n2210_, ori_ori_n2211_, ori_ori_n2212_, ori_ori_n2213_, ori_ori_n2214_, ori_ori_n2215_, ori_ori_n2216_, ori_ori_n2217_, ori_ori_n2218_, ori_ori_n2219_, ori_ori_n2220_, ori_ori_n2221_, ori_ori_n2222_, ori_ori_n2223_, ori_ori_n2224_, ori_ori_n2225_, ori_ori_n2226_, ori_ori_n2227_, ori_ori_n2228_, ori_ori_n2229_, ori_ori_n2230_, ori_ori_n2231_, ori_ori_n2232_, ori_ori_n2233_, ori_ori_n2234_, ori_ori_n2235_, ori_ori_n2236_, ori_ori_n2237_, ori_ori_n2238_, ori_ori_n2239_, ori_ori_n2240_, ori_ori_n2241_, ori_ori_n2242_, ori_ori_n2243_, ori_ori_n2244_, ori_ori_n2245_, ori_ori_n2246_, ori_ori_n2247_, ori_ori_n2248_, ori_ori_n2249_, ori_ori_n2250_, ori_ori_n2251_, ori_ori_n2252_, ori_ori_n2253_, ori_ori_n2254_, ori_ori_n2255_, ori_ori_n2256_, ori_ori_n2257_, ori_ori_n2258_, ori_ori_n2259_, ori_ori_n2260_, ori_ori_n2261_, ori_ori_n2262_, ori_ori_n2263_, ori_ori_n2264_, ori_ori_n2265_, ori_ori_n2266_, ori_ori_n2267_, ori_ori_n2268_, ori_ori_n2269_, ori_ori_n2270_, ori_ori_n2271_, ori_ori_n2272_, ori_ori_n2273_, ori_ori_n2274_, ori_ori_n2275_, ori_ori_n2276_, ori_ori_n2277_, ori_ori_n2279_, ori_ori_n2280_, ori_ori_n2281_, ori_ori_n2282_, ori_ori_n2283_, ori_ori_n2284_, ori_ori_n2285_, ori_ori_n2286_, ori_ori_n2287_, ori_ori_n2288_, ori_ori_n2289_, ori_ori_n2290_, ori_ori_n2291_, ori_ori_n2292_, ori_ori_n2293_, ori_ori_n2294_, ori_ori_n2295_, ori_ori_n2296_, ori_ori_n2297_, ori_ori_n2298_, ori_ori_n2299_, ori_ori_n2300_, ori_ori_n2301_, ori_ori_n2302_, ori_ori_n2303_, ori_ori_n2304_, ori_ori_n2305_, ori_ori_n2306_, ori_ori_n2307_, ori_ori_n2308_, ori_ori_n2309_, ori_ori_n2310_, ori_ori_n2311_, ori_ori_n2312_, ori_ori_n2313_, ori_ori_n2314_, ori_ori_n2315_, ori_ori_n2316_, ori_ori_n2317_, ori_ori_n2318_, ori_ori_n2319_, ori_ori_n2320_, ori_ori_n2321_, ori_ori_n2322_, ori_ori_n2323_, ori_ori_n2324_, ori_ori_n2325_, ori_ori_n2326_, ori_ori_n2327_, ori_ori_n2328_, ori_ori_n2329_, ori_ori_n2330_, ori_ori_n2331_, ori_ori_n2332_, ori_ori_n2333_, ori_ori_n2334_, ori_ori_n2335_, ori_ori_n2336_, ori_ori_n2337_, ori_ori_n2338_, ori_ori_n2339_, ori_ori_n2340_, ori_ori_n2341_, ori_ori_n2342_, ori_ori_n2343_, ori_ori_n2344_, ori_ori_n2345_, ori_ori_n2346_, ori_ori_n2347_, ori_ori_n2349_, ori_ori_n2350_, ori_ori_n2351_, ori_ori_n2352_, ori_ori_n2353_, ori_ori_n2354_, ori_ori_n2355_, ori_ori_n2356_, ori_ori_n2357_, ori_ori_n2358_, ori_ori_n2359_, ori_ori_n2360_, ori_ori_n2361_, ori_ori_n2362_, ori_ori_n2363_, ori_ori_n2364_, ori_ori_n2365_, ori_ori_n2366_, ori_ori_n2367_, ori_ori_n2368_, ori_ori_n2369_, ori_ori_n2370_, ori_ori_n2371_, ori_ori_n2372_, ori_ori_n2373_, ori_ori_n2374_, ori_ori_n2375_, ori_ori_n2376_, ori_ori_n2377_, ori_ori_n2378_, ori_ori_n2379_, ori_ori_n2380_, ori_ori_n2381_, ori_ori_n2382_, ori_ori_n2383_, ori_ori_n2384_, ori_ori_n2385_, ori_ori_n2386_, ori_ori_n2387_, ori_ori_n2388_, ori_ori_n2389_, ori_ori_n2390_, ori_ori_n2391_, ori_ori_n2392_, ori_ori_n2393_, ori_ori_n2394_, ori_ori_n2395_, ori_ori_n2396_, ori_ori_n2397_, ori_ori_n2398_, ori_ori_n2399_, ori_ori_n2400_, ori_ori_n2401_, ori_ori_n2402_, ori_ori_n2403_, ori_ori_n2404_, ori_ori_n2405_, ori_ori_n2406_, ori_ori_n2407_, ori_ori_n2408_, ori_ori_n2409_, ori_ori_n2411_, ori_ori_n2412_, ori_ori_n2413_, ori_ori_n2414_, ori_ori_n2415_, ori_ori_n2416_, ori_ori_n2417_, ori_ori_n2418_, ori_ori_n2419_, ori_ori_n2420_, ori_ori_n2421_, ori_ori_n2422_, ori_ori_n2423_, ori_ori_n2424_, ori_ori_n2425_, ori_ori_n2426_, ori_ori_n2427_, ori_ori_n2428_, ori_ori_n2429_, ori_ori_n2430_, ori_ori_n2431_, ori_ori_n2432_, ori_ori_n2433_, ori_ori_n2434_, ori_ori_n2435_, ori_ori_n2436_, ori_ori_n2437_, ori_ori_n2438_, ori_ori_n2439_, ori_ori_n2440_, ori_ori_n2441_, ori_ori_n2442_, ori_ori_n2443_, ori_ori_n2444_, ori_ori_n2445_, ori_ori_n2446_, ori_ori_n2447_, ori_ori_n2448_, ori_ori_n2449_, ori_ori_n2450_, ori_ori_n2451_, ori_ori_n2452_, ori_ori_n2453_, ori_ori_n2454_, ori_ori_n2455_, ori_ori_n2456_, ori_ori_n2457_, ori_ori_n2458_, ori_ori_n2459_, ori_ori_n2460_, ori_ori_n2461_, ori_ori_n2462_, ori_ori_n2463_, ori_ori_n2464_, ori_ori_n2465_, ori_ori_n2466_, ori_ori_n2467_, ori_ori_n2468_, ori_ori_n2469_, ori_ori_n2470_, ori_ori_n2471_, ori_ori_n2472_, ori_ori_n2473_, ori_ori_n2474_, ori_ori_n2475_, ori_ori_n2476_, ori_ori_n2477_, ori_ori_n2478_, ori_ori_n2479_, ori_ori_n2480_, ori_ori_n2481_, ori_ori_n2482_, ori_ori_n2483_, ori_ori_n2484_, ori_ori_n2485_, ori_ori_n2486_, ori_ori_n2487_, ori_ori_n2488_, ori_ori_n2490_, ori_ori_n2491_, ori_ori_n2492_, ori_ori_n2493_, ori_ori_n2494_, ori_ori_n2495_, ori_ori_n2496_, ori_ori_n2497_, ori_ori_n2498_, ori_ori_n2499_, ori_ori_n2500_, ori_ori_n2501_, ori_ori_n2502_, ori_ori_n2503_, ori_ori_n2504_, ori_ori_n2505_, ori_ori_n2506_, ori_ori_n2507_, ori_ori_n2508_, ori_ori_n2509_, ori_ori_n2510_, ori_ori_n2511_, ori_ori_n2512_, ori_ori_n2513_, ori_ori_n2514_, ori_ori_n2515_, ori_ori_n2516_, ori_ori_n2517_, ori_ori_n2518_, ori_ori_n2519_, ori_ori_n2520_, ori_ori_n2521_, ori_ori_n2522_, ori_ori_n2523_, ori_ori_n2524_, ori_ori_n2525_, ori_ori_n2526_, ori_ori_n2527_, ori_ori_n2528_, ori_ori_n2529_, ori_ori_n2530_, ori_ori_n2531_, ori_ori_n2532_, ori_ori_n2533_, ori_ori_n2534_, ori_ori_n2535_, ori_ori_n2536_, ori_ori_n2537_, ori_ori_n2538_, ori_ori_n2539_, ori_ori_n2540_, ori_ori_n2541_, ori_ori_n2542_, ori_ori_n2543_, ori_ori_n2544_, ori_ori_n2545_, ori_ori_n2546_, ori_ori_n2547_, ori_ori_n2548_, ori_ori_n2549_, ori_ori_n2550_, ori_ori_n2551_, ori_ori_n2552_, ori_ori_n2554_, ori_ori_n2555_, ori_ori_n2556_, ori_ori_n2557_, ori_ori_n2558_, ori_ori_n2559_, ori_ori_n2560_, ori_ori_n2561_, ori_ori_n2562_, ori_ori_n2563_, ori_ori_n2564_, ori_ori_n2565_, ori_ori_n2566_, ori_ori_n2567_, ori_ori_n2568_, ori_ori_n2569_, ori_ori_n2570_, ori_ori_n2571_, ori_ori_n2572_, ori_ori_n2573_, ori_ori_n2574_, ori_ori_n2575_, ori_ori_n2576_, ori_ori_n2577_, ori_ori_n2578_, ori_ori_n2579_, ori_ori_n2580_, ori_ori_n2581_, ori_ori_n2582_, ori_ori_n2583_, ori_ori_n2584_, ori_ori_n2585_, ori_ori_n2586_, ori_ori_n2587_, ori_ori_n2588_, ori_ori_n2589_, ori_ori_n2590_, ori_ori_n2591_, ori_ori_n2592_, ori_ori_n2593_, ori_ori_n2594_, ori_ori_n2595_, ori_ori_n2596_, ori_ori_n2597_, ori_ori_n2598_, ori_ori_n2599_, ori_ori_n2600_, ori_ori_n2601_, ori_ori_n2602_, ori_ori_n2603_, ori_ori_n2604_, ori_ori_n2605_, ori_ori_n2606_, ori_ori_n2607_, ori_ori_n2608_, ori_ori_n2609_, ori_ori_n2610_, ori_ori_n2611_, ori_ori_n2612_, ori_ori_n2613_, ori_ori_n2614_, ori_ori_n2615_, ori_ori_n2616_, ori_ori_n2617_, ori_ori_n2618_, ori_ori_n2619_, ori_ori_n2620_, ori_ori_n2621_, ori_ori_n2622_, ori_ori_n2623_, ori_ori_n2625_, ori_ori_n2626_, ori_ori_n2627_, ori_ori_n2628_, ori_ori_n2629_, ori_ori_n2630_, ori_ori_n2631_, ori_ori_n2632_, ori_ori_n2633_, ori_ori_n2634_, ori_ori_n2635_, ori_ori_n2636_, ori_ori_n2637_, ori_ori_n2638_, ori_ori_n2639_, ori_ori_n2640_, ori_ori_n2641_, ori_ori_n2642_, ori_ori_n2643_, ori_ori_n2644_, ori_ori_n2645_, ori_ori_n2646_, ori_ori_n2647_, ori_ori_n2648_, ori_ori_n2649_, ori_ori_n2650_, ori_ori_n2651_, ori_ori_n2652_, ori_ori_n2653_, ori_ori_n2654_, ori_ori_n2655_, ori_ori_n2656_, ori_ori_n2657_, ori_ori_n2658_, ori_ori_n2659_, ori_ori_n2660_, ori_ori_n2661_, ori_ori_n2662_, ori_ori_n2663_, ori_ori_n2664_, ori_ori_n2665_, ori_ori_n2666_, ori_ori_n2667_, ori_ori_n2668_, ori_ori_n2669_, ori_ori_n2670_, ori_ori_n2671_, ori_ori_n2672_, ori_ori_n2673_, ori_ori_n2674_, ori_ori_n2675_, ori_ori_n2676_, ori_ori_n2677_, ori_ori_n2678_, ori_ori_n2679_, ori_ori_n2680_, ori_ori_n2681_, ori_ori_n2682_, ori_ori_n2683_, ori_ori_n2684_, ori_ori_n2685_, ori_ori_n2686_, ori_ori_n2687_, ori_ori_n2688_, ori_ori_n2689_, ori_ori_n2690_, ori_ori_n2691_, ori_ori_n2692_, ori_ori_n2696_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, mai_mai_n1552_, mai_mai_n1553_, mai_mai_n1554_, mai_mai_n1555_, mai_mai_n1556_, mai_mai_n1557_, mai_mai_n1558_, mai_mai_n1559_, mai_mai_n1560_, mai_mai_n1561_, mai_mai_n1562_, mai_mai_n1563_, mai_mai_n1564_, mai_mai_n1565_, mai_mai_n1566_, mai_mai_n1567_, mai_mai_n1568_, mai_mai_n1569_, mai_mai_n1570_, mai_mai_n1571_, mai_mai_n1572_, mai_mai_n1573_, mai_mai_n1574_, mai_mai_n1575_, mai_mai_n1576_, mai_mai_n1577_, mai_mai_n1578_, mai_mai_n1579_, mai_mai_n1580_, mai_mai_n1581_, mai_mai_n1582_, mai_mai_n1583_, mai_mai_n1584_, mai_mai_n1585_, mai_mai_n1586_, mai_mai_n1587_, mai_mai_n1589_, mai_mai_n1590_, mai_mai_n1591_, mai_mai_n1592_, mai_mai_n1593_, mai_mai_n1594_, mai_mai_n1595_, mai_mai_n1596_, mai_mai_n1597_, mai_mai_n1598_, mai_mai_n1599_, mai_mai_n1600_, mai_mai_n1601_, mai_mai_n1602_, mai_mai_n1603_, mai_mai_n1604_, mai_mai_n1605_, mai_mai_n1606_, mai_mai_n1607_, mai_mai_n1608_, mai_mai_n1609_, mai_mai_n1610_, mai_mai_n1611_, mai_mai_n1612_, mai_mai_n1613_, mai_mai_n1614_, mai_mai_n1615_, mai_mai_n1616_, mai_mai_n1617_, mai_mai_n1618_, mai_mai_n1619_, mai_mai_n1620_, mai_mai_n1621_, mai_mai_n1622_, mai_mai_n1623_, mai_mai_n1624_, mai_mai_n1625_, mai_mai_n1626_, mai_mai_n1627_, mai_mai_n1628_, mai_mai_n1629_, mai_mai_n1630_, mai_mai_n1631_, mai_mai_n1632_, mai_mai_n1633_, mai_mai_n1634_, mai_mai_n1635_, mai_mai_n1636_, mai_mai_n1637_, mai_mai_n1638_, mai_mai_n1639_, mai_mai_n1640_, mai_mai_n1641_, mai_mai_n1642_, mai_mai_n1643_, mai_mai_n1644_, mai_mai_n1645_, mai_mai_n1646_, mai_mai_n1648_, mai_mai_n1649_, mai_mai_n1650_, mai_mai_n1651_, mai_mai_n1652_, mai_mai_n1653_, mai_mai_n1654_, mai_mai_n1655_, mai_mai_n1656_, mai_mai_n1657_, mai_mai_n1658_, mai_mai_n1659_, mai_mai_n1660_, mai_mai_n1661_, mai_mai_n1662_, mai_mai_n1663_, mai_mai_n1664_, mai_mai_n1665_, mai_mai_n1666_, mai_mai_n1667_, mai_mai_n1668_, mai_mai_n1669_, mai_mai_n1670_, mai_mai_n1671_, mai_mai_n1672_, mai_mai_n1674_, mai_mai_n1675_, mai_mai_n1676_, mai_mai_n1677_, mai_mai_n1678_, mai_mai_n1679_, mai_mai_n1680_, mai_mai_n1681_, mai_mai_n1682_, mai_mai_n1683_, mai_mai_n1684_, mai_mai_n1685_, mai_mai_n1686_, mai_mai_n1687_, mai_mai_n1688_, mai_mai_n1689_, mai_mai_n1690_, mai_mai_n1691_, mai_mai_n1692_, mai_mai_n1693_, mai_mai_n1694_, mai_mai_n1695_, mai_mai_n1696_, mai_mai_n1697_, mai_mai_n1698_, mai_mai_n1699_, mai_mai_n1700_, mai_mai_n1701_, mai_mai_n1702_, mai_mai_n1703_, mai_mai_n1704_, mai_mai_n1705_, mai_mai_n1706_, mai_mai_n1707_, mai_mai_n1708_, mai_mai_n1709_, mai_mai_n1710_, mai_mai_n1711_, mai_mai_n1712_, mai_mai_n1713_, mai_mai_n1714_, mai_mai_n1715_, mai_mai_n1716_, mai_mai_n1717_, mai_mai_n1718_, mai_mai_n1719_, mai_mai_n1720_, mai_mai_n1721_, mai_mai_n1722_, mai_mai_n1723_, mai_mai_n1724_, mai_mai_n1725_, mai_mai_n1726_, mai_mai_n1727_, mai_mai_n1728_, mai_mai_n1729_, mai_mai_n1730_, mai_mai_n1731_, mai_mai_n1732_, mai_mai_n1733_, mai_mai_n1734_, mai_mai_n1735_, mai_mai_n1736_, mai_mai_n1737_, mai_mai_n1738_, mai_mai_n1739_, mai_mai_n1740_, mai_mai_n1741_, mai_mai_n1742_, mai_mai_n1743_, mai_mai_n1744_, mai_mai_n1745_, mai_mai_n1746_, mai_mai_n1747_, mai_mai_n1748_, mai_mai_n1749_, mai_mai_n1750_, mai_mai_n1751_, mai_mai_n1752_, mai_mai_n1753_, mai_mai_n1754_, mai_mai_n1755_, mai_mai_n1756_, mai_mai_n1757_, mai_mai_n1758_, mai_mai_n1759_, mai_mai_n1760_, mai_mai_n1762_, mai_mai_n1763_, mai_mai_n1764_, mai_mai_n1765_, mai_mai_n1766_, mai_mai_n1767_, mai_mai_n1768_, mai_mai_n1769_, mai_mai_n1770_, mai_mai_n1771_, mai_mai_n1772_, mai_mai_n1773_, mai_mai_n1774_, mai_mai_n1775_, mai_mai_n1776_, mai_mai_n1777_, mai_mai_n1778_, mai_mai_n1779_, mai_mai_n1780_, mai_mai_n1781_, mai_mai_n1782_, mai_mai_n1783_, mai_mai_n1784_, mai_mai_n1785_, mai_mai_n1786_, mai_mai_n1787_, mai_mai_n1788_, mai_mai_n1789_, mai_mai_n1790_, mai_mai_n1791_, mai_mai_n1792_, mai_mai_n1793_, mai_mai_n1794_, mai_mai_n1795_, mai_mai_n1796_, mai_mai_n1797_, mai_mai_n1798_, mai_mai_n1799_, mai_mai_n1800_, mai_mai_n1801_, mai_mai_n1802_, mai_mai_n1803_, mai_mai_n1804_, mai_mai_n1805_, mai_mai_n1806_, mai_mai_n1807_, mai_mai_n1808_, mai_mai_n1809_, mai_mai_n1810_, mai_mai_n1811_, mai_mai_n1812_, mai_mai_n1813_, mai_mai_n1814_, mai_mai_n1815_, mai_mai_n1816_, mai_mai_n1817_, mai_mai_n1818_, mai_mai_n1820_, mai_mai_n1821_, mai_mai_n1822_, mai_mai_n1823_, mai_mai_n1824_, mai_mai_n1825_, mai_mai_n1826_, mai_mai_n1827_, mai_mai_n1828_, mai_mai_n1829_, mai_mai_n1830_, mai_mai_n1831_, mai_mai_n1832_, mai_mai_n1833_, mai_mai_n1834_, mai_mai_n1835_, mai_mai_n1836_, mai_mai_n1837_, mai_mai_n1838_, mai_mai_n1840_, mai_mai_n1841_, mai_mai_n1842_, mai_mai_n1843_, mai_mai_n1844_, mai_mai_n1845_, mai_mai_n1846_, mai_mai_n1847_, mai_mai_n1848_, mai_mai_n1849_, mai_mai_n1850_, mai_mai_n1851_, mai_mai_n1853_, mai_mai_n1854_, mai_mai_n1855_, mai_mai_n1856_, mai_mai_n1857_, mai_mai_n1858_, mai_mai_n1859_, mai_mai_n1860_, mai_mai_n1861_, mai_mai_n1862_, mai_mai_n1863_, mai_mai_n1864_, mai_mai_n1865_, mai_mai_n1866_, mai_mai_n1867_, mai_mai_n1868_, mai_mai_n1869_, mai_mai_n1871_, mai_mai_n1872_, mai_mai_n1873_, mai_mai_n1874_, mai_mai_n1875_, mai_mai_n1876_, mai_mai_n1877_, mai_mai_n1878_, mai_mai_n1879_, mai_mai_n1880_, mai_mai_n1881_, mai_mai_n1882_, mai_mai_n1883_, mai_mai_n1884_, mai_mai_n1885_, mai_mai_n1886_, mai_mai_n1887_, mai_mai_n1888_, mai_mai_n1889_, mai_mai_n1890_, mai_mai_n1891_, mai_mai_n1892_, mai_mai_n1893_, mai_mai_n1894_, mai_mai_n1895_, mai_mai_n1896_, mai_mai_n1897_, mai_mai_n1898_, mai_mai_n1899_, mai_mai_n1900_, mai_mai_n1901_, mai_mai_n1902_, mai_mai_n1903_, mai_mai_n1904_, mai_mai_n1905_, mai_mai_n1906_, mai_mai_n1907_, mai_mai_n1908_, mai_mai_n1909_, mai_mai_n1910_, mai_mai_n1911_, mai_mai_n1912_, mai_mai_n1913_, mai_mai_n1914_, mai_mai_n1916_, mai_mai_n1917_, mai_mai_n1918_, mai_mai_n1919_, mai_mai_n1920_, mai_mai_n1921_, mai_mai_n1922_, mai_mai_n1923_, mai_mai_n1924_, mai_mai_n1925_, mai_mai_n1926_, mai_mai_n1927_, mai_mai_n1928_, mai_mai_n1929_, mai_mai_n1930_, mai_mai_n1931_, mai_mai_n1933_, mai_mai_n1934_, mai_mai_n1935_, mai_mai_n1936_, mai_mai_n1937_, mai_mai_n1938_, mai_mai_n1939_, mai_mai_n1940_, mai_mai_n1941_, mai_mai_n1942_, mai_mai_n1943_, mai_mai_n1944_, mai_mai_n1945_, mai_mai_n1946_, mai_mai_n1947_, mai_mai_n1948_, mai_mai_n1949_, mai_mai_n1950_, mai_mai_n1951_, mai_mai_n1952_, mai_mai_n1953_, mai_mai_n1954_, mai_mai_n1955_, mai_mai_n1956_, mai_mai_n1957_, mai_mai_n1958_, mai_mai_n1959_, mai_mai_n1960_, mai_mai_n1961_, mai_mai_n1962_, mai_mai_n1963_, mai_mai_n1964_, mai_mai_n1965_, mai_mai_n1966_, mai_mai_n1967_, mai_mai_n1968_, mai_mai_n1969_, mai_mai_n1970_, mai_mai_n1971_, mai_mai_n1972_, mai_mai_n1973_, mai_mai_n1974_, mai_mai_n1975_, mai_mai_n1976_, mai_mai_n1977_, mai_mai_n1978_, mai_mai_n1979_, mai_mai_n1980_, mai_mai_n1981_, mai_mai_n1982_, mai_mai_n1983_, mai_mai_n1985_, mai_mai_n1986_, mai_mai_n1987_, mai_mai_n1988_, mai_mai_n1989_, mai_mai_n1990_, mai_mai_n1991_, mai_mai_n1992_, mai_mai_n1993_, mai_mai_n1994_, mai_mai_n1995_, mai_mai_n1996_, mai_mai_n1997_, mai_mai_n1998_, mai_mai_n1999_, mai_mai_n2000_, mai_mai_n2001_, mai_mai_n2002_, mai_mai_n2003_, mai_mai_n2004_, mai_mai_n2005_, mai_mai_n2006_, mai_mai_n2007_, mai_mai_n2008_, mai_mai_n2009_, mai_mai_n2010_, mai_mai_n2011_, mai_mai_n2012_, mai_mai_n2013_, mai_mai_n2014_, mai_mai_n2015_, mai_mai_n2016_, mai_mai_n2017_, mai_mai_n2018_, mai_mai_n2019_, mai_mai_n2020_, mai_mai_n2021_, mai_mai_n2022_, mai_mai_n2023_, mai_mai_n2024_, mai_mai_n2025_, mai_mai_n2026_, mai_mai_n2027_, mai_mai_n2028_, mai_mai_n2029_, mai_mai_n2030_, mai_mai_n2031_, mai_mai_n2032_, mai_mai_n2033_, mai_mai_n2034_, mai_mai_n2035_, mai_mai_n2036_, mai_mai_n2037_, mai_mai_n2038_, mai_mai_n2039_, mai_mai_n2040_, mai_mai_n2041_, mai_mai_n2042_, mai_mai_n2043_, mai_mai_n2044_, mai_mai_n2045_, mai_mai_n2046_, mai_mai_n2047_, mai_mai_n2048_, mai_mai_n2049_, mai_mai_n2050_, mai_mai_n2052_, mai_mai_n2053_, mai_mai_n2054_, mai_mai_n2055_, mai_mai_n2056_, mai_mai_n2057_, mai_mai_n2058_, mai_mai_n2059_, mai_mai_n2060_, mai_mai_n2061_, mai_mai_n2062_, mai_mai_n2063_, mai_mai_n2064_, mai_mai_n2065_, mai_mai_n2066_, mai_mai_n2067_, mai_mai_n2068_, mai_mai_n2069_, mai_mai_n2070_, mai_mai_n2071_, mai_mai_n2072_, mai_mai_n2073_, mai_mai_n2074_, mai_mai_n2075_, mai_mai_n2076_, mai_mai_n2077_, mai_mai_n2078_, mai_mai_n2079_, mai_mai_n2080_, mai_mai_n2081_, mai_mai_n2082_, mai_mai_n2083_, mai_mai_n2084_, mai_mai_n2085_, mai_mai_n2086_, mai_mai_n2087_, mai_mai_n2088_, mai_mai_n2089_, mai_mai_n2090_, mai_mai_n2091_, mai_mai_n2092_, mai_mai_n2093_, mai_mai_n2094_, mai_mai_n2095_, mai_mai_n2096_, mai_mai_n2097_, mai_mai_n2098_, mai_mai_n2099_, mai_mai_n2100_, mai_mai_n2101_, mai_mai_n2102_, mai_mai_n2103_, mai_mai_n2104_, mai_mai_n2105_, mai_mai_n2106_, mai_mai_n2107_, mai_mai_n2108_, mai_mai_n2109_, mai_mai_n2110_, mai_mai_n2111_, mai_mai_n2112_, mai_mai_n2113_, mai_mai_n2114_, mai_mai_n2115_, mai_mai_n2116_, mai_mai_n2117_, mai_mai_n2118_, mai_mai_n2119_, mai_mai_n2120_, mai_mai_n2121_, mai_mai_n2122_, mai_mai_n2123_, mai_mai_n2124_, mai_mai_n2125_, mai_mai_n2126_, mai_mai_n2127_, mai_mai_n2129_, mai_mai_n2130_, mai_mai_n2131_, mai_mai_n2132_, mai_mai_n2133_, mai_mai_n2134_, mai_mai_n2135_, mai_mai_n2136_, mai_mai_n2137_, mai_mai_n2138_, mai_mai_n2139_, mai_mai_n2140_, mai_mai_n2141_, mai_mai_n2142_, mai_mai_n2143_, mai_mai_n2144_, mai_mai_n2145_, mai_mai_n2146_, mai_mai_n2147_, mai_mai_n2148_, mai_mai_n2149_, mai_mai_n2150_, mai_mai_n2151_, mai_mai_n2152_, mai_mai_n2153_, mai_mai_n2154_, mai_mai_n2155_, mai_mai_n2156_, mai_mai_n2157_, mai_mai_n2158_, mai_mai_n2159_, mai_mai_n2160_, mai_mai_n2161_, mai_mai_n2162_, mai_mai_n2163_, mai_mai_n2164_, mai_mai_n2165_, mai_mai_n2166_, mai_mai_n2167_, mai_mai_n2168_, mai_mai_n2169_, mai_mai_n2170_, mai_mai_n2171_, mai_mai_n2172_, mai_mai_n2173_, mai_mai_n2174_, mai_mai_n2175_, mai_mai_n2176_, mai_mai_n2177_, mai_mai_n2178_, mai_mai_n2179_, mai_mai_n2180_, mai_mai_n2181_, mai_mai_n2182_, mai_mai_n2183_, mai_mai_n2184_, mai_mai_n2185_, mai_mai_n2186_, mai_mai_n2187_, mai_mai_n2188_, mai_mai_n2189_, mai_mai_n2190_, mai_mai_n2191_, mai_mai_n2192_, mai_mai_n2193_, mai_mai_n2194_, mai_mai_n2195_, mai_mai_n2196_, mai_mai_n2197_, mai_mai_n2198_, mai_mai_n2199_, mai_mai_n2200_, mai_mai_n2201_, mai_mai_n2203_, mai_mai_n2204_, mai_mai_n2205_, mai_mai_n2206_, mai_mai_n2207_, mai_mai_n2208_, mai_mai_n2209_, mai_mai_n2210_, mai_mai_n2211_, mai_mai_n2212_, mai_mai_n2213_, mai_mai_n2214_, mai_mai_n2215_, mai_mai_n2216_, mai_mai_n2217_, mai_mai_n2218_, mai_mai_n2219_, mai_mai_n2220_, mai_mai_n2221_, mai_mai_n2222_, mai_mai_n2223_, mai_mai_n2224_, mai_mai_n2225_, mai_mai_n2226_, mai_mai_n2227_, mai_mai_n2228_, mai_mai_n2229_, mai_mai_n2230_, mai_mai_n2231_, mai_mai_n2232_, mai_mai_n2233_, mai_mai_n2234_, mai_mai_n2235_, mai_mai_n2236_, mai_mai_n2237_, mai_mai_n2238_, mai_mai_n2239_, mai_mai_n2240_, mai_mai_n2241_, mai_mai_n2242_, mai_mai_n2243_, mai_mai_n2244_, mai_mai_n2245_, mai_mai_n2246_, mai_mai_n2247_, mai_mai_n2248_, mai_mai_n2249_, mai_mai_n2250_, mai_mai_n2251_, mai_mai_n2252_, mai_mai_n2253_, mai_mai_n2254_, mai_mai_n2255_, mai_mai_n2256_, mai_mai_n2257_, mai_mai_n2258_, mai_mai_n2259_, mai_mai_n2260_, mai_mai_n2261_, mai_mai_n2262_, mai_mai_n2263_, mai_mai_n2264_, mai_mai_n2265_, mai_mai_n2266_, mai_mai_n2267_, mai_mai_n2268_, mai_mai_n2269_, mai_mai_n2270_, mai_mai_n2271_, mai_mai_n2272_, mai_mai_n2273_, mai_mai_n2274_, mai_mai_n2275_, mai_mai_n2276_, mai_mai_n2277_, mai_mai_n2278_, mai_mai_n2279_, mai_mai_n2280_, mai_mai_n2282_, mai_mai_n2283_, mai_mai_n2284_, mai_mai_n2285_, mai_mai_n2286_, mai_mai_n2287_, mai_mai_n2288_, mai_mai_n2289_, mai_mai_n2290_, mai_mai_n2291_, mai_mai_n2292_, mai_mai_n2293_, mai_mai_n2294_, mai_mai_n2295_, mai_mai_n2296_, mai_mai_n2297_, mai_mai_n2298_, mai_mai_n2299_, mai_mai_n2300_, mai_mai_n2301_, mai_mai_n2302_, mai_mai_n2303_, mai_mai_n2304_, mai_mai_n2305_, mai_mai_n2306_, mai_mai_n2307_, mai_mai_n2308_, mai_mai_n2309_, mai_mai_n2310_, mai_mai_n2311_, mai_mai_n2312_, mai_mai_n2313_, mai_mai_n2314_, mai_mai_n2315_, mai_mai_n2316_, mai_mai_n2317_, mai_mai_n2318_, mai_mai_n2319_, mai_mai_n2320_, mai_mai_n2321_, mai_mai_n2322_, mai_mai_n2323_, mai_mai_n2324_, mai_mai_n2325_, mai_mai_n2326_, mai_mai_n2327_, mai_mai_n2328_, mai_mai_n2329_, mai_mai_n2330_, mai_mai_n2331_, mai_mai_n2332_, mai_mai_n2333_, mai_mai_n2334_, mai_mai_n2335_, mai_mai_n2336_, mai_mai_n2337_, mai_mai_n2338_, mai_mai_n2339_, mai_mai_n2340_, mai_mai_n2341_, mai_mai_n2342_, mai_mai_n2343_, mai_mai_n2344_, mai_mai_n2345_, mai_mai_n2346_, mai_mai_n2347_, mai_mai_n2348_, mai_mai_n2350_, mai_mai_n2351_, mai_mai_n2352_, mai_mai_n2353_, mai_mai_n2354_, mai_mai_n2355_, mai_mai_n2356_, mai_mai_n2357_, mai_mai_n2358_, mai_mai_n2359_, mai_mai_n2360_, mai_mai_n2361_, mai_mai_n2362_, mai_mai_n2363_, mai_mai_n2364_, mai_mai_n2365_, mai_mai_n2366_, mai_mai_n2367_, mai_mai_n2368_, mai_mai_n2369_, mai_mai_n2370_, mai_mai_n2371_, mai_mai_n2372_, mai_mai_n2373_, mai_mai_n2374_, mai_mai_n2375_, mai_mai_n2376_, mai_mai_n2377_, mai_mai_n2378_, mai_mai_n2379_, mai_mai_n2380_, mai_mai_n2381_, mai_mai_n2382_, mai_mai_n2383_, mai_mai_n2384_, mai_mai_n2385_, mai_mai_n2386_, mai_mai_n2387_, mai_mai_n2388_, mai_mai_n2389_, mai_mai_n2390_, mai_mai_n2391_, mai_mai_n2392_, mai_mai_n2393_, mai_mai_n2394_, mai_mai_n2395_, mai_mai_n2396_, mai_mai_n2397_, mai_mai_n2398_, mai_mai_n2399_, mai_mai_n2400_, mai_mai_n2401_, mai_mai_n2402_, mai_mai_n2403_, mai_mai_n2404_, mai_mai_n2405_, mai_mai_n2406_, mai_mai_n2407_, mai_mai_n2408_, mai_mai_n2409_, mai_mai_n2410_, mai_mai_n2411_, mai_mai_n2413_, mai_mai_n2414_, mai_mai_n2415_, mai_mai_n2416_, mai_mai_n2417_, mai_mai_n2418_, mai_mai_n2419_, mai_mai_n2420_, mai_mai_n2421_, mai_mai_n2422_, mai_mai_n2423_, mai_mai_n2424_, mai_mai_n2425_, mai_mai_n2426_, mai_mai_n2427_, mai_mai_n2428_, mai_mai_n2429_, mai_mai_n2430_, mai_mai_n2431_, mai_mai_n2432_, mai_mai_n2433_, mai_mai_n2434_, mai_mai_n2435_, mai_mai_n2436_, mai_mai_n2437_, mai_mai_n2438_, mai_mai_n2439_, mai_mai_n2440_, mai_mai_n2441_, mai_mai_n2442_, mai_mai_n2443_, mai_mai_n2444_, mai_mai_n2445_, mai_mai_n2446_, mai_mai_n2447_, mai_mai_n2448_, mai_mai_n2449_, mai_mai_n2450_, mai_mai_n2451_, mai_mai_n2452_, mai_mai_n2453_, mai_mai_n2454_, mai_mai_n2455_, mai_mai_n2456_, mai_mai_n2457_, mai_mai_n2458_, mai_mai_n2459_, mai_mai_n2460_, mai_mai_n2461_, mai_mai_n2462_, mai_mai_n2463_, mai_mai_n2464_, mai_mai_n2465_, mai_mai_n2466_, mai_mai_n2467_, mai_mai_n2468_, mai_mai_n2469_, mai_mai_n2470_, mai_mai_n2471_, mai_mai_n2472_, mai_mai_n2473_, mai_mai_n2474_, mai_mai_n2475_, mai_mai_n2476_, mai_mai_n2477_, mai_mai_n2478_, mai_mai_n2479_, mai_mai_n2480_, mai_mai_n2481_, mai_mai_n2482_, mai_mai_n2483_, mai_mai_n2484_, mai_mai_n2485_, mai_mai_n2486_, mai_mai_n2487_, mai_mai_n2488_, mai_mai_n2489_, mai_mai_n2490_, mai_mai_n2492_, mai_mai_n2493_, mai_mai_n2494_, mai_mai_n2495_, mai_mai_n2496_, mai_mai_n2497_, mai_mai_n2498_, mai_mai_n2499_, mai_mai_n2500_, mai_mai_n2501_, mai_mai_n2502_, mai_mai_n2503_, mai_mai_n2504_, mai_mai_n2505_, mai_mai_n2506_, mai_mai_n2507_, mai_mai_n2508_, mai_mai_n2509_, mai_mai_n2510_, mai_mai_n2511_, mai_mai_n2512_, mai_mai_n2513_, mai_mai_n2514_, mai_mai_n2515_, mai_mai_n2516_, mai_mai_n2517_, mai_mai_n2518_, mai_mai_n2519_, mai_mai_n2520_, mai_mai_n2521_, mai_mai_n2522_, mai_mai_n2523_, mai_mai_n2524_, mai_mai_n2525_, mai_mai_n2526_, mai_mai_n2527_, mai_mai_n2528_, mai_mai_n2529_, mai_mai_n2530_, mai_mai_n2531_, mai_mai_n2532_, mai_mai_n2533_, mai_mai_n2534_, mai_mai_n2535_, mai_mai_n2536_, mai_mai_n2537_, mai_mai_n2538_, mai_mai_n2539_, mai_mai_n2540_, mai_mai_n2541_, mai_mai_n2542_, mai_mai_n2543_, mai_mai_n2544_, mai_mai_n2545_, mai_mai_n2546_, mai_mai_n2547_, mai_mai_n2548_, mai_mai_n2549_, mai_mai_n2550_, mai_mai_n2551_, mai_mai_n2552_, mai_mai_n2553_, mai_mai_n2555_, mai_mai_n2556_, mai_mai_n2557_, mai_mai_n2558_, mai_mai_n2559_, mai_mai_n2560_, mai_mai_n2561_, mai_mai_n2562_, mai_mai_n2563_, mai_mai_n2564_, mai_mai_n2565_, mai_mai_n2566_, mai_mai_n2567_, mai_mai_n2568_, mai_mai_n2569_, mai_mai_n2570_, mai_mai_n2571_, mai_mai_n2572_, mai_mai_n2573_, mai_mai_n2574_, mai_mai_n2575_, mai_mai_n2576_, mai_mai_n2577_, mai_mai_n2578_, mai_mai_n2579_, mai_mai_n2580_, mai_mai_n2581_, mai_mai_n2582_, mai_mai_n2583_, mai_mai_n2584_, mai_mai_n2585_, mai_mai_n2586_, mai_mai_n2587_, mai_mai_n2588_, mai_mai_n2589_, mai_mai_n2590_, mai_mai_n2591_, mai_mai_n2592_, mai_mai_n2593_, mai_mai_n2594_, mai_mai_n2595_, mai_mai_n2596_, mai_mai_n2597_, mai_mai_n2598_, mai_mai_n2599_, mai_mai_n2600_, mai_mai_n2601_, mai_mai_n2602_, mai_mai_n2603_, mai_mai_n2604_, mai_mai_n2605_, mai_mai_n2606_, mai_mai_n2607_, mai_mai_n2608_, mai_mai_n2609_, mai_mai_n2610_, mai_mai_n2611_, mai_mai_n2612_, mai_mai_n2613_, mai_mai_n2614_, mai_mai_n2615_, mai_mai_n2616_, mai_mai_n2617_, mai_mai_n2618_, mai_mai_n2619_, mai_mai_n2620_, mai_mai_n2621_, mai_mai_n2622_, mai_mai_n2623_, mai_mai_n2624_, mai_mai_n2626_, mai_mai_n2627_, mai_mai_n2628_, mai_mai_n2629_, mai_mai_n2630_, mai_mai_n2631_, mai_mai_n2632_, mai_mai_n2633_, mai_mai_n2634_, mai_mai_n2635_, mai_mai_n2636_, mai_mai_n2637_, mai_mai_n2638_, mai_mai_n2639_, mai_mai_n2640_, mai_mai_n2641_, mai_mai_n2642_, mai_mai_n2643_, mai_mai_n2644_, mai_mai_n2645_, mai_mai_n2646_, mai_mai_n2647_, mai_mai_n2648_, mai_mai_n2649_, mai_mai_n2650_, mai_mai_n2651_, mai_mai_n2652_, mai_mai_n2653_, mai_mai_n2654_, mai_mai_n2655_, mai_mai_n2656_, mai_mai_n2657_, mai_mai_n2658_, mai_mai_n2659_, mai_mai_n2660_, mai_mai_n2661_, mai_mai_n2662_, mai_mai_n2663_, mai_mai_n2664_, mai_mai_n2665_, mai_mai_n2666_, mai_mai_n2667_, mai_mai_n2668_, mai_mai_n2669_, mai_mai_n2670_, mai_mai_n2671_, mai_mai_n2672_, mai_mai_n2673_, mai_mai_n2674_, mai_mai_n2675_, mai_mai_n2676_, mai_mai_n2677_, mai_mai_n2678_, mai_mai_n2679_, mai_mai_n2680_, mai_mai_n2681_, mai_mai_n2682_, mai_mai_n2683_, mai_mai_n2684_, mai_mai_n2685_, mai_mai_n2686_, mai_mai_n2687_, mai_mai_n2688_, mai_mai_n2689_, mai_mai_n2690_, mai_mai_n2691_, mai_mai_n2692_, mai_mai_n2696_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1618_, men_men_n1619_, men_men_n1620_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, men_men_n1632_, men_men_n1633_, men_men_n1634_, men_men_n1635_, men_men_n1636_, men_men_n1637_, men_men_n1638_, men_men_n1639_, men_men_n1640_, men_men_n1641_, men_men_n1642_, men_men_n1643_, men_men_n1644_, men_men_n1645_, men_men_n1646_, men_men_n1647_, men_men_n1649_, men_men_n1650_, men_men_n1651_, men_men_n1652_, men_men_n1653_, men_men_n1654_, men_men_n1655_, men_men_n1656_, men_men_n1657_, men_men_n1658_, men_men_n1659_, men_men_n1660_, men_men_n1661_, men_men_n1662_, men_men_n1663_, men_men_n1664_, men_men_n1665_, men_men_n1666_, men_men_n1667_, men_men_n1668_, men_men_n1669_, men_men_n1670_, men_men_n1671_, men_men_n1672_, men_men_n1673_, men_men_n1674_, men_men_n1676_, men_men_n1677_, men_men_n1678_, men_men_n1679_, men_men_n1680_, men_men_n1681_, men_men_n1682_, men_men_n1683_, men_men_n1684_, men_men_n1685_, men_men_n1686_, men_men_n1687_, men_men_n1688_, men_men_n1689_, men_men_n1690_, men_men_n1691_, men_men_n1692_, men_men_n1693_, men_men_n1694_, men_men_n1695_, men_men_n1696_, men_men_n1697_, men_men_n1698_, men_men_n1699_, men_men_n1700_, men_men_n1701_, men_men_n1702_, men_men_n1703_, men_men_n1704_, men_men_n1705_, men_men_n1706_, men_men_n1707_, men_men_n1708_, men_men_n1709_, men_men_n1710_, men_men_n1711_, men_men_n1712_, men_men_n1713_, men_men_n1714_, men_men_n1715_, men_men_n1716_, men_men_n1717_, men_men_n1718_, men_men_n1719_, men_men_n1720_, men_men_n1721_, men_men_n1722_, men_men_n1723_, men_men_n1724_, men_men_n1725_, men_men_n1726_, men_men_n1727_, men_men_n1728_, men_men_n1729_, men_men_n1730_, men_men_n1731_, men_men_n1732_, men_men_n1733_, men_men_n1734_, men_men_n1735_, men_men_n1736_, men_men_n1737_, men_men_n1738_, men_men_n1739_, men_men_n1740_, men_men_n1741_, men_men_n1742_, men_men_n1743_, men_men_n1744_, men_men_n1745_, men_men_n1746_, men_men_n1747_, men_men_n1748_, men_men_n1749_, men_men_n1750_, men_men_n1751_, men_men_n1752_, men_men_n1753_, men_men_n1754_, men_men_n1755_, men_men_n1756_, men_men_n1757_, men_men_n1758_, men_men_n1759_, men_men_n1760_, men_men_n1761_, men_men_n1762_, men_men_n1764_, men_men_n1765_, men_men_n1766_, men_men_n1767_, men_men_n1768_, men_men_n1769_, men_men_n1770_, men_men_n1771_, men_men_n1772_, men_men_n1773_, men_men_n1774_, men_men_n1775_, men_men_n1776_, men_men_n1777_, men_men_n1778_, men_men_n1779_, men_men_n1780_, men_men_n1781_, men_men_n1782_, men_men_n1783_, men_men_n1784_, men_men_n1785_, men_men_n1786_, men_men_n1787_, men_men_n1788_, men_men_n1789_, men_men_n1790_, men_men_n1791_, men_men_n1792_, men_men_n1793_, men_men_n1794_, men_men_n1795_, men_men_n1796_, men_men_n1797_, men_men_n1798_, men_men_n1799_, men_men_n1800_, men_men_n1801_, men_men_n1802_, men_men_n1803_, men_men_n1804_, men_men_n1805_, men_men_n1806_, men_men_n1807_, men_men_n1808_, men_men_n1809_, men_men_n1810_, men_men_n1811_, men_men_n1812_, men_men_n1813_, men_men_n1814_, men_men_n1815_, men_men_n1816_, men_men_n1817_, men_men_n1818_, men_men_n1819_, men_men_n1820_, men_men_n1822_, men_men_n1823_, men_men_n1824_, men_men_n1825_, men_men_n1826_, men_men_n1827_, men_men_n1828_, men_men_n1829_, men_men_n1830_, men_men_n1831_, men_men_n1832_, men_men_n1833_, men_men_n1834_, men_men_n1835_, men_men_n1836_, men_men_n1837_, men_men_n1838_, men_men_n1839_, men_men_n1840_, men_men_n1842_, men_men_n1843_, men_men_n1844_, men_men_n1845_, men_men_n1846_, men_men_n1847_, men_men_n1848_, men_men_n1849_, men_men_n1850_, men_men_n1851_, men_men_n1852_, men_men_n1853_, men_men_n1854_, men_men_n1856_, men_men_n1857_, men_men_n1858_, men_men_n1859_, men_men_n1860_, men_men_n1861_, men_men_n1862_, men_men_n1863_, men_men_n1864_, men_men_n1865_, men_men_n1866_, men_men_n1867_, men_men_n1868_, men_men_n1869_, men_men_n1870_, men_men_n1871_, men_men_n1872_, men_men_n1874_, men_men_n1875_, men_men_n1876_, men_men_n1877_, men_men_n1878_, men_men_n1879_, men_men_n1880_, men_men_n1881_, men_men_n1882_, men_men_n1883_, men_men_n1884_, men_men_n1885_, men_men_n1886_, men_men_n1887_, men_men_n1888_, men_men_n1889_, men_men_n1890_, men_men_n1891_, men_men_n1892_, men_men_n1893_, men_men_n1894_, men_men_n1895_, men_men_n1896_, men_men_n1897_, men_men_n1898_, men_men_n1899_, men_men_n1900_, men_men_n1901_, men_men_n1902_, men_men_n1903_, men_men_n1904_, men_men_n1905_, men_men_n1906_, men_men_n1907_, men_men_n1908_, men_men_n1909_, men_men_n1910_, men_men_n1911_, men_men_n1912_, men_men_n1913_, men_men_n1914_, men_men_n1915_, men_men_n1916_, men_men_n1917_, men_men_n1918_, men_men_n1919_, men_men_n1920_, men_men_n1922_, men_men_n1923_, men_men_n1924_, men_men_n1925_, men_men_n1926_, men_men_n1927_, men_men_n1928_, men_men_n1929_, men_men_n1930_, men_men_n1931_, men_men_n1932_, men_men_n1933_, men_men_n1934_, men_men_n1935_, men_men_n1936_, men_men_n1937_, men_men_n1939_, men_men_n1940_, men_men_n1941_, men_men_n1942_, men_men_n1943_, men_men_n1944_, men_men_n1945_, men_men_n1946_, men_men_n1947_, men_men_n1948_, men_men_n1949_, men_men_n1950_, men_men_n1951_, men_men_n1952_, men_men_n1953_, men_men_n1954_, men_men_n1955_, men_men_n1956_, men_men_n1957_, men_men_n1958_, men_men_n1959_, men_men_n1960_, men_men_n1961_, men_men_n1962_, men_men_n1963_, men_men_n1964_, men_men_n1965_, men_men_n1966_, men_men_n1967_, men_men_n1968_, men_men_n1969_, men_men_n1970_, men_men_n1971_, men_men_n1972_, men_men_n1973_, men_men_n1974_, men_men_n1975_, men_men_n1976_, men_men_n1977_, men_men_n1978_, men_men_n1979_, men_men_n1980_, men_men_n1981_, men_men_n1982_, men_men_n1983_, men_men_n1984_, men_men_n1985_, men_men_n1986_, men_men_n1987_, men_men_n1988_, men_men_n1989_, men_men_n1991_, men_men_n1992_, men_men_n1993_, men_men_n1994_, men_men_n1995_, men_men_n1996_, men_men_n1997_, men_men_n1998_, men_men_n1999_, men_men_n2000_, men_men_n2001_, men_men_n2002_, men_men_n2003_, men_men_n2004_, men_men_n2005_, men_men_n2006_, men_men_n2007_, men_men_n2008_, men_men_n2009_, men_men_n2010_, men_men_n2011_, men_men_n2012_, men_men_n2013_, men_men_n2014_, men_men_n2015_, men_men_n2016_, men_men_n2017_, men_men_n2018_, men_men_n2019_, men_men_n2020_, men_men_n2021_, men_men_n2022_, men_men_n2023_, men_men_n2024_, men_men_n2025_, men_men_n2026_, men_men_n2027_, men_men_n2028_, men_men_n2029_, men_men_n2030_, men_men_n2031_, men_men_n2032_, men_men_n2033_, men_men_n2034_, men_men_n2035_, men_men_n2036_, men_men_n2037_, men_men_n2038_, men_men_n2039_, men_men_n2040_, men_men_n2041_, men_men_n2042_, men_men_n2043_, men_men_n2044_, men_men_n2045_, men_men_n2046_, men_men_n2047_, men_men_n2048_, men_men_n2049_, men_men_n2050_, men_men_n2051_, men_men_n2052_, men_men_n2053_, men_men_n2054_, men_men_n2055_, men_men_n2056_, men_men_n2058_, men_men_n2059_, men_men_n2060_, men_men_n2061_, men_men_n2062_, men_men_n2063_, men_men_n2064_, men_men_n2065_, men_men_n2066_, men_men_n2067_, men_men_n2068_, men_men_n2069_, men_men_n2070_, men_men_n2071_, men_men_n2072_, men_men_n2073_, men_men_n2074_, men_men_n2075_, men_men_n2076_, men_men_n2077_, men_men_n2078_, men_men_n2079_, men_men_n2080_, men_men_n2081_, men_men_n2082_, men_men_n2083_, men_men_n2084_, men_men_n2085_, men_men_n2086_, men_men_n2087_, men_men_n2088_, men_men_n2089_, men_men_n2090_, men_men_n2091_, men_men_n2092_, men_men_n2093_, men_men_n2094_, men_men_n2095_, men_men_n2096_, men_men_n2097_, men_men_n2098_, men_men_n2099_, men_men_n2100_, men_men_n2101_, men_men_n2102_, men_men_n2103_, men_men_n2104_, men_men_n2105_, men_men_n2106_, men_men_n2107_, men_men_n2108_, men_men_n2109_, men_men_n2110_, men_men_n2111_, men_men_n2112_, men_men_n2113_, men_men_n2114_, men_men_n2115_, men_men_n2116_, men_men_n2117_, men_men_n2118_, men_men_n2119_, men_men_n2120_, men_men_n2121_, men_men_n2122_, men_men_n2123_, men_men_n2124_, men_men_n2125_, men_men_n2126_, men_men_n2127_, men_men_n2128_, men_men_n2129_, men_men_n2130_, men_men_n2131_, men_men_n2132_, men_men_n2134_, men_men_n2135_, men_men_n2136_, men_men_n2137_, men_men_n2138_, men_men_n2139_, men_men_n2140_, men_men_n2141_, men_men_n2142_, men_men_n2143_, men_men_n2144_, men_men_n2145_, men_men_n2146_, men_men_n2147_, men_men_n2148_, men_men_n2149_, men_men_n2150_, men_men_n2151_, men_men_n2152_, men_men_n2153_, men_men_n2154_, men_men_n2155_, men_men_n2156_, men_men_n2157_, men_men_n2158_, men_men_n2159_, men_men_n2160_, men_men_n2161_, men_men_n2162_, men_men_n2163_, men_men_n2164_, men_men_n2165_, men_men_n2166_, men_men_n2167_, men_men_n2168_, men_men_n2169_, men_men_n2170_, men_men_n2171_, men_men_n2172_, men_men_n2173_, men_men_n2174_, men_men_n2175_, men_men_n2176_, men_men_n2177_, men_men_n2178_, men_men_n2179_, men_men_n2180_, men_men_n2181_, men_men_n2182_, men_men_n2183_, men_men_n2184_, men_men_n2185_, men_men_n2186_, men_men_n2187_, men_men_n2188_, men_men_n2189_, men_men_n2190_, men_men_n2191_, men_men_n2192_, men_men_n2193_, men_men_n2194_, men_men_n2195_, men_men_n2196_, men_men_n2197_, men_men_n2198_, men_men_n2199_, men_men_n2200_, men_men_n2201_, men_men_n2202_, men_men_n2203_, men_men_n2204_, men_men_n2205_, men_men_n2206_, men_men_n2207_, men_men_n2208_, men_men_n2210_, men_men_n2211_, men_men_n2212_, men_men_n2213_, men_men_n2214_, men_men_n2215_, men_men_n2216_, men_men_n2217_, men_men_n2218_, men_men_n2219_, men_men_n2220_, men_men_n2221_, men_men_n2222_, men_men_n2223_, men_men_n2224_, men_men_n2225_, men_men_n2226_, men_men_n2227_, men_men_n2228_, men_men_n2229_, men_men_n2230_, men_men_n2231_, men_men_n2232_, men_men_n2233_, men_men_n2234_, men_men_n2235_, men_men_n2236_, men_men_n2237_, men_men_n2238_, men_men_n2239_, men_men_n2240_, men_men_n2241_, men_men_n2242_, men_men_n2243_, men_men_n2244_, men_men_n2245_, men_men_n2246_, men_men_n2247_, men_men_n2248_, men_men_n2249_, men_men_n2250_, men_men_n2251_, men_men_n2252_, men_men_n2253_, men_men_n2254_, men_men_n2255_, men_men_n2256_, men_men_n2257_, men_men_n2258_, men_men_n2259_, men_men_n2260_, men_men_n2261_, men_men_n2262_, men_men_n2263_, men_men_n2264_, men_men_n2265_, men_men_n2266_, men_men_n2267_, men_men_n2268_, men_men_n2269_, men_men_n2270_, men_men_n2271_, men_men_n2272_, men_men_n2273_, men_men_n2274_, men_men_n2275_, men_men_n2276_, men_men_n2277_, men_men_n2278_, men_men_n2279_, men_men_n2280_, men_men_n2281_, men_men_n2282_, men_men_n2283_, men_men_n2284_, men_men_n2285_, men_men_n2286_, men_men_n2287_, men_men_n2289_, men_men_n2290_, men_men_n2291_, men_men_n2292_, men_men_n2293_, men_men_n2294_, men_men_n2295_, men_men_n2296_, men_men_n2297_, men_men_n2298_, men_men_n2299_, men_men_n2300_, men_men_n2301_, men_men_n2302_, men_men_n2303_, men_men_n2304_, men_men_n2305_, men_men_n2306_, men_men_n2307_, men_men_n2308_, men_men_n2309_, men_men_n2310_, men_men_n2311_, men_men_n2312_, men_men_n2313_, men_men_n2314_, men_men_n2315_, men_men_n2316_, men_men_n2317_, men_men_n2318_, men_men_n2319_, men_men_n2320_, men_men_n2321_, men_men_n2322_, men_men_n2323_, men_men_n2324_, men_men_n2325_, men_men_n2326_, men_men_n2327_, men_men_n2328_, men_men_n2329_, men_men_n2330_, men_men_n2331_, men_men_n2332_, men_men_n2333_, men_men_n2334_, men_men_n2335_, men_men_n2336_, men_men_n2337_, men_men_n2338_, men_men_n2339_, men_men_n2340_, men_men_n2341_, men_men_n2342_, men_men_n2343_, men_men_n2344_, men_men_n2345_, men_men_n2346_, men_men_n2347_, men_men_n2348_, men_men_n2349_, men_men_n2350_, men_men_n2351_, men_men_n2352_, men_men_n2353_, men_men_n2354_, men_men_n2356_, men_men_n2357_, men_men_n2358_, men_men_n2359_, men_men_n2360_, men_men_n2361_, men_men_n2362_, men_men_n2363_, men_men_n2364_, men_men_n2365_, men_men_n2366_, men_men_n2367_, men_men_n2368_, men_men_n2369_, men_men_n2370_, men_men_n2371_, men_men_n2372_, men_men_n2373_, men_men_n2374_, men_men_n2375_, men_men_n2376_, men_men_n2377_, men_men_n2378_, men_men_n2379_, men_men_n2380_, men_men_n2381_, men_men_n2382_, men_men_n2383_, men_men_n2384_, men_men_n2385_, men_men_n2386_, men_men_n2387_, men_men_n2388_, men_men_n2389_, men_men_n2390_, men_men_n2391_, men_men_n2392_, men_men_n2393_, men_men_n2394_, men_men_n2395_, men_men_n2396_, men_men_n2397_, men_men_n2398_, men_men_n2399_, men_men_n2400_, men_men_n2401_, men_men_n2402_, men_men_n2403_, men_men_n2404_, men_men_n2405_, men_men_n2406_, men_men_n2407_, men_men_n2408_, men_men_n2409_, men_men_n2410_, men_men_n2411_, men_men_n2412_, men_men_n2413_, men_men_n2414_, men_men_n2415_, men_men_n2417_, men_men_n2418_, men_men_n2419_, men_men_n2420_, men_men_n2421_, men_men_n2422_, men_men_n2423_, men_men_n2424_, men_men_n2425_, men_men_n2426_, men_men_n2427_, men_men_n2428_, men_men_n2429_, men_men_n2430_, men_men_n2431_, men_men_n2432_, men_men_n2433_, men_men_n2434_, men_men_n2435_, men_men_n2436_, men_men_n2437_, men_men_n2438_, men_men_n2439_, men_men_n2440_, men_men_n2441_, men_men_n2442_, men_men_n2443_, men_men_n2444_, men_men_n2445_, men_men_n2446_, men_men_n2447_, men_men_n2448_, men_men_n2449_, men_men_n2450_, men_men_n2451_, men_men_n2452_, men_men_n2453_, men_men_n2454_, men_men_n2455_, men_men_n2456_, men_men_n2457_, men_men_n2458_, men_men_n2459_, men_men_n2460_, men_men_n2461_, men_men_n2462_, men_men_n2463_, men_men_n2464_, men_men_n2465_, men_men_n2466_, men_men_n2467_, men_men_n2468_, men_men_n2469_, men_men_n2470_, men_men_n2471_, men_men_n2472_, men_men_n2473_, men_men_n2474_, men_men_n2475_, men_men_n2476_, men_men_n2477_, men_men_n2478_, men_men_n2479_, men_men_n2480_, men_men_n2481_, men_men_n2482_, men_men_n2483_, men_men_n2484_, men_men_n2485_, men_men_n2486_, men_men_n2487_, men_men_n2488_, men_men_n2489_, men_men_n2490_, men_men_n2491_, men_men_n2492_, men_men_n2493_, men_men_n2495_, men_men_n2496_, men_men_n2497_, men_men_n2498_, men_men_n2499_, men_men_n2500_, men_men_n2501_, men_men_n2502_, men_men_n2503_, men_men_n2504_, men_men_n2505_, men_men_n2506_, men_men_n2507_, men_men_n2508_, men_men_n2509_, men_men_n2510_, men_men_n2511_, men_men_n2512_, men_men_n2513_, men_men_n2514_, men_men_n2515_, men_men_n2516_, men_men_n2517_, men_men_n2518_, men_men_n2519_, men_men_n2520_, men_men_n2521_, men_men_n2522_, men_men_n2523_, men_men_n2524_, men_men_n2525_, men_men_n2526_, men_men_n2527_, men_men_n2528_, men_men_n2529_, men_men_n2530_, men_men_n2531_, men_men_n2532_, men_men_n2533_, men_men_n2534_, men_men_n2535_, men_men_n2536_, men_men_n2537_, men_men_n2538_, men_men_n2539_, men_men_n2540_, men_men_n2541_, men_men_n2542_, men_men_n2543_, men_men_n2544_, men_men_n2545_, men_men_n2546_, men_men_n2547_, men_men_n2548_, men_men_n2549_, men_men_n2550_, men_men_n2551_, men_men_n2552_, men_men_n2553_, men_men_n2554_, men_men_n2555_, men_men_n2556_, men_men_n2557_, men_men_n2559_, men_men_n2560_, men_men_n2561_, men_men_n2562_, men_men_n2563_, men_men_n2564_, men_men_n2565_, men_men_n2566_, men_men_n2567_, men_men_n2568_, men_men_n2569_, men_men_n2570_, men_men_n2571_, men_men_n2572_, men_men_n2573_, men_men_n2574_, men_men_n2575_, men_men_n2576_, men_men_n2577_, men_men_n2578_, men_men_n2579_, men_men_n2580_, men_men_n2581_, men_men_n2582_, men_men_n2583_, men_men_n2584_, men_men_n2585_, men_men_n2586_, men_men_n2587_, men_men_n2588_, men_men_n2589_, men_men_n2590_, men_men_n2591_, men_men_n2592_, men_men_n2593_, men_men_n2594_, men_men_n2595_, men_men_n2596_, men_men_n2597_, men_men_n2598_, men_men_n2599_, men_men_n2600_, men_men_n2601_, men_men_n2602_, men_men_n2603_, men_men_n2604_, men_men_n2605_, men_men_n2606_, men_men_n2607_, men_men_n2608_, men_men_n2609_, men_men_n2610_, men_men_n2611_, men_men_n2612_, men_men_n2613_, men_men_n2614_, men_men_n2615_, men_men_n2616_, men_men_n2617_, men_men_n2618_, men_men_n2619_, men_men_n2620_, men_men_n2621_, men_men_n2622_, men_men_n2623_, men_men_n2624_, men_men_n2625_, men_men_n2627_, men_men_n2628_, men_men_n2629_, men_men_n2630_, men_men_n2631_, men_men_n2632_, men_men_n2633_, men_men_n2634_, men_men_n2635_, men_men_n2636_, men_men_n2637_, men_men_n2638_, men_men_n2639_, men_men_n2640_, men_men_n2641_, men_men_n2642_, men_men_n2643_, men_men_n2644_, men_men_n2645_, men_men_n2646_, men_men_n2647_, men_men_n2648_, men_men_n2649_, men_men_n2650_, men_men_n2651_, men_men_n2652_, men_men_n2653_, men_men_n2654_, men_men_n2655_, men_men_n2656_, men_men_n2657_, men_men_n2658_, men_men_n2659_, men_men_n2660_, men_men_n2661_, men_men_n2662_, men_men_n2663_, men_men_n2664_, men_men_n2665_, men_men_n2666_, men_men_n2667_, men_men_n2668_, men_men_n2669_, men_men_n2670_, men_men_n2671_, men_men_n2672_, men_men_n2673_, men_men_n2674_, men_men_n2675_, men_men_n2676_, men_men_n2677_, men_men_n2678_, men_men_n2679_, men_men_n2680_, men_men_n2681_, men_men_n2682_, men_men_n2683_, men_men_n2684_, men_men_n2685_, men_men_n2686_, men_men_n2687_, men_men_n2688_, men_men_n2689_, men_men_n2690_, men_men_n2691_, men_men_n2692_, men_men_n2696_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13, ori14, mai14, men14, ori15, mai15, men15, ori16, mai16, men16, ori17, mai17, men17, ori18, mai18, men18, ori19, mai19, men19, ori20, mai20, men20, ori21, mai21, men21, ori22, mai22, men22, ori23, mai23, men23, ori24, mai24, men24, ori25, mai25, men25, ori26, mai26, men26, ori27, mai27, men27, ori28, mai28, men28, ori29, mai29, men29, ori30, mai30, men30, ori31, mai31, men31, ori32, mai32, men32, ori33, mai33, men33, ori34, mai34, men34, ori35, mai35, men35, ori36, mai36, men36, ori37, mai37, men37, ori38, mai38, men38, ori39, mai39, men39;
  INV        o0000(.A(x3), .Y(ori_ori_n50_));
  NA2        o0001(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n51_));
  NA2        o0002(.A(x7), .B(x0), .Y(ori_ori_n52_));
  INV        o0003(.A(x1), .Y(ori_ori_n53_));
  NA2        o0004(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o0005(.A(x8), .Y(ori_ori_n55_));
  INV        o0006(.A(x4), .Y(ori_ori_n56_));
  INV        o0007(.A(x7), .Y(ori_ori_n57_));
  NA2        o0008(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0009(.A(x0), .Y(ori_ori_n59_));
  NA2        o0010(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NA4        o0011(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n55_), .D(x6), .Y(ori_ori_n61_));
  NA2        o0012(.A(ori_ori_n56_), .B(ori_ori_n59_), .Y(ori_ori_n62_));
  NO2        o0013(.A(ori_ori_n55_), .B(x6), .Y(ori_ori_n63_));
  NA2        o0014(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n64_));
  NA3        o0015(.A(ori_ori_n64_), .B(ori_ori_n63_), .C(ori_ori_n62_), .Y(ori_ori_n65_));
  AOI210     o0016(.A0(ori_ori_n65_), .A1(ori_ori_n61_), .B0(ori_ori_n54_), .Y(ori_ori_n66_));
  NO2        o0017(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n67_));
  NO2        o0018(.A(x7), .B(ori_ori_n59_), .Y(ori_ori_n68_));
  NO2        o0019(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  NAi21      o0020(.An(x5), .B(x1), .Y(ori_ori_n70_));
  INV        o0021(.A(x6), .Y(ori_ori_n71_));
  NA2        o0022(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NO3        o0023(.A(ori_ori_n72_), .B(ori_ori_n70_), .C(ori_ori_n69_), .Y(ori_ori_n73_));
  OAI210     o0024(.A0(ori_ori_n73_), .A1(ori_ori_n66_), .B0(ori_ori_n52_), .Y(ori_ori_n74_));
  NA2        o0025(.A(x7), .B(x4), .Y(ori_ori_n75_));
  NO2        o0026(.A(ori_ori_n75_), .B(x1), .Y(ori_ori_n76_));
  NO2        o0027(.A(ori_ori_n71_), .B(x5), .Y(ori_ori_n77_));
  NO2        o0028(.A(x8), .B(ori_ori_n59_), .Y(ori_ori_n78_));
  NA3        o0029(.A(ori_ori_n78_), .B(ori_ori_n77_), .C(ori_ori_n76_), .Y(ori_ori_n79_));
  AOI210     o0030(.A0(ori_ori_n79_), .A1(ori_ori_n74_), .B0(ori_ori_n51_), .Y(ori_ori_n80_));
  NA2        o0031(.A(x5), .B(x3), .Y(ori_ori_n81_));
  NO2        o0032(.A(x6), .B(x0), .Y(ori_ori_n82_));
  NO2        o0033(.A(ori_ori_n82_), .B(x4), .Y(ori_ori_n83_));
  NO2        o0034(.A(x4), .B(x2), .Y(ori_ori_n84_));
  NO2        o0035(.A(ori_ori_n71_), .B(ori_ori_n59_), .Y(ori_ori_n85_));
  NO2        o0036(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  NA2        o0037(.A(x8), .B(x1), .Y(ori_ori_n87_));
  NO2        o0038(.A(ori_ori_n87_), .B(x7), .Y(ori_ori_n88_));
  NO3        o0039(.A(x8), .B(ori_ori_n57_), .C(x6), .Y(ori_ori_n89_));
  NO2        o0040(.A(x1), .B(ori_ori_n59_), .Y(ori_ori_n90_));
  NO2        o0041(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n91_));
  XO2        o0042(.A(x7), .B(x1), .Y(ori_ori_n92_));
  INV        o0043(.A(ori_ori_n92_), .Y(ori_ori_n93_));
  NO2        o0044(.A(ori_ori_n93_), .B(x6), .Y(ori_ori_n94_));
  NO2        o0045(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n95_));
  NA2        o0046(.A(ori_ori_n95_), .B(ori_ori_n55_), .Y(ori_ori_n96_));
  NO2        o0047(.A(x6), .B(x5), .Y(ori_ori_n97_));
  NO2        o0048(.A(ori_ori_n57_), .B(x5), .Y(ori_ori_n98_));
  NO2        o0049(.A(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  NA2        o0050(.A(x6), .B(x1), .Y(ori_ori_n100_));
  NA2        o0051(.A(ori_ori_n100_), .B(ori_ori_n84_), .Y(ori_ori_n101_));
  NO4        o0052(.A(ori_ori_n101_), .B(ori_ori_n99_), .C(ori_ori_n96_), .D(ori_ori_n94_), .Y(ori_ori_n102_));
  NA2        o0053(.A(x3), .B(x0), .Y(ori_ori_n103_));
  INV        o0054(.A(x5), .Y(ori_ori_n104_));
  NA2        o0055(.A(ori_ori_n71_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  INV        o0056(.A(x2), .Y(ori_ori_n106_));
  NO2        o0057(.A(ori_ori_n56_), .B(ori_ori_n106_), .Y(ori_ori_n107_));
  NA2        o0058(.A(ori_ori_n57_), .B(ori_ori_n104_), .Y(ori_ori_n108_));
  NA3        o0059(.A(ori_ori_n108_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n109_));
  NO3        o0060(.A(ori_ori_n109_), .B(ori_ori_n103_), .C(ori_ori_n53_), .Y(ori_ori_n110_));
  NO3        o0061(.A(ori_ori_n110_), .B(ori_ori_n102_), .C(ori_ori_n80_), .Y(ori00));
  NO2        o0062(.A(x7), .B(x6), .Y(ori_ori_n112_));
  INV        o0063(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NO2        o0064(.A(ori_ori_n55_), .B(ori_ori_n53_), .Y(ori_ori_n114_));
  NA2        o0065(.A(ori_ori_n114_), .B(ori_ori_n56_), .Y(ori_ori_n115_));
  XN2        o0066(.A(x6), .B(x1), .Y(ori_ori_n116_));
  INV        o0067(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o0068(.A(x6), .B(x4), .Y(ori_ori_n118_));
  NA2        o0069(.A(x6), .B(x4), .Y(ori_ori_n119_));
  NAi21      o0070(.An(ori_ori_n118_), .B(ori_ori_n119_), .Y(ori_ori_n120_));
  XN2        o0071(.A(x7), .B(x6), .Y(ori_ori_n121_));
  NO2        o0072(.A(x3), .B(ori_ori_n106_), .Y(ori_ori_n122_));
  NA2        o0073(.A(ori_ori_n122_), .B(ori_ori_n104_), .Y(ori_ori_n123_));
  NA2        o0074(.A(x3), .B(ori_ori_n106_), .Y(ori_ori_n124_));
  NO2        o0075(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n125_));
  NA2        o0076(.A(ori_ori_n125_), .B(ori_ori_n56_), .Y(ori_ori_n126_));
  NA2        o0077(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n127_));
  NA2        o0078(.A(ori_ori_n127_), .B(x2), .Y(ori_ori_n128_));
  NA2        o0079(.A(x8), .B(x3), .Y(ori_ori_n129_));
  NA2        o0080(.A(ori_ori_n129_), .B(ori_ori_n75_), .Y(ori_ori_n130_));
  OAI220     o0081(.A0(ori_ori_n130_), .A1(ori_ori_n128_), .B0(ori_ori_n126_), .B1(ori_ori_n124_), .Y(ori_ori_n131_));
  NO2        o0082(.A(x5), .B(x0), .Y(ori_ori_n132_));
  NO2        o0083(.A(x6), .B(x1), .Y(ori_ori_n133_));
  NA3        o0084(.A(ori_ori_n133_), .B(ori_ori_n132_), .C(ori_ori_n131_), .Y(ori_ori_n134_));
  NA2        o0085(.A(x8), .B(ori_ori_n104_), .Y(ori_ori_n135_));
  NA2        o0086(.A(x4), .B(ori_ori_n50_), .Y(ori_ori_n136_));
  NO3        o0087(.A(ori_ori_n136_), .B(ori_ori_n135_), .C(ori_ori_n100_), .Y(ori_ori_n137_));
  NAi21      o0088(.An(x7), .B(x2), .Y(ori_ori_n138_));
  NO2        o0089(.A(ori_ori_n138_), .B(x0), .Y(ori_ori_n139_));
  XO2        o0090(.A(x8), .B(x7), .Y(ori_ori_n140_));
  NA2        o0091(.A(ori_ori_n140_), .B(ori_ori_n106_), .Y(ori_ori_n141_));
  NA2        o0092(.A(x6), .B(x5), .Y(ori_ori_n142_));
  NO2        o0093(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n143_));
  NO2        o0094(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n144_));
  NA2        o0095(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n145_));
  NO3        o0096(.A(ori_ori_n145_), .B(ori_ori_n142_), .C(ori_ori_n141_), .Y(ori_ori_n146_));
  AOI210     o0097(.A0(ori_ori_n139_), .A1(ori_ori_n137_), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NA2        o0098(.A(ori_ori_n147_), .B(ori_ori_n134_), .Y(ori01));
  NA2        o0099(.A(ori_ori_n57_), .B(ori_ori_n59_), .Y(ori_ori_n149_));
  NO2        o0100(.A(x2), .B(x1), .Y(ori_ori_n150_));
  NA2        o0101(.A(x2), .B(x1), .Y(ori_ori_n151_));
  NOi21      o0102(.An(ori_ori_n151_), .B(ori_ori_n150_), .Y(ori_ori_n152_));
  NA2        o0103(.A(ori_ori_n104_), .B(ori_ori_n53_), .Y(ori_ori_n153_));
  NO2        o0104(.A(ori_ori_n153_), .B(x8), .Y(ori_ori_n154_));
  NAi21      o0105(.An(x8), .B(x1), .Y(ori_ori_n155_));
  NO2        o0106(.A(ori_ori_n155_), .B(x3), .Y(ori_ori_n156_));
  OAI210     o0107(.A0(ori_ori_n156_), .A1(ori_ori_n154_), .B0(ori_ori_n152_), .Y(ori_ori_n157_));
  NO2        o0108(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n158_));
  NO2        o0109(.A(ori_ori_n106_), .B(x1), .Y(ori_ori_n159_));
  NA2        o0110(.A(ori_ori_n159_), .B(ori_ori_n158_), .Y(ori_ori_n160_));
  AOI210     o0111(.A0(ori_ori_n160_), .A1(ori_ori_n157_), .B0(ori_ori_n149_), .Y(ori_ori_n161_));
  NAi21      o0112(.An(x7), .B(x0), .Y(ori_ori_n162_));
  NO2        o0113(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n163_));
  NO2        o0114(.A(ori_ori_n81_), .B(x1), .Y(ori_ori_n164_));
  NA2        o0115(.A(ori_ori_n164_), .B(ori_ori_n163_), .Y(ori_ori_n165_));
  NA2        o0116(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n166_));
  NO2        o0117(.A(ori_ori_n166_), .B(ori_ori_n155_), .Y(ori_ori_n167_));
  NA2        o0118(.A(x8), .B(x5), .Y(ori_ori_n168_));
  NO3        o0119(.A(x3), .B(ori_ori_n106_), .C(ori_ori_n53_), .Y(ori_ori_n169_));
  NO2        o0120(.A(ori_ori_n169_), .B(ori_ori_n167_), .Y(ori_ori_n170_));
  AOI210     o0121(.A0(ori_ori_n170_), .A1(ori_ori_n165_), .B0(ori_ori_n162_), .Y(ori_ori_n171_));
  NO2        o0122(.A(ori_ori_n57_), .B(x3), .Y(ori_ori_n172_));
  NO2        o0123(.A(ori_ori_n55_), .B(x0), .Y(ori_ori_n173_));
  NA3        o0124(.A(ori_ori_n104_), .B(ori_ori_n106_), .C(x1), .Y(ori_ori_n174_));
  NO2        o0125(.A(ori_ori_n174_), .B(ori_ori_n173_), .Y(ori_ori_n175_));
  NO2        o0126(.A(ori_ori_n87_), .B(ori_ori_n50_), .Y(ori_ori_n176_));
  NA2        o0127(.A(ori_ori_n104_), .B(x0), .Y(ori_ori_n177_));
  NO2        o0128(.A(ori_ori_n177_), .B(x2), .Y(ori_ori_n178_));
  AOI220     o0129(.A0(ori_ori_n178_), .A1(ori_ori_n176_), .B0(ori_ori_n175_), .B1(ori_ori_n172_), .Y(ori_ori_n179_));
  NA2        o0130(.A(x7), .B(ori_ori_n106_), .Y(ori_ori_n180_));
  NA2        o0131(.A(ori_ori_n158_), .B(x8), .Y(ori_ori_n181_));
  NA4        o0132(.A(x5), .B(x3), .C(x1), .D(x0), .Y(ori_ori_n182_));
  AO210      o0133(.A0(ori_ori_n182_), .A1(ori_ori_n181_), .B0(ori_ori_n180_), .Y(ori_ori_n183_));
  NO2        o0134(.A(ori_ori_n151_), .B(ori_ori_n50_), .Y(ori_ori_n184_));
  NAi21      o0135(.An(x1), .B(x2), .Y(ori_ori_n185_));
  NO2        o0136(.A(ori_ori_n166_), .B(ori_ori_n185_), .Y(ori_ori_n186_));
  NA2        o0137(.A(x8), .B(x7), .Y(ori_ori_n187_));
  NO2        o0138(.A(ori_ori_n187_), .B(x0), .Y(ori_ori_n188_));
  OAI210     o0139(.A0(ori_ori_n186_), .A1(ori_ori_n184_), .B0(ori_ori_n188_), .Y(ori_ori_n189_));
  NA3        o0140(.A(ori_ori_n189_), .B(ori_ori_n183_), .C(ori_ori_n179_), .Y(ori_ori_n190_));
  NO3        o0141(.A(ori_ori_n190_), .B(ori_ori_n171_), .C(ori_ori_n161_), .Y(ori_ori_n191_));
  NA2        o0142(.A(x3), .B(x1), .Y(ori_ori_n192_));
  NA2        o0143(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n193_));
  NO2        o0144(.A(ori_ori_n193_), .B(ori_ori_n70_), .Y(ori_ori_n194_));
  OAI210     o0145(.A0(ori_ori_n194_), .A1(ori_ori_n186_), .B0(ori_ori_n67_), .Y(ori_ori_n195_));
  NA2        o0146(.A(ori_ori_n125_), .B(ori_ori_n106_), .Y(ori_ori_n196_));
  OAI210     o0147(.A0(ori_ori_n196_), .A1(ori_ori_n192_), .B0(ori_ori_n195_), .Y(ori_ori_n197_));
  XO2        o0148(.A(x5), .B(x3), .Y(ori_ori_n198_));
  NA2        o0149(.A(ori_ori_n198_), .B(x8), .Y(ori_ori_n199_));
  NA2        o0150(.A(x8), .B(ori_ori_n59_), .Y(ori_ori_n200_));
  NA2        o0151(.A(ori_ori_n200_), .B(ori_ori_n129_), .Y(ori_ori_n201_));
  NA2        o0152(.A(x7), .B(ori_ori_n71_), .Y(ori_ori_n202_));
  NO2        o0153(.A(ori_ori_n185_), .B(ori_ori_n202_), .Y(ori_ori_n203_));
  OA210      o0154(.A0(ori_ori_n201_), .A1(ori_ori_n198_), .B0(ori_ori_n203_), .Y(ori_ori_n204_));
  AOI220     o0155(.A0(ori_ori_n204_), .A1(ori_ori_n199_), .B0(ori_ori_n197_), .B1(x0), .Y(ori_ori_n205_));
  OAI210     o0156(.A0(ori_ori_n191_), .A1(ori_ori_n71_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  NO2        o0157(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n207_));
  NA4        o0158(.A(ori_ori_n55_), .B(x5), .C(x3), .D(x2), .Y(ori_ori_n208_));
  NA2        o0159(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n209_));
  NA2        o0160(.A(ori_ori_n209_), .B(x2), .Y(ori_ori_n210_));
  NA2        o0161(.A(ori_ori_n55_), .B(x3), .Y(ori_ori_n211_));
  NA4        o0162(.A(ori_ori_n211_), .B(ori_ori_n210_), .C(ori_ori_n198_), .D(ori_ori_n82_), .Y(ori_ori_n212_));
  AOI210     o0163(.A0(ori_ori_n212_), .A1(ori_ori_n208_), .B0(ori_ori_n53_), .Y(ori_ori_n213_));
  NO2        o0164(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n214_));
  NA2        o0165(.A(x5), .B(x1), .Y(ori_ori_n215_));
  NO2        o0166(.A(ori_ori_n215_), .B(x6), .Y(ori_ori_n216_));
  NO2        o0167(.A(x3), .B(x1), .Y(ori_ori_n217_));
  AOI210     o0168(.A0(ori_ori_n217_), .A1(ori_ori_n77_), .B0(ori_ori_n216_), .Y(ori_ori_n218_));
  NO2        o0169(.A(ori_ori_n81_), .B(ori_ori_n55_), .Y(ori_ori_n219_));
  NO2        o0170(.A(ori_ori_n100_), .B(ori_ori_n50_), .Y(ori_ori_n220_));
  NO2        o0171(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n221_));
  OAI210     o0172(.A0(ori_ori_n218_), .A1(x8), .B0(ori_ori_n221_), .Y(ori_ori_n222_));
  NO2        o0173(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n223_));
  NA2        o0174(.A(ori_ori_n223_), .B(ori_ori_n71_), .Y(ori_ori_n224_));
  NAi21      o0175(.An(x2), .B(x5), .Y(ori_ori_n225_));
  NA2        o0176(.A(x8), .B(x6), .Y(ori_ori_n226_));
  OAI210     o0177(.A0(ori_ori_n226_), .A1(ori_ori_n225_), .B0(ori_ori_n224_), .Y(ori_ori_n227_));
  NA2        o0178(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n228_));
  NO2        o0179(.A(ori_ori_n228_), .B(ori_ori_n59_), .Y(ori_ori_n229_));
  AO220      o0180(.A0(ori_ori_n229_), .A1(ori_ori_n227_), .B0(ori_ori_n222_), .B1(ori_ori_n214_), .Y(ori_ori_n230_));
  OAI210     o0181(.A0(ori_ori_n230_), .A1(ori_ori_n213_), .B0(ori_ori_n207_), .Y(ori_ori_n231_));
  NA2        o0182(.A(ori_ori_n71_), .B(ori_ori_n56_), .Y(ori_ori_n232_));
  NO2        o0183(.A(ori_ori_n232_), .B(x7), .Y(ori_ori_n233_));
  NO2        o0184(.A(ori_ori_n104_), .B(ori_ori_n53_), .Y(ori_ori_n234_));
  NA2        o0185(.A(ori_ori_n234_), .B(ori_ori_n106_), .Y(ori_ori_n235_));
  AOI210     o0186(.A0(ori_ori_n235_), .A1(ori_ori_n160_), .B0(ori_ori_n59_), .Y(ori_ori_n236_));
  NA2        o0187(.A(x3), .B(ori_ori_n59_), .Y(ori_ori_n237_));
  NO2        o0188(.A(ori_ori_n174_), .B(ori_ori_n237_), .Y(ori_ori_n238_));
  OA210      o0189(.A0(ori_ori_n238_), .A1(ori_ori_n236_), .B0(x8), .Y(ori_ori_n239_));
  NO2        o0190(.A(x1), .B(x0), .Y(ori_ori_n240_));
  NA2        o0191(.A(ori_ori_n240_), .B(ori_ori_n106_), .Y(ori_ori_n241_));
  NA2        o0192(.A(ori_ori_n104_), .B(ori_ori_n50_), .Y(ori_ori_n242_));
  XN2        o0193(.A(x3), .B(x2), .Y(ori_ori_n243_));
  NA2        o0194(.A(ori_ori_n243_), .B(ori_ori_n152_), .Y(ori_ori_n244_));
  NO2        o0195(.A(ori_ori_n104_), .B(x0), .Y(ori_ori_n245_));
  NA2        o0196(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n246_));
  NA2        o0197(.A(ori_ori_n246_), .B(ori_ori_n245_), .Y(ori_ori_n247_));
  OAI220     o0198(.A0(ori_ori_n247_), .A1(ori_ori_n244_), .B0(ori_ori_n242_), .B1(ori_ori_n241_), .Y(ori_ori_n248_));
  OAI210     o0199(.A0(ori_ori_n248_), .A1(ori_ori_n239_), .B0(ori_ori_n233_), .Y(ori_ori_n249_));
  NO2        o0200(.A(x7), .B(x1), .Y(ori_ori_n250_));
  NOi21      o0201(.An(x8), .B(x3), .Y(ori_ori_n251_));
  NA2        o0202(.A(ori_ori_n251_), .B(ori_ori_n59_), .Y(ori_ori_n252_));
  NA2        o0203(.A(x5), .B(x0), .Y(ori_ori_n253_));
  NAi21      o0204(.An(ori_ori_n132_), .B(ori_ori_n253_), .Y(ori_ori_n254_));
  NA2        o0205(.A(ori_ori_n71_), .B(ori_ori_n50_), .Y(ori_ori_n255_));
  OAI210     o0206(.A0(ori_ori_n255_), .A1(ori_ori_n254_), .B0(ori_ori_n252_), .Y(ori_ori_n256_));
  NA3        o0207(.A(ori_ori_n256_), .B(ori_ori_n135_), .C(ori_ori_n250_), .Y(ori_ori_n257_));
  NA2        o0208(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n258_));
  NO2        o0209(.A(ori_ori_n258_), .B(x5), .Y(ori_ori_n259_));
  NO2        o0210(.A(ori_ori_n144_), .B(ori_ori_n71_), .Y(ori_ori_n260_));
  NA2        o0211(.A(x1), .B(x0), .Y(ori_ori_n261_));
  NA2        o0212(.A(ori_ori_n50_), .B(ori_ori_n59_), .Y(ori_ori_n262_));
  NA4        o0213(.A(ori_ori_n262_), .B(ori_ori_n261_), .C(ori_ori_n260_), .D(ori_ori_n259_), .Y(ori_ori_n263_));
  NA3        o0214(.A(ori_ori_n263_), .B(ori_ori_n257_), .C(ori_ori_n182_), .Y(ori_ori_n264_));
  NO2        o0215(.A(ori_ori_n104_), .B(x3), .Y(ori_ori_n265_));
  NO2        o0216(.A(ori_ori_n106_), .B(x0), .Y(ori_ori_n266_));
  NA2        o0217(.A(ori_ori_n266_), .B(ori_ori_n265_), .Y(ori_ori_n267_));
  NO2        o0218(.A(ori_ori_n55_), .B(x7), .Y(ori_ori_n268_));
  NA2        o0219(.A(ori_ori_n268_), .B(ori_ori_n133_), .Y(ori_ori_n269_));
  NO3        o0220(.A(x8), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n270_));
  NAi21      o0221(.An(x8), .B(x0), .Y(ori_ori_n271_));
  NAi21      o0222(.An(x1), .B(x3), .Y(ori_ori_n272_));
  NO2        o0223(.A(ori_ori_n272_), .B(ori_ori_n271_), .Y(ori_ori_n273_));
  NO2        o0224(.A(x2), .B(ori_ori_n53_), .Y(ori_ori_n274_));
  AOI210     o0225(.A0(ori_ori_n274_), .A1(ori_ori_n270_), .B0(ori_ori_n273_), .Y(ori_ori_n275_));
  NOi21      o0226(.An(x5), .B(x6), .Y(ori_ori_n276_));
  NO2        o0227(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n277_));
  NA2        o0228(.A(ori_ori_n277_), .B(ori_ori_n276_), .Y(ori_ori_n278_));
  OAI220     o0229(.A0(ori_ori_n278_), .A1(ori_ori_n275_), .B0(ori_ori_n269_), .B1(ori_ori_n267_), .Y(ori_ori_n279_));
  AOI210     o0230(.A0(ori_ori_n264_), .A1(ori_ori_n107_), .B0(ori_ori_n279_), .Y(ori_ori_n280_));
  NA3        o0231(.A(ori_ori_n280_), .B(ori_ori_n249_), .C(ori_ori_n231_), .Y(ori_ori_n281_));
  AOI210     o0232(.A0(ori_ori_n206_), .A1(ori_ori_n56_), .B0(ori_ori_n281_), .Y(ori02));
  NO2        o0233(.A(x8), .B(ori_ori_n104_), .Y(ori_ori_n283_));
  XN2        o0234(.A(x7), .B(x3), .Y(ori_ori_n284_));
  INV        o0235(.A(ori_ori_n284_), .Y(ori_ori_n285_));
  NO2        o0236(.A(x2), .B(x0), .Y(ori_ori_n286_));
  NA2        o0237(.A(ori_ori_n286_), .B(ori_ori_n71_), .Y(ori_ori_n287_));
  NO2        o0238(.A(ori_ori_n57_), .B(x1), .Y(ori_ori_n288_));
  NO3        o0239(.A(ori_ori_n288_), .B(ori_ori_n287_), .C(ori_ori_n285_), .Y(ori_ori_n289_));
  NA2        o0240(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n290_));
  NO2        o0241(.A(ori_ori_n272_), .B(x6), .Y(ori_ori_n291_));
  XO2        o0242(.A(x7), .B(x0), .Y(ori_ori_n292_));
  NO2        o0243(.A(ori_ori_n292_), .B(ori_ori_n286_), .Y(ori_ori_n293_));
  NA2        o0244(.A(ori_ori_n293_), .B(ori_ori_n291_), .Y(ori_ori_n294_));
  AN2        o0245(.A(x7), .B(x2), .Y(ori_ori_n295_));
  NA2        o0246(.A(ori_ori_n295_), .B(ori_ori_n50_), .Y(ori_ori_n296_));
  OAI210     o0247(.A0(ori_ori_n296_), .A1(ori_ori_n290_), .B0(ori_ori_n294_), .Y(ori_ori_n297_));
  OAI210     o0248(.A0(ori_ori_n297_), .A1(ori_ori_n289_), .B0(ori_ori_n283_), .Y(ori_ori_n298_));
  NAi21      o0249(.An(x8), .B(x6), .Y(ori_ori_n299_));
  NO2        o0250(.A(ori_ori_n104_), .B(ori_ori_n59_), .Y(ori_ori_n300_));
  NA2        o0251(.A(x7), .B(x3), .Y(ori_ori_n301_));
  NO2        o0252(.A(ori_ori_n301_), .B(x2), .Y(ori_ori_n302_));
  NA2        o0253(.A(x2), .B(x0), .Y(ori_ori_n303_));
  NA2        o0254(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n304_));
  NA2        o0255(.A(ori_ori_n304_), .B(ori_ori_n303_), .Y(ori_ori_n305_));
  NAi21      o0256(.An(x7), .B(x1), .Y(ori_ori_n306_));
  NO2        o0257(.A(ori_ori_n306_), .B(x3), .Y(ori_ori_n307_));
  AOI220     o0258(.A0(ori_ori_n307_), .A1(ori_ori_n305_), .B0(ori_ori_n302_), .B1(ori_ori_n300_), .Y(ori_ori_n308_));
  NA2        o0259(.A(ori_ori_n274_), .B(ori_ori_n50_), .Y(ori_ori_n309_));
  NA3        o0260(.A(x7), .B(ori_ori_n104_), .C(x0), .Y(ori_ori_n310_));
  NA2        o0261(.A(ori_ori_n266_), .B(ori_ori_n53_), .Y(ori_ori_n311_));
  NA2        o0262(.A(ori_ori_n158_), .B(ori_ori_n57_), .Y(ori_ori_n312_));
  OA220      o0263(.A0(ori_ori_n312_), .A1(ori_ori_n311_), .B0(ori_ori_n310_), .B1(ori_ori_n309_), .Y(ori_ori_n313_));
  AOI210     o0264(.A0(ori_ori_n313_), .A1(ori_ori_n308_), .B0(ori_ori_n299_), .Y(ori_ori_n314_));
  INV        o0265(.A(ori_ori_n292_), .Y(ori_ori_n315_));
  NO2        o0266(.A(x7), .B(ori_ori_n71_), .Y(ori_ori_n316_));
  NA2        o0267(.A(ori_ori_n104_), .B(x3), .Y(ori_ori_n317_));
  NO2        o0268(.A(ori_ori_n317_), .B(ori_ori_n316_), .Y(ori_ori_n318_));
  NA2        o0269(.A(ori_ori_n318_), .B(ori_ori_n315_), .Y(ori_ori_n319_));
  NA2        o0270(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n320_));
  NO2        o0271(.A(ori_ori_n320_), .B(x7), .Y(ori_ori_n321_));
  NA2        o0272(.A(ori_ori_n321_), .B(ori_ori_n276_), .Y(ori_ori_n322_));
  NA2        o0273(.A(ori_ori_n163_), .B(x1), .Y(ori_ori_n323_));
  AOI210     o0274(.A0(ori_ori_n322_), .A1(ori_ori_n319_), .B0(ori_ori_n323_), .Y(ori_ori_n324_));
  NO2        o0275(.A(ori_ori_n57_), .B(ori_ori_n50_), .Y(ori_ori_n325_));
  NO2        o0276(.A(ori_ori_n55_), .B(ori_ori_n106_), .Y(ori_ori_n326_));
  NA3        o0277(.A(ori_ori_n326_), .B(ori_ori_n325_), .C(ori_ori_n59_), .Y(ori_ori_n327_));
  NO2        o0278(.A(ori_ori_n153_), .B(x6), .Y(ori_ori_n328_));
  NO2        o0279(.A(ori_ori_n100_), .B(ori_ori_n104_), .Y(ori_ori_n329_));
  NA2        o0280(.A(ori_ori_n57_), .B(ori_ori_n106_), .Y(ori_ori_n330_));
  NO2        o0281(.A(ori_ori_n330_), .B(ori_ori_n262_), .Y(ori_ori_n331_));
  OAI210     o0282(.A0(ori_ori_n329_), .A1(ori_ori_n328_), .B0(ori_ori_n331_), .Y(ori_ori_n332_));
  OAI210     o0283(.A0(ori_ori_n327_), .A1(ori_ori_n100_), .B0(ori_ori_n332_), .Y(ori_ori_n333_));
  NO3        o0284(.A(ori_ori_n333_), .B(ori_ori_n324_), .C(ori_ori_n314_), .Y(ori_ori_n334_));
  AOI210     o0285(.A0(ori_ori_n334_), .A1(ori_ori_n298_), .B0(x4), .Y(ori_ori_n335_));
  NA2        o0286(.A(x8), .B(ori_ori_n71_), .Y(ori_ori_n336_));
  NO2        o0287(.A(x3), .B(ori_ori_n59_), .Y(ori_ori_n337_));
  NA3        o0288(.A(ori_ori_n337_), .B(ori_ori_n104_), .C(ori_ori_n53_), .Y(ori_ori_n338_));
  NO2        o0289(.A(x3), .B(x0), .Y(ori_ori_n339_));
  NAi21      o0290(.An(ori_ori_n339_), .B(ori_ori_n103_), .Y(ori_ori_n340_));
  NA2        o0291(.A(x5), .B(x2), .Y(ori_ori_n341_));
  NO2        o0292(.A(ori_ori_n341_), .B(ori_ori_n217_), .Y(ori_ori_n342_));
  AOI210     o0293(.A0(ori_ori_n342_), .A1(ori_ori_n340_), .B0(ori_ori_n238_), .Y(ori_ori_n343_));
  AO210      o0294(.A0(ori_ori_n343_), .A1(ori_ori_n338_), .B0(ori_ori_n336_), .Y(ori_ori_n344_));
  NO2        o0295(.A(ori_ori_n106_), .B(ori_ori_n53_), .Y(ori_ori_n345_));
  NA2        o0296(.A(ori_ori_n345_), .B(x3), .Y(ori_ori_n346_));
  NO2        o0297(.A(ori_ori_n55_), .B(x1), .Y(ori_ori_n347_));
  NA2        o0298(.A(ori_ori_n347_), .B(ori_ori_n106_), .Y(ori_ori_n348_));
  OAI210     o0299(.A0(ori_ori_n348_), .A1(ori_ori_n166_), .B0(ori_ori_n346_), .Y(ori_ori_n349_));
  NAi32      o0300(.An(x3), .Bn(x0), .C(x2), .Y(ori_ori_n350_));
  NO2        o0301(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n351_));
  NAi21      o0302(.An(x6), .B(x5), .Y(ori_ori_n352_));
  NO2        o0303(.A(x2), .B(ori_ori_n59_), .Y(ori_ori_n353_));
  NO4        o0304(.A(ori_ori_n353_), .B(ori_ori_n352_), .C(ori_ori_n155_), .D(ori_ori_n351_), .Y(ori_ori_n354_));
  AOI220     o0305(.A0(ori_ori_n354_), .A1(ori_ori_n350_), .B0(ori_ori_n349_), .B1(ori_ori_n85_), .Y(ori_ori_n355_));
  AOI210     o0306(.A0(ori_ori_n355_), .A1(ori_ori_n344_), .B0(ori_ori_n75_), .Y(ori_ori_n356_));
  NA2        o0307(.A(ori_ori_n347_), .B(ori_ori_n56_), .Y(ori_ori_n357_));
  NO2        o0308(.A(ori_ori_n104_), .B(ori_ori_n50_), .Y(ori_ori_n358_));
  NO2        o0309(.A(ori_ori_n286_), .B(ori_ori_n214_), .Y(ori_ori_n359_));
  XO2        o0310(.A(x7), .B(x2), .Y(ori_ori_n360_));
  INV        o0311(.A(ori_ori_n360_), .Y(ori_ori_n361_));
  XO2        o0312(.A(x6), .B(x2), .Y(ori_ori_n362_));
  NA4        o0313(.A(ori_ori_n362_), .B(ori_ori_n361_), .C(ori_ori_n359_), .D(ori_ori_n358_), .Y(ori_ori_n363_));
  NAi21      o0314(.An(x0), .B(x6), .Y(ori_ori_n364_));
  AOI210     o0315(.A0(ori_ori_n364_), .A1(ori_ori_n138_), .B0(ori_ori_n266_), .Y(ori_ori_n365_));
  XN2        o0316(.A(x7), .B(x5), .Y(ori_ori_n366_));
  NA2        o0317(.A(ori_ori_n366_), .B(ori_ori_n71_), .Y(ori_ori_n367_));
  NA2        o0318(.A(x7), .B(x5), .Y(ori_ori_n368_));
  AOI210     o0319(.A0(ori_ori_n368_), .A1(x6), .B0(ori_ori_n350_), .Y(ori_ori_n369_));
  AOI220     o0320(.A0(ori_ori_n369_), .A1(ori_ori_n367_), .B0(ori_ori_n365_), .B1(ori_ori_n318_), .Y(ori_ori_n370_));
  AOI210     o0321(.A0(ori_ori_n370_), .A1(ori_ori_n363_), .B0(ori_ori_n357_), .Y(ori_ori_n371_));
  NO2        o0322(.A(x8), .B(x6), .Y(ori_ori_n372_));
  NAi21      o0323(.An(ori_ori_n372_), .B(ori_ori_n226_), .Y(ori_ori_n373_));
  AOI210     o0324(.A0(ori_ori_n373_), .A1(ori_ori_n90_), .B0(x3), .Y(ori_ori_n374_));
  NA2        o0325(.A(ori_ori_n104_), .B(x2), .Y(ori_ori_n375_));
  NO2        o0326(.A(ori_ori_n375_), .B(ori_ori_n64_), .Y(ori_ori_n376_));
  NA2        o0327(.A(x1), .B(ori_ori_n59_), .Y(ori_ori_n377_));
  NO2        o0328(.A(ori_ori_n377_), .B(ori_ori_n226_), .Y(ori_ori_n378_));
  OAI210     o0329(.A0(ori_ori_n378_), .A1(ori_ori_n50_), .B0(ori_ori_n376_), .Y(ori_ori_n379_));
  NA2        o0330(.A(x4), .B(x2), .Y(ori_ori_n380_));
  NO2        o0331(.A(ori_ori_n380_), .B(ori_ori_n104_), .Y(ori_ori_n381_));
  NAi21      o0332(.An(x1), .B(x6), .Y(ori_ori_n382_));
  NA2        o0333(.A(ori_ori_n339_), .B(ori_ori_n268_), .Y(ori_ori_n383_));
  OAI220     o0334(.A0(ori_ori_n383_), .A1(ori_ori_n382_), .B0(ori_ori_n103_), .B1(ori_ori_n53_), .Y(ori_ori_n384_));
  NA2        o0335(.A(x8), .B(x2), .Y(ori_ori_n385_));
  NO2        o0336(.A(ori_ori_n385_), .B(ori_ori_n50_), .Y(ori_ori_n386_));
  INV        o0337(.A(ori_ori_n216_), .Y(ori_ori_n387_));
  NO2        o0338(.A(ori_ori_n387_), .B(ori_ori_n52_), .Y(ori_ori_n388_));
  AOI220     o0339(.A0(ori_ori_n388_), .A1(ori_ori_n386_), .B0(ori_ori_n384_), .B1(ori_ori_n381_), .Y(ori_ori_n389_));
  OAI210     o0340(.A0(ori_ori_n379_), .A1(ori_ori_n374_), .B0(ori_ori_n389_), .Y(ori_ori_n390_));
  NO4        o0341(.A(ori_ori_n390_), .B(ori_ori_n371_), .C(ori_ori_n356_), .D(ori_ori_n335_), .Y(ori03));
  NAi21      o0342(.An(x2), .B(x0), .Y(ori_ori_n392_));
  NO3        o0343(.A(x8), .B(x6), .C(x4), .Y(ori_ori_n393_));
  INV        o0344(.A(ori_ori_n393_), .Y(ori_ori_n394_));
  NO2        o0345(.A(ori_ori_n394_), .B(ori_ori_n392_), .Y(ori_ori_n395_));
  NA2        o0346(.A(ori_ori_n107_), .B(ori_ori_n59_), .Y(ori_ori_n396_));
  NO2        o0347(.A(ori_ori_n396_), .B(ori_ori_n55_), .Y(ori_ori_n397_));
  OAI210     o0348(.A0(ori_ori_n397_), .A1(ori_ori_n395_), .B0(ori_ori_n158_), .Y(ori_ori_n398_));
  NA2        o0349(.A(x3), .B(x2), .Y(ori_ori_n399_));
  NO2        o0350(.A(ori_ori_n155_), .B(x0), .Y(ori_ori_n400_));
  NA2        o0351(.A(x8), .B(x0), .Y(ori_ori_n401_));
  NO2        o0352(.A(ori_ori_n401_), .B(x6), .Y(ori_ori_n402_));
  AOI210     o0353(.A0(ori_ori_n402_), .A1(x5), .B0(ori_ori_n400_), .Y(ori_ori_n403_));
  NO2        o0354(.A(ori_ori_n403_), .B(ori_ori_n399_), .Y(ori_ori_n404_));
  NO2        o0355(.A(x5), .B(ori_ori_n59_), .Y(ori_ori_n405_));
  NO2        o0356(.A(x3), .B(x2), .Y(ori_ori_n406_));
  NA2        o0357(.A(ori_ori_n406_), .B(ori_ori_n405_), .Y(ori_ori_n407_));
  NO2        o0358(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n408_));
  NA2        o0359(.A(ori_ori_n408_), .B(x5), .Y(ori_ori_n409_));
  AOI210     o0360(.A0(ori_ori_n409_), .A1(ori_ori_n407_), .B0(ori_ori_n299_), .Y(ori_ori_n410_));
  NA2        o0361(.A(ori_ori_n252_), .B(ori_ori_n168_), .Y(ori_ori_n411_));
  NO2        o0362(.A(ori_ori_n50_), .B(ori_ori_n59_), .Y(ori_ori_n412_));
  NO2        o0363(.A(ori_ori_n71_), .B(x0), .Y(ori_ori_n413_));
  NO4        o0364(.A(ori_ori_n413_), .B(ori_ori_n412_), .C(x2), .D(ori_ori_n53_), .Y(ori_ori_n414_));
  AO210      o0365(.A0(ori_ori_n414_), .A1(ori_ori_n411_), .B0(ori_ori_n410_), .Y(ori_ori_n415_));
  OAI210     o0366(.A0(ori_ori_n415_), .A1(ori_ori_n404_), .B0(x4), .Y(ori_ori_n416_));
  NO2        o0367(.A(x4), .B(ori_ori_n53_), .Y(ori_ori_n417_));
  NA2        o0368(.A(ori_ori_n417_), .B(ori_ori_n59_), .Y(ori_ori_n418_));
  NO3        o0369(.A(ori_ori_n418_), .B(ori_ori_n226_), .C(x5), .Y(ori_ori_n419_));
  NA2        o0370(.A(x7), .B(ori_ori_n104_), .Y(ori_ori_n420_));
  NO3        o0371(.A(x5), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n421_));
  INV        o0372(.A(ori_ori_n421_), .Y(ori_ori_n422_));
  NO2        o0373(.A(x6), .B(ori_ori_n56_), .Y(ori_ori_n423_));
  NO2        o0374(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n424_));
  NA2        o0375(.A(ori_ori_n424_), .B(ori_ori_n423_), .Y(ori_ori_n425_));
  OAI210     o0376(.A0(ori_ori_n425_), .A1(ori_ori_n422_), .B0(ori_ori_n420_), .Y(ori_ori_n426_));
  AOI210     o0377(.A0(ori_ori_n419_), .A1(x2), .B0(ori_ori_n426_), .Y(ori_ori_n427_));
  AOI220     o0378(.A0(ori_ori_n427_), .A1(ori_ori_n416_), .B0(ori_ori_n398_), .B1(x7), .Y(ori_ori_n428_));
  NA2        o0379(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n429_));
  NO2        o0380(.A(ori_ori_n251_), .B(ori_ori_n106_), .Y(ori_ori_n430_));
  NO2        o0381(.A(ori_ori_n55_), .B(ori_ori_n59_), .Y(ori_ori_n431_));
  NO3        o0382(.A(ori_ori_n431_), .B(ori_ori_n430_), .C(ori_ori_n142_), .Y(ori_ori_n432_));
  AOI210     o0383(.A0(ori_ori_n201_), .A1(ori_ori_n97_), .B0(ori_ori_n432_), .Y(ori_ori_n433_));
  NO2        o0384(.A(x5), .B(x2), .Y(ori_ori_n434_));
  NO2        o0385(.A(x8), .B(x3), .Y(ori_ori_n435_));
  NA2        o0386(.A(ori_ori_n435_), .B(ori_ori_n434_), .Y(ori_ori_n436_));
  NO2        o0387(.A(ori_ori_n436_), .B(x6), .Y(ori_ori_n437_));
  NA2        o0388(.A(ori_ori_n200_), .B(x2), .Y(ori_ori_n438_));
  NO3        o0389(.A(ori_ori_n435_), .B(ori_ori_n340_), .C(ori_ori_n352_), .Y(ori_ori_n439_));
  NA2        o0390(.A(ori_ori_n439_), .B(ori_ori_n438_), .Y(ori_ori_n440_));
  OAI210     o0391(.A0(ori_ori_n433_), .A1(ori_ori_n286_), .B0(ori_ori_n440_), .Y(ori_ori_n441_));
  NA2        o0392(.A(ori_ori_n441_), .B(x4), .Y(ori_ori_n442_));
  NA2        o0393(.A(ori_ori_n55_), .B(ori_ori_n59_), .Y(ori_ori_n443_));
  NO2        o0394(.A(ori_ori_n443_), .B(x5), .Y(ori_ori_n444_));
  NAi21      o0395(.An(x4), .B(x6), .Y(ori_ori_n445_));
  NO2        o0396(.A(ori_ori_n445_), .B(ori_ori_n51_), .Y(ori_ori_n446_));
  NO2        o0397(.A(ori_ori_n55_), .B(ori_ori_n71_), .Y(ori_ori_n447_));
  NO2        o0398(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n448_));
  NO2        o0399(.A(ori_ori_n226_), .B(x0), .Y(ori_ori_n449_));
  NO2        o0400(.A(ori_ori_n352_), .B(x8), .Y(ori_ori_n450_));
  OAI210     o0401(.A0(ori_ori_n450_), .A1(ori_ori_n449_), .B0(ori_ori_n448_), .Y(ori_ori_n451_));
  OAI210     o0402(.A0(ori_ori_n407_), .A1(ori_ori_n447_), .B0(ori_ori_n451_), .Y(ori_ori_n452_));
  AOI220     o0403(.A0(ori_ori_n452_), .A1(ori_ori_n56_), .B0(ori_ori_n446_), .B1(ori_ori_n444_), .Y(ori_ori_n453_));
  AOI210     o0404(.A0(ori_ori_n453_), .A1(ori_ori_n442_), .B0(ori_ori_n429_), .Y(ori_ori_n454_));
  NA2        o0405(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n455_));
  NO2        o0406(.A(ori_ori_n71_), .B(ori_ori_n56_), .Y(ori_ori_n456_));
  NA2        o0407(.A(ori_ori_n351_), .B(ori_ori_n59_), .Y(ori_ori_n457_));
  OAI220     o0408(.A0(ori_ori_n457_), .A1(ori_ori_n55_), .B0(ori_ori_n193_), .B1(ori_ori_n271_), .Y(ori_ori_n458_));
  NA2        o0409(.A(ori_ori_n458_), .B(ori_ori_n456_), .Y(ori_ori_n459_));
  NO3        o0410(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n460_));
  NA2        o0411(.A(ori_ori_n431_), .B(x5), .Y(ori_ori_n461_));
  NO2        o0412(.A(x8), .B(x5), .Y(ori_ori_n462_));
  NAi21      o0413(.An(ori_ori_n462_), .B(ori_ori_n168_), .Y(ori_ori_n463_));
  OAI210     o0414(.A0(ori_ori_n463_), .A1(ori_ori_n304_), .B0(ori_ori_n461_), .Y(ori_ori_n464_));
  NA2        o0415(.A(ori_ori_n359_), .B(ori_ori_n77_), .Y(ori_ori_n465_));
  NOi21      o0416(.An(x3), .B(x4), .Y(ori_ori_n466_));
  NA2        o0417(.A(ori_ori_n55_), .B(ori_ori_n106_), .Y(ori_ori_n467_));
  NA2        o0418(.A(ori_ori_n467_), .B(ori_ori_n466_), .Y(ori_ori_n468_));
  NO2        o0419(.A(ori_ori_n51_), .B(x6), .Y(ori_ori_n469_));
  NO2        o0420(.A(ori_ori_n142_), .B(ori_ori_n55_), .Y(ori_ori_n470_));
  NO3        o0421(.A(ori_ori_n56_), .B(x2), .C(x0), .Y(ori_ori_n471_));
  AOI220     o0422(.A0(ori_ori_n471_), .A1(ori_ori_n470_), .B0(ori_ori_n469_), .B1(ori_ori_n444_), .Y(ori_ori_n472_));
  OAI210     o0423(.A0(ori_ori_n468_), .A1(ori_ori_n465_), .B0(ori_ori_n472_), .Y(ori_ori_n473_));
  AOI210     o0424(.A0(ori_ori_n464_), .A1(ori_ori_n460_), .B0(ori_ori_n473_), .Y(ori_ori_n474_));
  AOI210     o0425(.A0(ori_ori_n474_), .A1(ori_ori_n459_), .B0(ori_ori_n455_), .Y(ori_ori_n475_));
  NA2        o0426(.A(x7), .B(x1), .Y(ori_ori_n476_));
  NO3        o0427(.A(x5), .B(x4), .C(x2), .Y(ori_ori_n477_));
  AN2        o0428(.A(ori_ori_n477_), .B(ori_ori_n372_), .Y(ori_ori_n478_));
  NO3        o0429(.A(ori_ori_n478_), .B(ori_ori_n470_), .C(ori_ori_n381_), .Y(ori_ori_n479_));
  OAI210     o0430(.A0(ori_ori_n372_), .A1(ori_ori_n84_), .B0(ori_ori_n339_), .Y(ori_ori_n480_));
  NO2        o0431(.A(ori_ori_n480_), .B(ori_ori_n479_), .Y(ori_ori_n481_));
  NO2        o0432(.A(x4), .B(ori_ori_n106_), .Y(ori_ori_n482_));
  NA2        o0433(.A(ori_ori_n482_), .B(x6), .Y(ori_ori_n483_));
  NA3        o0434(.A(ori_ori_n104_), .B(x4), .C(ori_ori_n106_), .Y(ori_ori_n484_));
  AOI210     o0435(.A0(ori_ori_n484_), .A1(ori_ori_n483_), .B0(ori_ori_n96_), .Y(ori_ori_n485_));
  NA2        o0436(.A(ori_ori_n466_), .B(ori_ori_n71_), .Y(ori_ori_n486_));
  NA2        o0437(.A(ori_ori_n163_), .B(ori_ori_n59_), .Y(ori_ori_n487_));
  NO2        o0438(.A(ori_ori_n487_), .B(ori_ori_n486_), .Y(ori_ori_n488_));
  NA2        o0439(.A(ori_ori_n448_), .B(x4), .Y(ori_ori_n489_));
  NO3        o0440(.A(ori_ori_n489_), .B(ori_ori_n372_), .C(ori_ori_n413_), .Y(ori_ori_n490_));
  NO4        o0441(.A(ori_ori_n490_), .B(ori_ori_n488_), .C(ori_ori_n485_), .D(ori_ori_n481_), .Y(ori_ori_n491_));
  NA2        o0442(.A(x5), .B(x4), .Y(ori_ori_n492_));
  NO2        o0443(.A(ori_ori_n71_), .B(ori_ori_n53_), .Y(ori_ori_n493_));
  NO3        o0444(.A(x8), .B(x3), .C(x2), .Y(ori_ori_n494_));
  NA3        o0445(.A(ori_ori_n494_), .B(ori_ori_n493_), .C(ori_ori_n59_), .Y(ori_ori_n495_));
  NO3        o0446(.A(x6), .B(x5), .C(x2), .Y(ori_ori_n496_));
  NA3        o0447(.A(ori_ori_n496_), .B(ori_ori_n288_), .C(ori_ori_n78_), .Y(ori_ori_n497_));
  OAI210     o0448(.A0(ori_ori_n495_), .A1(ori_ori_n492_), .B0(ori_ori_n497_), .Y(ori_ori_n498_));
  NA2        o0449(.A(ori_ori_n71_), .B(x2), .Y(ori_ori_n499_));
  NO3        o0450(.A(x4), .B(x3), .C(ori_ori_n59_), .Y(ori_ori_n500_));
  NA2        o0451(.A(ori_ori_n500_), .B(ori_ori_n223_), .Y(ori_ori_n501_));
  NO3        o0452(.A(ori_ori_n501_), .B(ori_ori_n499_), .C(ori_ori_n92_), .Y(ori_ori_n502_));
  XO2        o0453(.A(x4), .B(x0), .Y(ori_ori_n503_));
  NA2        o0454(.A(ori_ori_n262_), .B(x5), .Y(ori_ori_n504_));
  NO2        o0455(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n505_));
  NO2        o0456(.A(ori_ori_n505_), .B(ori_ori_n63_), .Y(ori_ori_n506_));
  NO4        o0457(.A(ori_ori_n506_), .B(ori_ori_n504_), .C(ori_ori_n503_), .D(ori_ori_n151_), .Y(ori_ori_n507_));
  NO3        o0458(.A(ori_ori_n507_), .B(ori_ori_n502_), .C(ori_ori_n498_), .Y(ori_ori_n508_));
  OAI210     o0459(.A0(ori_ori_n491_), .A1(ori_ori_n476_), .B0(ori_ori_n508_), .Y(ori_ori_n509_));
  NO4        o0460(.A(ori_ori_n509_), .B(ori_ori_n475_), .C(ori_ori_n454_), .D(ori_ori_n428_), .Y(ori04));
  NO2        o0461(.A(x7), .B(x2), .Y(ori_ori_n511_));
  NO2        o0462(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n512_));
  NO2        o0463(.A(ori_ori_n512_), .B(ori_ori_n144_), .Y(ori_ori_n513_));
  XN2        o0464(.A(x8), .B(x1), .Y(ori_ori_n514_));
  NO2        o0465(.A(ori_ori_n514_), .B(ori_ori_n142_), .Y(ori_ori_n515_));
  NA2        o0466(.A(ori_ori_n515_), .B(ori_ori_n513_), .Y(ori_ori_n516_));
  NA2        o0467(.A(x6), .B(x3), .Y(ori_ori_n517_));
  NO2        o0468(.A(ori_ori_n517_), .B(x5), .Y(ori_ori_n518_));
  NA2        o0469(.A(ori_ori_n71_), .B(x1), .Y(ori_ori_n519_));
  NO2        o0470(.A(ori_ori_n462_), .B(ori_ori_n251_), .Y(ori_ori_n520_));
  NO3        o0471(.A(ori_ori_n520_), .B(ori_ori_n435_), .C(ori_ori_n519_), .Y(ori_ori_n521_));
  AOI210     o0472(.A0(ori_ori_n518_), .A1(ori_ori_n347_), .B0(ori_ori_n521_), .Y(ori_ori_n522_));
  AOI210     o0473(.A0(ori_ori_n522_), .A1(ori_ori_n516_), .B0(x0), .Y(ori_ori_n523_));
  NOi21      o0474(.An(ori_ori_n168_), .B(ori_ori_n462_), .Y(ori_ori_n524_));
  NA2        o0475(.A(ori_ori_n105_), .B(x1), .Y(ori_ori_n525_));
  NO3        o0476(.A(ori_ori_n525_), .B(ori_ori_n524_), .C(ori_ori_n320_), .Y(ori_ori_n526_));
  OAI210     o0477(.A0(ori_ori_n526_), .A1(ori_ori_n523_), .B0(ori_ori_n511_), .Y(ori_ori_n527_));
  NA2        o0478(.A(ori_ori_n129_), .B(ori_ori_n237_), .Y(ori_ori_n528_));
  OR4        o0479(.A(ori_ori_n528_), .B(ori_ori_n373_), .C(ori_ori_n82_), .D(ori_ori_n54_), .Y(ori_ori_n529_));
  OR2        o0480(.A(x6), .B(x0), .Y(ori_ori_n530_));
  NO3        o0481(.A(ori_ori_n530_), .B(x3), .C(x1), .Y(ori_ori_n531_));
  AOI220     o0482(.A0(ori_ori_n531_), .A1(ori_ori_n104_), .B0(ori_ori_n276_), .B1(ori_ori_n270_), .Y(ori_ori_n532_));
  AOI210     o0483(.A0(ori_ori_n532_), .A1(ori_ori_n529_), .B0(ori_ori_n180_), .Y(ori_ori_n533_));
  NA2        o0484(.A(x7), .B(x2), .Y(ori_ori_n534_));
  INV        o0485(.A(ori_ori_n129_), .Y(ori_ori_n535_));
  OAI210     o0486(.A0(ori_ori_n167_), .A1(ori_ori_n535_), .B0(ori_ori_n82_), .Y(ori_ori_n536_));
  NO2        o0487(.A(ori_ori_n317_), .B(ori_ori_n55_), .Y(ori_ori_n537_));
  NO3        o0488(.A(x3), .B(x1), .C(x0), .Y(ori_ori_n538_));
  OR2        o0489(.A(x6), .B(x1), .Y(ori_ori_n539_));
  NA2        o0490(.A(ori_ori_n539_), .B(x0), .Y(ori_ori_n540_));
  AOI220     o0491(.A0(ori_ori_n540_), .A1(ori_ori_n537_), .B0(ori_ori_n538_), .B1(ori_ori_n470_), .Y(ori_ori_n541_));
  AOI210     o0492(.A0(ori_ori_n541_), .A1(ori_ori_n536_), .B0(ori_ori_n534_), .Y(ori_ori_n542_));
  NA2        o0493(.A(ori_ori_n71_), .B(x0), .Y(ori_ori_n543_));
  NOi31      o0494(.An(ori_ori_n342_), .B(ori_ori_n543_), .C(ori_ori_n258_), .Y(ori_ori_n544_));
  NO4        o0495(.A(ori_ori_n544_), .B(ori_ori_n542_), .C(ori_ori_n533_), .D(ori_ori_n56_), .Y(ori_ori_n545_));
  NA2        o0496(.A(ori_ori_n545_), .B(ori_ori_n527_), .Y(ori_ori_n546_));
  NA3        o0497(.A(x8), .B(x7), .C(x0), .Y(ori_ori_n547_));
  INV        o0498(.A(ori_ori_n547_), .Y(ori_ori_n548_));
  AOI210     o0499(.A0(ori_ori_n268_), .A1(ori_ori_n95_), .B0(ori_ori_n548_), .Y(ori_ori_n549_));
  NO2        o0500(.A(ori_ori_n549_), .B(ori_ori_n151_), .Y(ori_ori_n550_));
  NA2        o0501(.A(ori_ori_n431_), .B(ori_ori_n57_), .Y(ori_ori_n551_));
  NO2        o0502(.A(x8), .B(x0), .Y(ori_ori_n552_));
  NA2        o0503(.A(ori_ori_n552_), .B(ori_ori_n361_), .Y(ori_ori_n553_));
  AOI210     o0504(.A0(ori_ori_n553_), .A1(ori_ori_n551_), .B0(ori_ori_n272_), .Y(ori_ori_n554_));
  OAI210     o0505(.A0(ori_ori_n554_), .A1(ori_ori_n550_), .B0(ori_ori_n276_), .Y(ori_ori_n555_));
  NO2        o0506(.A(ori_ori_n71_), .B(ori_ori_n106_), .Y(ori_ori_n556_));
  NO2        o0507(.A(ori_ori_n368_), .B(x8), .Y(ori_ori_n557_));
  NO2        o0508(.A(ori_ori_n557_), .B(ori_ori_n259_), .Y(ori_ori_n558_));
  NO3        o0509(.A(ori_ori_n558_), .B(ori_ori_n377_), .C(ori_ori_n265_), .Y(ori_ori_n559_));
  NO2        o0510(.A(ori_ori_n285_), .B(x8), .Y(ori_ori_n560_));
  OAI210     o0511(.A0(ori_ori_n462_), .A1(ori_ori_n325_), .B0(ori_ori_n240_), .Y(ori_ori_n561_));
  NA2        o0512(.A(ori_ori_n347_), .B(ori_ori_n172_), .Y(ori_ori_n562_));
  OAI220     o0513(.A0(ori_ori_n562_), .A1(ori_ori_n59_), .B0(ori_ori_n561_), .B1(ori_ori_n560_), .Y(ori_ori_n563_));
  OAI210     o0514(.A0(ori_ori_n563_), .A1(ori_ori_n559_), .B0(ori_ori_n556_), .Y(ori_ori_n564_));
  NO2        o0515(.A(x8), .B(x2), .Y(ori_ori_n565_));
  NO2        o0516(.A(ori_ori_n217_), .B(ori_ori_n57_), .Y(ori_ori_n566_));
  NA3        o0517(.A(ori_ori_n566_), .B(ori_ori_n565_), .C(ori_ori_n340_), .Y(ori_ori_n567_));
  NO2        o0518(.A(ori_ori_n241_), .B(ori_ori_n129_), .Y(ori_ori_n568_));
  AOI210     o0519(.A0(ori_ori_n321_), .A1(ori_ori_n159_), .B0(ori_ori_n568_), .Y(ori_ori_n569_));
  AOI210     o0520(.A0(ori_ori_n569_), .A1(ori_ori_n567_), .B0(ori_ori_n105_), .Y(ori_ori_n570_));
  NA2        o0521(.A(ori_ori_n337_), .B(x2), .Y(ori_ori_n571_));
  NO2        o0522(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n572_));
  NA2        o0523(.A(ori_ori_n572_), .B(ori_ori_n63_), .Y(ori_ori_n573_));
  AOI210     o0524(.A0(ori_ori_n571_), .A1(ori_ori_n457_), .B0(ori_ori_n573_), .Y(ori_ori_n574_));
  NA2        o0525(.A(ori_ori_n106_), .B(ori_ori_n53_), .Y(ori_ori_n575_));
  NO2        o0526(.A(ori_ori_n575_), .B(x8), .Y(ori_ori_n576_));
  NA2        o0527(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n577_));
  NO2        o0528(.A(ori_ori_n177_), .B(ori_ori_n577_), .Y(ori_ori_n578_));
  AN2        o0529(.A(ori_ori_n578_), .B(ori_ori_n576_), .Y(ori_ori_n579_));
  NA2        o0530(.A(ori_ori_n405_), .B(ori_ori_n144_), .Y(ori_ori_n580_));
  NO2        o0531(.A(ori_ori_n71_), .B(x2), .Y(ori_ori_n581_));
  NA2        o0532(.A(ori_ori_n581_), .B(ori_ori_n268_), .Y(ori_ori_n582_));
  OAI210     o0533(.A0(ori_ori_n582_), .A1(ori_ori_n580_), .B0(ori_ori_n56_), .Y(ori_ori_n583_));
  NO4        o0534(.A(ori_ori_n583_), .B(ori_ori_n579_), .C(ori_ori_n574_), .D(ori_ori_n570_), .Y(ori_ori_n584_));
  NA3        o0535(.A(ori_ori_n584_), .B(ori_ori_n564_), .C(ori_ori_n555_), .Y(ori_ori_n585_));
  NA2        o0536(.A(ori_ori_n53_), .B(ori_ori_n59_), .Y(ori_ori_n586_));
  NOi21      o0537(.An(x2), .B(x7), .Y(ori_ori_n587_));
  NO2        o0538(.A(x6), .B(x3), .Y(ori_ori_n588_));
  NA2        o0539(.A(ori_ori_n588_), .B(ori_ori_n587_), .Y(ori_ori_n589_));
  NO2        o0540(.A(x6), .B(ori_ori_n59_), .Y(ori_ori_n590_));
  NO3        o0541(.A(ori_ori_n57_), .B(x2), .C(x1), .Y(ori_ori_n591_));
  NO3        o0542(.A(ori_ori_n57_), .B(x2), .C(x0), .Y(ori_ori_n592_));
  AOI220     o0543(.A0(ori_ori_n592_), .A1(ori_ori_n220_), .B0(ori_ori_n591_), .B1(ori_ori_n590_), .Y(ori_ori_n593_));
  OAI210     o0544(.A0(ori_ori_n589_), .A1(ori_ori_n586_), .B0(ori_ori_n593_), .Y(ori_ori_n594_));
  NO2        o0545(.A(ori_ori_n97_), .B(ori_ori_n53_), .Y(ori_ori_n595_));
  NA2        o0546(.A(ori_ori_n215_), .B(ori_ori_n57_), .Y(ori_ori_n596_));
  OAI210     o0547(.A0(ori_ori_n595_), .A1(ori_ori_n450_), .B0(ori_ori_n596_), .Y(ori_ori_n597_));
  NO3        o0548(.A(ori_ori_n597_), .B(ori_ori_n489_), .C(ori_ori_n59_), .Y(ori_ori_n598_));
  AO210      o0549(.A0(ori_ori_n594_), .A1(ori_ori_n462_), .B0(ori_ori_n598_), .Y(ori_ori_n599_));
  AOI210     o0550(.A0(ori_ori_n585_), .A1(ori_ori_n546_), .B0(ori_ori_n599_), .Y(ori05));
  AOI210     o0551(.A0(ori_ori_n158_), .A1(ori_ori_n55_), .B0(ori_ori_n505_), .Y(ori_ori_n601_));
  OR2        o0552(.A(ori_ori_n601_), .B(ori_ori_n57_), .Y(ori_ori_n602_));
  NO2        o0553(.A(x7), .B(ori_ori_n104_), .Y(ori_ori_n603_));
  NO2        o0554(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n604_));
  NA2        o0555(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n605_));
  NO2        o0556(.A(ori_ori_n605_), .B(ori_ori_n577_), .Y(ori_ori_n606_));
  AOI210     o0557(.A0(ori_ori_n604_), .A1(ori_ori_n603_), .B0(ori_ori_n606_), .Y(ori_ori_n607_));
  AOI210     o0558(.A0(ori_ori_n607_), .A1(ori_ori_n602_), .B0(ori_ori_n106_), .Y(ori_ori_n608_));
  NO2        o0559(.A(x7), .B(x4), .Y(ori_ori_n609_));
  NO2        o0560(.A(ori_ori_n64_), .B(ori_ori_n55_), .Y(ori_ori_n610_));
  NO2        o0561(.A(ori_ori_n193_), .B(x5), .Y(ori_ori_n611_));
  NA2        o0562(.A(ori_ori_n104_), .B(ori_ori_n106_), .Y(ori_ori_n612_));
  NO2        o0563(.A(ori_ori_n612_), .B(ori_ori_n211_), .Y(ori_ori_n613_));
  AO220      o0564(.A0(ori_ori_n613_), .A1(ori_ori_n609_), .B0(ori_ori_n611_), .B1(ori_ori_n610_), .Y(ori_ori_n614_));
  OAI210     o0565(.A0(ori_ori_n614_), .A1(ori_ori_n608_), .B0(ori_ori_n493_), .Y(ori_ori_n615_));
  NO2        o0566(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n616_));
  NA2        o0567(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n617_));
  NO2        o0568(.A(ori_ori_n104_), .B(ori_ori_n106_), .Y(ori_ori_n618_));
  NA2        o0569(.A(ori_ori_n618_), .B(x7), .Y(ori_ori_n619_));
  NA2        o0570(.A(ori_ori_n434_), .B(ori_ori_n250_), .Y(ori_ori_n620_));
  AOI210     o0571(.A0(ori_ori_n620_), .A1(ori_ori_n619_), .B0(ori_ori_n617_), .Y(ori_ori_n621_));
  NA2        o0572(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n622_));
  XO2        o0573(.A(x7), .B(x5), .Y(ori_ori_n623_));
  NO2        o0574(.A(ori_ori_n623_), .B(ori_ori_n53_), .Y(ori_ori_n624_));
  NA3        o0575(.A(ori_ori_n624_), .B(ori_ori_n622_), .C(ori_ori_n326_), .Y(ori_ori_n625_));
  NO2        o0576(.A(ori_ori_n104_), .B(x2), .Y(ori_ori_n626_));
  NO2        o0577(.A(ori_ori_n75_), .B(ori_ori_n55_), .Y(ori_ori_n627_));
  NA2        o0578(.A(ori_ori_n627_), .B(ori_ori_n626_), .Y(ori_ori_n628_));
  NA2        o0579(.A(ori_ori_n628_), .B(ori_ori_n625_), .Y(ori_ori_n629_));
  OAI210     o0580(.A0(ori_ori_n629_), .A1(ori_ori_n621_), .B0(ori_ori_n616_), .Y(ori_ori_n630_));
  NO2        o0581(.A(ori_ori_n71_), .B(ori_ori_n50_), .Y(ori_ori_n631_));
  NO2        o0582(.A(ori_ori_n187_), .B(x4), .Y(ori_ori_n632_));
  NO2        o0583(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n633_));
  XO2        o0584(.A(x5), .B(x2), .Y(ori_ori_n634_));
  NO3        o0585(.A(x8), .B(x7), .C(ori_ori_n106_), .Y(ori_ori_n635_));
  AO220      o0586(.A0(ori_ori_n635_), .A1(ori_ori_n633_), .B0(ori_ori_n634_), .B1(ori_ori_n632_), .Y(ori_ori_n636_));
  NA3        o0587(.A(ori_ori_n636_), .B(ori_ori_n631_), .C(ori_ori_n53_), .Y(ori_ori_n637_));
  NA2        o0588(.A(ori_ori_n265_), .B(ori_ori_n587_), .Y(ori_ori_n638_));
  NOi21      o0589(.An(x4), .B(x1), .Y(ori_ori_n639_));
  NA2        o0590(.A(ori_ori_n639_), .B(ori_ori_n63_), .Y(ori_ori_n640_));
  NA2        o0591(.A(x4), .B(x1), .Y(ori_ori_n641_));
  NO2        o0592(.A(ori_ori_n641_), .B(ori_ori_n50_), .Y(ori_ori_n642_));
  AOI210     o0593(.A0(ori_ori_n642_), .A1(ori_ori_n618_), .B0(ori_ori_n59_), .Y(ori_ori_n643_));
  OA210      o0594(.A0(ori_ori_n640_), .A1(ori_ori_n638_), .B0(ori_ori_n643_), .Y(ori_ori_n644_));
  NA4        o0595(.A(ori_ori_n644_), .B(ori_ori_n637_), .C(ori_ori_n630_), .D(ori_ori_n615_), .Y(ori_ori_n645_));
  NA2        o0596(.A(ori_ori_n631_), .B(ori_ori_n56_), .Y(ori_ori_n646_));
  NA2        o0597(.A(ori_ori_n565_), .B(ori_ori_n603_), .Y(ori_ori_n647_));
  NO2        o0598(.A(ori_ori_n647_), .B(ori_ori_n646_), .Y(ori_ori_n648_));
  NA2        o0599(.A(ori_ori_n268_), .B(ori_ori_n118_), .Y(ori_ori_n649_));
  OAI210     o0600(.A0(ori_ori_n649_), .A1(ori_ori_n160_), .B0(ori_ori_n59_), .Y(ori_ori_n650_));
  NA2        o0601(.A(ori_ori_n57_), .B(x6), .Y(ori_ori_n651_));
  NA2        o0602(.A(ori_ori_n651_), .B(x3), .Y(ori_ori_n652_));
  NA2        o0603(.A(ori_ori_n633_), .B(ori_ori_n150_), .Y(ori_ori_n653_));
  NO3        o0604(.A(ori_ori_n653_), .B(ori_ori_n652_), .C(ori_ori_n424_), .Y(ori_ori_n654_));
  NA2        o0605(.A(ori_ori_n277_), .B(ori_ori_n71_), .Y(ori_ori_n655_));
  NO2        o0606(.A(ori_ori_n385_), .B(x3), .Y(ori_ori_n656_));
  NA2        o0607(.A(ori_ori_n656_), .B(ori_ori_n234_), .Y(ori_ori_n657_));
  NO2        o0608(.A(ori_ori_n424_), .B(ori_ori_n632_), .Y(ori_ori_n658_));
  NO2        o0609(.A(ori_ori_n466_), .B(ori_ori_n104_), .Y(ori_ori_n659_));
  NO2        o0610(.A(ori_ori_n575_), .B(x6), .Y(ori_ori_n660_));
  NA2        o0611(.A(ori_ori_n660_), .B(ori_ori_n659_), .Y(ori_ori_n661_));
  OAI220     o0612(.A0(ori_ori_n661_), .A1(ori_ori_n658_), .B0(ori_ori_n657_), .B1(ori_ori_n655_), .Y(ori_ori_n662_));
  NO4        o0613(.A(ori_ori_n662_), .B(ori_ori_n654_), .C(ori_ori_n650_), .D(ori_ori_n648_), .Y(ori_ori_n663_));
  NA2        o0614(.A(ori_ori_n57_), .B(x5), .Y(ori_ori_n664_));
  NO2        o0615(.A(ori_ori_n664_), .B(x1), .Y(ori_ori_n665_));
  NA2        o0616(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n666_));
  NO2        o0617(.A(ori_ori_n666_), .B(ori_ori_n124_), .Y(ori_ori_n667_));
  NA2        o0618(.A(x8), .B(x4), .Y(ori_ori_n668_));
  NO2        o0619(.A(x8), .B(x4), .Y(ori_ori_n669_));
  NAi21      o0620(.An(ori_ori_n669_), .B(ori_ori_n668_), .Y(ori_ori_n670_));
  NAi21      o0621(.An(ori_ori_n565_), .B(ori_ori_n385_), .Y(ori_ori_n671_));
  NO4        o0622(.A(ori_ori_n671_), .B(ori_ori_n670_), .C(ori_ori_n424_), .D(ori_ori_n71_), .Y(ori_ori_n672_));
  OAI210     o0623(.A0(ori_ori_n672_), .A1(ori_ori_n667_), .B0(ori_ori_n665_), .Y(ori_ori_n673_));
  NO3        o0624(.A(x8), .B(ori_ori_n104_), .C(x4), .Y(ori_ori_n674_));
  INV        o0625(.A(ori_ori_n674_), .Y(ori_ori_n675_));
  NO2        o0626(.A(ori_ori_n675_), .B(ori_ori_n106_), .Y(ori_ori_n676_));
  NO2        o0627(.A(x5), .B(x4), .Y(ori_ori_n677_));
  NA3        o0628(.A(ori_ori_n677_), .B(ori_ori_n63_), .C(ori_ori_n106_), .Y(ori_ori_n678_));
  NO2        o0629(.A(x6), .B(ori_ori_n106_), .Y(ori_ori_n679_));
  NA2        o0630(.A(ori_ori_n666_), .B(ori_ori_n679_), .Y(ori_ori_n680_));
  OAI210     o0631(.A0(ori_ori_n680_), .A1(ori_ori_n524_), .B0(ori_ori_n678_), .Y(ori_ori_n681_));
  OAI210     o0632(.A0(ori_ori_n681_), .A1(ori_ori_n676_), .B0(ori_ori_n307_), .Y(ori_ori_n682_));
  NA3        o0633(.A(ori_ori_n682_), .B(ori_ori_n673_), .C(ori_ori_n663_), .Y(ori_ori_n683_));
  OR2        o0634(.A(x4), .B(x1), .Y(ori_ori_n684_));
  NO2        o0635(.A(ori_ori_n684_), .B(x3), .Y(ori_ori_n685_));
  NA2        o0636(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n686_));
  NO3        o0637(.A(ori_ori_n366_), .B(ori_ori_n686_), .C(x6), .Y(ori_ori_n687_));
  AOI220     o0638(.A0(ori_ori_n687_), .A1(ori_ori_n685_), .B0(ori_ori_n683_), .B1(ori_ori_n645_), .Y(ori06));
  NA2        o0639(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n689_));
  NA2        o0640(.A(x6), .B(ori_ori_n106_), .Y(ori_ori_n690_));
  NA2        o0641(.A(ori_ori_n690_), .B(ori_ori_n55_), .Y(ori_ori_n691_));
  NA2        o0642(.A(x5), .B(ori_ori_n59_), .Y(ori_ori_n692_));
  NO2        o0643(.A(ori_ori_n692_), .B(ori_ori_n114_), .Y(ori_ori_n693_));
  NA3        o0644(.A(ori_ori_n693_), .B(ori_ori_n691_), .C(ori_ori_n499_), .Y(ori_ori_n694_));
  NO2        o0645(.A(ori_ori_n385_), .B(x0), .Y(ori_ori_n695_));
  NA2        o0646(.A(ori_ori_n336_), .B(x2), .Y(ori_ori_n696_));
  NOi21      o0647(.An(x6), .B(x8), .Y(ori_ori_n697_));
  NO2        o0648(.A(ori_ori_n697_), .B(x2), .Y(ori_ori_n698_));
  NO3        o0649(.A(ori_ori_n698_), .B(ori_ori_n70_), .C(ori_ori_n59_), .Y(ori_ori_n699_));
  AOI220     o0650(.A0(ori_ori_n699_), .A1(ori_ori_n696_), .B0(ori_ori_n695_), .B1(ori_ori_n328_), .Y(ori_ori_n700_));
  AOI210     o0651(.A0(ori_ori_n700_), .A1(ori_ori_n694_), .B0(ori_ori_n689_), .Y(ori_ori_n701_));
  NA2        o0652(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n702_));
  NA2        o0653(.A(ori_ori_n364_), .B(ori_ori_n352_), .Y(ori_ori_n703_));
  NO2        o0654(.A(ori_ori_n71_), .B(ori_ori_n104_), .Y(ori_ori_n704_));
  NO2        o0655(.A(ori_ori_n53_), .B(ori_ori_n59_), .Y(ori_ori_n705_));
  NO4        o0656(.A(ori_ori_n705_), .B(ori_ori_n686_), .C(ori_ori_n704_), .D(ori_ori_n493_), .Y(ori_ori_n706_));
  AOI220     o0657(.A0(ori_ori_n706_), .A1(ori_ori_n703_), .B0(ori_ori_n421_), .B1(ori_ori_n63_), .Y(ori_ori_n707_));
  NO2        o0658(.A(ori_ori_n707_), .B(ori_ori_n702_), .Y(ori_ori_n708_));
  NO2        o0659(.A(ori_ori_n54_), .B(x0), .Y(ori_ori_n709_));
  NA2        o0660(.A(x4), .B(x3), .Y(ori_ori_n710_));
  OAI210     o0661(.A0(ori_ori_n710_), .A1(x8), .B0(ori_ori_n517_), .Y(ori_ori_n711_));
  NA2        o0662(.A(ori_ori_n711_), .B(ori_ori_n709_), .Y(ori_ori_n712_));
  NO2        o0663(.A(ori_ori_n100_), .B(ori_ori_n56_), .Y(ori_ori_n713_));
  NA3        o0664(.A(ori_ori_n713_), .B(ori_ori_n251_), .C(ori_ori_n405_), .Y(ori_ori_n714_));
  AOI210     o0665(.A0(ori_ori_n714_), .A1(ori_ori_n712_), .B0(x2), .Y(ori_ori_n715_));
  INV        o0666(.A(ori_ori_n381_), .Y(ori_ori_n716_));
  NO2        o0667(.A(ori_ori_n408_), .B(x8), .Y(ori_ori_n717_));
  NO2        o0668(.A(ori_ori_n252_), .B(ori_ori_n519_), .Y(ori_ori_n718_));
  AOI210     o0669(.A0(ori_ori_n717_), .A1(ori_ori_n260_), .B0(ori_ori_n718_), .Y(ori_ori_n719_));
  NO2        o0670(.A(x5), .B(x3), .Y(ori_ori_n720_));
  NA3        o0671(.A(ori_ori_n552_), .B(ori_ori_n720_), .C(x1), .Y(ori_ori_n721_));
  NA2        o0672(.A(ori_ori_n604_), .B(ori_ori_n556_), .Y(ori_ori_n722_));
  OA220      o0673(.A0(ori_ori_n722_), .A1(ori_ori_n580_), .B0(ori_ori_n721_), .B1(ori_ori_n499_), .Y(ori_ori_n723_));
  OAI210     o0674(.A0(ori_ori_n719_), .A1(ori_ori_n716_), .B0(ori_ori_n723_), .Y(ori_ori_n724_));
  OR4        o0675(.A(ori_ori_n724_), .B(ori_ori_n715_), .C(ori_ori_n708_), .D(ori_ori_n701_), .Y(ori_ori_n725_));
  NA2        o0676(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n726_));
  NO2        o0677(.A(ori_ori_n618_), .B(ori_ori_n59_), .Y(ori_ori_n727_));
  NA2        o0678(.A(ori_ori_n727_), .B(ori_ori_n631_), .Y(ori_ori_n728_));
  NO2        o0679(.A(ori_ori_n166_), .B(x6), .Y(ori_ori_n729_));
  NA2        o0680(.A(ori_ori_n729_), .B(ori_ori_n286_), .Y(ori_ori_n730_));
  AOI210     o0681(.A0(ori_ori_n730_), .A1(ori_ori_n728_), .B0(ori_ori_n726_), .Y(ori_ori_n731_));
  AN2        o0682(.A(ori_ori_n471_), .B(ori_ori_n318_), .Y(ori_ori_n732_));
  OAI210     o0683(.A0(ori_ori_n732_), .A1(ori_ori_n731_), .B0(ori_ori_n347_), .Y(ori_ori_n733_));
  NO2        o0684(.A(ori_ori_n303_), .B(ori_ori_n104_), .Y(ori_ori_n734_));
  NO2        o0685(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n735_));
  NA2        o0686(.A(ori_ori_n735_), .B(ori_ori_n71_), .Y(ori_ori_n736_));
  NO2        o0687(.A(ori_ori_n736_), .B(ori_ori_n246_), .Y(ori_ori_n737_));
  NO2        o0688(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n738_));
  NA3        o0689(.A(ori_ori_n738_), .B(ori_ori_n572_), .C(ori_ori_n56_), .Y(ori_ori_n739_));
  NO2        o0690(.A(ori_ori_n57_), .B(x6), .Y(ori_ori_n740_));
  NA2        o0691(.A(ori_ori_n176_), .B(ori_ori_n740_), .Y(ori_ori_n741_));
  NA3        o0692(.A(ori_ori_n604_), .B(ori_ori_n325_), .C(ori_ori_n71_), .Y(ori_ori_n742_));
  NA3        o0693(.A(ori_ori_n742_), .B(ori_ori_n741_), .C(ori_ori_n739_), .Y(ori_ori_n743_));
  OR3        o0694(.A(ori_ori_n743_), .B(ori_ori_n737_), .C(ori_ori_n642_), .Y(ori_ori_n744_));
  NA2        o0695(.A(ori_ori_n744_), .B(ori_ori_n734_), .Y(ori_ori_n745_));
  NA2        o0696(.A(ori_ori_n709_), .B(ori_ori_n631_), .Y(ori_ori_n746_));
  NA4        o0697(.A(ori_ori_n261_), .B(ori_ori_n588_), .C(ori_ori_n215_), .D(ori_ori_n253_), .Y(ori_ori_n747_));
  NA2        o0698(.A(ori_ori_n482_), .B(ori_ori_n67_), .Y(ori_ori_n748_));
  AOI210     o0699(.A0(ori_ori_n747_), .A1(ori_ori_n746_), .B0(ori_ori_n748_), .Y(ori_ori_n749_));
  NA2        o0700(.A(x7), .B(x6), .Y(ori_ori_n750_));
  NA3        o0701(.A(x2), .B(x1), .C(x0), .Y(ori_ori_n751_));
  NO3        o0702(.A(ori_ori_n751_), .B(ori_ori_n750_), .C(ori_ori_n601_), .Y(ori_ori_n752_));
  NA2        o0703(.A(ori_ori_n494_), .B(ori_ori_n143_), .Y(ori_ori_n753_));
  NO2        o0704(.A(x5), .B(x1), .Y(ori_ori_n754_));
  NA2        o0705(.A(ori_ori_n754_), .B(ori_ori_n740_), .Y(ori_ori_n755_));
  NA2        o0706(.A(x4), .B(x0), .Y(ori_ori_n756_));
  NO3        o0707(.A(ori_ori_n57_), .B(x6), .C(x2), .Y(ori_ori_n757_));
  NA2        o0708(.A(ori_ori_n757_), .B(ori_ori_n219_), .Y(ori_ori_n758_));
  NO2        o0709(.A(ori_ori_n758_), .B(ori_ori_n756_), .Y(ori_ori_n759_));
  NO3        o0710(.A(ori_ori_n759_), .B(ori_ori_n752_), .C(ori_ori_n749_), .Y(ori_ori_n760_));
  NA3        o0711(.A(ori_ori_n760_), .B(ori_ori_n745_), .C(ori_ori_n733_), .Y(ori_ori_n761_));
  AOI210     o0712(.A0(ori_ori_n725_), .A1(ori_ori_n57_), .B0(ori_ori_n761_), .Y(ori07));
  NA2        o0713(.A(ori_ori_n104_), .B(ori_ori_n59_), .Y(ori_ori_n763_));
  NOi21      o0714(.An(ori_ori_n750_), .B(ori_ori_n112_), .Y(ori_ori_n764_));
  NO4        o0715(.A(ori_ori_n764_), .B(ori_ori_n631_), .C(ori_ori_n246_), .D(ori_ori_n763_), .Y(ori_ori_n765_));
  NO3        o0716(.A(ori_ori_n57_), .B(x5), .C(x1), .Y(ori_ori_n766_));
  NA2        o0717(.A(ori_ori_n766_), .B(ori_ori_n372_), .Y(ori_ori_n767_));
  NO2        o0718(.A(ori_ori_n57_), .B(ori_ori_n71_), .Y(ori_ori_n768_));
  NO2        o0719(.A(ori_ori_n149_), .B(ori_ori_n105_), .Y(ori_ori_n769_));
  AOI210     o0720(.A0(ori_ori_n768_), .A1(ori_ori_n90_), .B0(ori_ori_n769_), .Y(ori_ori_n770_));
  OAI220     o0721(.A0(ori_ori_n770_), .A1(ori_ori_n129_), .B0(ori_ori_n767_), .B1(ori_ori_n320_), .Y(ori_ori_n771_));
  OAI210     o0722(.A0(ori_ori_n771_), .A1(ori_ori_n765_), .B0(x2), .Y(ori_ori_n772_));
  NAi21      o0723(.An(ori_ori_n150_), .B(ori_ori_n151_), .Y(ori_ori_n773_));
  NA3        o0724(.A(ori_ori_n773_), .B(ori_ori_n89_), .C(x3), .Y(ori_ori_n774_));
  NO3        o0725(.A(ori_ori_n55_), .B(x3), .C(x1), .Y(ori_ori_n775_));
  NO2        o0726(.A(ori_ori_n512_), .B(x2), .Y(ori_ori_n776_));
  AOI210     o0727(.A0(ori_ori_n776_), .A1(ori_ori_n514_), .B0(ori_ori_n775_), .Y(ori_ori_n777_));
  OAI210     o0728(.A0(ori_ori_n777_), .A1(ori_ori_n651_), .B0(ori_ori_n774_), .Y(ori_ori_n778_));
  NO2        o0729(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n779_));
  NA2        o0730(.A(ori_ori_n779_), .B(ori_ori_n59_), .Y(ori_ori_n780_));
  NA2        o0731(.A(ori_ori_n353_), .B(ori_ori_n347_), .Y(ori_ori_n781_));
  NO2        o0732(.A(x7), .B(x3), .Y(ori_ori_n782_));
  NA2        o0733(.A(ori_ori_n782_), .B(ori_ori_n97_), .Y(ori_ori_n783_));
  AOI210     o0734(.A0(ori_ori_n781_), .A1(ori_ori_n780_), .B0(ori_ori_n783_), .Y(ori_ori_n784_));
  AOI210     o0735(.A0(ori_ori_n778_), .A1(ori_ori_n245_), .B0(ori_ori_n784_), .Y(ori_ori_n785_));
  AOI210     o0736(.A0(ori_ori_n785_), .A1(ori_ori_n772_), .B0(x4), .Y(ori_ori_n786_));
  NA3        o0737(.A(ori_ori_n754_), .B(ori_ori_n316_), .C(ori_ori_n55_), .Y(ori_ori_n787_));
  AOI210     o0738(.A0(ori_ori_n787_), .A1(ori_ori_n597_), .B0(ori_ori_n106_), .Y(ori_ori_n788_));
  XO2        o0739(.A(x5), .B(x1), .Y(ori_ori_n789_));
  NO4        o0740(.A(ori_ori_n789_), .B(ori_ori_n159_), .C(ori_ori_n202_), .D(ori_ori_n55_), .Y(ori_ori_n790_));
  OAI210     o0741(.A0(ori_ori_n790_), .A1(ori_ori_n788_), .B0(ori_ori_n412_), .Y(ori_ori_n791_));
  NO3        o0742(.A(ori_ori_n50_), .B(x2), .C(x0), .Y(ori_ori_n792_));
  NO2        o0743(.A(ori_ori_n306_), .B(ori_ori_n104_), .Y(ori_ori_n793_));
  NA2        o0744(.A(x6), .B(x0), .Y(ori_ori_n794_));
  NO2        o0745(.A(ori_ori_n686_), .B(ori_ori_n794_), .Y(ori_ori_n795_));
  NO2        o0746(.A(ori_ori_n789_), .B(ori_ori_n697_), .Y(ori_ori_n796_));
  OAI210     o0747(.A0(ori_ori_n754_), .A1(ori_ori_n63_), .B0(ori_ori_n57_), .Y(ori_ori_n797_));
  OAI210     o0748(.A0(ori_ori_n797_), .A1(ori_ori_n796_), .B0(ori_ori_n767_), .Y(ori_ori_n798_));
  AOI220     o0749(.A0(ori_ori_n798_), .A1(ori_ori_n792_), .B0(ori_ori_n795_), .B1(ori_ori_n793_), .Y(ori_ori_n799_));
  AOI210     o0750(.A0(ori_ori_n799_), .A1(ori_ori_n791_), .B0(ori_ori_n56_), .Y(ori_ori_n800_));
  NOi21      o0751(.An(ori_ori_n226_), .B(ori_ori_n372_), .Y(ori_ori_n801_));
  NO3        o0752(.A(ori_ori_n801_), .B(ori_ori_n235_), .C(ori_ori_n67_), .Y(ori_ori_n802_));
  NO2        o0753(.A(ori_ori_n185_), .B(ori_ori_n71_), .Y(ori_ori_n803_));
  NO2        o0754(.A(ori_ori_n306_), .B(x6), .Y(ori_ori_n804_));
  AO220      o0755(.A0(ori_ori_n804_), .A1(ori_ori_n326_), .B0(ori_ori_n803_), .B1(ori_ori_n557_), .Y(ori_ori_n805_));
  OAI210     o0756(.A0(ori_ori_n805_), .A1(ori_ori_n802_), .B0(ori_ori_n59_), .Y(ori_ori_n806_));
  NA2        o0757(.A(ori_ori_n90_), .B(ori_ori_n71_), .Y(ori_ori_n807_));
  NO2        o0758(.A(ori_ori_n807_), .B(ori_ori_n647_), .Y(ori_ori_n808_));
  NAi21      o0759(.An(x8), .B(x7), .Y(ori_ori_n809_));
  NA2        o0760(.A(ori_ori_n801_), .B(ori_ori_n809_), .Y(ori_ori_n810_));
  NA2        o0761(.A(ori_ori_n405_), .B(ori_ori_n106_), .Y(ori_ori_n811_));
  NO2        o0762(.A(ori_ori_n697_), .B(x1), .Y(ori_ori_n812_));
  NO3        o0763(.A(ori_ori_n812_), .B(ori_ori_n811_), .C(ori_ori_n572_), .Y(ori_ori_n813_));
  AOI210     o0764(.A0(ori_ori_n813_), .A1(ori_ori_n810_), .B0(ori_ori_n808_), .Y(ori_ori_n814_));
  AOI210     o0765(.A0(ori_ori_n814_), .A1(ori_ori_n806_), .B0(ori_ori_n136_), .Y(ori_ori_n815_));
  NO2        o0766(.A(x8), .B(x7), .Y(ori_ori_n816_));
  NO2        o0767(.A(ori_ori_n816_), .B(x3), .Y(ori_ori_n817_));
  NA3        o0768(.A(ori_ori_n817_), .B(ori_ori_n361_), .C(x1), .Y(ori_ori_n818_));
  NO2        o0769(.A(x8), .B(ori_ori_n106_), .Y(ori_ori_n819_));
  AOI220     o0770(.A0(ori_ori_n325_), .A1(ori_ori_n347_), .B0(ori_ori_n819_), .B1(ori_ori_n250_), .Y(ori_ori_n820_));
  NO2        o0771(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n821_));
  NA2        o0772(.A(ori_ori_n821_), .B(ori_ori_n300_), .Y(ori_ori_n822_));
  AOI210     o0773(.A0(ori_ori_n820_), .A1(ori_ori_n818_), .B0(ori_ori_n822_), .Y(ori_ori_n823_));
  NO4        o0774(.A(ori_ori_n823_), .B(ori_ori_n815_), .C(ori_ori_n800_), .D(ori_ori_n786_), .Y(ori08));
  NA2        o0775(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n825_));
  XN2        o0776(.A(x5), .B(x4), .Y(ori_ori_n826_));
  INV        o0777(.A(ori_ori_n826_), .Y(ori_ori_n827_));
  AOI220     o0778(.A0(ori_ori_n827_), .A1(ori_ori_n353_), .B0(ori_ori_n132_), .B1(ori_ori_n56_), .Y(ori_ori_n828_));
  NO2        o0779(.A(ori_ori_n237_), .B(ori_ori_n104_), .Y(ori_ori_n829_));
  AOI210     o0780(.A0(ori_ori_n829_), .A1(ori_ori_n274_), .B0(ori_ori_n186_), .Y(ori_ori_n830_));
  OAI220     o0781(.A0(ori_ori_n830_), .A1(x4), .B0(ori_ori_n828_), .B1(ori_ori_n825_), .Y(ori_ori_n831_));
  NA2        o0782(.A(ori_ori_n831_), .B(ori_ori_n268_), .Y(ori_ori_n832_));
  AOI210     o0783(.A0(ori_ori_n267_), .A1(ori_ori_n811_), .B0(ori_ori_n617_), .Y(ori_ori_n833_));
  NA2        o0784(.A(ori_ori_n612_), .B(ori_ori_n166_), .Y(ori_ori_n834_));
  OAI220     o0785(.A0(ori_ori_n834_), .A1(ori_ori_n666_), .B0(ori_ori_n484_), .B1(ori_ori_n50_), .Y(ori_ori_n835_));
  AO210      o0786(.A0(ori_ori_n835_), .A1(ori_ori_n340_), .B0(ori_ori_n833_), .Y(ori_ori_n836_));
  NA2        o0787(.A(ori_ori_n274_), .B(ori_ori_n143_), .Y(ori_ori_n837_));
  NA2        o0788(.A(ori_ori_n136_), .B(x7), .Y(ori_ori_n838_));
  OR3        o0789(.A(ori_ori_n751_), .B(ori_ori_n466_), .C(ori_ori_n720_), .Y(ori_ori_n839_));
  OAI220     o0790(.A0(ori_ori_n839_), .A1(ori_ori_n838_), .B0(ori_ori_n837_), .B1(ori_ori_n199_), .Y(ori_ori_n840_));
  AOI210     o0791(.A0(ori_ori_n836_), .A1(ori_ori_n288_), .B0(ori_ori_n840_), .Y(ori_ori_n841_));
  AOI210     o0792(.A0(ori_ori_n841_), .A1(ori_ori_n832_), .B0(ori_ori_n71_), .Y(ori_ori_n842_));
  NO2        o0793(.A(ori_ori_n816_), .B(ori_ori_n106_), .Y(ori_ori_n843_));
  NA2        o0794(.A(ori_ori_n843_), .B(ori_ori_n187_), .Y(ori_ori_n844_));
  OAI210     o0795(.A0(ori_ori_n408_), .A1(ori_ori_n300_), .B0(ori_ori_n340_), .Y(ori_ori_n845_));
  NA2        o0796(.A(ori_ori_n434_), .B(ori_ori_n228_), .Y(ori_ori_n846_));
  NA2        o0797(.A(ori_ori_n717_), .B(ori_ori_n103_), .Y(ori_ori_n847_));
  OAI220     o0798(.A0(ori_ori_n847_), .A1(ori_ori_n846_), .B0(ori_ori_n845_), .B1(ori_ori_n844_), .Y(ori_ori_n848_));
  NA2        o0799(.A(ori_ori_n848_), .B(ori_ori_n284_), .Y(ori_ori_n849_));
  NA2        o0800(.A(ori_ori_n330_), .B(ori_ori_n53_), .Y(ori_ori_n850_));
  NO3        o0801(.A(ori_ori_n408_), .B(ori_ori_n129_), .C(ori_ori_n68_), .Y(ori_ori_n851_));
  NO2        o0802(.A(ori_ori_n705_), .B(ori_ori_n240_), .Y(ori_ori_n852_));
  NO3        o0803(.A(ori_ori_n566_), .B(ori_ori_n467_), .C(ori_ori_n95_), .Y(ori_ori_n853_));
  AO220      o0804(.A0(ori_ori_n853_), .A1(ori_ori_n852_), .B0(ori_ori_n851_), .B1(ori_ori_n850_), .Y(ori_ori_n854_));
  NA2        o0805(.A(x7), .B(ori_ori_n59_), .Y(ori_ori_n855_));
  NO3        o0806(.A(ori_ori_n309_), .B(ori_ori_n855_), .C(ori_ori_n283_), .Y(ori_ori_n856_));
  AOI210     o0807(.A0(ori_ori_n854_), .A1(x5), .B0(ori_ori_n856_), .Y(ori_ori_n857_));
  AOI210     o0808(.A0(ori_ori_n857_), .A1(ori_ori_n849_), .B0(ori_ori_n72_), .Y(ori_ori_n858_));
  NO2        o0809(.A(ori_ori_n70_), .B(x3), .Y(ori_ori_n859_));
  OAI210     o0810(.A0(ori_ori_n859_), .A1(ori_ori_n259_), .B0(ori_ori_n141_), .Y(ori_ori_n860_));
  MUX2       o0811(.S(x3), .A(ori_ori_n159_), .B(ori_ori_n773_), .Y(ori_ori_n861_));
  NA2        o0812(.A(ori_ori_n861_), .B(ori_ori_n557_), .Y(ori_ori_n862_));
  NO3        o0813(.A(x6), .B(x4), .C(x0), .Y(ori_ori_n863_));
  INV        o0814(.A(ori_ori_n863_), .Y(ori_ori_n864_));
  AOI210     o0815(.A0(ori_ori_n862_), .A1(ori_ori_n860_), .B0(ori_ori_n864_), .Y(ori_ori_n865_));
  NO3        o0816(.A(x5), .B(x3), .C(ori_ori_n106_), .Y(ori_ori_n866_));
  AOI220     o0817(.A0(ori_ori_n827_), .A1(ori_ori_n305_), .B0(ori_ori_n866_), .B1(ori_ori_n59_), .Y(ori_ori_n867_));
  OR2        o0818(.A(x8), .B(x1), .Y(ori_ori_n868_));
  NO3        o0819(.A(ori_ori_n868_), .B(ori_ori_n867_), .C(ori_ori_n735_), .Y(ori_ori_n869_));
  NAi21      o0820(.An(x4), .B(x1), .Y(ori_ori_n870_));
  NO2        o0821(.A(ori_ori_n870_), .B(x0), .Y(ori_ori_n871_));
  NA2        o0822(.A(ori_ori_n611_), .B(ori_ori_n871_), .Y(ori_ori_n872_));
  NA3        o0823(.A(ori_ori_n55_), .B(x1), .C(x0), .Y(ori_ori_n873_));
  OAI210     o0824(.A0(ori_ori_n873_), .A1(ori_ori_n716_), .B0(ori_ori_n872_), .Y(ori_ori_n874_));
  OAI210     o0825(.A0(ori_ori_n874_), .A1(ori_ori_n869_), .B0(ori_ori_n316_), .Y(ori_ori_n875_));
  AO210      o0826(.A0(ori_ori_n286_), .A1(ori_ori_n259_), .B0(ori_ori_n734_), .Y(ori_ori_n876_));
  NA2        o0827(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n877_));
  NO2        o0828(.A(ori_ori_n877_), .B(ori_ori_n255_), .Y(ori_ori_n878_));
  NO2        o0829(.A(ori_ori_n57_), .B(x2), .Y(ori_ori_n879_));
  NO4        o0830(.A(ori_ori_n326_), .B(ori_ori_n879_), .C(ori_ori_n816_), .D(ori_ori_n290_), .Y(ori_ori_n880_));
  AOI220     o0831(.A0(ori_ori_n880_), .A1(ori_ori_n878_), .B0(ori_ori_n876_), .B1(ori_ori_n642_), .Y(ori_ori_n881_));
  NA2        o0832(.A(ori_ori_n881_), .B(ori_ori_n875_), .Y(ori_ori_n882_));
  NO4        o0833(.A(ori_ori_n882_), .B(ori_ori_n865_), .C(ori_ori_n858_), .D(ori_ori_n842_), .Y(ori09));
  NO3        o0834(.A(ori_ori_n789_), .B(ori_ori_n116_), .C(ori_ori_n92_), .Y(ori_ori_n884_));
  AOI220     o0835(.A0(ori_ori_n295_), .A1(ori_ori_n70_), .B0(ori_ori_n587_), .B1(ori_ori_n539_), .Y(ori_ori_n885_));
  OAI210     o0836(.A0(ori_ori_n884_), .A1(x2), .B0(ori_ori_n885_), .Y(ori_ori_n886_));
  AOI210     o0837(.A0(ori_ori_n886_), .A1(ori_ori_n755_), .B0(ori_ori_n443_), .Y(ori_ori_n887_));
  NO2        o0838(.A(ori_ori_n586_), .B(ori_ori_n258_), .Y(ori_ori_n888_));
  NO2        o0839(.A(ori_ori_n754_), .B(ori_ori_n336_), .Y(ori_ori_n889_));
  NO3        o0840(.A(ori_ori_n603_), .B(ori_ori_n98_), .C(ori_ori_n106_), .Y(ori_ori_n890_));
  AO220      o0841(.A0(ori_ori_n890_), .A1(ori_ori_n889_), .B0(ori_ori_n888_), .B1(ori_ori_n618_), .Y(ori_ori_n891_));
  OAI210     o0842(.A0(ori_ori_n891_), .A1(ori_ori_n887_), .B0(x4), .Y(ori_ori_n892_));
  OAI220     o0843(.A0(ori_ori_n364_), .A1(ori_ori_n138_), .B0(ori_ori_n392_), .B1(ori_ori_n276_), .Y(ori_ori_n893_));
  NO2        o0844(.A(ori_ori_n185_), .B(ori_ori_n104_), .Y(ori_ori_n894_));
  AOI220     o0845(.A0(ori_ori_n894_), .A1(ori_ori_n121_), .B0(ori_ori_n893_), .B1(ori_ori_n624_), .Y(ori_ori_n895_));
  NO2        o0846(.A(ori_ori_n789_), .B(ori_ori_n92_), .Y(ori_ori_n896_));
  NAi21      o0847(.An(x0), .B(x2), .Y(ori_ori_n897_));
  NO2        o0848(.A(ori_ori_n299_), .B(ori_ori_n897_), .Y(ori_ori_n898_));
  OAI210     o0849(.A0(ori_ori_n476_), .A1(ori_ori_n271_), .B0(ori_ori_n185_), .Y(ori_ori_n899_));
  AOI210     o0850(.A0(ori_ori_n162_), .A1(ori_ori_n809_), .B0(ori_ori_n352_), .Y(ori_ori_n900_));
  AOI220     o0851(.A0(ori_ori_n900_), .A1(ori_ori_n899_), .B0(ori_ori_n898_), .B1(ori_ori_n896_), .Y(ori_ori_n901_));
  OAI210     o0852(.A0(ori_ori_n895_), .A1(ori_ori_n55_), .B0(ori_ori_n901_), .Y(ori_ori_n902_));
  NA2        o0853(.A(ori_ori_n902_), .B(ori_ori_n56_), .Y(ori_ori_n903_));
  NO2        o0854(.A(ori_ori_n56_), .B(ori_ori_n59_), .Y(ori_ori_n904_));
  INV        o0855(.A(ori_ori_n121_), .Y(ori_ori_n905_));
  NA2        o0856(.A(ori_ori_n754_), .B(ori_ori_n55_), .Y(ori_ori_n906_));
  AOI210     o0857(.A0(x6), .A1(x1), .B0(x5), .Y(ori_ori_n907_));
  OAI210     o0858(.A0(ori_ori_n907_), .A1(ori_ori_n329_), .B0(x2), .Y(ori_ori_n908_));
  AOI210     o0859(.A0(ori_ori_n908_), .A1(ori_ori_n906_), .B0(ori_ori_n905_), .Y(ori_ori_n909_));
  NA2        o0860(.A(ori_ori_n556_), .B(ori_ori_n55_), .Y(ori_ori_n910_));
  NO2        o0861(.A(ori_ori_n225_), .B(ori_ori_n382_), .Y(ori_ori_n911_));
  NO2        o0862(.A(ori_ori_n306_), .B(ori_ori_n142_), .Y(ori_ori_n912_));
  NO2        o0863(.A(ori_ori_n912_), .B(ori_ori_n911_), .Y(ori_ori_n913_));
  OAI220     o0864(.A0(ori_ori_n913_), .A1(ori_ori_n55_), .B0(ori_ori_n910_), .B1(ori_ori_n455_), .Y(ori_ori_n914_));
  OAI210     o0865(.A0(ori_ori_n914_), .A1(ori_ori_n909_), .B0(ori_ori_n904_), .Y(ori_ori_n915_));
  NO2        o0866(.A(ori_ori_n401_), .B(ori_ori_n104_), .Y(ori_ori_n916_));
  NO2        o0867(.A(ori_ori_n330_), .B(ori_ori_n493_), .Y(ori_ori_n917_));
  AOI220     o0868(.A0(ori_ori_n917_), .A1(ori_ori_n916_), .B0(ori_ori_n203_), .B1(ori_ori_n223_), .Y(ori_ori_n918_));
  NA4        o0869(.A(ori_ori_n918_), .B(ori_ori_n915_), .C(ori_ori_n903_), .D(ori_ori_n892_), .Y(ori_ori_n919_));
  NA2        o0870(.A(ori_ori_n919_), .B(ori_ori_n50_), .Y(ori_ori_n920_));
  NO2        o0871(.A(ori_ori_n375_), .B(ori_ori_n155_), .Y(ori_ori_n921_));
  NA2        o0872(.A(ori_ori_n234_), .B(ori_ori_n587_), .Y(ori_ori_n922_));
  OAI210     o0873(.A0(ori_ori_n429_), .A1(ori_ori_n819_), .B0(ori_ori_n922_), .Y(ori_ori_n923_));
  OAI210     o0874(.A0(ori_ori_n923_), .A1(ori_ori_n921_), .B0(x0), .Y(ori_ori_n924_));
  NO3        o0875(.A(x8), .B(x7), .C(x2), .Y(ori_ori_n925_));
  NO3        o0876(.A(ori_ori_n57_), .B(x5), .C(x2), .Y(ori_ori_n926_));
  OAI210     o0877(.A0(ori_ori_n926_), .A1(ori_ori_n925_), .B0(ori_ori_n514_), .Y(ori_ori_n927_));
  AOI210     o0878(.A0(ori_ori_n927_), .A1(ori_ori_n924_), .B0(x4), .Y(ori_ori_n928_));
  NO2        o0879(.A(ori_ori_n422_), .B(ori_ori_n141_), .Y(ori_ori_n929_));
  NO2        o0880(.A(ori_ori_n52_), .B(x2), .Y(ori_ori_n930_));
  NO2        o0881(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n931_));
  NA2        o0882(.A(ori_ori_n931_), .B(x8), .Y(ori_ori_n932_));
  NA2        o0883(.A(ori_ori_n932_), .B(ori_ori_n906_), .Y(ori_ori_n933_));
  AO210      o0884(.A0(ori_ori_n933_), .A1(ori_ori_n930_), .B0(ori_ori_n929_), .Y(ori_ori_n934_));
  OAI210     o0885(.A0(ori_ori_n934_), .A1(ori_ori_n928_), .B0(ori_ori_n616_), .Y(ori_ori_n935_));
  NO2        o0886(.A(ori_ori_n254_), .B(ori_ori_n115_), .Y(ori_ori_n936_));
  OAI210     o0887(.A0(x4), .A1(x2), .B0(x0), .Y(ori_ori_n937_));
  NA3        o0888(.A(ori_ori_n605_), .B(ori_ori_n617_), .C(ori_ori_n341_), .Y(ori_ori_n938_));
  OAI210     o0889(.A0(ori_ori_n937_), .A1(ori_ori_n283_), .B0(ori_ori_n53_), .Y(ori_ori_n939_));
  AOI210     o0890(.A0(ori_ori_n938_), .A1(ori_ori_n937_), .B0(ori_ori_n939_), .Y(ori_ori_n940_));
  OAI210     o0891(.A0(ori_ori_n940_), .A1(ori_ori_n936_), .B0(ori_ori_n325_), .Y(ori_ori_n941_));
  AOI220     o0892(.A0(ori_ori_n668_), .A1(ori_ori_n345_), .B0(ori_ori_n347_), .B1(ori_ori_n91_), .Y(ori_ori_n942_));
  NA2        o0893(.A(ori_ori_n91_), .B(x5), .Y(ori_ori_n943_));
  OAI220     o0894(.A0(ori_ori_n943_), .A1(ori_ori_n868_), .B0(ori_ori_n942_), .B1(ori_ori_n317_), .Y(ori_ori_n944_));
  NA2        o0895(.A(ori_ori_n944_), .B(ori_ori_n68_), .Y(ori_ori_n945_));
  NA2        o0896(.A(ori_ori_n405_), .B(ori_ori_n773_), .Y(ori_ori_n946_));
  NA2        o0897(.A(ori_ori_n245_), .B(ori_ori_n159_), .Y(ori_ori_n947_));
  AO210      o0898(.A0(ori_ori_n947_), .A1(ori_ori_n946_), .B0(ori_ori_n126_), .Y(ori_ori_n948_));
  NO2        o0899(.A(ori_ori_n435_), .B(x2), .Y(ori_ori_n949_));
  NO2        o0900(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n950_));
  NA2        o0901(.A(ori_ori_n950_), .B(x5), .Y(ori_ori_n951_));
  NO2        o0902(.A(ori_ori_n951_), .B(ori_ori_n60_), .Y(ori_ori_n952_));
  AOI220     o0903(.A0(ori_ori_n952_), .A1(ori_ori_n949_), .B0(ori_ori_n669_), .B1(ori_ori_n238_), .Y(ori_ori_n953_));
  NA4        o0904(.A(ori_ori_n953_), .B(ori_ori_n948_), .C(ori_ori_n945_), .D(ori_ori_n941_), .Y(ori_ori_n954_));
  NO4        o0905(.A(ori_ori_n938_), .B(ori_ori_n633_), .C(ori_ori_n455_), .D(ori_ori_n50_), .Y(ori_ori_n955_));
  AOI220     o0906(.A0(ori_ori_n604_), .A1(ori_ori_n603_), .B0(ori_ori_n277_), .B1(x5), .Y(ori_ori_n956_));
  NO2        o0907(.A(ori_ori_n677_), .B(ori_ori_n185_), .Y(ori_ori_n957_));
  NA3        o0908(.A(ori_ori_n957_), .B(ori_ori_n670_), .C(x7), .Y(ori_ori_n958_));
  OAI210     o0909(.A0(ori_ori_n956_), .A1(ori_ori_n346_), .B0(ori_ori_n958_), .Y(ori_ori_n959_));
  OAI210     o0910(.A0(ori_ori_n959_), .A1(ori_ori_n955_), .B0(ori_ori_n82_), .Y(ori_ori_n960_));
  NA2        o0911(.A(ori_ori_n779_), .B(x2), .Y(ori_ori_n961_));
  NO2        o0912(.A(ori_ori_n961_), .B(ori_ori_n58_), .Y(ori_ori_n962_));
  NO2        o0913(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n963_));
  NAi21      o0914(.An(x1), .B(x4), .Y(ori_ori_n964_));
  NA2        o0915(.A(ori_ori_n964_), .B(ori_ori_n870_), .Y(ori_ori_n965_));
  NO3        o0916(.A(ori_ori_n965_), .B(ori_ori_n196_), .C(ori_ori_n963_), .Y(ori_ori_n966_));
  OAI210     o0917(.A0(ori_ori_n966_), .A1(ori_ori_n962_), .B0(ori_ori_n412_), .Y(ori_ori_n967_));
  NA3        o0918(.A(ori_ori_n395_), .B(ori_ori_n754_), .C(ori_ori_n57_), .Y(ori_ori_n968_));
  NA3        o0919(.A(ori_ori_n968_), .B(ori_ori_n967_), .C(ori_ori_n960_), .Y(ori_ori_n969_));
  AOI210     o0920(.A0(ori_ori_n954_), .A1(x6), .B0(ori_ori_n969_), .Y(ori_ori_n970_));
  NA3        o0921(.A(ori_ori_n970_), .B(ori_ori_n935_), .C(ori_ori_n920_), .Y(ori10));
  NO2        o0922(.A(x4), .B(x1), .Y(ori_ori_n972_));
  NO2        o0923(.A(ori_ori_n972_), .B(ori_ori_n143_), .Y(ori_ori_n973_));
  NA3        o0924(.A(x5), .B(x4), .C(x0), .Y(ori_ori_n974_));
  OAI220     o0925(.A0(ori_ori_n974_), .A1(ori_ori_n272_), .B0(ori_ori_n705_), .B1(ori_ori_n242_), .Y(ori_ori_n975_));
  NA2        o0926(.A(ori_ori_n975_), .B(ori_ori_n973_), .Y(ori_ori_n976_));
  NO3        o0927(.A(ori_ori_n353_), .B(ori_ori_n317_), .C(ori_ori_n90_), .Y(ori_ori_n977_));
  NA3        o0928(.A(ori_ori_n977_), .B(ori_ori_n380_), .C(ori_ori_n62_), .Y(ori_ori_n978_));
  AOI210     o0929(.A0(ori_ori_n978_), .A1(ori_ori_n976_), .B0(ori_ori_n299_), .Y(ori_ori_n979_));
  NOi21      o0930(.An(ori_ori_n253_), .B(ori_ori_n132_), .Y(ori_ori_n980_));
  AOI210     o0931(.A0(ori_ori_n500_), .A1(ori_ori_n618_), .B0(ori_ori_n326_), .Y(ori_ori_n981_));
  NO2        o0932(.A(ori_ori_n904_), .B(ori_ori_n339_), .Y(ori_ori_n982_));
  NOi31      o0933(.An(ori_ori_n982_), .B(ori_ori_n981_), .C(ori_ori_n980_), .Y(ori_ori_n983_));
  NA2        o0934(.A(x4), .B(ori_ori_n106_), .Y(ori_ori_n984_));
  NO2        o0935(.A(ori_ori_n320_), .B(ori_ori_n984_), .Y(ori_ori_n985_));
  NA2        o0936(.A(ori_ori_n95_), .B(x5), .Y(ori_ori_n986_));
  NO3        o0937(.A(ori_ori_n986_), .B(ori_ori_n107_), .C(ori_ori_n55_), .Y(ori_ori_n987_));
  NO3        o0938(.A(ori_ori_n987_), .B(ori_ori_n985_), .C(ori_ori_n983_), .Y(ori_ori_n988_));
  NA2        o0939(.A(ori_ori_n963_), .B(ori_ori_n50_), .Y(ori_ori_n989_));
  NA2        o0940(.A(ori_ori_n604_), .B(ori_ori_n266_), .Y(ori_ori_n990_));
  NO2        o0941(.A(ori_ori_n990_), .B(ori_ori_n989_), .Y(ori_ori_n991_));
  OAI220     o0942(.A0(ori_ori_n932_), .A1(ori_ori_n103_), .B0(ori_ori_n877_), .B1(ori_ori_n443_), .Y(ori_ori_n992_));
  AOI210     o0943(.A0(ori_ori_n992_), .A1(ori_ori_n274_), .B0(ori_ori_n991_), .Y(ori_ori_n993_));
  OAI210     o0944(.A0(ori_ori_n988_), .A1(ori_ori_n382_), .B0(ori_ori_n993_), .Y(ori_ori_n994_));
  OAI210     o0945(.A0(ori_ori_n994_), .A1(ori_ori_n979_), .B0(x7), .Y(ori_ori_n995_));
  NA2        o0946(.A(ori_ori_n55_), .B(ori_ori_n71_), .Y(ori_ori_n996_));
  AOI210     o0947(.A0(ori_ori_n443_), .A1(ori_ori_n352_), .B0(ori_ori_n984_), .Y(ori_ori_n997_));
  NO3        o0948(.A(ori_ori_n445_), .B(ori_ori_n897_), .C(x5), .Y(ori_ori_n998_));
  OAI210     o0949(.A0(ori_ori_n998_), .A1(ori_ori_n997_), .B0(ori_ori_n996_), .Y(ori_ori_n999_));
  NO2        o0950(.A(ori_ori_n353_), .B(ori_ori_n135_), .Y(ori_ori_n1000_));
  NA2        o0951(.A(ori_ori_n1000_), .B(ori_ori_n423_), .Y(ori_ori_n1001_));
  AOI210     o0952(.A0(ori_ori_n1001_), .A1(ori_ori_n999_), .B0(x3), .Y(ori_ori_n1002_));
  NA2        o0953(.A(ori_ori_n697_), .B(ori_ori_n245_), .Y(ori_ori_n1003_));
  NO2        o0954(.A(x5), .B(ori_ori_n106_), .Y(ori_ori_n1004_));
  OAI210     o0955(.A0(ori_ori_n1004_), .A1(ori_ori_n232_), .B0(ori_ori_n943_), .Y(ori_ori_n1005_));
  NA3        o0956(.A(ori_ori_n462_), .B(ori_ori_n124_), .C(ori_ori_n423_), .Y(ori_ori_n1006_));
  OAI210     o0957(.A0(ori_ori_n445_), .A1(ori_ori_n208_), .B0(ori_ori_n1006_), .Y(ori_ori_n1007_));
  AOI210     o0958(.A0(ori_ori_n1005_), .A1(ori_ori_n251_), .B0(ori_ori_n1007_), .Y(ori_ori_n1008_));
  OAI220     o0959(.A0(ori_ori_n1008_), .A1(ori_ori_n59_), .B0(ori_ori_n1003_), .B1(ori_ori_n710_), .Y(ori_ori_n1009_));
  OAI210     o0960(.A0(ori_ori_n1009_), .A1(ori_ori_n1002_), .B0(ori_ori_n950_), .Y(ori_ori_n1010_));
  NO2        o0961(.A(x4), .B(x3), .Y(ori_ori_n1011_));
  NO3        o0962(.A(ori_ori_n1011_), .B(ori_ori_n340_), .C(ori_ori_n87_), .Y(ori_ori_n1012_));
  OAI210     o0963(.A0(ori_ori_n1012_), .A1(ori_ori_n273_), .B0(ori_ori_n434_), .Y(ori_ori_n1013_));
  AOI210     o0964(.A0(ori_ori_n396_), .A1(ori_ori_n123_), .B0(ori_ori_n246_), .Y(ori_ori_n1014_));
  NA2        o0965(.A(ori_ori_n972_), .B(ori_ori_n55_), .Y(ori_ori_n1015_));
  NO2        o0966(.A(ori_ori_n1015_), .B(ori_ori_n986_), .Y(ori_ori_n1016_));
  NO2        o0967(.A(ori_ori_n524_), .B(ori_ori_n358_), .Y(ori_ori_n1017_));
  NO3        o0968(.A(x4), .B(ori_ori_n106_), .C(ori_ori_n59_), .Y(ori_ori_n1018_));
  NO2        o0969(.A(ori_ori_n435_), .B(x1), .Y(ori_ori_n1019_));
  NOi31      o0970(.An(ori_ori_n1018_), .B(ori_ori_n1019_), .C(ori_ori_n1017_), .Y(ori_ori_n1020_));
  NA2        o0971(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n1021_));
  NO4        o0972(.A(ori_ori_n973_), .B(ori_ori_n513_), .C(ori_ori_n1021_), .D(x2), .Y(ori_ori_n1022_));
  NO4        o0973(.A(ori_ori_n1022_), .B(ori_ori_n1020_), .C(ori_ori_n1016_), .D(ori_ori_n1014_), .Y(ori_ori_n1023_));
  AOI210     o0974(.A0(ori_ori_n1023_), .A1(ori_ori_n1013_), .B0(ori_ori_n202_), .Y(ori_ori_n1024_));
  NO2        o0975(.A(ori_ori_n666_), .B(ori_ori_n499_), .Y(ori_ori_n1025_));
  NO2        o0976(.A(x6), .B(x2), .Y(ori_ori_n1026_));
  NO3        o0977(.A(ori_ori_n1026_), .B(ori_ori_n697_), .C(ori_ori_n60_), .Y(ori_ori_n1027_));
  OAI210     o0978(.A0(ori_ori_n1027_), .A1(ori_ori_n1025_), .B0(ori_ori_n265_), .Y(ori_ori_n1028_));
  NO2        o0979(.A(ori_ori_n877_), .B(ori_ori_n443_), .Y(ori_ori_n1029_));
  NA3        o0980(.A(x4), .B(x3), .C(ori_ori_n106_), .Y(ori_ori_n1030_));
  NO3        o0981(.A(ori_ori_n1030_), .B(ori_ori_n703_), .C(ori_ori_n462_), .Y(ori_ori_n1031_));
  AOI210     o0982(.A0(ori_ori_n1029_), .A1(ori_ori_n469_), .B0(ori_ori_n1031_), .Y(ori_ori_n1032_));
  AOI210     o0983(.A0(ori_ori_n1032_), .A1(ori_ori_n1028_), .B0(ori_ori_n455_), .Y(ori_ori_n1033_));
  NO2        o0984(.A(ori_ori_n55_), .B(ori_ori_n56_), .Y(ori_ori_n1034_));
  OAI220     o0985(.A0(ori_ori_n827_), .A1(ori_ori_n457_), .B0(ori_ori_n756_), .B1(ori_ori_n123_), .Y(ori_ori_n1035_));
  NOi21      o0986(.An(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n1036_));
  NO3        o0987(.A(ori_ori_n341_), .B(ori_ori_n320_), .C(ori_ori_n1036_), .Y(ori_ori_n1037_));
  AOI220     o0988(.A0(ori_ori_n1037_), .A1(ori_ori_n250_), .B0(ori_ori_n1035_), .B1(ori_ori_n112_), .Y(ori_ori_n1038_));
  NO2        o0989(.A(ori_ori_n1038_), .B(ori_ori_n1034_), .Y(ori_ori_n1039_));
  NA2        o0990(.A(ori_ori_n517_), .B(ori_ori_n255_), .Y(ori_ori_n1040_));
  NO2        o0991(.A(ori_ori_n484_), .B(ori_ori_n586_), .Y(ori_ori_n1041_));
  NA3        o0992(.A(ori_ori_n1041_), .B(ori_ori_n1040_), .C(ori_ori_n55_), .Y(ori_ori_n1042_));
  NO2        o0993(.A(ori_ori_n177_), .B(ori_ori_n106_), .Y(ori_ori_n1043_));
  NA3        o0994(.A(ori_ori_n1043_), .B(ori_ori_n176_), .C(ori_ori_n118_), .Y(ori_ori_n1044_));
  NA2        o0995(.A(ori_ori_n1044_), .B(ori_ori_n1042_), .Y(ori_ori_n1045_));
  NO4        o0996(.A(ori_ori_n1045_), .B(ori_ori_n1039_), .C(ori_ori_n1033_), .D(ori_ori_n1024_), .Y(ori_ori_n1046_));
  NA3        o0997(.A(ori_ori_n1046_), .B(ori_ori_n1010_), .C(ori_ori_n995_), .Y(ori11));
  NA2        o0998(.A(ori_ori_n373_), .B(ori_ori_n90_), .Y(ori_ori_n1048_));
  INV        o0999(.A(ori_ori_n898_), .Y(ori_ori_n1049_));
  OAI220     o1000(.A0(ori_ori_n1049_), .A1(ori_ori_n53_), .B0(ori_ori_n1048_), .B1(ori_ori_n362_), .Y(ori_ori_n1050_));
  NO2        o1001(.A(ori_ori_n773_), .B(x5), .Y(ori_ori_n1051_));
  NO2        o1002(.A(ori_ori_n163_), .B(ori_ori_n530_), .Y(ori_ori_n1052_));
  AOI220     o1003(.A0(ori_ori_n1052_), .A1(ori_ori_n1051_), .B0(ori_ori_n1050_), .B1(x5), .Y(ori_ori_n1053_));
  OAI220     o1004(.A0(ori_ori_n980_), .A1(ori_ori_n211_), .B0(ori_ori_n209_), .B1(ori_ori_n177_), .Y(ori_ori_n1054_));
  NO2        o1005(.A(ori_ori_n337_), .B(ori_ori_n424_), .Y(ori_ori_n1055_));
  AOI220     o1006(.A0(ori_ori_n1055_), .A1(ori_ori_n175_), .B0(ori_ori_n1054_), .B1(ori_ori_n159_), .Y(ori_ori_n1056_));
  NO2        o1007(.A(ori_ori_n1056_), .B(ori_ori_n445_), .Y(ori_ori_n1057_));
  NO2        o1008(.A(ori_ori_n246_), .B(x2), .Y(ori_ori_n1058_));
  OAI210     o1009(.A0(ori_ori_n921_), .A1(ori_ori_n1058_), .B0(ori_ori_n413_), .Y(ori_ori_n1059_));
  NO2        o1010(.A(ori_ori_n55_), .B(ori_ori_n104_), .Y(ori_ori_n1060_));
  NA2        o1011(.A(ori_ori_n274_), .B(ori_ori_n1060_), .Y(ori_ori_n1061_));
  NO2        o1012(.A(ori_ori_n71_), .B(x1), .Y(ori_ori_n1062_));
  NA2        o1013(.A(ori_ori_n1062_), .B(ori_ori_n78_), .Y(ori_ori_n1063_));
  OA220      o1014(.A0(ori_ori_n1063_), .A1(ori_ori_n612_), .B0(ori_ori_n1061_), .B1(ori_ori_n530_), .Y(ori_ori_n1064_));
  AOI210     o1015(.A0(ori_ori_n1064_), .A1(ori_ori_n1059_), .B0(ori_ori_n710_), .Y(ori_ori_n1065_));
  NO2        o1016(.A(ori_ori_n300_), .B(ori_ori_n53_), .Y(ori_ori_n1066_));
  NO2        o1017(.A(ori_ori_n434_), .B(x3), .Y(ori_ori_n1067_));
  NA3        o1018(.A(ori_ori_n1067_), .B(ori_ori_n1066_), .C(ori_ori_n897_), .Y(ori_ori_n1068_));
  AOI210     o1019(.A0(ori_ori_n1068_), .A1(ori_ori_n947_), .B0(ori_ori_n394_), .Y(ori_ori_n1069_));
  NA2        o1020(.A(ori_ori_n106_), .B(x1), .Y(ori_ori_n1070_));
  NO2        o1021(.A(ori_ori_n618_), .B(ori_ori_n214_), .Y(ori_ori_n1071_));
  NA4        o1022(.A(ori_ori_n1071_), .B(ori_ori_n889_), .C(ori_ori_n466_), .D(ori_ori_n1070_), .Y(ori_ori_n1072_));
  NA3        o1023(.A(x6), .B(x5), .C(ori_ori_n106_), .Y(ori_ori_n1073_));
  NO2        o1024(.A(ori_ori_n1073_), .B(ori_ori_n272_), .Y(ori_ori_n1074_));
  NO2        o1025(.A(ori_ori_n445_), .B(x0), .Y(ori_ori_n1075_));
  NOi31      o1026(.An(ori_ori_n1075_), .B(ori_ori_n168_), .C(ori_ori_n51_), .Y(ori_ori_n1076_));
  AOI210     o1027(.A0(ori_ori_n1074_), .A1(ori_ori_n173_), .B0(ori_ori_n1076_), .Y(ori_ori_n1077_));
  NA2        o1028(.A(ori_ori_n1077_), .B(ori_ori_n1072_), .Y(ori_ori_n1078_));
  NO4        o1029(.A(ori_ori_n1078_), .B(ori_ori_n1069_), .C(ori_ori_n1065_), .D(ori_ori_n1057_), .Y(ori_ori_n1079_));
  OAI210     o1030(.A0(ori_ori_n1053_), .A1(ori_ori_n136_), .B0(ori_ori_n1079_), .Y(ori_ori_n1080_));
  NA2        o1031(.A(ori_ori_n868_), .B(ori_ori_n87_), .Y(ori_ori_n1081_));
  NO3        o1032(.A(ori_ori_n463_), .B(ori_ori_n779_), .C(ori_ori_n119_), .Y(ori_ori_n1082_));
  AOI210     o1033(.A0(ori_ori_n1081_), .A1(ori_ori_n97_), .B0(ori_ori_n1082_), .Y(ori_ori_n1083_));
  NO2        o1034(.A(x8), .B(x1), .Y(ori_ori_n1084_));
  NO3        o1035(.A(ori_ori_n1084_), .B(ori_ori_n689_), .C(ori_ori_n447_), .Y(ori_ori_n1085_));
  OAI210     o1036(.A0(ori_ori_n77_), .A1(ori_ori_n53_), .B0(ori_ori_n1085_), .Y(ori_ori_n1086_));
  OAI210     o1037(.A0(ori_ori_n1083_), .A1(x3), .B0(ori_ori_n1086_), .Y(ori_ori_n1087_));
  NO2        o1038(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n1088_));
  OAI210     o1039(.A0(ori_ori_n1088_), .A1(x2), .B0(ori_ori_n228_), .Y(ori_ori_n1089_));
  NO2        o1040(.A(ori_ori_n605_), .B(ori_ori_n226_), .Y(ori_ori_n1090_));
  NA2        o1041(.A(ori_ori_n1090_), .B(ori_ori_n1089_), .Y(ori_ori_n1091_));
  NO2        o1042(.A(ori_ori_n517_), .B(x4), .Y(ori_ori_n1092_));
  NO3        o1043(.A(ori_ori_n55_), .B(x6), .C(x1), .Y(ori_ori_n1093_));
  NOi21      o1044(.An(ori_ori_n1093_), .B(ori_ori_n484_), .Y(ori_ori_n1094_));
  AOI210     o1045(.A0(ori_ori_n1092_), .A1(ori_ori_n576_), .B0(ori_ori_n1094_), .Y(ori_ori_n1095_));
  NA2        o1046(.A(ori_ori_n1095_), .B(ori_ori_n1091_), .Y(ori_ori_n1096_));
  AOI210     o1047(.A0(ori_ori_n1087_), .A1(x2), .B0(ori_ori_n1096_), .Y(ori_ori_n1097_));
  NO2        o1048(.A(ori_ori_n226_), .B(x2), .Y(ori_ori_n1098_));
  NA2        o1049(.A(ori_ori_n1098_), .B(ori_ori_n1011_), .Y(ori_ori_n1099_));
  NOi21      o1050(.An(ori_ori_n385_), .B(ori_ori_n565_), .Y(ori_ori_n1100_));
  NO3        o1051(.A(ori_ori_n1100_), .B(ori_ori_n604_), .C(ori_ori_n320_), .Y(ori_ori_n1101_));
  NA2        o1052(.A(x8), .B(ori_ori_n106_), .Y(ori_ori_n1102_));
  OAI220     o1053(.A0(ori_ori_n710_), .A1(ori_ori_n1102_), .B0(ori_ori_n320_), .B1(ori_ori_n380_), .Y(ori_ori_n1103_));
  OAI210     o1054(.A0(ori_ori_n1103_), .A1(ori_ori_n1101_), .B0(ori_ori_n71_), .Y(ori_ori_n1104_));
  NO2        o1055(.A(ori_ori_n104_), .B(x1), .Y(ori_ori_n1105_));
  NA2        o1056(.A(ori_ori_n1105_), .B(x7), .Y(ori_ori_n1106_));
  AOI210     o1057(.A0(ori_ori_n1104_), .A1(ori_ori_n1099_), .B0(ori_ori_n1106_), .Y(ori_ori_n1107_));
  NA2        o1058(.A(ori_ori_n84_), .B(ori_ori_n71_), .Y(ori_ori_n1108_));
  INV        o1059(.A(ori_ori_n243_), .Y(ori_ori_n1109_));
  NA2        o1060(.A(ori_ori_n1109_), .B(ori_ori_n143_), .Y(ori_ori_n1110_));
  OAI220     o1061(.A0(ori_ori_n1110_), .A1(ori_ori_n362_), .B0(ori_ori_n1108_), .B1(ori_ori_n320_), .Y(ori_ori_n1111_));
  NO2        o1062(.A(ori_ori_n153_), .B(ori_ori_n55_), .Y(ori_ori_n1112_));
  AOI210     o1063(.A0(ori_ori_n1112_), .A1(ori_ori_n1111_), .B0(ori_ori_n1107_), .Y(ori_ori_n1113_));
  OAI210     o1064(.A0(ori_ori_n1097_), .A1(ori_ori_n855_), .B0(ori_ori_n1113_), .Y(ori_ori_n1114_));
  AO210      o1065(.A0(ori_ori_n1080_), .A1(ori_ori_n57_), .B0(ori_ori_n1114_), .Y(ori12));
  NA2        o1066(.A(ori_ori_n888_), .B(ori_ori_n242_), .Y(ori_ori_n1116_));
  NO2        o1067(.A(ori_ori_n622_), .B(x7), .Y(ori_ori_n1117_));
  NA2        o1068(.A(ori_ori_n1117_), .B(ori_ori_n273_), .Y(ori_ori_n1118_));
  NA2        o1069(.A(ori_ori_n702_), .B(ori_ori_n877_), .Y(ori_ori_n1119_));
  AOI210     o1070(.A0(ori_ori_n1118_), .A1(ori_ori_n1116_), .B0(ori_ori_n1119_), .Y(ori_ori_n1120_));
  NOi21      o1071(.An(ori_ori_n401_), .B(ori_ori_n552_), .Y(ori_ori_n1121_));
  NO2        o1072(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n1122_));
  NO2        o1073(.A(ori_ori_n605_), .B(ori_ori_n1122_), .Y(ori_ori_n1123_));
  NO3        o1074(.A(ori_ori_n870_), .B(ori_ori_n108_), .C(ori_ori_n95_), .Y(ori_ori_n1124_));
  AOI210     o1075(.A0(ori_ori_n1123_), .A1(ori_ori_n1019_), .B0(ori_ori_n1124_), .Y(ori_ori_n1125_));
  NA2        o1076(.A(ori_ori_n1060_), .B(ori_ori_n56_), .Y(ori_ori_n1126_));
  OAI220     o1077(.A0(ori_ori_n1126_), .A1(ori_ori_n577_), .B0(ori_ori_n1125_), .B1(ori_ori_n1121_), .Y(ori_ori_n1127_));
  OAI210     o1078(.A0(ori_ori_n1127_), .A1(ori_ori_n1120_), .B0(ori_ori_n581_), .Y(ori_ori_n1128_));
  NA2        o1079(.A(ori_ori_n87_), .B(x5), .Y(ori_ori_n1129_));
  OAI210     o1080(.A0(ori_ori_n1129_), .A1(ori_ori_n320_), .B0(ori_ori_n721_), .Y(ori_ori_n1130_));
  AOI210     o1081(.A0(ori_ori_n829_), .A1(ori_ori_n114_), .B0(ori_ori_n1130_), .Y(ori_ori_n1131_));
  NA2        o1082(.A(ori_ori_n603_), .B(ori_ori_n53_), .Y(ori_ori_n1132_));
  NA2        o1083(.A(ori_ori_n283_), .B(ori_ori_n50_), .Y(ori_ori_n1133_));
  OAI220     o1084(.A0(ori_ori_n1133_), .A1(ori_ori_n306_), .B0(ori_ori_n1132_), .B1(ori_ori_n129_), .Y(ori_ori_n1134_));
  NO2        o1085(.A(ori_ori_n1081_), .B(ori_ori_n512_), .Y(ori_ori_n1135_));
  NO4        o1086(.A(ori_ori_n234_), .B(ori_ori_n265_), .C(ori_ori_n60_), .D(ori_ori_n57_), .Y(ori_ori_n1136_));
  AOI220     o1087(.A0(ori_ori_n1136_), .A1(ori_ori_n1135_), .B0(ori_ori_n1134_), .B1(ori_ori_n56_), .Y(ori_ori_n1137_));
  OAI210     o1088(.A0(ori_ori_n1131_), .A1(ori_ori_n64_), .B0(ori_ori_n1137_), .Y(ori_ori_n1138_));
  NO2        o1089(.A(ori_ori_n57_), .B(x0), .Y(ori_ori_n1139_));
  NO2        o1090(.A(ori_ori_n666_), .B(ori_ori_n317_), .Y(ori_ori_n1140_));
  NO2        o1091(.A(ori_ori_n756_), .B(x3), .Y(ori_ori_n1141_));
  NO2        o1092(.A(ori_ori_n664_), .B(x8), .Y(ori_ori_n1142_));
  AOI220     o1093(.A0(ori_ori_n1142_), .A1(ori_ori_n1141_), .B0(ori_ori_n1140_), .B1(ori_ori_n1139_), .Y(ori_ori_n1143_));
  AOI210     o1094(.A0(ori_ori_n689_), .A1(ori_ori_n242_), .B0(x7), .Y(ori_ori_n1144_));
  NO3        o1095(.A(ori_ori_n1144_), .B(ori_ori_n606_), .C(x8), .Y(ori_ori_n1145_));
  NA4        o1096(.A(ori_ori_n668_), .B(ori_ori_n660_), .C(ori_ori_n199_), .D(x0), .Y(ori_ori_n1146_));
  OAI220     o1097(.A0(ori_ori_n1146_), .A1(ori_ori_n1145_), .B0(ori_ori_n1143_), .B1(ori_ori_n575_), .Y(ori_ori_n1147_));
  AOI210     o1098(.A0(ori_ori_n1138_), .A1(ori_ori_n1026_), .B0(ori_ori_n1147_), .Y(ori_ori_n1148_));
  NO2        o1099(.A(ori_ori_n242_), .B(ori_ori_n55_), .Y(ori_ori_n1149_));
  NO2        o1100(.A(ori_ori_n250_), .B(x8), .Y(ori_ori_n1150_));
  NOi32      o1101(.An(ori_ori_n1150_), .Bn(ori_ori_n198_), .C(ori_ori_n566_), .Y(ori_ori_n1151_));
  NO2        o1102(.A(ori_ori_n88_), .B(ori_ori_n60_), .Y(ori_ori_n1152_));
  OAI210     o1103(.A0(ori_ori_n1151_), .A1(ori_ori_n1149_), .B0(ori_ori_n1152_), .Y(ori_ori_n1153_));
  NO2        o1104(.A(ori_ori_n950_), .B(ori_ori_n96_), .Y(ori_ori_n1154_));
  NO2        o1105(.A(ori_ori_n162_), .B(ori_ori_n53_), .Y(ori_ori_n1155_));
  AOI210     o1106(.A0(ori_ori_n337_), .A1(x8), .B0(ori_ori_n1155_), .Y(ori_ori_n1156_));
  AOI210     o1107(.A0(ori_ori_n211_), .A1(ori_ori_n92_), .B0(ori_ori_n1156_), .Y(ori_ori_n1157_));
  OAI210     o1108(.A0(ori_ori_n1157_), .A1(ori_ori_n1154_), .B0(ori_ori_n677_), .Y(ori_ori_n1158_));
  NO2        o1109(.A(x7), .B(x0), .Y(ori_ori_n1159_));
  NO3        o1110(.A(ori_ori_n153_), .B(ori_ori_n1159_), .C(ori_ori_n140_), .Y(ori_ori_n1160_));
  XN2        o1111(.A(x8), .B(x7), .Y(ori_ori_n1161_));
  NO3        o1112(.A(ori_ori_n1084_), .B(ori_ori_n253_), .C(ori_ori_n1161_), .Y(ori_ori_n1162_));
  OAI210     o1113(.A0(ori_ori_n1162_), .A1(ori_ori_n1160_), .B0(ori_ori_n735_), .Y(ori_ori_n1163_));
  NO2        o1114(.A(ori_ori_n262_), .B(ori_ori_n258_), .Y(ori_ori_n1164_));
  NO2        o1115(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n1165_));
  OAI210     o1116(.A0(ori_ori_n1164_), .A1(ori_ori_n273_), .B0(ori_ori_n1165_), .Y(ori_ori_n1166_));
  NA4        o1117(.A(ori_ori_n1166_), .B(ori_ori_n1163_), .C(ori_ori_n1158_), .D(ori_ori_n1153_), .Y(ori_ori_n1167_));
  NA2        o1118(.A(ori_ori_n1167_), .B(ori_ori_n556_), .Y(ori_ori_n1168_));
  NO2        o1119(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n1169_));
  NA2        o1120(.A(ori_ori_n1169_), .B(ori_ori_n158_), .Y(ori_ori_n1170_));
  NO2        o1121(.A(ori_ori_n670_), .B(ori_ori_n253_), .Y(ori_ori_n1171_));
  OAI210     o1122(.A0(ori_ori_n1171_), .A1(ori_ori_n1029_), .B0(ori_ori_n50_), .Y(ori_ori_n1172_));
  AOI210     o1123(.A0(ori_ori_n1172_), .A1(ori_ori_n1170_), .B0(ori_ori_n429_), .Y(ori_ori_n1173_));
  OAI220     o1124(.A0(ori_ori_n285_), .A1(ori_ori_n271_), .B0(ori_ori_n258_), .B1(ori_ori_n237_), .Y(ori_ori_n1174_));
  NA3        o1125(.A(ori_ori_n1174_), .B(ori_ori_n677_), .C(x1), .Y(ori_ori_n1175_));
  OAI210     o1126(.A0(x8), .A1(x0), .B0(x4), .Y(ori_ori_n1176_));
  NO2        o1127(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n1177_));
  NO2        o1128(.A(ori_ori_n68_), .B(ori_ori_n1177_), .Y(ori_ori_n1178_));
  NOi21      o1129(.An(ori_ori_n1176_), .B(ori_ori_n1178_), .Y(ori_ori_n1179_));
  NO2        o1130(.A(ori_ori_n668_), .B(ori_ori_n320_), .Y(ori_ori_n1180_));
  NO2        o1131(.A(ori_ori_n782_), .B(ori_ori_n215_), .Y(ori_ori_n1181_));
  OAI210     o1132(.A0(ori_ori_n1180_), .A1(ori_ori_n1179_), .B0(ori_ori_n1181_), .Y(ori_ori_n1182_));
  NO2        o1133(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n1183_));
  NO2        o1134(.A(ori_ori_n605_), .B(ori_ori_n443_), .Y(ori_ori_n1184_));
  OAI210     o1135(.A0(ori_ori_n1184_), .A1(ori_ori_n1183_), .B0(ori_ori_n250_), .Y(ori_ori_n1185_));
  NO2        o1136(.A(ori_ori_n825_), .B(ori_ori_n420_), .Y(ori_ori_n1186_));
  NA2        o1137(.A(ori_ori_n325_), .B(ori_ori_n59_), .Y(ori_ori_n1187_));
  NO2        o1138(.A(ori_ori_n1126_), .B(ori_ori_n1187_), .Y(ori_ori_n1188_));
  AOI210     o1139(.A0(ori_ori_n1186_), .A1(ori_ori_n173_), .B0(ori_ori_n1188_), .Y(ori_ori_n1189_));
  NA4        o1140(.A(ori_ori_n1189_), .B(ori_ori_n1185_), .C(ori_ori_n1182_), .D(ori_ori_n1175_), .Y(ori_ori_n1190_));
  OAI210     o1141(.A0(ori_ori_n1190_), .A1(ori_ori_n1173_), .B0(ori_ori_n679_), .Y(ori_ori_n1191_));
  NA4        o1142(.A(ori_ori_n1191_), .B(ori_ori_n1168_), .C(ori_ori_n1148_), .D(ori_ori_n1128_), .Y(ori13));
  NO2        o1143(.A(ori_ori_n462_), .B(ori_ori_n347_), .Y(ori_ori_n1193_));
  NOi41      o1144(.An(ori_ori_n1193_), .B(ori_ori_n677_), .C(ori_ori_n287_), .D(ori_ori_n234_), .Y(ori_ori_n1194_));
  NO2        o1145(.A(ori_ori_n870_), .B(ori_ori_n177_), .Y(ori_ori_n1195_));
  NO2        o1146(.A(ori_ori_n152_), .B(ori_ori_n71_), .Y(ori_ori_n1196_));
  XN2        o1147(.A(x4), .B(x0), .Y(ori_ori_n1197_));
  NO3        o1148(.A(ori_ori_n1197_), .B(ori_ori_n107_), .C(ori_ori_n420_), .Y(ori_ori_n1198_));
  AO220      o1149(.A0(ori_ori_n1198_), .A1(ori_ori_n1196_), .B0(ori_ori_n1195_), .B1(ori_ori_n326_), .Y(ori_ori_n1199_));
  OAI210     o1150(.A0(ori_ori_n1199_), .A1(ori_ori_n1194_), .B0(x3), .Y(ori_ori_n1200_));
  NO2        o1151(.A(ori_ori_n870_), .B(x6), .Y(ori_ori_n1201_));
  NO2        o1152(.A(ori_ori_n1133_), .B(ori_ori_n392_), .Y(ori_ori_n1202_));
  NO3        o1153(.A(x8), .B(x5), .C(ori_ori_n106_), .Y(ori_ori_n1203_));
  NA2        o1154(.A(ori_ori_n1203_), .B(ori_ori_n642_), .Y(ori_ori_n1204_));
  NO2        o1155(.A(ori_ori_n605_), .B(ori_ori_n193_), .Y(ori_ori_n1205_));
  NA2        o1156(.A(ori_ori_n1205_), .B(ori_ori_n1093_), .Y(ori_ori_n1206_));
  NA2        o1157(.A(ori_ori_n447_), .B(ori_ori_n53_), .Y(ori_ori_n1207_));
  NO2        o1158(.A(ori_ori_n1207_), .B(ori_ori_n943_), .Y(ori_ori_n1208_));
  NA2        o1159(.A(ori_ori_n1126_), .B(ori_ori_n467_), .Y(ori_ori_n1209_));
  NA2        o1160(.A(ori_ori_n56_), .B(ori_ori_n106_), .Y(ori_ori_n1210_));
  NA2        o1161(.A(ori_ori_n1210_), .B(x1), .Y(ori_ori_n1211_));
  NO2        o1162(.A(ori_ori_n1211_), .B(ori_ori_n255_), .Y(ori_ori_n1212_));
  NO2        o1163(.A(ori_ori_n317_), .B(x6), .Y(ori_ori_n1213_));
  OAI210     o1164(.A0(ori_ori_n246_), .A1(ori_ori_n984_), .B0(ori_ori_n961_), .Y(ori_ori_n1214_));
  AOI220     o1165(.A0(ori_ori_n1214_), .A1(ori_ori_n1213_), .B0(ori_ori_n1212_), .B1(ori_ori_n1209_), .Y(ori_ori_n1215_));
  NAi41      o1166(.An(ori_ori_n1208_), .B(ori_ori_n1215_), .C(ori_ori_n1206_), .D(ori_ori_n1204_), .Y(ori_ori_n1216_));
  AOI220     o1167(.A0(ori_ori_n1216_), .A1(ori_ori_n68_), .B0(ori_ori_n1202_), .B1(ori_ori_n1201_), .Y(ori_ori_n1217_));
  NA2        o1168(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n1218_));
  NA2        o1169(.A(ori_ori_n1218_), .B(ori_ori_n906_), .Y(ori_ori_n1219_));
  OAI220     o1170(.A0(ori_ori_n299_), .A1(ori_ori_n825_), .B0(ori_ori_n87_), .B1(ori_ori_n77_), .Y(ori_ori_n1220_));
  AOI210     o1171(.A0(ori_ori_n1129_), .A1(ori_ori_n616_), .B0(ori_ori_n984_), .Y(ori_ori_n1221_));
  OA210      o1172(.A0(ori_ori_n1220_), .A1(ori_ori_n1219_), .B0(ori_ori_n1221_), .Y(ori_ori_n1222_));
  NA2        o1173(.A(ori_ori_n618_), .B(ori_ori_n55_), .Y(ori_ori_n1223_));
  NA2        o1174(.A(ori_ori_n505_), .B(ori_ori_n493_), .Y(ori_ori_n1224_));
  NA2        o1175(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n1225_));
  NA2        o1176(.A(ori_ori_n1225_), .B(ori_ori_n539_), .Y(ori_ori_n1226_));
  NO2        o1177(.A(ori_ori_n155_), .B(ori_ori_n124_), .Y(ori_ori_n1227_));
  AOI210     o1178(.A0(ori_ori_n1226_), .A1(ori_ori_n430_), .B0(ori_ori_n1227_), .Y(ori_ori_n1228_));
  OAI220     o1179(.A0(ori_ori_n1228_), .A1(ori_ori_n877_), .B0(ori_ori_n1224_), .B1(ori_ori_n1223_), .Y(ori_ori_n1229_));
  OAI210     o1180(.A0(ori_ori_n1229_), .A1(ori_ori_n1222_), .B0(ori_ori_n1159_), .Y(ori_ori_n1230_));
  NAi21      o1181(.An(ori_ori_n84_), .B(ori_ori_n380_), .Y(ori_ori_n1231_));
  NO2        o1182(.A(ori_ori_n1231_), .B(ori_ori_n71_), .Y(ori_ori_n1232_));
  AOI210     o1183(.A0(ori_ori_n158_), .A1(x4), .B0(ori_ori_n169_), .Y(ori_ori_n1233_));
  NO2        o1184(.A(ori_ori_n1233_), .B(x0), .Y(ori_ori_n1234_));
  NO2        o1185(.A(ori_ori_n166_), .B(ori_ori_n290_), .Y(ori_ori_n1235_));
  OAI210     o1186(.A0(ori_ori_n1235_), .A1(ori_ori_n1234_), .B0(ori_ori_n1232_), .Y(ori_ori_n1236_));
  NA3        o1187(.A(ori_ori_n1165_), .B(ori_ori_n184_), .C(ori_ori_n71_), .Y(ori_ori_n1237_));
  NO2        o1188(.A(x4), .B(x0), .Y(ori_ori_n1238_));
  NO3        o1189(.A(ori_ori_n1004_), .B(ori_ori_n243_), .C(ori_ori_n539_), .Y(ori_ori_n1239_));
  OAI210     o1190(.A0(ori_ori_n1239_), .A1(ori_ori_n194_), .B0(ori_ori_n1238_), .Y(ori_ori_n1240_));
  NA3        o1191(.A(ori_ori_n1240_), .B(ori_ori_n1237_), .C(ori_ori_n1236_), .Y(ori_ori_n1241_));
  NA2        o1192(.A(ori_ori_n245_), .B(ori_ori_n735_), .Y(ori_ori_n1242_));
  NO2        o1193(.A(ori_ori_n1242_), .B(ori_ori_n519_), .Y(ori_ori_n1243_));
  NA2        o1194(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n1244_));
  NO3        o1195(.A(ori_ori_n1244_), .B(ori_ori_n493_), .C(ori_ori_n81_), .Y(ori_ori_n1245_));
  OAI210     o1196(.A0(ori_ori_n1245_), .A1(ori_ori_n1243_), .B0(x2), .Y(ori_ori_n1246_));
  NO2        o1197(.A(ori_ori_n320_), .B(ori_ori_n380_), .Y(ori_ori_n1247_));
  NO2        o1198(.A(ori_ori_n689_), .B(x0), .Y(ori_ori_n1248_));
  OAI210     o1199(.A0(ori_ori_n1248_), .A1(ori_ori_n1247_), .B0(ori_ori_n329_), .Y(ori_ori_n1249_));
  NO2        o1200(.A(ori_ori_n794_), .B(x1), .Y(ori_ori_n1250_));
  AOI220     o1201(.A0(ori_ori_n1250_), .A1(ori_ori_n611_), .B0(ori_ori_n477_), .B1(ori_ori_n291_), .Y(ori_ori_n1251_));
  NA2        o1202(.A(ori_ori_n499_), .B(ori_ori_n50_), .Y(ori_ori_n1252_));
  AOI220     o1203(.A0(ori_ori_n1252_), .A1(ori_ori_n1195_), .B0(ori_ori_n985_), .B1(ori_ori_n97_), .Y(ori_ori_n1253_));
  NA4        o1204(.A(ori_ori_n1253_), .B(ori_ori_n1251_), .C(ori_ori_n1249_), .D(ori_ori_n1246_), .Y(ori_ori_n1254_));
  AOI220     o1205(.A0(ori_ori_n1254_), .A1(ori_ori_n125_), .B0(ori_ori_n1241_), .B1(ori_ori_n67_), .Y(ori_ori_n1255_));
  NA4        o1206(.A(ori_ori_n1255_), .B(ori_ori_n1230_), .C(ori_ori_n1217_), .D(ori_ori_n1200_), .Y(ori14));
  NO2        o1207(.A(ori_ori_n368_), .B(ori_ori_n71_), .Y(ori_ori_n1257_));
  NO3        o1208(.A(x7), .B(x6), .C(x0), .Y(ori_ori_n1258_));
  OAI210     o1209(.A0(ori_ori_n1258_), .A1(ori_ori_n1257_), .B0(x8), .Y(ori_ori_n1259_));
  NA2        o1210(.A(ori_ori_n1142_), .B(ori_ori_n85_), .Y(ori_ori_n1260_));
  AOI210     o1211(.A0(ori_ori_n1260_), .A1(ori_ori_n1259_), .B0(ori_ori_n151_), .Y(ori_ori_n1261_));
  AOI220     o1212(.A0(ori_ori_n372_), .A1(ori_ori_n855_), .B0(ori_ori_n447_), .B1(ori_ori_n420_), .Y(ori_ori_n1262_));
  NA2        o1213(.A(ori_ori_n274_), .B(ori_ori_n980_), .Y(ori_ori_n1263_));
  OAI220     o1214(.A0(ori_ori_n1263_), .A1(ori_ori_n1262_), .B0(ori_ori_n465_), .B1(ori_ori_n809_), .Y(ori_ori_n1264_));
  OA210      o1215(.A0(ori_ori_n1264_), .A1(ori_ori_n1261_), .B0(x4), .Y(ori_ori_n1265_));
  NO2        o1216(.A(ori_ori_n135_), .B(ori_ori_n609_), .Y(ori_ori_n1266_));
  NA2        o1217(.A(x6), .B(x2), .Y(ori_ori_n1267_));
  NO2        o1218(.A(ori_ori_n627_), .B(ori_ori_n1267_), .Y(ori_ori_n1268_));
  OA210      o1219(.A0(ori_ori_n1266_), .A1(ori_ori_n207_), .B0(ori_ori_n1268_), .Y(ori_ori_n1269_));
  NO4        o1220(.A(ori_ori_n605_), .B(ori_ori_n373_), .C(ori_ori_n295_), .D(ori_ori_n112_), .Y(ori_ori_n1270_));
  OAI210     o1221(.A0(ori_ori_n1270_), .A1(ori_ori_n1269_), .B0(ori_ori_n59_), .Y(ori_ori_n1271_));
  NA2        o1222(.A(x6), .B(ori_ori_n104_), .Y(ori_ori_n1272_));
  NO2        o1223(.A(ori_ori_n666_), .B(ori_ori_n1272_), .Y(ori_ori_n1273_));
  NA2        o1224(.A(ori_ori_n1273_), .B(ori_ori_n930_), .Y(ori_ori_n1274_));
  AOI210     o1225(.A0(ori_ori_n1142_), .A1(ori_ori_n1018_), .B0(x1), .Y(ori_ori_n1275_));
  NO2        o1226(.A(ori_ori_n534_), .B(x5), .Y(ori_ori_n1276_));
  NA3        o1227(.A(ori_ori_n1276_), .B(ori_ori_n118_), .C(x0), .Y(ori_ori_n1277_));
  NA4        o1228(.A(ori_ori_n696_), .B(ori_ori_n931_), .C(ori_ori_n299_), .D(ori_ori_n68_), .Y(ori_ori_n1278_));
  AN4        o1229(.A(ori_ori_n1278_), .B(ori_ori_n1277_), .C(ori_ori_n1275_), .D(ori_ori_n1274_), .Y(ori_ori_n1279_));
  NO2        o1230(.A(ori_ori_n703_), .B(ori_ori_n1102_), .Y(ori_ori_n1280_));
  NO2        o1231(.A(ori_ori_n77_), .B(ori_ori_n58_), .Y(ori_ori_n1281_));
  OAI210     o1232(.A0(ori_ori_n1280_), .A1(ori_ori_n444_), .B0(ori_ori_n1281_), .Y(ori_ori_n1282_));
  AO210      o1233(.A0(ori_ori_n1257_), .A1(ori_ori_n1018_), .B0(ori_ori_n53_), .Y(ori_ori_n1283_));
  AOI210     o1234(.A0(ori_ori_n769_), .A1(ori_ori_n819_), .B0(ori_ori_n1283_), .Y(ori_ori_n1284_));
  AOI220     o1235(.A0(ori_ori_n1284_), .A1(ori_ori_n1282_), .B0(ori_ori_n1279_), .B1(ori_ori_n1271_), .Y(ori_ori_n1285_));
  NO2        o1236(.A(ori_ori_n678_), .B(ori_ori_n162_), .Y(ori_ori_n1286_));
  NO3        o1237(.A(ori_ori_n1286_), .B(ori_ori_n1285_), .C(ori_ori_n1265_), .Y(ori_ori_n1287_));
  NO2        o1238(.A(ori_ori_n317_), .B(x2), .Y(ori_ori_n1288_));
  XN2        o1239(.A(x4), .B(x1), .Y(ori_ori_n1289_));
  NO2        o1240(.A(ori_ori_n1289_), .B(ori_ori_n299_), .Y(ori_ori_n1290_));
  NOi21      o1241(.An(ori_ori_n1290_), .B(ori_ori_n408_), .Y(ori_ori_n1291_));
  NO2        o1242(.A(ori_ori_n336_), .B(ori_ori_n60_), .Y(ori_ori_n1292_));
  OAI210     o1243(.A0(ori_ori_n1292_), .A1(ori_ori_n1291_), .B0(ori_ori_n1288_), .Y(ori_ori_n1293_));
  NA2        o1244(.A(ori_ori_n690_), .B(ori_ori_n56_), .Y(ori_ori_n1294_));
  OAI220     o1245(.A0(ori_ori_n1294_), .A1(ori_ori_n152_), .B0(ori_ori_n185_), .B1(ori_ori_n71_), .Y(ori_ori_n1295_));
  NO2        o1246(.A(ori_ori_n211_), .B(ori_ori_n253_), .Y(ori_ori_n1296_));
  AOI220     o1247(.A0(ori_ori_n132_), .A1(ori_ori_n56_), .B0(ori_ori_n91_), .B1(x5), .Y(ori_ori_n1297_));
  NA2        o1248(.A(ori_ori_n1093_), .B(ori_ori_n304_), .Y(ori_ori_n1298_));
  NA2        o1249(.A(ori_ori_n245_), .B(ori_ori_n351_), .Y(ori_ori_n1299_));
  NA2        o1250(.A(ori_ori_n641_), .B(ori_ori_n1036_), .Y(ori_ori_n1300_));
  OAI220     o1251(.A0(ori_ori_n1300_), .A1(ori_ori_n1299_), .B0(ori_ori_n1298_), .B1(ori_ori_n1297_), .Y(ori_ori_n1301_));
  AOI210     o1252(.A0(ori_ori_n1296_), .A1(ori_ori_n1295_), .B0(ori_ori_n1301_), .Y(ori_ori_n1302_));
  AOI210     o1253(.A0(ori_ori_n1302_), .A1(ori_ori_n1293_), .B0(x7), .Y(ori_ori_n1303_));
  NO2        o1254(.A(ori_ori_n492_), .B(x6), .Y(ori_ori_n1304_));
  AOI210     o1255(.A0(ori_ori_n821_), .A1(ori_ori_n963_), .B0(ori_ori_n1304_), .Y(ori_ori_n1305_));
  OAI220     o1256(.A0(ori_ori_n1305_), .A1(ori_ori_n55_), .B0(ori_ori_n492_), .B1(ori_ori_n100_), .Y(ori_ori_n1306_));
  NA2        o1257(.A(ori_ori_n1306_), .B(ori_ori_n353_), .Y(ori_ori_n1307_));
  NA3        o1258(.A(ori_ori_n612_), .B(ori_ori_n1070_), .C(ori_ori_n70_), .Y(ori_ori_n1308_));
  NO4        o1259(.A(ori_ori_n1308_), .B(ori_ori_n1244_), .C(ori_ori_n116_), .D(ori_ori_n55_), .Y(ori_ori_n1309_));
  NO3        o1260(.A(ori_ori_n1063_), .B(ori_ori_n827_), .C(ori_ori_n482_), .Y(ori_ori_n1310_));
  NO3        o1261(.A(ori_ori_n756_), .B(ori_ori_n499_), .C(ori_ori_n54_), .Y(ori_ori_n1311_));
  NO4        o1262(.A(ori_ori_n1311_), .B(ori_ori_n1310_), .C(ori_ori_n1309_), .D(ori_ori_n1041_), .Y(ori_ori_n1312_));
  AOI210     o1263(.A0(ori_ori_n1312_), .A1(ori_ori_n1307_), .B0(ori_ori_n301_), .Y(ori_ori_n1313_));
  NA2        o1264(.A(ori_ori_n904_), .B(ori_ori_n53_), .Y(ori_ori_n1314_));
  OAI210     o1265(.A0(ori_ori_n240_), .A1(ori_ori_n114_), .B0(x2), .Y(ori_ori_n1315_));
  NA2        o1266(.A(ori_ori_n364_), .B(ori_ori_n56_), .Y(ori_ori_n1316_));
  OA220      o1267(.A0(ori_ori_n1316_), .A1(ori_ori_n1315_), .B0(ori_ori_n1314_), .B1(ori_ori_n372_), .Y(ori_ori_n1317_));
  NA2        o1268(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n1318_));
  NO2        o1269(.A(ori_ori_n1318_), .B(ori_ori_n192_), .Y(ori_ori_n1319_));
  NA4        o1270(.A(ori_ori_n1319_), .B(ori_ori_n364_), .C(ori_ori_n253_), .D(ori_ori_n67_), .Y(ori_ori_n1320_));
  OAI210     o1271(.A0(ori_ori_n1317_), .A1(ori_ori_n312_), .B0(ori_ori_n1320_), .Y(ori_ori_n1321_));
  NO3        o1272(.A(ori_ori_n1321_), .B(ori_ori_n1313_), .C(ori_ori_n1303_), .Y(ori_ori_n1322_));
  OAI210     o1273(.A0(ori_ori_n1287_), .A1(x3), .B0(ori_ori_n1322_), .Y(ori15));
  NA2        o1274(.A(ori_ori_n587_), .B(ori_ori_n59_), .Y(ori_ori_n1324_));
  NAi41      o1275(.An(x2), .B(x7), .C(x6), .D(x0), .Y(ori_ori_n1325_));
  AOI210     o1276(.A0(ori_ori_n1325_), .A1(ori_ori_n1324_), .B0(ori_ori_n53_), .Y(ori_ori_n1326_));
  NA3        o1277(.A(ori_ori_n57_), .B(x6), .C(ori_ori_n106_), .Y(ori_ori_n1327_));
  NO2        o1278(.A(ori_ori_n1327_), .B(ori_ori_n290_), .Y(ori_ori_n1328_));
  OAI210     o1279(.A0(ori_ori_n1328_), .A1(ori_ori_n1326_), .B0(ori_ori_n1165_), .Y(ori_ori_n1329_));
  NA2        o1280(.A(ori_ori_n108_), .B(ori_ori_n106_), .Y(ori_ori_n1330_));
  NA4        o1281(.A(ori_ori_n1330_), .B(ori_ori_n639_), .C(ori_ori_n305_), .D(x6), .Y(ori_ori_n1331_));
  AOI210     o1282(.A0(ori_ori_n734_), .A1(ori_ori_n76_), .B0(x3), .Y(ori_ori_n1332_));
  NA3        o1283(.A(ori_ori_n1332_), .B(ori_ori_n1331_), .C(ori_ori_n1329_), .Y(ori_ori_n1333_));
  AOI210     o1284(.A0(ori_ori_n1075_), .A1(ori_ori_n591_), .B0(ori_ori_n50_), .Y(ori_ori_n1334_));
  NO2        o1285(.A(ori_ori_n290_), .B(ori_ori_n106_), .Y(ori_ori_n1335_));
  NO2        o1286(.A(ori_ori_n232_), .B(x5), .Y(ori_ori_n1336_));
  NA2        o1287(.A(ori_ori_n1336_), .B(ori_ori_n1335_), .Y(ori_ori_n1337_));
  NA3        o1288(.A(ori_ori_n1250_), .B(ori_ori_n626_), .C(ori_ori_n1177_), .Y(ori_ori_n1338_));
  NA4        o1289(.A(ori_ori_n1338_), .B(ori_ori_n1337_), .C(ori_ori_n1334_), .D(ori_ori_n1277_), .Y(ori_ori_n1339_));
  NA2        o1290(.A(ori_ori_n330_), .B(ori_ori_n339_), .Y(ori_ori_n1340_));
  AOI210     o1291(.A0(ori_ori_n1211_), .A1(ori_ori_n58_), .B0(ori_ori_n1340_), .Y(ori_ori_n1341_));
  NA4        o1292(.A(ori_ori_n1211_), .B(ori_ori_n702_), .C(ori_ori_n1139_), .D(ori_ori_n380_), .Y(ori_ori_n1342_));
  NA2        o1293(.A(ori_ori_n591_), .B(ori_ori_n466_), .Y(ori_ori_n1343_));
  NO2        o1294(.A(ori_ori_n756_), .B(ori_ori_n53_), .Y(ori_ori_n1344_));
  NO2        o1295(.A(ori_ori_n782_), .B(ori_ori_n295_), .Y(ori_ori_n1345_));
  NA2        o1296(.A(ori_ori_n1345_), .B(ori_ori_n1344_), .Y(ori_ori_n1346_));
  NA3        o1297(.A(ori_ori_n1346_), .B(ori_ori_n1343_), .C(ori_ori_n1342_), .Y(ori_ori_n1347_));
  OAI210     o1298(.A0(ori_ori_n1347_), .A1(ori_ori_n1341_), .B0(ori_ori_n77_), .Y(ori_ori_n1348_));
  NA2        o1299(.A(ori_ori_n366_), .B(ori_ori_n705_), .Y(ori_ori_n1349_));
  NA2        o1300(.A(ori_ori_n572_), .B(ori_ori_n56_), .Y(ori_ori_n1350_));
  NA3        o1301(.A(ori_ori_n1350_), .B(ori_ori_n339_), .C(ori_ori_n108_), .Y(ori_ori_n1351_));
  AOI210     o1302(.A0(ori_ori_n1351_), .A1(ori_ori_n1349_), .B0(ori_ori_n499_), .Y(ori_ori_n1352_));
  NO3        o1303(.A(ori_ori_n807_), .B(ori_ori_n623_), .C(ori_ori_n193_), .Y(ori_ori_n1353_));
  OAI210     o1304(.A0(ori_ori_n1353_), .A1(ori_ori_n1352_), .B0(ori_ori_n492_), .Y(ori_ori_n1354_));
  NO2        o1305(.A(ori_ori_n877_), .B(ori_ori_n50_), .Y(ori_ori_n1355_));
  NO2        o1306(.A(ori_ori_n242_), .B(ori_ori_n64_), .Y(ori_ori_n1356_));
  OA210      o1307(.A0(ori_ori_n1356_), .A1(ori_ori_n1355_), .B0(ori_ori_n408_), .Y(ori_ori_n1357_));
  NA2        o1308(.A(ori_ori_n57_), .B(x3), .Y(ori_ori_n1358_));
  AOI210     o1309(.A0(ori_ori_n986_), .A1(ori_ori_n1358_), .B0(ori_ori_n684_), .Y(ori_ori_n1359_));
  OAI210     o1310(.A0(ori_ori_n1359_), .A1(ori_ori_n1357_), .B0(ori_ori_n1026_), .Y(ori_ori_n1360_));
  NA2        o1311(.A(ori_ori_n1319_), .B(ori_ori_n68_), .Y(ori_ori_n1361_));
  NO2        o1312(.A(ori_ori_n1267_), .B(x0), .Y(ori_ori_n1362_));
  AOI210     o1313(.A0(ori_ori_n1362_), .A1(ori_ori_n606_), .B0(x8), .Y(ori_ori_n1363_));
  NO2        o1314(.A(ori_ori_n429_), .B(ori_ori_n81_), .Y(ori_ori_n1364_));
  NO2        o1315(.A(ori_ori_n937_), .B(ori_ori_n71_), .Y(ori_ori_n1365_));
  NA2        o1316(.A(ori_ori_n1365_), .B(ori_ori_n1364_), .Y(ori_ori_n1366_));
  NO2        o1317(.A(ori_ori_n984_), .B(x6), .Y(ori_ori_n1367_));
  NA4        o1318(.A(ori_ori_n1367_), .B(ori_ori_n596_), .C(ori_ori_n153_), .D(ori_ori_n412_), .Y(ori_ori_n1368_));
  AN4        o1319(.A(ori_ori_n1368_), .B(ori_ori_n1366_), .C(ori_ori_n1363_), .D(ori_ori_n1361_), .Y(ori_ori_n1369_));
  NA4        o1320(.A(ori_ori_n1369_), .B(ori_ori_n1360_), .C(ori_ori_n1354_), .D(ori_ori_n1348_), .Y(ori_ori_n1370_));
  NA2        o1321(.A(ori_ori_n159_), .B(ori_ori_n740_), .Y(ori_ori_n1371_));
  NO2        o1322(.A(ori_ori_n651_), .B(x2), .Y(ori_ori_n1372_));
  OAI210     o1323(.A0(ori_ori_n68_), .A1(ori_ori_n53_), .B0(ori_ori_n138_), .Y(ori_ori_n1373_));
  OAI210     o1324(.A0(ori_ori_n1372_), .A1(ori_ori_n85_), .B0(ori_ori_n1373_), .Y(ori_ori_n1374_));
  AOI210     o1325(.A0(ori_ori_n1374_), .A1(ori_ori_n1371_), .B0(ori_ori_n317_), .Y(ori_ori_n1375_));
  NO3        o1326(.A(ori_ori_n1327_), .B(ori_ori_n261_), .C(ori_ori_n242_), .Y(ori_ori_n1376_));
  NA3        o1327(.A(ori_ori_n57_), .B(x1), .C(x0), .Y(ori_ori_n1377_));
  NA3        o1328(.A(ori_ori_n71_), .B(x5), .C(x2), .Y(ori_ori_n1378_));
  NA4        o1329(.A(x7), .B(x3), .C(ori_ori_n53_), .D(x0), .Y(ori_ori_n1379_));
  OAI220     o1330(.A0(ori_ori_n1379_), .A1(x6), .B0(ori_ori_n1378_), .B1(ori_ori_n1377_), .Y(ori_ori_n1380_));
  NO2        o1331(.A(ori_ori_n1380_), .B(ori_ori_n1376_), .Y(ori_ori_n1381_));
  NAi21      o1332(.An(ori_ori_n112_), .B(ori_ori_n750_), .Y(ori_ori_n1382_));
  NA4        o1333(.A(ori_ori_n1382_), .B(ori_ori_n315_), .C(ori_ori_n285_), .D(ori_ori_n626_), .Y(ori_ori_n1383_));
  OAI220     o1334(.A0(ori_ori_n320_), .A1(x7), .B0(ori_ori_n124_), .B1(ori_ori_n71_), .Y(ori_ori_n1384_));
  NA3        o1335(.A(ori_ori_n1384_), .B(ori_ori_n794_), .C(ori_ori_n1105_), .Y(ori_ori_n1385_));
  NA2        o1336(.A(ori_ori_n82_), .B(ori_ori_n50_), .Y(ori_ori_n1386_));
  AO210      o1337(.A0(ori_ori_n1386_), .A1(ori_ori_n310_), .B0(ori_ori_n151_), .Y(ori_ori_n1387_));
  NA4        o1338(.A(ori_ori_n1387_), .B(ori_ori_n1385_), .C(ori_ori_n1383_), .D(ori_ori_n1381_), .Y(ori_ori_n1388_));
  OAI210     o1339(.A0(ori_ori_n1388_), .A1(ori_ori_n1375_), .B0(ori_ori_n56_), .Y(ori_ori_n1389_));
  AOI210     o1340(.A0(ori_ori_n692_), .A1(x4), .B0(ori_ori_n963_), .Y(ori_ori_n1390_));
  OAI220     o1341(.A0(ori_ori_n1390_), .A1(ori_ori_n296_), .B0(ori_ori_n1030_), .B1(ori_ori_n951_), .Y(ori_ori_n1391_));
  NA2        o1342(.A(ori_ori_n838_), .B(ori_ori_n405_), .Y(ori_ori_n1392_));
  OAI210     o1343(.A0(ori_ori_n1364_), .A1(ori_ori_n1356_), .B0(ori_ori_n286_), .Y(ori_ori_n1393_));
  OAI210     o1344(.A0(ori_ori_n1392_), .A1(ori_ori_n850_), .B0(ori_ori_n1393_), .Y(ori_ori_n1394_));
  OAI210     o1345(.A0(ori_ori_n1394_), .A1(ori_ori_n1391_), .B0(x6), .Y(ori_ori_n1395_));
  NO2        o1346(.A(ori_ori_n57_), .B(ori_ori_n59_), .Y(ori_ori_n1396_));
  NO2        o1347(.A(x7), .B(x5), .Y(ori_ori_n1397_));
  AOI220     o1348(.A0(ori_ori_n859_), .A1(ori_ori_n1396_), .B0(ori_ori_n538_), .B1(ori_ori_n1397_), .Y(ori_ori_n1398_));
  NA2        o1349(.A(ori_ori_n766_), .B(ori_ori_n286_), .Y(ori_ori_n1399_));
  NA3        o1350(.A(ori_ori_n618_), .B(ori_ori_n288_), .C(ori_ori_n237_), .Y(ori_ori_n1400_));
  NA3        o1351(.A(ori_ori_n1400_), .B(ori_ori_n1399_), .C(ori_ori_n1398_), .Y(ori_ori_n1401_));
  NA2        o1352(.A(ori_ori_n1401_), .B(ori_ori_n423_), .Y(ori_ori_n1402_));
  AOI210     o1353(.A0(ori_ori_n376_), .A1(ori_ori_n337_), .B0(ori_ori_n55_), .Y(ori_ori_n1403_));
  NA4        o1354(.A(ori_ori_n1403_), .B(ori_ori_n1402_), .C(ori_ori_n1395_), .D(ori_ori_n1389_), .Y(ori_ori_n1404_));
  AO220      o1355(.A0(ori_ori_n1404_), .A1(ori_ori_n1370_), .B0(ori_ori_n1339_), .B1(ori_ori_n1333_), .Y(ori16));
  NO2        o1356(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n1406_));
  NA2        o1357(.A(ori_ori_n665_), .B(ori_ori_n535_), .Y(ori_ori_n1407_));
  NA3        o1358(.A(ori_ori_n226_), .B(ori_ori_n430_), .C(ori_ori_n963_), .Y(ori_ori_n1408_));
  NA2        o1359(.A(ori_ori_n127_), .B(ori_ori_n202_), .Y(ori_ori_n1409_));
  AOI210     o1360(.A0(ori_ori_n1408_), .A1(ori_ori_n1407_), .B0(ori_ori_n1409_), .Y(ori_ori_n1410_));
  NO3        o1361(.A(x8), .B(x6), .C(ori_ori_n50_), .Y(ori_ori_n1411_));
  NO2        o1362(.A(ori_ori_n738_), .B(ori_ori_n180_), .Y(ori_ori_n1412_));
  OAI210     o1363(.A0(ori_ori_n1411_), .A1(ori_ori_n234_), .B0(ori_ori_n1412_), .Y(ori_ori_n1413_));
  NO2        o1364(.A(ori_ori_n155_), .B(x5), .Y(ori_ori_n1414_));
  NA2        o1365(.A(ori_ori_n1414_), .B(ori_ori_n1372_), .Y(ori_ori_n1415_));
  NA3        o1366(.A(ori_ori_n581_), .B(ori_ori_n537_), .C(ori_ori_n476_), .Y(ori_ori_n1416_));
  NA3        o1367(.A(ori_ori_n1416_), .B(ori_ori_n1415_), .C(ori_ori_n1413_), .Y(ori_ori_n1417_));
  OAI210     o1368(.A0(ori_ori_n1417_), .A1(ori_ori_n1410_), .B0(ori_ori_n1406_), .Y(ori_ori_n1418_));
  OAI210     o1369(.A0(ori_ori_n1288_), .A1(ori_ori_n930_), .B0(ori_ori_n420_), .Y(ori_ori_n1419_));
  NO2        o1370(.A(ori_ori_n317_), .B(x7), .Y(ori_ori_n1420_));
  NO2        o1371(.A(ori_ori_n1419_), .B(ori_ori_n640_), .Y(ori_ori_n1421_));
  NA2        o1372(.A(ori_ori_n1084_), .B(ori_ori_n193_), .Y(ori_ori_n1422_));
  NA2        o1373(.A(ori_ori_n55_), .B(ori_ori_n104_), .Y(ori_ori_n1423_));
  NA2        o1374(.A(ori_ori_n1423_), .B(ori_ori_n686_), .Y(ori_ori_n1424_));
  NA2        o1375(.A(ori_ori_n375_), .B(ori_ori_n1088_), .Y(ori_ori_n1425_));
  OA220      o1376(.A0(ori_ori_n1425_), .A1(ori_ori_n1424_), .B0(ori_ori_n1422_), .B1(ori_ori_n634_), .Y(ori_ori_n1426_));
  OAI210     o1377(.A0(ori_ori_n1426_), .A1(ori_ori_n655_), .B0(ori_ori_n497_), .Y(ori_ori_n1427_));
  INV        o1378(.A(ori_ori_n1026_), .Y(ori_ori_n1428_));
  NO2        o1379(.A(ori_ori_n1428_), .B(ori_ori_n62_), .Y(ori_ori_n1429_));
  AOI220     o1380(.A0(ori_ori_n1429_), .A1(ori_ori_n265_), .B0(ori_ori_n1273_), .B1(ori_ori_n122_), .Y(ori_ori_n1430_));
  AOI220     o1381(.A0(ori_ori_n639_), .A1(ori_ori_n360_), .B0(ori_ori_n626_), .B1(ori_ori_n88_), .Y(ori_ori_n1431_));
  NA3        o1382(.A(ori_ori_n463_), .B(ori_ori_n588_), .C(ori_ori_n187_), .Y(ori_ori_n1432_));
  OAI220     o1383(.A0(ori_ori_n1432_), .A1(ori_ori_n1431_), .B0(ori_ori_n1430_), .B1(ori_ori_n306_), .Y(ori_ori_n1433_));
  NO3        o1384(.A(ori_ori_n1433_), .B(ori_ori_n1427_), .C(ori_ori_n1421_), .Y(ori_ori_n1434_));
  NO3        o1385(.A(x6), .B(x4), .C(x3), .Y(ori_ori_n1435_));
  NA2        o1386(.A(ori_ori_n1435_), .B(ori_ori_n534_), .Y(ori_ori_n1436_));
  NA4        o1387(.A(ori_ori_n710_), .B(ori_ori_n180_), .C(ori_ori_n58_), .D(x6), .Y(ori_ori_n1437_));
  AOI210     o1388(.A0(ori_ori_n1437_), .A1(ori_ori_n1436_), .B0(ori_ori_n54_), .Y(ori_ori_n1438_));
  NO2        o1389(.A(ori_ori_n726_), .B(x3), .Y(ori_ori_n1439_));
  AOI210     o1390(.A0(ori_ori_n664_), .A1(ori_ori_n142_), .B0(ori_ori_n1070_), .Y(ori_ori_n1440_));
  OA210      o1391(.A0(ori_ori_n1439_), .A1(ori_ori_n423_), .B0(ori_ori_n1440_), .Y(ori_ori_n1441_));
  NO3        o1392(.A(ori_ori_n499_), .B(ori_ori_n215_), .C(ori_ori_n75_), .Y(ori_ori_n1442_));
  NO2        o1393(.A(ori_ori_n766_), .B(ori_ori_n511_), .Y(ori_ori_n1443_));
  NO3        o1394(.A(ori_ori_n1443_), .B(ori_ori_n255_), .C(ori_ori_n150_), .Y(ori_ori_n1444_));
  NO4        o1395(.A(ori_ori_n1444_), .B(ori_ori_n1442_), .C(ori_ori_n1441_), .D(ori_ori_n1438_), .Y(ori_ori_n1445_));
  NA2        o1396(.A(ori_ori_n406_), .B(ori_ori_n963_), .Y(ori_ori_n1446_));
  NA4        o1397(.A(ori_ori_n482_), .B(ori_ori_n368_), .C(ori_ori_n217_), .D(x6), .Y(ori_ori_n1447_));
  OAI210     o1398(.A0(ori_ori_n726_), .A1(ori_ori_n1446_), .B0(ori_ori_n1447_), .Y(ori_ori_n1448_));
  NA2        o1399(.A(ori_ori_n912_), .B(ori_ori_n1318_), .Y(ori_ori_n1449_));
  NA2        o1400(.A(ori_ori_n735_), .B(x7), .Y(ori_ori_n1450_));
  OAI210     o1401(.A0(ori_ori_n1450_), .A1(ori_ori_n387_), .B0(ori_ori_n1449_), .Y(ori_ori_n1451_));
  NA2        o1402(.A(ori_ori_n272_), .B(x2), .Y(ori_ori_n1452_));
  NO3        o1403(.A(ori_ori_n1452_), .B(ori_ori_n596_), .C(ori_ori_n72_), .Y(ori_ori_n1453_));
  OA210      o1404(.A0(ori_ori_n1272_), .A1(ori_ori_n58_), .B0(ori_ori_n783_), .Y(ori_ori_n1454_));
  AOI210     o1405(.A0(ori_ori_n581_), .A1(ori_ori_n50_), .B0(ori_ori_n591_), .Y(ori_ori_n1455_));
  OAI210     o1406(.A0(ori_ori_n931_), .A1(ori_ori_n950_), .B0(ori_ori_n382_), .Y(ori_ori_n1456_));
  OAI220     o1407(.A0(ori_ori_n1456_), .A1(ori_ori_n1455_), .B0(ori_ori_n1454_), .B1(ori_ori_n185_), .Y(ori_ori_n1457_));
  NO4        o1408(.A(ori_ori_n1457_), .B(ori_ori_n1453_), .C(ori_ori_n1451_), .D(ori_ori_n1448_), .Y(ori_ori_n1458_));
  OA220      o1409(.A0(ori_ori_n1458_), .A1(ori_ori_n443_), .B0(ori_ori_n1445_), .B1(ori_ori_n200_), .Y(ori_ori_n1459_));
  NO2        o1410(.A(ori_ori_n926_), .B(ori_ori_n55_), .Y(ori_ori_n1460_));
  NA2        o1411(.A(ori_ori_n417_), .B(ori_ori_n809_), .Y(ori_ori_n1461_));
  NO2        o1412(.A(ori_ori_n1461_), .B(ori_ori_n1460_), .Y(ori_ori_n1462_));
  NO3        o1413(.A(ori_ori_n964_), .B(ori_ori_n330_), .C(x8), .Y(ori_ori_n1463_));
  OAI210     o1414(.A0(ori_ori_n1463_), .A1(ori_ori_n1462_), .B0(x6), .Y(ori_ori_n1464_));
  NO2        o1415(.A(ori_ori_n1100_), .B(ori_ori_n1062_), .Y(ori_ori_n1465_));
  NA2        o1416(.A(ori_ori_n185_), .B(x7), .Y(ori_ori_n1466_));
  OAI220     o1417(.A0(ori_ori_n1466_), .A1(ori_ori_n1465_), .B0(ori_ori_n768_), .B1(ori_ori_n87_), .Y(ori_ori_n1467_));
  NA2        o1418(.A(ori_ori_n1467_), .B(ori_ori_n931_), .Y(ori_ori_n1468_));
  NA2        o1419(.A(ori_ori_n879_), .B(ori_ori_n71_), .Y(ori_ori_n1469_));
  INV        o1420(.A(ori_ori_n1015_), .Y(ori_ori_n1470_));
  AOI210     o1421(.A0(ori_ori_n499_), .A1(ori_ori_n57_), .B0(ori_ori_n634_), .Y(ori_ori_n1471_));
  NA3        o1422(.A(ori_ori_n223_), .B(ori_ori_n76_), .C(ori_ori_n71_), .Y(ori_ori_n1472_));
  OAI210     o1423(.A0(ori_ori_n922_), .A1(ori_ori_n226_), .B0(ori_ori_n1472_), .Y(ori_ori_n1473_));
  AOI210     o1424(.A0(ori_ori_n1471_), .A1(ori_ori_n1470_), .B0(ori_ori_n1473_), .Y(ori_ori_n1474_));
  NA3        o1425(.A(ori_ori_n1474_), .B(ori_ori_n1468_), .C(ori_ori_n1464_), .Y(ori_ori_n1475_));
  NO2        o1426(.A(ori_ori_n641_), .B(x6), .Y(ori_ori_n1476_));
  OAI210     o1427(.A0(ori_ori_n382_), .A1(ori_ori_n84_), .B0(ori_ori_n380_), .Y(ori_ori_n1477_));
  OA210      o1428(.A0(ori_ori_n1477_), .A1(ori_ori_n1476_), .B0(ori_ori_n125_), .Y(ori_ori_n1478_));
  NO3        o1429(.A(ori_ori_n445_), .B(ori_ori_n385_), .C(x7), .Y(ori_ori_n1479_));
  NO3        o1430(.A(ori_ori_n155_), .B(ori_ori_n75_), .C(x2), .Y(ori_ori_n1480_));
  NO3        o1431(.A(ori_ori_n1480_), .B(ori_ori_n1479_), .C(ori_ori_n1478_), .Y(ori_ori_n1481_));
  NO2        o1432(.A(ori_ori_n226_), .B(x1), .Y(ori_ori_n1482_));
  OAI210     o1433(.A0(ori_ori_n1482_), .A1(ori_ori_n450_), .B0(ori_ori_n511_), .Y(ori_ori_n1483_));
  NO2        o1434(.A(ori_ori_n57_), .B(ori_ori_n104_), .Y(ori_ori_n1484_));
  NA2        o1435(.A(ori_ori_n1093_), .B(ori_ori_n1484_), .Y(ori_ori_n1485_));
  AOI210     o1436(.A0(ori_ori_n1485_), .A1(ori_ori_n1483_), .B0(ori_ori_n56_), .Y(ori_ori_n1486_));
  AOI220     o1437(.A0(ori_ori_n768_), .A1(ori_ori_n779_), .B0(ori_ori_n514_), .B1(ori_ori_n276_), .Y(ori_ori_n1487_));
  NO2        o1438(.A(ori_ori_n1487_), .B(ori_ori_n1318_), .Y(ori_ori_n1488_));
  NO3        o1439(.A(ori_ori_n534_), .B(ori_ori_n168_), .C(ori_ori_n1062_), .Y(ori_ori_n1489_));
  NA2        o1440(.A(ori_ori_n950_), .B(x4), .Y(ori_ori_n1490_));
  OAI220     o1441(.A0(ori_ori_n1490_), .A1(ori_ori_n691_), .B0(ori_ori_n649_), .B1(ori_ori_n612_), .Y(ori_ori_n1491_));
  NO4        o1442(.A(ori_ori_n1491_), .B(ori_ori_n1489_), .C(ori_ori_n1488_), .D(ori_ori_n1486_), .Y(ori_ori_n1492_));
  OAI210     o1443(.A0(ori_ori_n1481_), .A1(x5), .B0(ori_ori_n1492_), .Y(ori_ori_n1493_));
  AOI220     o1444(.A0(ori_ori_n1493_), .A1(ori_ori_n95_), .B0(ori_ori_n1475_), .B1(ori_ori_n337_), .Y(ori_ori_n1494_));
  NA4        o1445(.A(ori_ori_n1494_), .B(ori_ori_n1459_), .C(ori_ori_n1434_), .D(ori_ori_n1418_), .Y(ori17));
  NO4        o1446(.A(ori_ori_n603_), .B(ori_ori_n704_), .C(ori_ori_n98_), .D(ori_ori_n97_), .Y(ori_ori_n1496_));
  NO2        o1447(.A(ori_ori_n121_), .B(ori_ori_n1177_), .Y(ori_ori_n1497_));
  AOI220     o1448(.A0(ori_ori_n1497_), .A1(ori_ori_n720_), .B0(ori_ori_n1496_), .B1(ori_ori_n505_), .Y(ori_ori_n1498_));
  NA2        o1449(.A(ori_ori_n159_), .B(ori_ori_n78_), .Y(ori_ori_n1499_));
  NOi21      o1450(.An(ori_ori_n380_), .B(ori_ori_n84_), .Y(ori_ori_n1500_));
  OAI210     o1451(.A0(ori_ori_n626_), .A1(ori_ori_n55_), .B0(ori_ori_n1500_), .Y(ori_ori_n1501_));
  NA2        o1452(.A(ori_ori_n1231_), .B(ori_ori_n1021_), .Y(ori_ori_n1502_));
  NA4        o1453(.A(ori_ori_n1502_), .B(ori_ori_n1501_), .C(ori_ori_n738_), .D(ori_ori_n57_), .Y(ori_ori_n1503_));
  OAI210     o1454(.A0(ori_ori_n710_), .A1(x8), .B0(ori_ori_n1318_), .Y(ori_ori_n1504_));
  NA3        o1455(.A(ori_ori_n1504_), .B(ori_ori_n1257_), .C(ori_ori_n399_), .Y(ori_ori_n1505_));
  NA3        o1456(.A(ori_ori_n393_), .B(ori_ori_n265_), .C(ori_ori_n587_), .Y(ori_ori_n1506_));
  OA210      o1457(.A0(ori_ori_n1327_), .A1(ori_ori_n1170_), .B0(ori_ori_n758_), .Y(ori_ori_n1507_));
  NA4        o1458(.A(ori_ori_n1507_), .B(ori_ori_n1506_), .C(ori_ori_n1505_), .D(ori_ori_n1503_), .Y(ori_ori_n1508_));
  NA3        o1459(.A(ori_ori_n158_), .B(ori_ori_n632_), .C(ori_ori_n1062_), .Y(ori_ori_n1509_));
  AOI210     o1460(.A0(ori_ori_n1090_), .A1(ori_ori_n302_), .B0(ori_ori_n59_), .Y(ori_ori_n1510_));
  NA2        o1461(.A(ori_ori_n1510_), .B(ori_ori_n1509_), .Y(ori_ori_n1511_));
  AOI210     o1462(.A0(ori_ori_n1508_), .A1(x1), .B0(ori_ori_n1511_), .Y(ori_ori_n1512_));
  NO2        o1463(.A(ori_ori_n989_), .B(ori_ori_n499_), .Y(ori_ori_n1513_));
  OAI210     o1464(.A0(ori_ori_n1513_), .A1(ori_ori_n1074_), .B0(ori_ori_n609_), .Y(ori_ori_n1514_));
  NO3        o1465(.A(ori_ori_n634_), .B(ori_ori_n556_), .C(ori_ori_n525_), .Y(ori_ori_n1515_));
  OAI210     o1466(.A0(ori_ori_n1515_), .A1(ori_ori_n911_), .B0(ori_ori_n1439_), .Y(ori_ori_n1516_));
  AOI210     o1467(.A0(ori_ori_n1516_), .A1(ori_ori_n1514_), .B0(x8), .Y(ori_ori_n1517_));
  NA3        o1468(.A(ori_ori_n634_), .B(ori_ori_n268_), .C(ori_ori_n118_), .Y(ori_ori_n1518_));
  NO2        o1469(.A(ori_ori_n138_), .B(ori_ori_n136_), .Y(ori_ori_n1519_));
  NO3        o1470(.A(ori_ori_n907_), .B(ori_ori_n779_), .C(ori_ori_n704_), .Y(ori_ori_n1520_));
  AOI210     o1471(.A0(ori_ori_n1520_), .A1(ori_ori_n1519_), .B0(x0), .Y(ori_ori_n1521_));
  OAI210     o1472(.A0(ori_ori_n1518_), .A1(ori_ori_n244_), .B0(ori_ori_n1521_), .Y(ori_ori_n1522_));
  NO2        o1473(.A(ori_ori_n1522_), .B(ori_ori_n1517_), .Y(ori_ori_n1523_));
  OAI220     o1474(.A0(ori_ori_n1523_), .A1(ori_ori_n1512_), .B0(ori_ori_n1499_), .B1(ori_ori_n1498_), .Y(ori18));
  AOI210     o1475(.A0(x8), .A1(x0), .B0(x5), .Y(ori_ori_n1525_));
  NOi31      o1476(.An(ori_ori_n302_), .B(ori_ori_n1525_), .C(ori_ori_n1060_), .Y(ori_ori_n1526_));
  NA2        o1477(.A(ori_ori_n603_), .B(ori_ori_n59_), .Y(ori_ori_n1527_));
  AOI210     o1478(.A0(ori_ori_n1422_), .A1(ori_ori_n348_), .B0(ori_ori_n1527_), .Y(ori_ori_n1528_));
  NO2        o1479(.A(ori_ori_n619_), .B(ori_ori_n780_), .Y(ori_ori_n1529_));
  NO4        o1480(.A(ori_ori_n251_), .B(ori_ori_n819_), .C(ori_ori_n149_), .D(ori_ori_n70_), .Y(ori_ori_n1530_));
  NO4        o1481(.A(ori_ori_n1530_), .B(ori_ori_n1529_), .C(ori_ori_n1528_), .D(ori_ori_n1526_), .Y(ori_ori_n1531_));
  NA3        o1482(.A(ori_ori_n520_), .B(ori_ori_n211_), .C(x0), .Y(ori_ori_n1532_));
  NAi21      o1483(.An(ori_ori_n386_), .B(ori_ori_n1532_), .Y(ori_ori_n1533_));
  NO2        o1484(.A(ori_ori_n897_), .B(x5), .Y(ori_ori_n1534_));
  AOI210     o1485(.A0(ori_ori_n1155_), .A1(x5), .B0(ori_ori_n1534_), .Y(ori_ori_n1535_));
  OA220      o1486(.A0(ori_ori_n520_), .A1(ori_ori_n330_), .B0(ori_ori_n399_), .B1(x5), .Y(ori_ori_n1536_));
  OAI220     o1487(.A0(ori_ori_n1536_), .A1(ori_ori_n290_), .B0(ori_ori_n1535_), .B1(ori_ori_n209_), .Y(ori_ori_n1537_));
  AOI210     o1488(.A0(ori_ori_n1533_), .A1(ori_ori_n288_), .B0(ori_ori_n1537_), .Y(ori_ori_n1538_));
  AOI210     o1489(.A0(ori_ori_n1538_), .A1(ori_ori_n1531_), .B0(x6), .Y(ori_ori_n1539_));
  NA3        o1490(.A(ori_ori_n524_), .B(ori_ori_n420_), .C(x2), .Y(ori_ori_n1540_));
  NA3        o1491(.A(ori_ori_n1060_), .B(ori_ori_n51_), .C(ori_ori_n57_), .Y(ori_ori_n1541_));
  AOI210     o1492(.A0(ori_ori_n1541_), .A1(ori_ori_n1540_), .B0(ori_ori_n794_), .Y(ori_ori_n1542_));
  AOI210     o1493(.A0(ori_ori_n424_), .A1(ori_ori_n132_), .B0(ori_ori_n792_), .Y(ori_ori_n1543_));
  NA2        o1494(.A(ori_ori_n265_), .B(x6), .Y(ori_ori_n1544_));
  OAI210     o1495(.A0(ori_ori_n173_), .A1(ori_ori_n106_), .B0(ori_ori_n1161_), .Y(ori_ori_n1545_));
  OAI220     o1496(.A0(ori_ori_n1545_), .A1(ori_ori_n1544_), .B0(ori_ori_n1543_), .B1(ori_ori_n750_), .Y(ori_ori_n1546_));
  OAI210     o1497(.A0(ori_ori_n1546_), .A1(ori_ori_n1542_), .B0(ori_ori_n53_), .Y(ori_ori_n1547_));
  NO2        o1498(.A(ori_ori_n690_), .B(ori_ori_n258_), .Y(ori_ori_n1548_));
  NO2        o1499(.A(ori_ori_n261_), .B(x3), .Y(ori_ori_n1549_));
  NO3        o1500(.A(ori_ori_n434_), .B(ori_ori_n603_), .C(ori_ori_n843_), .Y(ori_ori_n1550_));
  OAI210     o1501(.A0(ori_ori_n1550_), .A1(ori_ori_n1548_), .B0(ori_ori_n1549_), .Y(ori_ori_n1551_));
  AOI210     o1502(.A0(ori_ori_n1164_), .A1(ori_ori_n618_), .B0(x4), .Y(ori_ori_n1552_));
  OAI210     o1503(.A0(ori_ori_n556_), .A1(ori_ori_n603_), .B0(ori_ori_n59_), .Y(ori_ori_n1553_));
  OAI210     o1504(.A0(ori_ori_n626_), .A1(ori_ori_n651_), .B0(ori_ori_n1553_), .Y(ori_ori_n1554_));
  AO220      o1505(.A0(ori_ori_n1276_), .A1(ori_ori_n738_), .B0(ori_ori_n557_), .B1(ori_ori_n353_), .Y(ori_ori_n1555_));
  AOI220     o1506(.A0(ori_ori_n1555_), .A1(x1), .B0(ori_ori_n1554_), .B1(ori_ori_n156_), .Y(ori_ori_n1556_));
  NA4        o1507(.A(ori_ori_n1556_), .B(ori_ori_n1552_), .C(ori_ori_n1551_), .D(ori_ori_n1547_), .Y(ori_ori_n1557_));
  NO3        o1508(.A(ori_ori_n1081_), .B(ori_ori_n125_), .C(ori_ori_n124_), .Y(ori_ori_n1558_));
  OAI210     o1509(.A0(ori_ori_n1558_), .A1(ori_ori_n656_), .B0(ori_ori_n104_), .Y(ori_ori_n1559_));
  AOI210     o1510(.A0(ori_ori_n1559_), .A1(ori_ori_n562_), .B0(ori_ori_n794_), .Y(ori_ori_n1560_));
  NA3        o1511(.A(ori_ori_n1223_), .B(ori_ori_n185_), .C(ori_ori_n135_), .Y(ori_ori_n1561_));
  NA3        o1512(.A(ori_ori_n1084_), .B(ori_ori_n782_), .C(ori_ori_n341_), .Y(ori_ori_n1562_));
  NA2        o1513(.A(ori_ori_n166_), .B(ori_ori_n779_), .Y(ori_ori_n1563_));
  OAI210     o1514(.A0(ori_ori_n1563_), .A1(ori_ori_n1330_), .B0(ori_ori_n1562_), .Y(ori_ori_n1564_));
  AOI210     o1515(.A0(ori_ori_n1561_), .A1(ori_ori_n172_), .B0(ori_ori_n1564_), .Y(ori_ori_n1565_));
  OAI210     o1516(.A0(ori_ori_n1565_), .A1(ori_ori_n543_), .B0(x4), .Y(ori_ori_n1566_));
  OAI220     o1517(.A0(ori_ori_n1566_), .A1(ori_ori_n1560_), .B0(ori_ori_n1557_), .B1(ori_ori_n1539_), .Y(ori_ori_n1567_));
  NO2        o1518(.A(ori_ori_n141_), .B(ori_ori_n119_), .Y(ori_ori_n1568_));
  NO2        o1519(.A(ori_ori_n185_), .B(ori_ori_n809_), .Y(ori_ori_n1569_));
  AOI210     o1520(.A0(ori_ori_n604_), .A1(ori_ori_n511_), .B0(ori_ori_n1569_), .Y(ori_ori_n1570_));
  NO2        o1521(.A(ori_ori_n1570_), .B(x6), .Y(ori_ori_n1571_));
  NO2        o1522(.A(ori_ori_n385_), .B(ori_ori_n250_), .Y(ori_ori_n1572_));
  NO2        o1523(.A(ori_ori_n125_), .B(ori_ori_n740_), .Y(ori_ori_n1573_));
  NO2        o1524(.A(ori_ori_n964_), .B(ori_ori_n587_), .Y(ori_ori_n1574_));
  AO220      o1525(.A0(ori_ori_n1574_), .A1(ori_ori_n1573_), .B0(ori_ori_n1572_), .B1(ori_ori_n121_), .Y(ori_ori_n1575_));
  NO3        o1526(.A(ori_ori_n1575_), .B(ori_ori_n1571_), .C(ori_ori_n1568_), .Y(ori_ori_n1576_));
  NA2        o1527(.A(ori_ori_n1081_), .B(x3), .Y(ori_ori_n1577_));
  NA2        o1528(.A(ori_ori_n1367_), .B(ori_ori_n127_), .Y(ori_ori_n1578_));
  OAI220     o1529(.A0(ori_ori_n1578_), .A1(ori_ori_n1577_), .B0(ori_ori_n1576_), .B1(x3), .Y(ori_ori_n1579_));
  NO3        o1530(.A(ori_ori_n1011_), .B(ori_ori_n690_), .C(ori_ori_n325_), .Y(ori_ori_n1580_));
  AO210      o1531(.A0(ori_ori_n1040_), .A1(ori_ori_n295_), .B0(ori_ori_n1580_), .Y(ori_ori_n1581_));
  AOI220     o1532(.A0(ori_ori_n1581_), .A1(x8), .B0(ori_ori_n1367_), .B1(ori_ori_n435_), .Y(ori_ori_n1582_));
  NA2        o1533(.A(ori_ori_n754_), .B(ori_ori_n316_), .Y(ori_ori_n1583_));
  NO4        o1534(.A(ori_ori_n366_), .B(ori_ori_n198_), .C(ori_ori_n336_), .D(x2), .Y(ori_ori_n1584_));
  NA2        o1535(.A(ori_ori_n1423_), .B(ori_ori_n106_), .Y(ori_ori_n1585_));
  NO3        o1536(.A(ori_ori_n1225_), .B(ori_ori_n1004_), .C(ori_ori_n1161_), .Y(ori_ori_n1586_));
  AOI210     o1537(.A0(ori_ori_n1586_), .A1(ori_ori_n1585_), .B0(ori_ori_n1584_), .Y(ori_ori_n1587_));
  OA220      o1538(.A0(ori_ori_n1587_), .A1(ori_ori_n964_), .B0(ori_ori_n1583_), .B1(ori_ori_n571_), .Y(ori_ori_n1588_));
  OAI210     o1539(.A0(ori_ori_n1582_), .A1(ori_ori_n409_), .B0(ori_ori_n1588_), .Y(ori_ori_n1589_));
  AOI210     o1540(.A0(ori_ori_n1579_), .A1(ori_ori_n132_), .B0(ori_ori_n1589_), .Y(ori_ori_n1590_));
  NA2        o1541(.A(ori_ori_n1590_), .B(ori_ori_n1567_), .Y(ori19));
  NO2        o1542(.A(ori_ori_n1469_), .B(ori_ori_n254_), .Y(ori_ori_n1592_));
  NA2        o1543(.A(ori_ori_n651_), .B(x3), .Y(ori_ori_n1593_));
  OAI210     o1544(.A0(ori_ori_n149_), .A1(ori_ori_n105_), .B0(ori_ori_n81_), .Y(ori_ori_n1594_));
  NA3        o1545(.A(ori_ori_n1594_), .B(ori_ori_n1593_), .C(ori_ori_n237_), .Y(ori_ori_n1595_));
  NO2        o1546(.A(ori_ori_n1325_), .B(ori_ori_n166_), .Y(ori_ori_n1596_));
  AOI210     o1547(.A0(ori_ori_n1496_), .A1(ori_ori_n351_), .B0(ori_ori_n1596_), .Y(ori_ori_n1597_));
  AOI210     o1548(.A0(ori_ori_n1597_), .A1(ori_ori_n1595_), .B0(ori_ori_n56_), .Y(ori_ori_n1598_));
  NO2        o1549(.A(ori_ori_n868_), .B(ori_ori_n1238_), .Y(ori_ori_n1599_));
  OAI210     o1550(.A0(ori_ori_n1598_), .A1(ori_ori_n1592_), .B0(ori_ori_n1599_), .Y(ori_ori_n1600_));
  NOi21      o1551(.An(ori_ori_n613_), .B(ori_ori_n655_), .Y(ori_ori_n1601_));
  AOI210     o1552(.A0(ori_ori_n351_), .A1(x6), .B0(ori_ori_n118_), .Y(ori_ori_n1602_));
  NO3        o1553(.A(ori_ori_n1602_), .B(ori_ori_n763_), .C(ori_ori_n122_), .Y(ori_ori_n1603_));
  NA2        o1554(.A(ori_ori_n1218_), .B(ori_ori_n119_), .Y(ori_ori_n1604_));
  NO4        o1555(.A(ori_ori_n1604_), .B(ori_ori_n1011_), .C(ori_ori_n897_), .D(ori_ori_n77_), .Y(ori_ori_n1605_));
  NO3        o1556(.A(ori_ori_n1605_), .B(ori_ori_n1603_), .C(ori_ori_n1037_), .Y(ori_ori_n1606_));
  NO2        o1557(.A(ori_ori_n543_), .B(ori_ori_n622_), .Y(ori_ori_n1607_));
  NA2        o1558(.A(ori_ori_n1272_), .B(ori_ori_n50_), .Y(ori_ori_n1608_));
  NO3        o1559(.A(ori_ori_n518_), .B(ori_ori_n304_), .C(ori_ori_n64_), .Y(ori_ori_n1609_));
  AOI220     o1560(.A0(ori_ori_n1609_), .A1(ori_ori_n1608_), .B0(ori_ori_n1607_), .B1(ori_ori_n782_), .Y(ori_ori_n1610_));
  OAI210     o1561(.A0(ori_ori_n1606_), .A1(ori_ori_n57_), .B0(ori_ori_n1610_), .Y(ori_ori_n1611_));
  AOI210     o1562(.A0(ori_ori_n1611_), .A1(ori_ori_n779_), .B0(ori_ori_n1601_), .Y(ori_ori_n1612_));
  AOI210     o1563(.A0(ori_ori_n829_), .A1(ori_ori_n740_), .B0(ori_ori_n769_), .Y(ori_ori_n1613_));
  NO2        o1564(.A(ori_ori_n1613_), .B(x4), .Y(ori_ori_n1614_));
  NA3        o1565(.A(ori_ori_n738_), .B(ori_ori_n253_), .C(x7), .Y(ori_ori_n1615_));
  AOI220     o1566(.A0(ori_ori_n1420_), .A1(ori_ori_n794_), .B0(ori_ori_n704_), .B1(ori_ori_n1177_), .Y(ori_ori_n1616_));
  AOI210     o1567(.A0(ori_ori_n1616_), .A1(ori_ori_n1615_), .B0(ori_ori_n503_), .Y(ori_ori_n1617_));
  OAI210     o1568(.A0(ori_ori_n1617_), .A1(ori_ori_n1614_), .B0(ori_ori_n819_), .Y(ori_ori_n1618_));
  NO2        o1569(.A(ori_ori_n750_), .B(ori_ori_n320_), .Y(ori_ori_n1619_));
  NO2        o1570(.A(ori_ori_n149_), .B(ori_ori_n1036_), .Y(ori_ori_n1620_));
  AOI220     o1571(.A0(ori_ori_n1620_), .A1(ori_ori_n1288_), .B0(ori_ori_n1619_), .B1(ori_ori_n477_), .Y(ori_ori_n1621_));
  AO210      o1572(.A0(ori_ori_n1621_), .A1(ori_ori_n1618_), .B0(x1), .Y(ori_ori_n1622_));
  NA2        o1573(.A(ori_ori_n634_), .B(ori_ori_n1062_), .Y(ori_ori_n1623_));
  NA2        o1574(.A(ori_ori_n142_), .B(ori_ori_n107_), .Y(ori_ori_n1624_));
  NOi21      o1575(.An(x1), .B(x6), .Y(ori_ori_n1625_));
  NA2        o1576(.A(ori_ori_n1625_), .B(ori_ori_n84_), .Y(ori_ori_n1626_));
  NA3        o1577(.A(ori_ori_n1626_), .B(ori_ori_n1624_), .C(ori_ori_n1623_), .Y(ori_ori_n1627_));
  AOI220     o1578(.A0(ori_ori_n1627_), .A1(x3), .B0(ori_ori_n1226_), .B1(ori_ori_n381_), .Y(ori_ori_n1628_));
  NA3        o1579(.A(ori_ori_n1231_), .B(ori_ori_n804_), .C(ori_ori_n605_), .Y(ori_ori_n1629_));
  AOI220     o1580(.A0(ori_ori_n1276_), .A1(ori_ori_n118_), .B0(ori_ori_n926_), .B1(ori_ori_n821_), .Y(ori_ori_n1630_));
  AOI210     o1581(.A0(ori_ori_n1630_), .A1(ori_ori_n1629_), .B0(ori_ori_n320_), .Y(ori_ori_n1631_));
  NA3        o1582(.A(ori_ori_n1218_), .B(ori_ori_n382_), .C(ori_ori_n106_), .Y(ori_ori_n1632_));
  NO2        o1583(.A(ori_ori_n1632_), .B(ori_ori_n974_), .Y(ori_ori_n1633_));
  NO3        o1584(.A(ori_ori_n620_), .B(ori_ori_n517_), .C(ori_ori_n1244_), .Y(ori_ori_n1634_));
  NO3        o1585(.A(ori_ori_n1634_), .B(ori_ori_n1633_), .C(ori_ori_n1631_), .Y(ori_ori_n1635_));
  OAI210     o1586(.A0(ori_ori_n1628_), .A1(ori_ori_n855_), .B0(ori_ori_n1635_), .Y(ori_ori_n1636_));
  NO2        o1587(.A(ori_ori_n556_), .B(ori_ori_n68_), .Y(ori_ori_n1637_));
  OAI220     o1588(.A0(ori_ori_n1637_), .A1(ori_ori_n1593_), .B0(ori_ori_n303_), .B1(ori_ori_n905_), .Y(ori_ori_n1638_));
  AOI220     o1589(.A0(ori_ori_n1638_), .A1(ori_ori_n56_), .B0(ori_ori_n1372_), .B1(ori_ori_n735_), .Y(ori_ori_n1639_));
  NO2        o1590(.A(ori_ori_n54_), .B(ori_ori_n71_), .Y(ori_ori_n1640_));
  AO220      o1591(.A0(ori_ori_n1640_), .A1(ori_ori_n1011_), .B0(ori_ori_n821_), .B1(ori_ori_n963_), .Y(ori_ori_n1641_));
  NA2        o1592(.A(ori_ori_n1201_), .B(ori_ori_n358_), .Y(ori_ori_n1642_));
  NO2        o1593(.A(ori_ori_n1004_), .B(ori_ori_n1625_), .Y(ori_ori_n1643_));
  NA2        o1594(.A(ori_ori_n499_), .B(ori_ori_n735_), .Y(ori_ori_n1644_));
  OAI210     o1595(.A0(ori_ori_n1644_), .A1(ori_ori_n1643_), .B0(ori_ori_n1642_), .Y(ori_ori_n1645_));
  AOI210     o1596(.A0(ori_ori_n1641_), .A1(x2), .B0(ori_ori_n1645_), .Y(ori_ori_n1646_));
  OAI220     o1597(.A0(ori_ori_n1646_), .A1(ori_ori_n149_), .B0(ori_ori_n1639_), .B1(ori_ori_n54_), .Y(ori_ori_n1647_));
  OAI210     o1598(.A0(ori_ori_n1647_), .A1(ori_ori_n1636_), .B0(x8), .Y(ori_ori_n1648_));
  NA4        o1599(.A(ori_ori_n1648_), .B(ori_ori_n1622_), .C(ori_ori_n1612_), .D(ori_ori_n1600_), .Y(ori20));
  NA4        o1600(.A(ori_ori_n392_), .B(ori_ori_n276_), .C(ori_ori_n380_), .D(ori_ori_n62_), .Y(ori_ori_n1650_));
  NA2        o1601(.A(ori_ori_n477_), .B(ori_ori_n413_), .Y(ori_ori_n1651_));
  AOI210     o1602(.A0(ori_ori_n1651_), .A1(ori_ori_n1650_), .B0(ori_ori_n87_), .Y(ori_ori_n1652_));
  AOI210     o1603(.A0(ori_ori_n1066_), .A1(ori_ori_n62_), .B0(ori_ori_n1607_), .Y(ori_ori_n1653_));
  AOI210     o1604(.A0(ori_ori_n998_), .A1(ori_ori_n347_), .B0(ori_ori_n1208_), .Y(ori_ori_n1654_));
  OAI210     o1605(.A0(ori_ori_n1653_), .A1(ori_ori_n686_), .B0(ori_ori_n1654_), .Y(ori_ori_n1655_));
  OAI210     o1606(.A0(ori_ori_n1655_), .A1(ori_ori_n1652_), .B0(ori_ori_n1122_), .Y(ori_ori_n1656_));
  NAi21      o1607(.An(ori_ori_n552_), .B(ori_ori_n401_), .Y(ori_ori_n1657_));
  NA3        o1608(.A(ori_ori_n1657_), .B(ori_ori_n996_), .C(ori_ori_n963_), .Y(ori_ori_n1658_));
  NA3        o1609(.A(ori_ori_n1121_), .B(ori_ori_n276_), .C(ori_ori_n586_), .Y(ori_ori_n1659_));
  AOI210     o1610(.A0(ori_ori_n1659_), .A1(ori_ori_n1658_), .B0(ori_ori_n1318_), .Y(ori_ori_n1660_));
  NO2        o1611(.A(ori_ori_n754_), .B(ori_ori_n984_), .Y(ori_ori_n1661_));
  NOi31      o1612(.An(ori_ori_n1661_), .B(ori_ori_n1193_), .C(ori_ori_n530_), .Y(ori_ori_n1662_));
  OAI210     o1613(.A0(ori_ori_n1662_), .A1(ori_ori_n1660_), .B0(ori_ori_n325_), .Y(ori_ori_n1663_));
  NA2        o1614(.A(ori_ori_n316_), .B(ori_ori_n91_), .Y(ori_ori_n1664_));
  NA2        o1615(.A(ori_ori_n326_), .B(ori_ori_n104_), .Y(ori_ori_n1665_));
  NA2        o1616(.A(ori_ori_n423_), .B(ori_ori_n52_), .Y(ori_ori_n1666_));
  OAI220     o1617(.A0(ori_ori_n1666_), .A1(ori_ori_n1665_), .B0(ori_ori_n1664_), .B1(ori_ori_n271_), .Y(ori_ori_n1667_));
  NA2        o1618(.A(ori_ori_n1667_), .B(ori_ori_n217_), .Y(ori_ori_n1668_));
  NO2        o1619(.A(ori_ori_n670_), .B(ori_ori_n609_), .Y(ori_ori_n1669_));
  NA2        o1620(.A(ori_ori_n964_), .B(ori_ori_n50_), .Y(ori_ori_n1670_));
  NO3        o1621(.A(ori_ori_n1670_), .B(ori_ori_n364_), .C(ori_ori_n225_), .Y(ori_ori_n1671_));
  NA4        o1622(.A(ori_ori_n337_), .B(ori_ori_n234_), .C(ori_ori_n809_), .D(ori_ori_n64_), .Y(ori_ori_n1672_));
  OAI220     o1623(.A0(ori_ori_n1672_), .A1(ori_ori_n680_), .B0(ori_ori_n1490_), .B1(ori_ori_n1049_), .Y(ori_ori_n1673_));
  AOI210     o1624(.A0(ori_ori_n1671_), .A1(ori_ori_n1669_), .B0(ori_ori_n1673_), .Y(ori_ori_n1674_));
  NA4        o1625(.A(ori_ori_n1674_), .B(ori_ori_n1668_), .C(ori_ori_n1663_), .D(ori_ori_n1656_), .Y(ori21));
  OAI210     o1626(.A0(ori_ori_n406_), .A1(ori_ori_n54_), .B0(x7), .Y(ori_ori_n1676_));
  OAI220     o1627(.A0(ori_ori_n1676_), .A1(ori_ori_n1308_), .B0(ori_ori_n1067_), .B1(ori_ori_n92_), .Y(ori_ori_n1677_));
  NA2        o1628(.A(ori_ori_n1677_), .B(ori_ori_n78_), .Y(ori_ori_n1678_));
  NA2        o1629(.A(ori_ori_n288_), .B(ori_ori_n866_), .Y(ori_ori_n1679_));
  AOI220     o1630(.A0(ori_ori_n1679_), .A1(ori_ori_n306_), .B0(ori_ori_n571_), .B1(ori_ori_n461_), .Y(ori_ori_n1680_));
  NA2        o1631(.A(ori_ori_n950_), .B(ori_ori_n270_), .Y(ori_ori_n1681_));
  NA2        o1632(.A(ori_ori_n538_), .B(ori_ori_n462_), .Y(ori_ori_n1682_));
  NA4        o1633(.A(ori_ori_n1682_), .B(ori_ori_n1681_), .C(ori_ori_n1399_), .D(ori_ori_n56_), .Y(ori_ori_n1683_));
  NO2        o1634(.A(ori_ori_n782_), .B(ori_ori_n434_), .Y(ori_ori_n1684_));
  NO3        o1635(.A(ori_ori_n1684_), .B(ori_ori_n727_), .C(ori_ori_n246_), .Y(ori_ori_n1685_));
  NOi31      o1636(.An(ori_ori_n188_), .B(ori_ori_n634_), .C(ori_ori_n1105_), .Y(ori_ori_n1686_));
  NO4        o1637(.A(ori_ori_n1686_), .B(ori_ori_n1685_), .C(ori_ori_n1683_), .D(ori_ori_n1680_), .Y(ori_ori_n1687_));
  NO3        o1638(.A(ori_ori_n434_), .B(ori_ori_n274_), .C(ori_ori_n52_), .Y(ori_ori_n1688_));
  OA210      o1639(.A0(ori_ori_n1688_), .A1(ori_ori_n894_), .B0(x3), .Y(ori_ori_n1689_));
  OAI210     o1640(.A0(ori_ori_n793_), .A1(ori_ori_n591_), .B0(ori_ori_n339_), .Y(ori_ori_n1690_));
  NO2        o1641(.A(ori_ori_n70_), .B(x2), .Y(ori_ori_n1691_));
  OAI210     o1642(.A0(ori_ori_n172_), .A1(x0), .B0(ori_ori_n1691_), .Y(ori_ori_n1692_));
  NA2        o1643(.A(ori_ori_n139_), .B(ori_ori_n104_), .Y(ori_ori_n1693_));
  NA3        o1644(.A(ori_ori_n1693_), .B(ori_ori_n1692_), .C(ori_ori_n1690_), .Y(ori_ori_n1694_));
  OAI210     o1645(.A0(ori_ori_n1694_), .A1(ori_ori_n1689_), .B0(x8), .Y(ori_ori_n1695_));
  NO3        o1646(.A(ori_ori_n780_), .B(ori_ori_n623_), .C(ori_ori_n587_), .Y(ori_ori_n1696_));
  NA2        o1647(.A(ori_ori_n55_), .B(ori_ori_n50_), .Y(ori_ori_n1697_));
  MUX2       o1648(.S(ori_ori_n603_), .A(ori_ori_n1697_), .B(ori_ori_n103_), .Y(ori_ori_n1698_));
  AOI210     o1649(.A0(ori_ori_n1377_), .A1(ori_ori_n235_), .B0(ori_ori_n1698_), .Y(ori_ori_n1699_));
  OAI210     o1650(.A0(ori_ori_n647_), .A1(ori_ori_n586_), .B0(x4), .Y(ori_ori_n1700_));
  NO3        o1651(.A(ori_ori_n1700_), .B(ori_ori_n1699_), .C(ori_ori_n1696_), .Y(ori_ori_n1701_));
  AO220      o1652(.A0(ori_ori_n1701_), .A1(ori_ori_n1695_), .B0(ori_ori_n1687_), .B1(ori_ori_n1678_), .Y(ori_ori_n1702_));
  AO220      o1653(.A0(ori_ori_n635_), .A1(ori_ori_n320_), .B0(ori_ori_n592_), .B1(x8), .Y(ori_ori_n1703_));
  NO2        o1654(.A(ori_ori_n868_), .B(x0), .Y(ori_ori_n1704_));
  NO3        o1655(.A(ori_ori_n1704_), .B(ori_ori_n548_), .C(ori_ori_n88_), .Y(ori_ori_n1705_));
  NO2        o1656(.A(ori_ori_n155_), .B(x2), .Y(ori_ori_n1706_));
  NO3        o1657(.A(ori_ori_n377_), .B(ori_ori_n251_), .C(ori_ori_n180_), .Y(ori_ori_n1707_));
  AOI210     o1658(.A0(ori_ori_n1706_), .A1(ori_ori_n68_), .B0(ori_ori_n1707_), .Y(ori_ori_n1708_));
  OAI210     o1659(.A0(ori_ori_n1705_), .A1(ori_ori_n399_), .B0(ori_ori_n1708_), .Y(ori_ori_n1709_));
  AOI220     o1660(.A0(ori_ori_n1709_), .A1(x5), .B0(ori_ori_n1703_), .B1(ori_ori_n754_), .Y(ori_ori_n1710_));
  AOI210     o1661(.A0(ori_ori_n1710_), .A1(ori_ori_n1702_), .B0(ori_ori_n71_), .Y(ori_ori_n1711_));
  NO2        o1662(.A(ori_ori_n916_), .B(ori_ori_n164_), .Y(ori_ori_n1712_));
  NOi41      o1663(.An(ori_ori_n1452_), .B(ori_ori_n1525_), .C(ori_ori_n1176_), .D(ori_ori_n859_), .Y(ori_ori_n1713_));
  NA2        o1664(.A(ori_ori_n1713_), .B(ori_ori_n1712_), .Y(ori_ori_n1714_));
  NO2        o1665(.A(ori_ori_n78_), .B(x4), .Y(ori_ori_n1715_));
  OAI210     o1666(.A0(ori_ori_n286_), .A1(ori_ori_n153_), .B0(ori_ori_n1715_), .Y(ori_ori_n1716_));
  OAI210     o1667(.A0(ori_ori_n408_), .A1(ori_ori_n424_), .B0(ori_ori_n225_), .Y(ori_ori_n1717_));
  NO2        o1668(.A(ori_ori_n253_), .B(ori_ori_n50_), .Y(ori_ori_n1718_));
  NO2        o1669(.A(ori_ori_n1718_), .B(ori_ori_n57_), .Y(ori_ori_n1719_));
  NA2        o1670(.A(ori_ori_n1719_), .B(ori_ori_n1717_), .Y(ori_ori_n1720_));
  AOI210     o1671(.A0(ori_ori_n1716_), .A1(ori_ori_n1714_), .B0(ori_ori_n1720_), .Y(ori_ori_n1721_));
  NA2        o1672(.A(ori_ori_n766_), .B(ori_ori_n552_), .Y(ori_ori_n1722_));
  AO210      o1673(.A0(ori_ori_n1722_), .A1(ori_ori_n974_), .B0(ori_ori_n50_), .Y(ori_ori_n1723_));
  NO2        o1674(.A(ori_ori_n1657_), .B(ori_ori_n1238_), .Y(ori_ori_n1724_));
  AOI220     o1675(.A0(ori_ori_n1724_), .A1(ori_ori_n1186_), .B0(ori_ori_n1344_), .B1(ori_ori_n1060_), .Y(ori_ori_n1725_));
  AOI210     o1676(.A0(ori_ori_n1725_), .A1(ori_ori_n1723_), .B0(ori_ori_n106_), .Y(ori_ori_n1726_));
  NA2        o1677(.A(ori_ori_n295_), .B(ori_ori_n104_), .Y(ori_ori_n1727_));
  NA2        o1678(.A(ori_ori_n904_), .B(ori_ori_n55_), .Y(ori_ori_n1728_));
  NO2        o1679(.A(ori_ori_n675_), .B(ori_ori_n1070_), .Y(ori_ori_n1729_));
  NO3        o1680(.A(ori_ori_n1729_), .B(ori_ori_n1726_), .C(ori_ori_n1721_), .Y(ori_ori_n1730_));
  NO2        o1681(.A(ori_ori_n1730_), .B(x6), .Y(ori_ori_n1731_));
  AOI210     o1682(.A0(ori_ori_n612_), .A1(ori_ori_n1070_), .B0(ori_ori_n1525_), .Y(ori_ori_n1732_));
  OAI210     o1683(.A0(ori_ori_n1732_), .A1(ori_ori_n693_), .B0(ori_ori_n56_), .Y(ori_ori_n1733_));
  NO2        o1684(.A(ori_ori_n756_), .B(ori_ori_n54_), .Y(ori_ori_n1734_));
  NO4        o1685(.A(ori_ori_n972_), .B(ori_ori_n274_), .C(ori_ori_n779_), .D(ori_ori_n763_), .Y(ori_ori_n1735_));
  NO2        o1686(.A(ori_ori_n873_), .B(x5), .Y(ori_ori_n1736_));
  NO4        o1687(.A(ori_ori_n1736_), .B(ori_ori_n1735_), .C(ori_ori_n1734_), .D(ori_ori_n957_), .Y(ori_ori_n1737_));
  AOI210     o1688(.A0(ori_ori_n1737_), .A1(ori_ori_n1733_), .B0(ori_ori_n50_), .Y(ori_ori_n1738_));
  NA2        o1689(.A(ori_ori_n155_), .B(ori_ori_n104_), .Y(ori_ori_n1739_));
  OA220      o1690(.A0(ori_ori_n1739_), .A1(ori_ori_n438_), .B0(ori_ori_n467_), .B1(ori_ori_n754_), .Y(ori_ori_n1740_));
  NA3        o1691(.A(ori_ori_n55_), .B(x2), .C(x0), .Y(ori_ori_n1741_));
  AOI220     o1692(.A0(ori_ori_n1741_), .A1(ori_ori_n166_), .B0(ori_ori_n873_), .B1(ori_ori_n151_), .Y(ori_ori_n1742_));
  NO2        o1693(.A(ori_ori_n686_), .B(ori_ori_n253_), .Y(ori_ori_n1743_));
  NO3        o1694(.A(ori_ori_n241_), .B(ori_ori_n223_), .C(ori_ori_n358_), .Y(ori_ori_n1744_));
  NO3        o1695(.A(ori_ori_n1744_), .B(ori_ori_n1743_), .C(ori_ori_n1742_), .Y(ori_ori_n1745_));
  OAI220     o1696(.A0(ori_ori_n1745_), .A1(ori_ori_n56_), .B0(ori_ori_n1740_), .B1(ori_ori_n702_), .Y(ori_ori_n1746_));
  OAI210     o1697(.A0(ori_ori_n1746_), .A1(ori_ori_n1738_), .B0(ori_ori_n112_), .Y(ori_ori_n1747_));
  NO2        o1698(.A(ori_ori_n617_), .B(ori_ori_n301_), .Y(ori_ori_n1748_));
  AOI210     o1699(.A0(ori_ori_n610_), .A1(x5), .B0(ori_ori_n1748_), .Y(ori_ori_n1749_));
  NO2        o1700(.A(ori_ori_n1749_), .B(ori_ori_n106_), .Y(ori_ori_n1750_));
  NA2        o1701(.A(ori_ori_n710_), .B(ori_ori_n81_), .Y(ori_ori_n1751_));
  NA3        o1702(.A(ori_ori_n1751_), .B(ori_ori_n431_), .C(ori_ori_n57_), .Y(ori_ori_n1752_));
  OAI210     o1703(.A0(ori_ori_n1728_), .A1(ori_ori_n1727_), .B0(ori_ori_n1752_), .Y(ori_ori_n1753_));
  OAI210     o1704(.A0(ori_ori_n1753_), .A1(ori_ori_n1750_), .B0(x1), .Y(ori_ori_n1754_));
  NO4        o1705(.A(ori_ori_n417_), .B(ori_ori_n78_), .C(ori_ori_n143_), .D(x3), .Y(ori_ori_n1755_));
  NO2        o1706(.A(ori_ori_n326_), .B(ori_ori_n108_), .Y(ori_ori_n1756_));
  OAI210     o1707(.A0(ori_ori_n1755_), .A1(ori_ori_n1319_), .B0(ori_ori_n1756_), .Y(ori_ori_n1757_));
  NO2        o1708(.A(ori_ori_n60_), .B(ori_ori_n104_), .Y(ori_ori_n1758_));
  NO4        o1709(.A(ori_ori_n1727_), .B(ori_ori_n972_), .C(ori_ori_n670_), .D(ori_ori_n50_), .Y(ori_ori_n1759_));
  AOI210     o1710(.A0(ori_ori_n1758_), .A1(ori_ori_n1569_), .B0(ori_ori_n1759_), .Y(ori_ori_n1760_));
  NA4        o1711(.A(ori_ori_n1760_), .B(ori_ori_n1757_), .C(ori_ori_n1754_), .D(ori_ori_n1747_), .Y(ori_ori_n1761_));
  NO3        o1712(.A(ori_ori_n1761_), .B(ori_ori_n1731_), .C(ori_ori_n1711_), .Y(ori22));
  AOI210     o1713(.A0(ori_ori_n524_), .A1(ori_ori_n71_), .B0(ori_ori_n470_), .Y(ori_ori_n1763_));
  NO3        o1714(.A(ori_ori_n1213_), .B(ori_ori_n556_), .C(ori_ori_n704_), .Y(ori_ori_n1764_));
  AOI210     o1715(.A0(x5), .A1(x2), .B0(x8), .Y(ori_ori_n1765_));
  NA2        o1716(.A(ori_ori_n1765_), .B(ori_ori_n59_), .Y(ori_ori_n1766_));
  OAI220     o1717(.A0(ori_ori_n1766_), .A1(ori_ori_n1764_), .B0(ori_ori_n1763_), .B1(ori_ori_n399_), .Y(ori_ori_n1767_));
  NA2        o1718(.A(ori_ori_n586_), .B(ori_ori_n87_), .Y(ori_ori_n1768_));
  NA2        o1719(.A(ori_ori_n271_), .B(ori_ori_n77_), .Y(ori_ori_n1769_));
  OA220      o1720(.A0(ori_ori_n1769_), .A1(ori_ori_n1768_), .B0(ori_ori_n852_), .B1(ori_ori_n1021_), .Y(ori_ori_n1770_));
  NO3        o1721(.A(ori_ori_n1267_), .B(ori_ori_n87_), .C(x0), .Y(ori_ori_n1771_));
  OAI210     o1722(.A0(ori_ori_n399_), .A1(ori_ori_n200_), .B0(x4), .Y(ori_ori_n1772_));
  NO2        o1723(.A(ori_ori_n1772_), .B(ori_ori_n1771_), .Y(ori_ori_n1773_));
  OAI210     o1724(.A0(ori_ori_n1770_), .A1(ori_ori_n193_), .B0(ori_ori_n1773_), .Y(ori_ori_n1774_));
  AOI210     o1725(.A0(ori_ori_n1767_), .A1(ori_ori_n53_), .B0(ori_ori_n1774_), .Y(ori_ori_n1775_));
  NA2        o1726(.A(ori_ori_n299_), .B(ori_ori_n304_), .Y(ori_ori_n1776_));
  NA3        o1727(.A(ori_ori_n1776_), .B(ori_ori_n217_), .C(ori_ori_n303_), .Y(ori_ori_n1777_));
  NA2        o1728(.A(ori_ori_n581_), .B(ori_ori_n240_), .Y(ori_ori_n1778_));
  NA2        o1729(.A(ori_ori_n1778_), .B(ori_ori_n1777_), .Y(ori_ori_n1779_));
  NO2        o1730(.A(ori_ori_n467_), .B(ori_ori_n255_), .Y(ori_ori_n1780_));
  INV        o1731(.A(ori_ori_n1780_), .Y(ori_ori_n1781_));
  OAI210     o1732(.A0(ori_ori_n1100_), .A1(ori_ori_n182_), .B0(ori_ori_n56_), .Y(ori_ori_n1782_));
  NA3        o1733(.A(ori_ori_n55_), .B(ori_ori_n71_), .C(x0), .Y(ori_ori_n1783_));
  OAI220     o1734(.A0(ori_ori_n1783_), .A1(ori_ori_n1070_), .B0(ori_ori_n364_), .B1(ori_ori_n208_), .Y(ori_ori_n1784_));
  NO2        o1735(.A(ori_ori_n1784_), .B(ori_ori_n1782_), .Y(ori_ori_n1785_));
  OAI210     o1736(.A0(ori_ori_n1781_), .A1(ori_ori_n253_), .B0(ori_ori_n1785_), .Y(ori_ori_n1786_));
  AOI210     o1737(.A0(ori_ori_n1779_), .A1(ori_ori_n104_), .B0(ori_ori_n1786_), .Y(ori_ori_n1787_));
  AOI210     o1738(.A0(ori_ori_n961_), .A1(ori_ori_n781_), .B0(ori_ori_n877_), .Y(ori_ori_n1788_));
  OAI210     o1739(.A0(ori_ori_n811_), .A1(ori_ori_n155_), .B0(ori_ori_n947_), .Y(ori_ori_n1789_));
  OAI210     o1740(.A0(ori_ori_n1789_), .A1(ori_ori_n1788_), .B0(ori_ori_n616_), .Y(ori_ori_n1790_));
  OA210      o1741(.A0(ori_ori_n1787_), .A1(ori_ori_n1775_), .B0(ori_ori_n1790_), .Y(ori_ori_n1791_));
  OAI210     o1742(.A0(ori_ori_n1195_), .A1(ori_ori_n709_), .B0(ori_ori_n697_), .Y(ori_ori_n1792_));
  NO2        o1743(.A(ori_ori_n352_), .B(x0), .Y(ori_ori_n1793_));
  NA3        o1744(.A(ori_ori_n1793_), .B(ori_ori_n347_), .C(ori_ori_n56_), .Y(ori_ori_n1794_));
  AOI210     o1745(.A0(ori_ori_n1794_), .A1(ori_ori_n1792_), .B0(ori_ori_n399_), .Y(ori_ori_n1795_));
  NO3        o1746(.A(ori_ori_n166_), .B(ori_ori_n155_), .C(ori_ori_n62_), .Y(ori_ori_n1796_));
  OAI210     o1747(.A0(ori_ori_n1796_), .A1(ori_ori_n419_), .B0(ori_ori_n106_), .Y(ori_ori_n1797_));
  NA2        o1748(.A(ori_ori_n135_), .B(ori_ori_n794_), .Y(ori_ori_n1798_));
  NA2        o1749(.A(ori_ori_n417_), .B(x3), .Y(ori_ori_n1799_));
  NAi31      o1750(.An(ori_ori_n1799_), .B(ori_ori_n1798_), .C(ori_ori_n1585_), .Y(ori_ori_n1800_));
  NO3        o1751(.A(ori_ori_n868_), .B(ori_ori_n466_), .C(ori_ori_n106_), .Y(ori_ori_n1801_));
  NO2        o1752(.A(ori_ori_n1102_), .B(ori_ori_n136_), .Y(ori_ori_n1802_));
  NO3        o1753(.A(ori_ori_n907_), .B(ori_ori_n413_), .C(ori_ori_n300_), .Y(ori_ori_n1803_));
  AOI220     o1754(.A0(ori_ori_n1803_), .A1(ori_ori_n1802_), .B0(ori_ori_n1801_), .B1(ori_ori_n1793_), .Y(ori_ori_n1804_));
  NA3        o1755(.A(ori_ori_n413_), .B(ori_ori_n91_), .C(ori_ori_n81_), .Y(ori_ori_n1805_));
  AOI210     o1756(.A0(ori_ori_n612_), .A1(ori_ori_n456_), .B0(ori_ori_n496_), .Y(ori_ori_n1806_));
  NA2        o1757(.A(ori_ori_n1197_), .B(x3), .Y(ori_ori_n1807_));
  OAI210     o1758(.A0(ori_ori_n1807_), .A1(ori_ori_n1806_), .B0(ori_ori_n1805_), .Y(ori_ori_n1808_));
  NA3        o1759(.A(ori_ori_n56_), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n1809_));
  NOi21      o1760(.An(ori_ori_n83_), .B(ori_ori_n738_), .Y(ori_ori_n1810_));
  NA3        o1761(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n1811_));
  NA3        o1762(.A(ori_ori_n1811_), .B(ori_ori_n1004_), .C(ori_ori_n262_), .Y(ori_ori_n1812_));
  OAI220     o1763(.A0(ori_ori_n1812_), .A1(ori_ori_n1810_), .B0(ori_ori_n1073_), .B1(ori_ori_n1809_), .Y(ori_ori_n1813_));
  AOI220     o1764(.A0(ori_ori_n1813_), .A1(ori_ori_n1084_), .B0(ori_ori_n1808_), .B1(ori_ori_n347_), .Y(ori_ori_n1814_));
  NA4        o1765(.A(ori_ori_n1814_), .B(ori_ori_n1804_), .C(ori_ori_n1800_), .D(ori_ori_n1797_), .Y(ori_ori_n1815_));
  AOI210     o1766(.A0(ori_ori_n1815_), .A1(x7), .B0(ori_ori_n1795_), .Y(ori_ori_n1816_));
  OAI210     o1767(.A0(ori_ori_n1791_), .A1(x7), .B0(ori_ori_n1816_), .Y(ori23));
  OR2        o1768(.A(ori_ori_n518_), .B(ori_ori_n217_), .Y(ori_ori_n1818_));
  AOI220     o1769(.A0(ori_ori_n1818_), .A1(ori_ori_n1661_), .B0(ori_ori_n618_), .B1(ori_ori_n291_), .Y(ori_ori_n1819_));
  NO3        o1770(.A(ori_ori_n852_), .B(ori_ori_n595_), .C(ori_ori_n489_), .Y(ori_ori_n1820_));
  NO3        o1771(.A(ori_ori_n965_), .B(ori_ori_n144_), .C(ori_ori_n113_), .Y(ori_ori_n1821_));
  AOI210     o1772(.A0(ori_ori_n1821_), .A1(ori_ori_n1043_), .B0(ori_ori_n1820_), .Y(ori_ori_n1822_));
  OAI210     o1773(.A0(ori_ori_n1819_), .A1(ori_ori_n149_), .B0(ori_ori_n1822_), .Y(ori_ori_n1823_));
  NA2        o1774(.A(ori_ori_n1823_), .B(ori_ori_n55_), .Y(ori_ori_n1824_));
  NO2        o1775(.A(ori_ori_n972_), .B(ori_ori_n516_), .Y(ori_ori_n1825_));
  AO220      o1776(.A0(ori_ori_n1304_), .A1(ori_ori_n176_), .B0(ori_ori_n1011_), .B1(ori_ori_n754_), .Y(ori_ori_n1826_));
  OAI210     o1777(.A0(ori_ori_n1826_), .A1(ori_ori_n1825_), .B0(ori_ori_n592_), .Y(ori_ori_n1827_));
  NA2        o1778(.A(ori_ori_n173_), .B(ori_ori_n164_), .Y(ori_ori_n1828_));
  NA2        o1779(.A(ori_ori_n405_), .B(ori_ori_n156_), .Y(ori_ori_n1829_));
  AOI210     o1780(.A0(ori_ori_n1829_), .A1(ori_ori_n1828_), .B0(ori_ori_n232_), .Y(ori_ori_n1830_));
  NA3        o1781(.A(ori_ori_n877_), .B(ori_ori_n424_), .C(ori_ori_n253_), .Y(ori_ori_n1831_));
  AOI210     o1782(.A0(ori_ori_n1831_), .A1(ori_ori_n501_), .B0(ori_ori_n382_), .Y(ori_ori_n1832_));
  OAI210     o1783(.A0(ori_ori_n1832_), .A1(ori_ori_n1830_), .B0(ori_ori_n295_), .Y(ori_ori_n1833_));
  NA3        o1784(.A(ori_ori_n57_), .B(x4), .C(x3), .Y(ori_ori_n1834_));
  NO3        o1785(.A(ori_ori_n1834_), .B(ori_ori_n751_), .C(ori_ori_n135_), .Y(ori_ori_n1835_));
  AOI210     o1786(.A0(ori_ori_n930_), .A1(ori_ori_n137_), .B0(ori_ori_n1835_), .Y(ori_ori_n1836_));
  NA4        o1787(.A(ori_ori_n1836_), .B(ori_ori_n1833_), .C(ori_ori_n1827_), .D(ori_ori_n1824_), .Y(ori24));
  NO2        o1788(.A(ori_ori_n237_), .B(x1), .Y(ori_ori_n1838_));
  NA2        o1789(.A(ori_ori_n337_), .B(ori_ori_n493_), .Y(ori_ori_n1839_));
  NAi21      o1790(.An(ori_ori_n1838_), .B(ori_ori_n1839_), .Y(ori_ori_n1840_));
  NO3        o1791(.A(ori_ori_n543_), .B(ori_ori_n689_), .C(ori_ori_n151_), .Y(ori_ori_n1841_));
  AOI210     o1792(.A0(ori_ori_n1840_), .A1(ori_ori_n91_), .B0(ori_ori_n1841_), .Y(ori_ori_n1842_));
  NA2        o1793(.A(ori_ori_n98_), .B(x8), .Y(ori_ori_n1843_));
  NO3        o1794(.A(ori_ori_n1081_), .B(ori_ori_n1358_), .C(ori_ori_n1062_), .Y(ori_ori_n1844_));
  AOI210     o1795(.A0(ori_ori_n996_), .A1(ori_ori_n56_), .B0(ori_ori_n1476_), .Y(ori_ori_n1845_));
  AO220      o1796(.A0(ori_ori_n1845_), .A1(ori_ori_n1844_), .B0(ori_ori_n1290_), .B1(ori_ori_n325_), .Y(ori_ori_n1846_));
  NA2        o1797(.A(ori_ori_n456_), .B(x8), .Y(ori_ori_n1847_));
  NA2        o1798(.A(ori_ori_n671_), .B(ori_ori_n121_), .Y(ori_ori_n1848_));
  OAI220     o1799(.A0(ori_ori_n1848_), .A1(ori_ori_n1461_), .B0(ori_ori_n1847_), .B1(ori_ori_n850_), .Y(ori_ori_n1849_));
  AOI220     o1800(.A0(ori_ori_n1849_), .A1(ori_ori_n1718_), .B0(ori_ori_n1846_), .B1(ori_ori_n1043_), .Y(ori_ori_n1850_));
  OAI210     o1801(.A0(ori_ori_n1843_), .A1(ori_ori_n1842_), .B0(ori_ori_n1850_), .Y(ori25));
  NA2        o1802(.A(ori_ori_n326_), .B(ori_ori_n59_), .Y(ori_ori_n1852_));
  NO2        o1803(.A(ori_ori_n1852_), .B(ori_ori_n317_), .Y(ori_ori_n1853_));
  OAI210     o1804(.A0(ori_ori_n1853_), .A1(ori_ori_n1202_), .B0(ori_ori_n112_), .Y(ori_ori_n1854_));
  NA2        o1805(.A(ori_ori_n1619_), .B(ori_ori_n1203_), .Y(ori_ori_n1855_));
  AOI210     o1806(.A0(ori_ori_n1855_), .A1(ori_ori_n1854_), .B0(ori_ori_n684_), .Y(ori_ori_n1856_));
  NO3        o1807(.A(ori_ori_n1055_), .B(ori_ori_n138_), .C(ori_ori_n78_), .Y(ori_ori_n1857_));
  OAI210     o1808(.A0(ori_ori_n193_), .A1(ori_ori_n271_), .B0(ori_ori_n327_), .Y(ori_ori_n1858_));
  OAI210     o1809(.A0(ori_ori_n1858_), .A1(ori_ori_n1857_), .B0(ori_ori_n1201_), .Y(ori_ori_n1859_));
  NO2        o1810(.A(ori_ori_n1411_), .B(ori_ori_n449_), .Y(ori_ori_n1860_));
  NO3        o1811(.A(ori_ori_n1860_), .B(ori_ori_n534_), .C(ori_ori_n95_), .Y(ori_ori_n1861_));
  NA2        o1812(.A(ori_ori_n511_), .B(ori_ori_n55_), .Y(ori_ori_n1862_));
  OAI220     o1813(.A0(ori_ori_n1862_), .A1(ori_ori_n237_), .B0(ori_ori_n589_), .B1(ori_ori_n271_), .Y(ori_ori_n1863_));
  OAI210     o1814(.A0(ori_ori_n1863_), .A1(ori_ori_n1861_), .B0(ori_ori_n639_), .Y(ori_ori_n1864_));
  AOI220     o1815(.A0(ori_ori_n1780_), .A1(ori_ori_n1155_), .B0(ori_ori_n1519_), .B1(ori_ori_n378_), .Y(ori_ori_n1865_));
  NA3        o1816(.A(ori_ori_n1865_), .B(ori_ori_n1864_), .C(ori_ori_n1859_), .Y(ori_ori_n1866_));
  AO210      o1817(.A0(ori_ori_n1866_), .A1(ori_ori_n104_), .B0(ori_ori_n1856_), .Y(ori26));
  NA2        o1818(.A(ori_ori_n779_), .B(ori_ori_n50_), .Y(ori_ori_n1868_));
  OAI220     o1819(.A0(ori_ori_n301_), .A1(ori_ori_n246_), .B0(ori_ori_n1868_), .B1(x7), .Y(ori_ori_n1869_));
  AOI220     o1820(.A0(ori_ori_n1869_), .A1(ori_ori_n91_), .B0(ori_ori_n1319_), .B1(ori_ori_n1161_), .Y(ori_ori_n1870_));
  NA2        o1821(.A(ori_ori_n627_), .B(ori_ori_n581_), .Y(ori_ori_n1871_));
  OAI210     o1822(.A0(ori_ori_n635_), .A1(ori_ori_n627_), .B0(ori_ori_n754_), .Y(ori_ori_n1872_));
  AOI210     o1823(.A0(ori_ori_n1871_), .A1(ori_ori_n1225_), .B0(ori_ori_n1872_), .Y(ori_ori_n1873_));
  NA2        o1824(.A(ori_ori_n1034_), .B(ori_ori_n587_), .Y(ori_ori_n1874_));
  NO2        o1825(.A(ori_ori_n1874_), .B(ori_ori_n1272_), .Y(ori_ori_n1875_));
  AOI210     o1826(.A0(ori_ori_n1802_), .A1(ori_ori_n1484_), .B0(ori_ori_n1875_), .Y(ori_ori_n1876_));
  NO2        o1827(.A(ori_ori_n1102_), .B(ori_ori_n75_), .Y(ori_ori_n1877_));
  NA2        o1828(.A(ori_ori_n819_), .B(ori_ori_n172_), .Y(ori_ori_n1878_));
  NO2        o1829(.A(ori_ori_n1878_), .B(ori_ori_n539_), .Y(ori_ori_n1879_));
  AOI210     o1830(.A0(ori_ori_n1877_), .A1(ori_ori_n588_), .B0(ori_ori_n1879_), .Y(ori_ori_n1880_));
  OAI220     o1831(.A0(ori_ori_n1880_), .A1(ori_ori_n104_), .B0(ori_ori_n1876_), .B1(ori_ori_n53_), .Y(ori_ori_n1881_));
  NA2        o1832(.A(ori_ori_n604_), .B(ori_ori_n511_), .Y(ori_ori_n1882_));
  NO2        o1833(.A(ori_ori_n128_), .B(ori_ori_n125_), .Y(ori_ori_n1883_));
  NA2        o1834(.A(ori_ori_n1883_), .B(ori_ori_n118_), .Y(ori_ori_n1884_));
  NA2        o1835(.A(ori_ori_n754_), .B(x3), .Y(ori_ori_n1885_));
  AOI210     o1836(.A0(ori_ori_n1884_), .A1(ori_ori_n1882_), .B0(ori_ori_n1885_), .Y(ori_ori_n1886_));
  NO2        o1837(.A(ori_ori_n1021_), .B(x3), .Y(ori_ori_n1887_));
  AOI210     o1838(.A0(ori_ori_n447_), .A1(ori_ori_n104_), .B0(ori_ori_n1887_), .Y(ori_ori_n1888_));
  NA3        o1839(.A(ori_ori_n572_), .B(ori_ori_n51_), .C(ori_ori_n56_), .Y(ori_ori_n1889_));
  AOI210     o1840(.A0(ori_ori_n1669_), .A1(ori_ori_n1074_), .B0(x0), .Y(ori_ori_n1890_));
  OAI210     o1841(.A0(ori_ori_n1889_), .A1(ori_ori_n1888_), .B0(ori_ori_n1890_), .Y(ori_ori_n1891_));
  NO4        o1842(.A(ori_ori_n1891_), .B(ori_ori_n1886_), .C(ori_ori_n1881_), .D(ori_ori_n1873_), .Y(ori_ori_n1892_));
  AOI210     o1843(.A0(x8), .A1(x6), .B0(x5), .Y(ori_ori_n1893_));
  AO220      o1844(.A0(ori_ori_n1893_), .A1(ori_ori_n140_), .B0(ori_ori_n595_), .B1(ori_ori_n135_), .Y(ori_ori_n1894_));
  NA2        o1845(.A(ori_ori_n1894_), .B(ori_ori_n448_), .Y(ori_ori_n1895_));
  NO2        o1846(.A(ori_ori_n764_), .B(ori_ori_n140_), .Y(ori_ori_n1896_));
  NA3        o1847(.A(ori_ori_n1896_), .B(ori_ori_n1691_), .C(ori_ori_n129_), .Y(ori_ori_n1897_));
  NO2        o1848(.A(ori_ori_n399_), .B(ori_ori_n1397_), .Y(ori_ori_n1898_));
  OAI210     o1849(.A0(ori_ori_n1898_), .A1(ori_ori_n1364_), .B0(ori_ori_n447_), .Y(ori_ori_n1899_));
  NA3        o1850(.A(ori_ori_n372_), .B(ori_ori_n866_), .C(ori_ori_n250_), .Y(ori_ori_n1900_));
  NA4        o1851(.A(ori_ori_n1900_), .B(ori_ori_n1899_), .C(ori_ori_n1897_), .D(ori_ori_n1895_), .Y(ori_ori_n1901_));
  AOI210     o1852(.A0(ori_ori_n219_), .A1(x2), .B0(ori_ori_n494_), .Y(ori_ori_n1902_));
  NO2        o1853(.A(ori_ori_n1902_), .B(ori_ori_n113_), .Y(ori_ori_n1903_));
  NA3        o1854(.A(ori_ori_n821_), .B(ori_ori_n1021_), .C(x7), .Y(ori_ori_n1904_));
  AOI210     o1855(.A0(ori_ori_n341_), .A1(ori_ori_n211_), .B0(ori_ori_n1904_), .Y(ori_ori_n1905_));
  OAI220     o1856(.A0(ori_ori_n910_), .A1(ori_ori_n301_), .B0(ori_ori_n647_), .B1(ori_ori_n689_), .Y(ori_ori_n1906_));
  NO3        o1857(.A(ori_ori_n1906_), .B(ori_ori_n1905_), .C(ori_ori_n1903_), .Y(ori_ori_n1907_));
  NA3        o1858(.A(ori_ori_n671_), .B(ori_ori_n187_), .C(ori_ori_n963_), .Y(ori_ori_n1908_));
  NA2        o1859(.A(ori_ori_n1908_), .B(ori_ori_n647_), .Y(ori_ori_n1909_));
  NA2        o1860(.A(ori_ori_n135_), .B(ori_ori_n127_), .Y(ori_ori_n1910_));
  OAI210     o1861(.A0(ori_ori_n1910_), .A1(ori_ori_n1447_), .B0(x0), .Y(ori_ori_n1911_));
  AOI210     o1862(.A0(ori_ori_n1909_), .A1(ori_ori_n1435_), .B0(ori_ori_n1911_), .Y(ori_ori_n1912_));
  OAI210     o1863(.A0(ori_ori_n1907_), .A1(ori_ori_n53_), .B0(ori_ori_n1912_), .Y(ori_ori_n1913_));
  AOI210     o1864(.A0(ori_ori_n1901_), .A1(x4), .B0(ori_ori_n1913_), .Y(ori_ori_n1914_));
  OA220      o1865(.A0(ori_ori_n1914_), .A1(ori_ori_n1892_), .B0(ori_ori_n1870_), .B1(ori_ori_n105_), .Y(ori27));
  NA2        o1866(.A(ori_ori_n1165_), .B(ori_ori_n447_), .Y(ori_ori_n1916_));
  NO2        o1867(.A(ori_ori_n1916_), .B(ori_ori_n296_), .Y(ori_ori_n1917_));
  NA2        o1868(.A(ori_ori_n926_), .B(ori_ori_n821_), .Y(ori_ori_n1918_));
  NA3        o1869(.A(ori_ori_n827_), .B(ori_ori_n361_), .C(ori_ori_n1036_), .Y(ori_ori_n1919_));
  AOI210     o1870(.A0(ori_ori_n1919_), .A1(ori_ori_n1918_), .B0(ori_ori_n211_), .Y(ori_ori_n1920_));
  OAI210     o1871(.A0(ori_ori_n1920_), .A1(ori_ori_n1917_), .B0(ori_ori_n705_), .Y(ori_ori_n1921_));
  XO2        o1872(.A(x8), .B(x4), .Y(ori_ori_n1922_));
  NO3        o1873(.A(ori_ori_n1922_), .B(ori_ori_n447_), .C(ori_ori_n166_), .Y(ori_ori_n1923_));
  OA210      o1874(.A0(ori_ori_n1923_), .A1(ori_ori_n1273_), .B0(ori_ori_n274_), .Y(ori_ori_n1924_));
  NO2        o1875(.A(ori_ori_n394_), .B(ori_ori_n160_), .Y(ori_ori_n1925_));
  OAI210     o1876(.A0(ori_ori_n1925_), .A1(ori_ori_n1924_), .B0(ori_ori_n1139_), .Y(ori_ori_n1926_));
  AOI210     o1877(.A0(ori_ori_n635_), .A1(ori_ori_n56_), .B0(ori_ori_n1877_), .Y(ori_ori_n1927_));
  OAI220     o1878(.A0(ori_ori_n1927_), .A1(ori_ori_n1272_), .B0(ori_ori_n1223_), .B1(ori_ori_n202_), .Y(ori_ori_n1928_));
  NA2        o1879(.A(ori_ori_n1928_), .B(ori_ori_n538_), .Y(ori_ori_n1929_));
  NA3        o1880(.A(ori_ori_n1929_), .B(ori_ori_n1926_), .C(ori_ori_n1921_), .Y(ori28));
  NO3        o1881(.A(ori_ori_n1922_), .B(ori_ori_n1406_), .C(ori_ori_n142_), .Y(ori_ori_n1931_));
  OAI210     o1882(.A0(ori_ori_n1931_), .A1(ori_ori_n1292_), .B0(ori_ori_n587_), .Y(ori_ori_n1932_));
  NA3        o1883(.A(ori_ori_n1203_), .B(ori_ori_n904_), .C(x7), .Y(ori_ori_n1933_));
  NA3        o1884(.A(ori_ori_n496_), .B(ori_ori_n78_), .C(ori_ori_n609_), .Y(ori_ori_n1934_));
  NA3        o1885(.A(ori_ori_n1934_), .B(ori_ori_n1933_), .C(ori_ori_n1932_), .Y(ori_ori_n1935_));
  NA2        o1886(.A(ori_ori_n1267_), .B(ori_ori_n445_), .Y(ori_ori_n1936_));
  NA3        o1887(.A(ori_ori_n1936_), .B(ori_ori_n1424_), .C(ori_ori_n412_), .Y(ori_ori_n1937_));
  NO2        o1888(.A(ori_ori_n304_), .B(x4), .Y(ori_ori_n1938_));
  AOI220     o1889(.A0(ori_ori_n1938_), .A1(ori_ori_n1887_), .B0(ori_ori_n1140_), .B1(ori_ori_n679_), .Y(ori_ori_n1939_));
  NA2        o1890(.A(ori_ori_n1939_), .B(ori_ori_n1937_), .Y(ori_ori_n1940_));
  NO2        o1891(.A(ori_ori_n1267_), .B(ori_ori_n1244_), .Y(ori_ori_n1941_));
  NO4        o1892(.A(x6), .B(ori_ori_n56_), .C(x2), .D(x0), .Y(ori_ori_n1942_));
  OAI210     o1893(.A0(ori_ori_n1942_), .A1(ori_ori_n1941_), .B0(ori_ori_n1060_), .Y(ori_ori_n1943_));
  NA2        o1894(.A(ori_ori_n1197_), .B(ori_ori_n104_), .Y(ori_ori_n1944_));
  NA2        o1895(.A(ori_ori_n1098_), .B(ori_ori_n103_), .Y(ori_ori_n1945_));
  OAI210     o1896(.A0(ori_ori_n1945_), .A1(ori_ori_n1944_), .B0(ori_ori_n1943_), .Y(ori_ori_n1946_));
  OAI210     o1897(.A0(ori_ori_n1946_), .A1(ori_ori_n1940_), .B0(x7), .Y(ori_ori_n1947_));
  NO2        o1898(.A(ori_ori_n385_), .B(x7), .Y(ori_ori_n1948_));
  NO3        o1899(.A(ori_ori_n399_), .B(ori_ori_n268_), .C(ori_ori_n119_), .Y(ori_ori_n1949_));
  OAI220     o1900(.A0(ori_ori_n2696_), .A1(ori_ori_n1949_), .B0(ori_ori_n1948_), .B1(ori_ori_n107_), .Y(ori_ori_n1950_));
  NA2        o1901(.A(ori_ori_n1811_), .B(ori_ori_n659_), .Y(ori_ori_n1951_));
  NO2        o1902(.A(ori_ori_n1862_), .B(ori_ori_n77_), .Y(ori_ori_n1952_));
  AOI220     o1903(.A0(ori_ori_n1952_), .A1(ori_ori_n1951_), .B0(ori_ori_n478_), .B1(ori_ori_n50_), .Y(ori_ori_n1953_));
  AOI210     o1904(.A0(ori_ori_n1953_), .A1(ori_ori_n1950_), .B0(ori_ori_n59_), .Y(ori_ori_n1954_));
  AOI220     o1905(.A0(ori_ori_n1411_), .A1(ori_ori_n677_), .B0(ori_ori_n411_), .B1(ori_ori_n456_), .Y(ori_ori_n1955_));
  OAI210     o1906(.A0(ori_ori_n1955_), .A1(ori_ori_n138_), .B0(x1), .Y(ori_ori_n1956_));
  NO2        o1907(.A(ori_ori_n1956_), .B(ori_ori_n1954_), .Y(ori_ori_n1957_));
  AOI210     o1908(.A0(ori_ori_n1604_), .A1(ori_ori_n399_), .B0(ori_ori_n669_), .Y(ori_ori_n1958_));
  NO2        o1909(.A(ori_ori_n399_), .B(x5), .Y(ori_ori_n1959_));
  NO2        o1910(.A(ori_ori_n1959_), .B(ori_ori_n223_), .Y(ori_ori_n1960_));
  NO2        o1911(.A(ori_ori_n1960_), .B(ori_ori_n1958_), .Y(ori_ori_n1961_));
  NOi21      o1912(.An(ori_ori_n710_), .B(ori_ori_n1011_), .Y(ori_ori_n1962_));
  NA3        o1913(.A(ori_ori_n1962_), .B(ori_ori_n1098_), .C(ori_ori_n877_), .Y(ori_ori_n1963_));
  OAI210     o1914(.A0(ori_ori_n1378_), .A1(ori_ori_n1697_), .B0(ori_ori_n1963_), .Y(ori_ori_n1964_));
  OAI210     o1915(.A0(ori_ori_n1964_), .A1(ori_ori_n1961_), .B0(ori_ori_n1139_), .Y(ori_ori_n1965_));
  OAI210     o1916(.A0(ori_ori_n445_), .A1(ori_ori_n51_), .B0(ori_ori_n1030_), .Y(ori_ori_n1966_));
  AOI220     o1917(.A0(ori_ori_n1966_), .A1(ori_ori_n462_), .B0(ori_ori_n445_), .B1(ori_ori_n386_), .Y(ori_ori_n1967_));
  NO2        o1918(.A(ori_ori_n1967_), .B(ori_ori_n149_), .Y(ori_ori_n1968_));
  OAI220     o1919(.A0(ori_ori_n690_), .A1(ori_ori_n258_), .B0(ori_ori_n686_), .B1(x6), .Y(ori_ori_n1969_));
  NO2        o1920(.A(ori_ori_n299_), .B(x4), .Y(ori_ori_n1970_));
  AOI220     o1921(.A0(ori_ori_n1970_), .A1(ori_ori_n361_), .B0(ori_ori_n1969_), .B1(x4), .Y(ori_ori_n1971_));
  NO3        o1922(.A(ori_ori_n1971_), .B(ori_ori_n320_), .C(x5), .Y(ori_ori_n1972_));
  NO2        o1923(.A(ori_ori_n710_), .B(ori_ori_n57_), .Y(ori_ori_n1973_));
  NA2        o1924(.A(ori_ori_n1973_), .B(ori_ori_n447_), .Y(ori_ori_n1974_));
  AOI220     o1925(.A0(ori_ori_n667_), .A1(ori_ori_n740_), .B0(ori_ori_n494_), .B1(ori_ori_n233_), .Y(ori_ori_n1975_));
  AOI210     o1926(.A0(ori_ori_n1975_), .A1(ori_ori_n1974_), .B0(ori_ori_n253_), .Y(ori_ori_n1976_));
  NO4        o1927(.A(ori_ori_n1976_), .B(ori_ori_n1972_), .C(x1), .D(ori_ori_n1968_), .Y(ori_ori_n1977_));
  AOI220     o1928(.A0(ori_ori_n1977_), .A1(ori_ori_n1965_), .B0(ori_ori_n1957_), .B1(ori_ori_n1947_), .Y(ori_ori_n1978_));
  AOI210     o1929(.A0(ori_ori_n1935_), .A1(x3), .B0(ori_ori_n1978_), .Y(ori29));
  OAI210     o1930(.A0(ori_ori_n557_), .A1(ori_ori_n259_), .B0(ori_ori_n735_), .Y(ori_ori_n1980_));
  NA2        o1931(.A(ori_ori_n756_), .B(ori_ori_n1060_), .Y(ori_ori_n1981_));
  AO210      o1932(.A0(ori_ori_n1178_), .A1(ori_ori_n1187_), .B0(ori_ori_n1981_), .Y(ori_ori_n1982_));
  AOI210     o1933(.A0(ori_ori_n177_), .A1(ori_ori_n162_), .B0(ori_ori_n710_), .Y(ori_ori_n1983_));
  AOI210     o1934(.A0(ori_ori_n1439_), .A1(ori_ori_n78_), .B0(ori_ori_n1983_), .Y(ori_ori_n1984_));
  NA3        o1935(.A(ori_ori_n1984_), .B(ori_ori_n1982_), .C(ori_ori_n1980_), .Y(ori_ori_n1985_));
  NO3        o1936(.A(ori_ori_n669_), .B(ori_ori_n1161_), .C(ori_ori_n50_), .Y(ori_ori_n1986_));
  NO3        o1937(.A(ori_ori_n1986_), .B(ori_ori_n1266_), .C(ori_ori_n557_), .Y(ori_ori_n1987_));
  NO2        o1938(.A(ori_ori_n443_), .B(ori_ori_n58_), .Y(ori_ori_n1988_));
  AOI220     o1939(.A0(ori_ori_n1988_), .A1(ori_ori_n1225_), .B0(ori_ori_n674_), .B1(ori_ori_n1396_), .Y(ori_ori_n1989_));
  OAI210     o1940(.A0(ori_ori_n1987_), .A1(ori_ori_n543_), .B0(ori_ori_n1989_), .Y(ori_ori_n1990_));
  AOI210     o1941(.A0(ori_ori_n1985_), .A1(x6), .B0(ori_ori_n1990_), .Y(ori_ori_n1991_));
  OAI210     o1942(.A0(x8), .A1(x4), .B0(x5), .Y(ori_ori_n1992_));
  NA2        o1943(.A(ori_ori_n1992_), .B(ori_ori_n108_), .Y(ori_ori_n1993_));
  NA2        o1944(.A(ori_ori_n299_), .B(ori_ori_n142_), .Y(ori_ori_n1994_));
  NA4        o1945(.A(ori_ori_n1994_), .B(ori_ori_n1993_), .C(ori_ori_n668_), .D(ori_ori_n64_), .Y(ori_ori_n1995_));
  AOI210     o1946(.A0(ori_ori_n1336_), .A1(ori_ori_n268_), .B0(ori_ori_n1748_), .Y(ori_ori_n1996_));
  AOI210     o1947(.A0(ori_ori_n1996_), .A1(ori_ori_n1995_), .B0(ori_ori_n897_), .Y(ori_ori_n1997_));
  NA4        o1948(.A(ori_ori_n669_), .B(ori_ori_n304_), .C(ori_ori_n177_), .D(ori_ori_n162_), .Y(ori_ori_n1998_));
  NA3        o1949(.A(ori_ori_n633_), .B(ori_ori_n292_), .C(ori_ori_n809_), .Y(ori_ori_n1999_));
  AOI210     o1950(.A0(ori_ori_n1999_), .A1(ori_ori_n1998_), .B0(ori_ori_n1225_), .Y(ori_ori_n2000_));
  OAI210     o1951(.A0(ori_ori_n904_), .A1(x8), .B0(x7), .Y(ori_ori_n2001_));
  NO2        o1952(.A(ori_ori_n2001_), .B(ori_ori_n123_), .Y(ori_ori_n2002_));
  OA210      o1953(.A0(ori_ori_n877_), .A1(ori_ori_n271_), .B0(ori_ori_n1992_), .Y(ori_ori_n2003_));
  OAI220     o1954(.A0(ori_ori_n2003_), .A1(ori_ori_n589_), .B0(ori_ori_n1527_), .B1(ori_ori_n394_), .Y(ori_ori_n2004_));
  NO4        o1955(.A(ori_ori_n2004_), .B(ori_ori_n2002_), .C(ori_ori_n2000_), .D(ori_ori_n1997_), .Y(ori_ori_n2005_));
  OAI210     o1956(.A0(ori_ori_n1991_), .A1(x2), .B0(ori_ori_n2005_), .Y(ori_ori_n2006_));
  NA3        o1957(.A(x6), .B(ori_ori_n50_), .C(x2), .Y(ori_ori_n2007_));
  OAI210     o1958(.A0(ori_ori_n1244_), .A1(ori_ori_n351_), .B0(ori_ori_n2007_), .Y(ori_ori_n2008_));
  NO3        o1959(.A(ori_ori_n445_), .B(x3), .C(x0), .Y(ori_ori_n2009_));
  AO220      o1960(.A0(ori_ori_n2009_), .A1(x5), .B0(ori_ori_n1942_), .B1(ori_ori_n81_), .Y(ori_ori_n2010_));
  AOI210     o1961(.A0(ori_ori_n2008_), .A1(ori_ori_n341_), .B0(ori_ori_n2010_), .Y(ori_ori_n2011_));
  NO3        o1962(.A(ori_ori_n703_), .B(ori_ori_n362_), .C(ori_ori_n136_), .Y(ori_ori_n2012_));
  AOI210     o1963(.A0(ori_ori_n734_), .A1(ori_ori_n616_), .B0(ori_ori_n2012_), .Y(ori_ori_n2013_));
  OAI210     o1964(.A0(ori_ori_n2011_), .A1(x7), .B0(ori_ori_n2013_), .Y(ori_ori_n2014_));
  AOI210     o1965(.A0(ori_ori_n1108_), .A1(ori_ori_n399_), .B0(ori_ori_n1423_), .Y(ori_ori_n2015_));
  NO2        o1966(.A(ori_ori_n142_), .B(x2), .Y(ori_ori_n2016_));
  OA210      o1967(.A0(ori_ori_n2016_), .A1(ori_ori_n631_), .B0(ori_ori_n669_), .Y(ori_ori_n2017_));
  OAI210     o1968(.A0(ori_ori_n2017_), .A1(ori_ori_n2015_), .B0(ori_ori_n68_), .Y(ori_ori_n2018_));
  NO2        o1969(.A(ori_ori_n193_), .B(ori_ori_n85_), .Y(ori_ori_n2019_));
  OAI210     o1970(.A0(ori_ori_n2019_), .A1(ori_ori_n795_), .B0(ori_ori_n1117_), .Y(ori_ori_n2020_));
  NA3        o1971(.A(ori_ori_n1959_), .B(ori_ori_n226_), .C(ori_ori_n83_), .Y(ori_ori_n2021_));
  NA3        o1972(.A(ori_ori_n2021_), .B(ori_ori_n2020_), .C(ori_ori_n2018_), .Y(ori_ori_n2022_));
  AOI210     o1973(.A0(ori_ori_n2014_), .A1(x8), .B0(ori_ori_n2022_), .Y(ori_ori_n2023_));
  OAI210     o1974(.A0(ori_ori_n443_), .A1(ori_ori_n242_), .B0(ori_ori_n974_), .Y(ori_ori_n2024_));
  OAI210     o1975(.A0(ori_ori_n2024_), .A1(ori_ori_n1140_), .B0(ori_ori_n679_), .Y(ori_ori_n2025_));
  NO3        o1976(.A(ori_ori_n1034_), .B(ori_ori_n352_), .C(ori_ori_n143_), .Y(ori_ori_n2026_));
  NA3        o1977(.A(ori_ori_n2026_), .B(ori_ori_n1318_), .C(ori_ori_n50_), .Y(ori_ori_n2027_));
  NO2        o1978(.A(ori_ori_n129_), .B(ori_ori_n91_), .Y(ori_ori_n2028_));
  AOI220     o1979(.A0(ori_ori_n2028_), .A1(ori_ori_n590_), .B0(ori_ori_n1941_), .B1(ori_ori_n358_), .Y(ori_ori_n2029_));
  NOi31      o1980(.An(ori_ori_n1141_), .B(ori_ori_n1893_), .C(ori_ori_n626_), .Y(ori_ori_n2030_));
  NA2        o1981(.A(ori_ori_n168_), .B(x4), .Y(ori_ori_n2031_));
  NO3        o1982(.A(ori_ori_n1500_), .B(ori_ori_n237_), .C(ori_ori_n71_), .Y(ori_ori_n2032_));
  AOI210     o1983(.A0(ori_ori_n2032_), .A1(ori_ori_n2031_), .B0(ori_ori_n2030_), .Y(ori_ori_n2033_));
  NA4        o1984(.A(ori_ori_n2033_), .B(ori_ori_n2029_), .C(ori_ori_n2027_), .D(ori_ori_n2025_), .Y(ori_ori_n2034_));
  NO4        o1985(.A(ori_ori_n1244_), .B(ori_ori_n166_), .C(ori_ori_n55_), .D(ori_ori_n71_), .Y(ori_ori_n2035_));
  NO4        o1986(.A(ori_ori_n1218_), .B(ori_ori_n503_), .C(ori_ori_n1396_), .D(ori_ori_n104_), .Y(ori_ori_n2036_));
  OAI210     o1987(.A0(ori_ori_n2036_), .A1(ori_ori_n2035_), .B0(ori_ori_n106_), .Y(ori_ori_n2037_));
  AOI210     o1988(.A0(ori_ori_n303_), .A1(x4), .B0(ori_ori_n187_), .Y(ori_ori_n2038_));
  OAI210     o1989(.A0(ori_ori_n2038_), .A1(ori_ori_n1988_), .B0(ori_ori_n729_), .Y(ori_ori_n2039_));
  OR3        o1990(.A(ori_ori_n1769_), .B(ori_ori_n1450_), .C(ori_ori_n1100_), .Y(ori_ori_n2040_));
  NA2        o1991(.A(ori_ori_n1942_), .B(ori_ori_n816_), .Y(ori_ori_n2041_));
  OA220      o1992(.A0(ori_ori_n2041_), .A1(ori_ori_n242_), .B0(ori_ori_n582_), .B1(ori_ori_n1809_), .Y(ori_ori_n2042_));
  NA4        o1993(.A(ori_ori_n2042_), .B(ori_ori_n2040_), .C(ori_ori_n2039_), .D(ori_ori_n2037_), .Y(ori_ori_n2043_));
  AOI210     o1994(.A0(ori_ori_n2034_), .A1(ori_ori_n288_), .B0(ori_ori_n2043_), .Y(ori_ori_n2044_));
  OAI210     o1995(.A0(ori_ori_n2023_), .A1(x1), .B0(ori_ori_n2044_), .Y(ori_ori_n2045_));
  AO210      o1996(.A0(ori_ori_n2006_), .A1(x1), .B0(ori_ori_n2045_), .Y(ori30));
  NO3        o1997(.A(ori_ori_n1793_), .B(ori_ori_n578_), .C(ori_ori_n95_), .Y(ori_ori_n2047_));
  NO3        o1998(.A(ori_ori_n1159_), .B(ori_ori_n132_), .C(ori_ori_n382_), .Y(ori_ori_n2048_));
  AOI210     o1999(.A0(ori_ori_n729_), .A1(ori_ori_n250_), .B0(ori_ori_n2048_), .Y(ori_ori_n2049_));
  AOI210     o2000(.A0(ori_ori_n2049_), .A1(ori_ori_n2047_), .B0(ori_ori_n56_), .Y(ori_ori_n2050_));
  NA2        o2001(.A(ori_ori_n821_), .B(ori_ori_n339_), .Y(ori_ori_n2051_));
  NA2        o2002(.A(ori_ori_n2051_), .B(ori_ori_n1379_), .Y(ori_ori_n2052_));
  OAI210     o2003(.A0(ori_ori_n2052_), .A1(ori_ori_n2050_), .B0(ori_ori_n106_), .Y(ori_ori_n2053_));
  OAI210     o2004(.A0(ori_ori_n1011_), .A1(ori_ori_n572_), .B0(ori_ori_n679_), .Y(ori_ori_n2054_));
  AOI220     o2005(.A0(ori_ori_n448_), .A1(ori_ori_n950_), .B0(ori_ori_n325_), .B1(ori_ori_n456_), .Y(ori_ori_n2055_));
  AOI210     o2006(.A0(ori_ori_n2055_), .A1(ori_ori_n2054_), .B0(ori_ori_n253_), .Y(ori_ori_n2056_));
  NO3        o2007(.A(ori_ori_n277_), .B(ori_ori_n120_), .C(x0), .Y(ori_ori_n2057_));
  AOI210     o2008(.A0(ori_ori_n505_), .A1(x6), .B0(ori_ori_n2057_), .Y(ori_ori_n2058_));
  AOI220     o2009(.A0(ori_ori_n1155_), .A1(ori_ori_n423_), .B0(ori_ori_n768_), .B1(ori_ori_n90_), .Y(ori_ori_n2059_));
  OAI220     o2010(.A0(ori_ori_n2059_), .A1(ori_ori_n242_), .B0(ori_ori_n2058_), .B1(ori_ori_n54_), .Y(ori_ori_n2060_));
  NA3        o2011(.A(ori_ori_n321_), .B(ori_ori_n159_), .C(ori_ori_n71_), .Y(ori_ori_n2061_));
  AO210      o2012(.A0(ori_ori_n571_), .A1(ori_ori_n519_), .B0(x5), .Y(ori_ori_n2062_));
  AOI210     o2013(.A0(ori_ori_n2061_), .A1(ori_ori_n726_), .B0(ori_ori_n2062_), .Y(ori_ori_n2063_));
  AOI210     o2014(.A0(ori_ori_n1625_), .A1(ori_ori_n50_), .B0(ori_ori_n456_), .Y(ori_ori_n2064_));
  NA2        o2015(.A(ori_ori_n192_), .B(x2), .Y(ori_ori_n2065_));
  OA220      o2016(.A0(ori_ori_n2065_), .A1(ori_ori_n2064_), .B0(ori_ori_n272_), .B1(x6), .Y(ori_ori_n2066_));
  OAI210     o2017(.A0(x7), .A1(x6), .B0(x1), .Y(ori_ori_n2067_));
  NA3        o2018(.A(ori_ori_n57_), .B(x4), .C(ori_ori_n59_), .Y(ori_ori_n2068_));
  AOI220     o2019(.A0(ori_ori_n2068_), .A1(ori_ori_n1386_), .B0(ori_ori_n2067_), .B1(ori_ori_n1834_), .Y(ori_ori_n2069_));
  NO3        o2020(.A(ori_ori_n1382_), .B(ori_ori_n341_), .C(ori_ori_n1036_), .Y(ori_ori_n2070_));
  NO2        o2021(.A(ori_ori_n517_), .B(ori_ori_n870_), .Y(ori_ori_n2071_));
  NOi21      o2022(.An(ori_ori_n2071_), .B(ori_ori_n855_), .Y(ori_ori_n2072_));
  NO3        o2023(.A(ori_ori_n1318_), .B(ori_ori_n228_), .C(ori_ori_n651_), .Y(ori_ori_n2073_));
  NO4        o2024(.A(ori_ori_n2073_), .B(ori_ori_n2072_), .C(ori_ori_n2070_), .D(ori_ori_n2069_), .Y(ori_ori_n2074_));
  OAI210     o2025(.A0(ori_ori_n2066_), .A1(ori_ori_n763_), .B0(ori_ori_n2074_), .Y(ori_ori_n2075_));
  NO4        o2026(.A(ori_ori_n2075_), .B(ori_ori_n2063_), .C(ori_ori_n2060_), .D(ori_ori_n2056_), .Y(ori_ori_n2076_));
  AOI210     o2027(.A0(ori_ori_n2076_), .A1(ori_ori_n2053_), .B0(x8), .Y(ori_ori_n2077_));
  NO3        o2028(.A(ori_ori_n492_), .B(ori_ori_n792_), .C(ori_ori_n53_), .Y(ori_ori_n2078_));
  OAI220     o2029(.A0(ori_ori_n1809_), .A1(ori_ori_n341_), .B0(ori_ori_n484_), .B1(ori_ori_n586_), .Y(ori_ori_n2079_));
  OAI210     o2030(.A0(ori_ori_n2079_), .A1(ori_ori_n2078_), .B0(x6), .Y(ori_ori_n2080_));
  OAI210     o2031(.A0(ori_ori_n1051_), .A1(ori_ori_n538_), .B0(ori_ori_n821_), .Y(ori_ori_n2081_));
  OAI210     o2032(.A0(ori_ori_n1758_), .A1(ori_ori_n328_), .B0(ori_ori_n122_), .Y(ori_ori_n2082_));
  AOI210     o2033(.A0(ori_ori_n377_), .A1(ori_ori_n225_), .B0(ori_ori_n72_), .Y(ori_ori_n2083_));
  AOI210     o2034(.A0(ori_ori_n1011_), .A1(ori_ori_n754_), .B0(ori_ori_n2083_), .Y(ori_ori_n2084_));
  NA4        o2035(.A(ori_ori_n2084_), .B(ori_ori_n2082_), .C(ori_ori_n2081_), .D(ori_ori_n2080_), .Y(ori_ori_n2085_));
  NA2        o2036(.A(ori_ori_n1105_), .B(ori_ori_n59_), .Y(ori_ori_n2086_));
  AOI210     o2037(.A0(ori_ori_n931_), .A1(ori_ori_n493_), .B0(ori_ori_n685_), .Y(ori_ori_n2087_));
  OAI220     o2038(.A0(ori_ori_n2087_), .A1(ori_ori_n303_), .B0(ori_ori_n2086_), .B1(ori_ori_n483_), .Y(ori_ori_n2088_));
  AOI210     o2039(.A0(ori_ori_n2085_), .A1(x8), .B0(ori_ori_n2088_), .Y(ori_ori_n2089_));
  NO2        o2040(.A(ori_ori_n2089_), .B(ori_ori_n57_), .Y(ori_ori_n2090_));
  NA2        o2041(.A(ori_ori_n434_), .B(ori_ori_n855_), .Y(ori_ori_n2091_));
  NO2        o2042(.A(ori_ori_n930_), .B(ori_ori_n665_), .Y(ori_ori_n2092_));
  AOI210     o2043(.A0(ori_ori_n2092_), .A1(ori_ori_n2091_), .B0(ori_ori_n445_), .Y(ori_ori_n2093_));
  NO3        o2044(.A(ori_ori_n639_), .B(ori_ori_n408_), .C(ori_ori_n1159_), .Y(ori_ori_n2094_));
  NO3        o2045(.A(ori_ori_n2094_), .B(ori_ori_n1272_), .C(ori_ori_n1396_), .Y(ori_ori_n2095_));
  AOI210     o2046(.A0(ori_ori_n300_), .A1(x1), .B0(ori_ori_n143_), .Y(ori_ori_n2096_));
  NO2        o2047(.A(ori_ori_n306_), .B(x5), .Y(ori_ori_n2097_));
  NO2        o2048(.A(ori_ori_n2097_), .B(ori_ori_n863_), .Y(ori_ori_n2098_));
  OAI220     o2049(.A0(ori_ori_n2098_), .A1(ori_ori_n1071_), .B0(ori_ori_n2096_), .B1(ori_ori_n202_), .Y(ori_ori_n2099_));
  NO3        o2050(.A(ori_ori_n2099_), .B(ori_ori_n2095_), .C(ori_ori_n2093_), .Y(ori_ori_n2100_));
  NA2        o2051(.A(ori_ori_n972_), .B(ori_ori_n82_), .Y(ori_ori_n2101_));
  AO210      o2052(.A0(ori_ori_n2101_), .A1(ori_ori_n1626_), .B0(x3), .Y(ori_ori_n2102_));
  NO2        o2053(.A(ori_ori_n214_), .B(ori_ori_n56_), .Y(ori_ori_n2103_));
  OAI220     o2054(.A0(ori_ori_n377_), .A1(ori_ori_n1272_), .B0(ori_ori_n352_), .B1(ori_ori_n228_), .Y(ori_ori_n2104_));
  AOI220     o2055(.A0(ori_ori_n2104_), .A1(x2), .B0(ori_ori_n2103_), .B1(ori_ori_n1640_), .Y(ori_ori_n2105_));
  AOI210     o2056(.A0(ori_ori_n2105_), .A1(ori_ori_n2102_), .B0(ori_ori_n258_), .Y(ori_ori_n2106_));
  NO2        o2057(.A(ori_ori_n300_), .B(ori_ori_n119_), .Y(ori_ori_n2107_));
  NO3        o2058(.A(ori_ori_n826_), .B(ori_ori_n704_), .C(ori_ori_n162_), .Y(ori_ori_n2108_));
  OAI210     o2059(.A0(ori_ori_n2108_), .A1(ori_ori_n2107_), .B0(ori_ori_n150_), .Y(ori_ori_n2109_));
  NA3        o2060(.A(x5), .B(x4), .C(ori_ori_n59_), .Y(ori_ori_n2110_));
  AOI210     o2061(.A0(ori_ori_n2110_), .A1(ori_ori_n1324_), .B0(ori_ori_n539_), .Y(ori_ori_n2111_));
  AOI210     o2062(.A0(ori_ori_n1344_), .A1(x2), .B0(ori_ori_n2111_), .Y(ori_ori_n2112_));
  AOI210     o2063(.A0(ori_ori_n2112_), .A1(ori_ori_n2109_), .B0(ori_ori_n50_), .Y(ori_ori_n2113_));
  NA3        o2064(.A(ori_ori_n1497_), .B(ori_ori_n1150_), .C(ori_ori_n476_), .Y(ori_ori_n2114_));
  AOI210     o2065(.A0(ori_ori_n2114_), .A1(ori_ori_n2101_), .B0(ori_ori_n612_), .Y(ori_ori_n2115_));
  AOI210     o2066(.A0(ori_ori_n1036_), .A1(x1), .B0(ori_ori_n1336_), .Y(ori_ori_n2116_));
  OAI220     o2067(.A0(ori_ori_n304_), .A1(x4), .B0(ori_ori_n51_), .B1(x6), .Y(ori_ori_n2117_));
  NO2        o2068(.A(ori_ori_n118_), .B(ori_ori_n108_), .Y(ori_ori_n2118_));
  AOI220     o2069(.A0(ori_ori_n2118_), .A1(ori_ori_n2117_), .B0(ori_ori_n1180_), .B1(ori_ori_n626_), .Y(ori_ori_n2119_));
  OAI210     o2070(.A0(ori_ori_n2116_), .A1(ori_ori_n487_), .B0(ori_ori_n2119_), .Y(ori_ori_n2120_));
  NO4        o2071(.A(ori_ori_n2120_), .B(ori_ori_n2115_), .C(ori_ori_n2113_), .D(ori_ori_n2106_), .Y(ori_ori_n2121_));
  OAI210     o2072(.A0(ori_ori_n2100_), .A1(ori_ori_n129_), .B0(ori_ori_n2121_), .Y(ori_ori_n2122_));
  NO3        o2073(.A(ori_ori_n2122_), .B(ori_ori_n2090_), .C(ori_ori_n2077_), .Y(ori31));
  NA2        o2074(.A(ori_ori_n996_), .B(ori_ori_n353_), .Y(ori_ori_n2124_));
  NO2        o2075(.A(ori_ori_n449_), .B(ori_ori_n679_), .Y(ori_ori_n2125_));
  AOI210     o2076(.A0(ori_ori_n2125_), .A1(ori_ori_n2124_), .B0(ori_ori_n58_), .Y(ori_ori_n2126_));
  NO2        o2077(.A(ori_ori_n794_), .B(ori_ori_n56_), .Y(ori_ori_n2127_));
  AOI220     o2078(.A0(ori_ori_n2127_), .A1(x2), .B0(ori_ori_n89_), .B1(x0), .Y(ori_ori_n2128_));
  NA3        o2079(.A(ori_ori_n2128_), .B(ori_ori_n2041_), .C(ori_ori_n1871_), .Y(ori_ori_n2129_));
  OAI210     o2080(.A0(ori_ori_n2129_), .A1(ori_ori_n2126_), .B0(ori_ori_n53_), .Y(ori_ori_n2130_));
  INV        o2081(.A(ori_ori_n679_), .Y(ori_ori_n2131_));
  NO3        o2082(.A(ori_ori_n1970_), .B(ori_ori_n1942_), .C(ori_ori_n898_), .Y(ori_ori_n2132_));
  OA220      o2083(.A0(ori_ori_n2132_), .A1(ori_ori_n476_), .B0(ori_ori_n2131_), .B1(ori_ori_n1490_), .Y(ori_ori_n2133_));
  AOI210     o2084(.A0(ori_ori_n2133_), .A1(ori_ori_n2130_), .B0(ori_ori_n104_), .Y(ori_ori_n2134_));
  NO2        o2085(.A(ori_ori_n499_), .B(ori_ori_n75_), .Y(ori_ori_n2135_));
  NA2        o2086(.A(ori_ori_n445_), .B(ori_ori_n57_), .Y(ori_ori_n2136_));
  AOI210     o2087(.A0(ori_ori_n303_), .A1(ori_ori_n86_), .B0(ori_ori_n2136_), .Y(ori_ori_n2137_));
  OAI210     o2088(.A0(ori_ori_n2137_), .A1(ori_ori_n2135_), .B0(ori_ori_n779_), .Y(ori_ori_n2138_));
  NO4        o2089(.A(ori_ori_n1176_), .B(ori_ori_n362_), .C(ori_ori_n1625_), .D(ori_ori_n67_), .Y(ori_ori_n2139_));
  AOI210     o2090(.A0(ori_ori_n1664_), .A1(ori_ori_n1371_), .B0(ori_ori_n443_), .Y(ori_ori_n2140_));
  OAI220     o2091(.A0(ori_ori_n1325_), .A1(ori_ori_n964_), .B0(ori_ori_n781_), .B1(ori_ori_n113_), .Y(ori_ori_n2141_));
  NO3        o2092(.A(ori_ori_n2141_), .B(ori_ori_n2140_), .C(ori_ori_n2139_), .Y(ori_ori_n2142_));
  AOI210     o2093(.A0(ori_ori_n2142_), .A1(ori_ori_n2138_), .B0(x5), .Y(ori_ori_n2143_));
  AOI220     o2094(.A0(ori_ori_n447_), .A1(ori_ori_n626_), .B0(ori_ori_n572_), .B1(ori_ori_n63_), .Y(ori_ori_n2144_));
  AOI210     o2095(.A0(ori_ori_n2144_), .A1(ori_ori_n582_), .B0(ori_ori_n1244_), .Y(ori_ori_n2145_));
  AOI220     o2096(.A0(ori_ori_n973_), .A1(ori_ori_n740_), .B0(ori_ori_n1159_), .B1(ori_ori_n117_), .Y(ori_ori_n2146_));
  OAI220     o2097(.A0(ori_ori_n2146_), .A1(ori_ori_n385_), .B0(ori_ori_n483_), .B1(ori_ori_n780_), .Y(ori_ori_n2147_));
  NO4        o2098(.A(ori_ori_n2147_), .B(ori_ori_n2145_), .C(ori_ori_n2143_), .D(ori_ori_n2134_), .Y(ori_ori_n2148_));
  NA2        o2099(.A(ori_ori_n493_), .B(ori_ori_n59_), .Y(ori_ori_n2149_));
  AOI210     o2100(.A0(ori_ori_n543_), .A1(ori_ori_n2149_), .B0(ori_ori_n135_), .Y(ori_ori_n2150_));
  OAI210     o2101(.A0(ori_ori_n100_), .A1(ori_ori_n271_), .B0(ori_ori_n2086_), .Y(ori_ori_n2151_));
  OAI210     o2102(.A0(ori_ori_n2151_), .A1(ori_ori_n2150_), .B0(x7), .Y(ori_ori_n2152_));
  NO3        o2103(.A(ori_ori_n377_), .B(ori_ori_n55_), .C(x7), .Y(ori_ori_n2153_));
  OA210      o2104(.A0(ori_ori_n2153_), .A1(ori_ori_n1335_), .B0(ori_ori_n97_), .Y(ori_ori_n2154_));
  NA2        o2105(.A(ori_ori_n1102_), .B(ori_ori_n90_), .Y(ori_ori_n2155_));
  AOI210     o2106(.A0(ori_ori_n910_), .A1(ori_ori_n108_), .B0(ori_ori_n2155_), .Y(ori_ori_n2156_));
  NA2        o2107(.A(ori_ori_n1572_), .B(x6), .Y(ori_ori_n2157_));
  AOI210     o2108(.A0(ori_ori_n2157_), .A1(ori_ori_n287_), .B0(ori_ori_n104_), .Y(ori_ori_n2158_));
  NA2        o2109(.A(ori_ori_n1203_), .B(ori_ori_n316_), .Y(ori_ori_n2159_));
  AOI210     o2110(.A0(ori_ori_n2159_), .A1(ori_ori_n647_), .B0(ori_ori_n53_), .Y(ori_ori_n2160_));
  NO4        o2111(.A(ori_ori_n2160_), .B(ori_ori_n2158_), .C(ori_ori_n2156_), .D(ori_ori_n2154_), .Y(ori_ori_n2161_));
  AOI210     o2112(.A0(ori_ori_n2161_), .A1(ori_ori_n2152_), .B0(ori_ori_n689_), .Y(ori_ori_n2162_));
  NOi21      o2113(.An(ori_ori_n1783_), .B(ori_ori_n1075_), .Y(ori_ori_n2163_));
  OAI220     o2114(.A0(ori_ori_n2163_), .A1(ori_ori_n1944_), .B0(ori_ori_n932_), .B1(ori_ori_n2149_), .Y(ori_ori_n2164_));
  NA2        o2115(.A(ori_ori_n2164_), .B(x3), .Y(ori_ori_n2165_));
  AOI220     o2116(.A0(ori_ori_n1406_), .A1(x8), .B0(ori_ori_n60_), .B1(x1), .Y(ori_ori_n2166_));
  NO3        o2117(.A(ori_ori_n2166_), .B(ori_ori_n1129_), .C(x6), .Y(ori_ori_n2167_));
  AOI220     o2118(.A0(ori_ori_n616_), .A1(ori_ori_n408_), .B0(ori_ori_n493_), .B1(ori_ori_n78_), .Y(ori_ori_n2168_));
  NA2        o2119(.A(ori_ori_n114_), .B(ori_ori_n530_), .Y(ori_ori_n2169_));
  OAI220     o2120(.A0(ori_ori_n2169_), .A1(ori_ori_n1944_), .B0(ori_ori_n2168_), .B1(x4), .Y(ori_ori_n2170_));
  NO2        o2121(.A(ori_ori_n2170_), .B(ori_ori_n2167_), .Y(ori_ori_n2171_));
  AOI210     o2122(.A0(ori_ori_n2171_), .A1(ori_ori_n2165_), .B0(ori_ori_n180_), .Y(ori_ori_n2172_));
  NO4        o2123(.A(ori_ori_n617_), .B(ori_ori_n590_), .C(ori_ori_n705_), .D(ori_ori_n704_), .Y(ori_ori_n2173_));
  OAI210     o2124(.A0(ori_ori_n2173_), .A1(ori_ori_n1093_), .B0(x3), .Y(ori_ori_n2174_));
  NO4        o2125(.A(ori_ori_n812_), .B(ori_ori_n1244_), .C(ori_ori_n779_), .D(x5), .Y(ori_ori_n2175_));
  NO3        o2126(.A(x6), .B(ori_ori_n56_), .C(x1), .Y(ori_ori_n2176_));
  NA2        o2127(.A(ori_ori_n2176_), .B(ori_ori_n283_), .Y(ori_ori_n2177_));
  OAI210     o2128(.A0(ori_ori_n1916_), .A1(ori_ori_n377_), .B0(ori_ori_n2177_), .Y(ori_ori_n2178_));
  NA4        o2129(.A(ori_ori_n639_), .B(ori_ori_n173_), .C(x6), .D(ori_ori_n104_), .Y(ori_ori_n2179_));
  NO2        o2130(.A(ori_ori_n864_), .B(ori_ori_n246_), .Y(ori_ori_n2180_));
  NOi41      o2131(.An(ori_ori_n2179_), .B(ori_ori_n2180_), .C(ori_ori_n2178_), .D(ori_ori_n2175_), .Y(ori_ori_n2181_));
  AOI210     o2132(.A0(ori_ori_n2181_), .A1(ori_ori_n2174_), .B0(ori_ori_n534_), .Y(ori_ori_n2182_));
  OAI210     o2133(.A0(ori_ori_n616_), .A1(ori_ori_n470_), .B0(ori_ori_n950_), .Y(ori_ori_n2183_));
  NO3        o2134(.A(ori_ori_n372_), .B(ori_ori_n77_), .C(ori_ori_n53_), .Y(ori_ori_n2184_));
  NO3        o2135(.A(ori_ori_n462_), .B(ori_ori_n347_), .C(ori_ori_n50_), .Y(ori_ori_n2185_));
  OAI210     o2136(.A0(ori_ori_n2185_), .A1(ori_ori_n2184_), .B0(ori_ori_n1177_), .Y(ori_ori_n2186_));
  AOI210     o2137(.A0(ori_ori_n2186_), .A1(ori_ori_n2183_), .B0(ori_ori_n392_), .Y(ori_ori_n2187_));
  NO2        o2138(.A(ori_ori_n211_), .B(ori_ori_n539_), .Y(ori_ori_n2188_));
  OAI210     o2139(.A0(ori_ori_n132_), .A1(x2), .B0(ori_ori_n2188_), .Y(ori_ori_n2189_));
  NA3        o2140(.A(ori_ori_n408_), .B(ori_ori_n326_), .C(ori_ori_n77_), .Y(ori_ori_n2190_));
  OA210      o2141(.A0(ori_ori_n241_), .A1(ori_ori_n224_), .B0(ori_ori_n2190_), .Y(ori_ori_n2191_));
  AOI210     o2142(.A0(ori_ori_n2191_), .A1(ori_ori_n2189_), .B0(ori_ori_n64_), .Y(ori_ori_n2192_));
  NA2        o2143(.A(ori_ori_n118_), .B(ori_ori_n57_), .Y(ori_ori_n2193_));
  AOI220     o2144(.A0(ori_ori_n1604_), .A1(ori_ori_n916_), .B0(ori_ori_n270_), .B1(x4), .Y(ori_ori_n2194_));
  AOI220     o2145(.A0(ori_ori_n1657_), .A1(ori_ori_n618_), .B0(ori_ori_n727_), .B1(ori_ori_n779_), .Y(ori_ori_n2195_));
  OAI220     o2146(.A0(ori_ori_n2195_), .A1(ori_ori_n2193_), .B0(ori_ori_n2194_), .B1(ori_ori_n185_), .Y(ori_ori_n2196_));
  OR3        o2147(.A(ori_ori_n2196_), .B(ori_ori_n2192_), .C(ori_ori_n2187_), .Y(ori_ori_n2197_));
  NO4        o2148(.A(ori_ori_n2197_), .B(ori_ori_n2182_), .C(ori_ori_n2172_), .D(ori_ori_n2162_), .Y(ori_ori_n2198_));
  OAI210     o2149(.A0(ori_ori_n2148_), .A1(x3), .B0(ori_ori_n2198_), .Y(ori32));
  OAI210     o2150(.A0(ori_ori_n565_), .A1(ori_ori_n53_), .B0(ori_ori_n413_), .Y(ori_ori_n2200_));
  NA2        o2151(.A(ori_ori_n514_), .B(x2), .Y(ori_ori_n2201_));
  AOI210     o2152(.A0(ori_ori_n2201_), .A1(ori_ori_n2200_), .B0(ori_ori_n57_), .Y(ori_ori_n2202_));
  OAI210     o2153(.A0(ori_ori_n2202_), .A1(ori_ori_n795_), .B0(ori_ori_n56_), .Y(ori_ori_n2203_));
  OAI210     o2154(.A0(ori_ori_n1728_), .A1(ori_ori_n1469_), .B0(ori_ori_n1499_), .Y(ori_ori_n2204_));
  AOI210     o2155(.A0(ori_ori_n2127_), .A1(ori_ori_n274_), .B0(ori_ori_n2204_), .Y(ori_ori_n2205_));
  AOI210     o2156(.A0(ori_ori_n2205_), .A1(ori_ori_n2203_), .B0(ori_ori_n50_), .Y(ori_ori_n2206_));
  NA3        o2157(.A(ori_ori_n1573_), .B(ori_ori_n810_), .C(ori_ori_n286_), .Y(ori_ori_n2207_));
  NA2        o2158(.A(ori_ori_n751_), .B(ori_ori_n547_), .Y(ori_ori_n2208_));
  OAI220     o2159(.A0(ori_ori_n1070_), .A1(ori_ori_n226_), .B0(ori_ori_n686_), .B1(ori_ori_n202_), .Y(ori_ori_n2209_));
  NO3        o2160(.A(ori_ori_n373_), .B(ori_ori_n575_), .C(ori_ori_n816_), .Y(ori_ori_n2210_));
  NO3        o2161(.A(ori_ori_n1382_), .B(ori_ori_n586_), .C(ori_ori_n268_), .Y(ori_ori_n2211_));
  NO4        o2162(.A(ori_ori_n2211_), .B(ori_ori_n2210_), .C(ori_ori_n2209_), .D(ori_ori_n2208_), .Y(ori_ori_n2212_));
  AOI210     o2163(.A0(ori_ori_n2212_), .A1(ori_ori_n2207_), .B0(ori_ori_n136_), .Y(ori_ori_n2213_));
  OAI220     o2164(.A0(ori_ori_n401_), .A1(x7), .B0(ori_ori_n299_), .B1(ori_ori_n292_), .Y(ori_ori_n2214_));
  NA2        o2165(.A(ori_ori_n2214_), .B(ori_ori_n972_), .Y(ori_ori_n2215_));
  NO2        o2166(.A(ori_ori_n552_), .B(ori_ori_n870_), .Y(ori_ori_n2216_));
  AOI220     o2167(.A0(ori_ori_n2216_), .A1(ori_ori_n1896_), .B0(ori_ori_n531_), .B1(ori_ori_n125_), .Y(ori_ori_n2217_));
  AOI210     o2168(.A0(ori_ori_n2217_), .A1(ori_ori_n2215_), .B0(ori_ori_n106_), .Y(ori_ori_n2218_));
  NA3        o2169(.A(ori_ori_n1335_), .B(ori_ori_n1161_), .C(ori_ori_n113_), .Y(ori_ori_n2219_));
  AOI220     o2170(.A0(ori_ori_n1372_), .A1(ori_ori_n705_), .B0(ori_ori_n1258_), .B1(ori_ori_n1058_), .Y(ori_ori_n2220_));
  AOI210     o2171(.A0(ori_ori_n2220_), .A1(ori_ori_n2219_), .B0(ori_ori_n56_), .Y(ori_ori_n2221_));
  NA2        o2172(.A(ori_ori_n972_), .B(ori_ori_n57_), .Y(ori_ori_n2222_));
  NOi21      o2173(.An(ori_ori_n2222_), .B(ori_ori_n125_), .Y(ori_ori_n2223_));
  NA2        o2174(.A(ori_ori_n1026_), .B(ori_ori_n246_), .Y(ori_ori_n2224_));
  NO3        o2175(.A(ori_ori_n2224_), .B(ori_ori_n2223_), .C(ori_ori_n59_), .Y(ori_ori_n2225_));
  OR4        o2176(.A(ori_ori_n2225_), .B(ori_ori_n2221_), .C(ori_ori_n2218_), .D(ori_ori_n2213_), .Y(ori_ori_n2226_));
  OAI210     o2177(.A0(ori_ori_n2226_), .A1(ori_ori_n2206_), .B0(ori_ori_n104_), .Y(ori_ori_n2227_));
  NO3        o2178(.A(ori_ori_n1244_), .B(ori_ori_n140_), .C(ori_ori_n121_), .Y(ori_ori_n2228_));
  NO2        o2179(.A(ori_ori_n380_), .B(ori_ori_n55_), .Y(ori_ori_n2229_));
  NA2        o2180(.A(ori_ori_n2229_), .B(ori_ori_n112_), .Y(ori_ori_n2230_));
  OAI210     o2181(.A0(ori_ori_n635_), .A1(ori_ori_n592_), .B0(ori_ori_n821_), .Y(ori_ori_n2231_));
  NA2        o2182(.A(ori_ori_n2231_), .B(ori_ori_n2230_), .Y(ori_ori_n2232_));
  OAI210     o2183(.A0(ori_ori_n2232_), .A1(ori_ori_n2228_), .B0(x3), .Y(ori_ori_n2233_));
  OAI210     o2184(.A0(ori_ori_n904_), .A1(ori_ori_n268_), .B0(ori_ori_n50_), .Y(ori_ori_n2234_));
  AOI210     o2185(.A0(ori_ori_n62_), .A1(ori_ori_n106_), .B0(ori_ori_n2234_), .Y(ori_ori_n2235_));
  OAI210     o2186(.A0(ori_ori_n2235_), .A1(ori_ori_n1877_), .B0(ori_ori_n704_), .Y(ori_ori_n2236_));
  NO3        o2187(.A(ori_ori_n301_), .B(ori_ori_n168_), .C(ori_ori_n119_), .Y(ori_ori_n2237_));
  NO3        o2188(.A(ori_ori_n810_), .B(ori_ori_n360_), .C(ori_ori_n136_), .Y(ori_ori_n2238_));
  OAI210     o2189(.A0(ori_ori_n2238_), .A1(ori_ori_n2237_), .B0(ori_ori_n59_), .Y(ori_ori_n2239_));
  NA2        o2190(.A(ori_ori_n1165_), .B(ori_ori_n71_), .Y(ori_ori_n2240_));
  NO2        o2191(.A(ori_ori_n1948_), .B(ori_ori_n592_), .Y(ori_ori_n2241_));
  AOI210     o2192(.A0(ori_ori_n2241_), .A1(ori_ori_n1878_), .B0(ori_ori_n2240_), .Y(ori_ori_n2242_));
  NO2        o2193(.A(ori_ori_n271_), .B(ori_ori_n57_), .Y(ori_ori_n2243_));
  NO2        o2194(.A(ori_ori_n2243_), .B(ori_ori_n1018_), .Y(ori_ori_n2244_));
  NOi31      o2195(.An(ori_ori_n729_), .B(ori_ori_n2244_), .C(ori_ori_n277_), .Y(ori_ori_n2245_));
  NO3        o2196(.A(ori_ori_n1327_), .B(ori_ori_n211_), .C(ori_ori_n253_), .Y(ori_ori_n2246_));
  NO4        o2197(.A(ori_ori_n2246_), .B(ori_ori_n2245_), .C(ori_ori_n2242_), .D(x1), .Y(ori_ori_n2247_));
  NA4        o2198(.A(ori_ori_n2247_), .B(ori_ori_n2239_), .C(ori_ori_n2236_), .D(ori_ori_n2233_), .Y(ori_ori_n2248_));
  AO210      o2199(.A0(ori_ori_n1108_), .A1(ori_ori_n396_), .B0(ori_ori_n1021_), .Y(ori_ori_n2249_));
  NA3        o2200(.A(ori_ori_n1922_), .B(ori_ori_n556_), .C(ori_ori_n271_), .Y(ori_ori_n2250_));
  AOI210     o2201(.A0(ori_ori_n2250_), .A1(ori_ori_n2249_), .B0(ori_ori_n301_), .Y(ori_ori_n2251_));
  NA4        o2202(.A(ori_ori_n1281_), .B(ori_ori_n528_), .C(ori_ori_n385_), .D(ori_ori_n226_), .Y(ori_ori_n2252_));
  NO3        o2203(.A(ori_ori_n1450_), .B(ori_ori_n1021_), .C(x2), .Y(ori_ori_n2253_));
  NO2        o2204(.A(ori_ori_n1267_), .B(ori_ori_n383_), .Y(ori_ori_n2254_));
  NO2        o2205(.A(ori_ori_n1852_), .B(ori_ori_n64_), .Y(ori_ori_n2255_));
  NO4        o2206(.A(ori_ori_n2255_), .B(ori_ori_n2254_), .C(ori_ori_n2253_), .D(ori_ori_n53_), .Y(ori_ori_n2256_));
  NO3        o2207(.A(ori_ori_n466_), .B(ori_ori_n1102_), .C(ori_ori_n118_), .Y(ori_ori_n2257_));
  OAI220     o2208(.A0(ori_ori_n689_), .A1(ori_ori_n168_), .B0(ori_ori_n352_), .B1(ori_ori_n136_), .Y(ori_ori_n2258_));
  OAI210     o2209(.A0(ori_ori_n2258_), .A1(ori_ori_n2257_), .B0(ori_ori_n68_), .Y(ori_ori_n2259_));
  NO2        o2210(.A(ori_ori_n1992_), .B(ori_ori_n364_), .Y(ori_ori_n2260_));
  OAI210     o2211(.A0(ori_ori_n1883_), .A1(ori_ori_n610_), .B0(ori_ori_n2260_), .Y(ori_ori_n2261_));
  NA4        o2212(.A(ori_ori_n2261_), .B(ori_ori_n2259_), .C(ori_ori_n2256_), .D(ori_ori_n2252_), .Y(ori_ori_n2262_));
  OAI210     o2213(.A0(ori_ori_n2262_), .A1(ori_ori_n2251_), .B0(ori_ori_n2248_), .Y(ori_ori_n2263_));
  NO3        o2214(.A(ori_ori_n1231_), .B(ori_ori_n103_), .C(ori_ori_n71_), .Y(ori_ori_n2264_));
  NO2        o2215(.A(ori_ori_n565_), .B(ori_ori_n368_), .Y(ori_ori_n2265_));
  OAI210     o2216(.A0(ori_ori_n2264_), .A1(ori_ori_n1429_), .B0(ori_ori_n2265_), .Y(ori_ori_n2266_));
  NO3        o2217(.A(x8), .B(ori_ori_n71_), .C(x2), .Y(ori_ori_n2267_));
  OAI220     o2218(.A0(ori_ori_n2267_), .A1(ori_ori_n626_), .B0(ori_ori_n1439_), .B1(ori_ori_n89_), .Y(ori_ori_n2268_));
  AOI220     o2219(.A0(ori_ori_n557_), .A1(ori_ori_n821_), .B0(ori_ori_n679_), .B1(ori_ori_n251_), .Y(ori_ori_n2269_));
  AOI210     o2220(.A0(ori_ori_n2269_), .A1(ori_ori_n2268_), .B0(ori_ori_n261_), .Y(ori_ori_n2270_));
  NA2        o2221(.A(ori_ori_n1026_), .B(ori_ori_n1159_), .Y(ori_ori_n2271_));
  AOI210     o2222(.A0(ori_ori_n675_), .A1(ori_ori_n689_), .B0(ori_ori_n2271_), .Y(ori_ori_n2272_));
  AOI210     o2223(.A0(ori_ori_n590_), .A1(ori_ori_n626_), .B0(ori_ori_n695_), .Y(ori_ori_n2273_));
  NO2        o2224(.A(ori_ori_n2273_), .B(ori_ori_n1834_), .Y(ori_ori_n2274_));
  NO2        o2225(.A(ori_ori_n450_), .B(ori_ori_n431_), .Y(ori_ori_n2275_));
  NOi31      o2226(.An(ori_ori_n1519_), .B(ori_ori_n2275_), .C(ori_ori_n590_), .Y(ori_ori_n2276_));
  NO4        o2227(.A(ori_ori_n2276_), .B(ori_ori_n2274_), .C(ori_ori_n2272_), .D(ori_ori_n2270_), .Y(ori_ori_n2277_));
  NA4        o2228(.A(ori_ori_n2277_), .B(ori_ori_n2266_), .C(ori_ori_n2263_), .D(ori_ori_n2227_), .Y(ori33));
  OAI210     o2229(.A0(ori_ori_n817_), .A1(x1), .B0(ori_ori_n196_), .Y(ori_ori_n2279_));
  OAI210     o2230(.A0(ori_ori_n2097_), .A1(ori_ori_n172_), .B0(ori_ori_n326_), .Y(ori_ori_n2280_));
  OAI220     o2231(.A0(ori_ori_n1088_), .A1(ori_ori_n816_), .B0(ori_ori_n1691_), .B1(ori_ori_n351_), .Y(ori_ori_n2281_));
  NA3        o2232(.A(ori_ori_n2281_), .B(ori_ori_n2280_), .C(ori_ori_n638_), .Y(ori_ori_n2282_));
  AOI210     o2233(.A0(ori_ori_n2279_), .A1(x5), .B0(ori_ori_n2282_), .Y(ori_ori_n2283_));
  NA2        o2234(.A(ori_ori_n225_), .B(ori_ori_n76_), .Y(ori_ori_n2284_));
  NA4        o2235(.A(ori_ori_n1765_), .B(ori_ori_n566_), .C(ori_ori_n242_), .D(x4), .Y(ori_ori_n2285_));
  AOI210     o2236(.A0(ori_ori_n2285_), .A1(ori_ori_n2284_), .B0(ori_ori_n351_), .Y(ori_ori_n2286_));
  OAI210     o2237(.A0(ori_ori_n434_), .A1(ori_ori_n265_), .B0(ori_ori_n53_), .Y(ori_ori_n2287_));
  AOI210     o2238(.A0(ori_ori_n2287_), .A1(ori_ori_n436_), .B0(ori_ori_n64_), .Y(ori_ori_n2288_));
  NA2        o2239(.A(ori_ori_n1679_), .B(ori_ori_n71_), .Y(ori_ori_n2289_));
  NO3        o2240(.A(ori_ori_n2289_), .B(ori_ori_n2288_), .C(ori_ori_n2286_), .Y(ori_ori_n2290_));
  OAI210     o2241(.A0(ori_ori_n2283_), .A1(x4), .B0(ori_ori_n2290_), .Y(ori_ori_n2291_));
  OAI210     o2242(.A0(ori_ori_n138_), .A1(x5), .B0(ori_ori_n235_), .Y(ori_ori_n2292_));
  NA2        o2243(.A(ori_ori_n180_), .B(x4), .Y(ori_ori_n2293_));
  NA2        o2244(.A(ori_ori_n306_), .B(ori_ori_n283_), .Y(ori_ori_n2294_));
  NO2        o2245(.A(ori_ori_n972_), .B(ori_ori_n223_), .Y(ori_ori_n2295_));
  NA2        o2246(.A(ori_ori_n641_), .B(x7), .Y(ori_ori_n2296_));
  OAI220     o2247(.A0(ori_ori_n2296_), .A1(ori_ori_n2295_), .B0(ori_ori_n2294_), .B1(ori_ori_n2293_), .Y(ori_ori_n2297_));
  AOI210     o2248(.A0(ori_ori_n2292_), .A1(ori_ori_n1034_), .B0(ori_ori_n2297_), .Y(ori_ori_n2298_));
  NA2        o2249(.A(ori_ori_n207_), .B(ori_ori_n963_), .Y(ori_ori_n2299_));
  AOI210     o2250(.A0(ori_ori_n2299_), .A1(ori_ori_n2222_), .B0(ori_ori_n209_), .Y(ori_ori_n2300_));
  NO2        o2251(.A(ori_ori_n1665_), .B(ori_ori_n964_), .Y(ori_ori_n2301_));
  OAI210     o2252(.A0(ori_ori_n870_), .A1(ori_ori_n51_), .B0(x6), .Y(ori_ori_n2302_));
  NA3        o2253(.A(ori_ori_n926_), .B(ori_ori_n735_), .C(ori_ori_n55_), .Y(ori_ori_n2303_));
  OAI210     o2254(.A0(ori_ori_n620_), .A1(ori_ori_n505_), .B0(ori_ori_n2303_), .Y(ori_ori_n2304_));
  NO4        o2255(.A(ori_ori_n2304_), .B(ori_ori_n2302_), .C(ori_ori_n2301_), .D(ori_ori_n2300_), .Y(ori_ori_n2305_));
  OAI210     o2256(.A0(ori_ori_n2298_), .A1(ori_ori_n50_), .B0(ori_ori_n2305_), .Y(ori_ori_n2306_));
  NA3        o2257(.A(ori_ori_n2306_), .B(ori_ori_n2291_), .C(ori_ori_n59_), .Y(ori_ori_n2307_));
  NA2        o2258(.A(ori_ori_n535_), .B(ori_ori_n105_), .Y(ori_ori_n2308_));
  NO3        o2259(.A(ori_ori_n1585_), .B(ori_ori_n372_), .C(x4), .Y(ori_ori_n2309_));
  AOI210     o2260(.A0(ori_ori_n2309_), .A1(ori_ori_n2308_), .B0(ori_ori_n437_), .Y(ori_ori_n2310_));
  NA2        o2261(.A(ori_ori_n819_), .B(ori_ori_n104_), .Y(ori_ori_n2311_));
  NA2        o2262(.A(ori_ori_n2311_), .B(ori_ori_n461_), .Y(ori_ori_n2312_));
  NO2        o2263(.A(ori_ori_n710_), .B(ori_ori_n373_), .Y(ori_ori_n2313_));
  NA2        o2264(.A(ori_ori_n501_), .B(ori_ori_n53_), .Y(ori_ori_n2314_));
  AOI210     o2265(.A0(ori_ori_n2313_), .A1(ori_ori_n2312_), .B0(ori_ori_n2314_), .Y(ori_ori_n2315_));
  OAI210     o2266(.A0(ori_ori_n2310_), .A1(ori_ori_n59_), .B0(ori_ori_n2315_), .Y(ori_ori_n2316_));
  AOI220     o2267(.A0(ori_ori_n689_), .A1(ori_ori_n232_), .B0(ori_ori_n385_), .B1(ori_ori_n226_), .Y(ori_ori_n2317_));
  NA2        o2268(.A(ori_ori_n736_), .B(ori_ori_n984_), .Y(ori_ori_n2318_));
  OAI210     o2269(.A0(ori_ori_n2318_), .A1(ori_ori_n2317_), .B0(ori_ori_n300_), .Y(ori_ori_n2319_));
  AOI210     o2270(.A0(ori_ori_n2127_), .A1(ori_ori_n210_), .B0(ori_ori_n53_), .Y(ori_ori_n2320_));
  NO2        o2271(.A(ori_ori_n136_), .B(ori_ori_n336_), .Y(ori_ori_n2321_));
  AOI220     o2272(.A0(ori_ori_n2321_), .A1(ori_ori_n1004_), .B0(ori_ori_n674_), .B1(ori_ori_n351_), .Y(ori_ori_n2322_));
  NA2        o2273(.A(ori_ori_n445_), .B(ori_ori_n499_), .Y(ori_ori_n2323_));
  NO3        o2274(.A(ori_ori_n2323_), .B(ori_ori_n1040_), .C(ori_ori_n177_), .Y(ori_ori_n2324_));
  AOI210     o2275(.A0(ori_ori_n1810_), .A1(ori_ori_n1203_), .B0(ori_ori_n2324_), .Y(ori_ori_n2325_));
  NA4        o2276(.A(ori_ori_n2325_), .B(ori_ori_n2322_), .C(ori_ori_n2320_), .D(ori_ori_n2319_), .Y(ori_ori_n2326_));
  NA3        o2277(.A(ori_ori_n2326_), .B(ori_ori_n2316_), .C(ori_ori_n57_), .Y(ori_ori_n2327_));
  NAi21      o2278(.An(ori_ori_n1205_), .B(ori_ori_n489_), .Y(ori_ori_n2328_));
  NA4        o2279(.A(ori_ori_n641_), .B(ori_ori_n1318_), .C(ori_ori_n470_), .D(ori_ori_n50_), .Y(ori_ori_n2329_));
  OAI210     o2280(.A0(ori_ori_n2321_), .A1(ori_ori_n2071_), .B0(x2), .Y(ori_ori_n2330_));
  NA4        o2281(.A(ori_ori_n283_), .B(ori_ori_n151_), .C(ori_ori_n272_), .D(ori_ori_n118_), .Y(ori_ori_n2331_));
  NA3        o2282(.A(ori_ori_n2331_), .B(ori_ori_n2330_), .C(ori_ori_n2329_), .Y(ori_ori_n2332_));
  AO220      o2283(.A0(ori_ori_n2332_), .A1(x0), .B0(ori_ori_n2328_), .B1(ori_ori_n133_), .Y(ori_ori_n2333_));
  NA3        o2284(.A(ori_ori_n779_), .B(ori_ori_n351_), .C(ori_ori_n60_), .Y(ori_ori_n2334_));
  NO2        o2285(.A(ori_ori_n2267_), .B(ori_ori_n412_), .Y(ori_ori_n2335_));
  NA2        o2286(.A(ori_ori_n639_), .B(ori_ori_n517_), .Y(ori_ori_n2336_));
  OAI220     o2287(.A0(ori_ori_n2336_), .A1(ori_ori_n2335_), .B0(ori_ori_n2334_), .B1(ori_ori_n71_), .Y(ori_ori_n2337_));
  OAI210     o2288(.A0(ori_ori_n1549_), .A1(ori_ori_n347_), .B0(ori_ori_n107_), .Y(ori_ori_n2338_));
  AOI210     o2289(.A0(ori_ori_n590_), .A1(ori_ori_n466_), .B0(ori_ori_n133_), .Y(ori_ori_n2339_));
  OAI210     o2290(.A0(ori_ori_n2339_), .A1(ori_ori_n385_), .B0(ori_ori_n2338_), .Y(ori_ori_n2340_));
  OAI210     o2291(.A0(ori_ori_n2340_), .A1(ori_ori_n2337_), .B0(ori_ori_n98_), .Y(ori_ori_n2341_));
  NA3        o2292(.A(ori_ori_n1223_), .B(ori_ori_n126_), .C(ori_ori_n380_), .Y(ori_ori_n2342_));
  NA2        o2293(.A(ori_ori_n2342_), .B(ori_ori_n1838_), .Y(ori_ori_n2343_));
  NA2        o2294(.A(ori_ori_n1202_), .B(ori_ori_n713_), .Y(ori_ori_n2344_));
  NA2        o2295(.A(ori_ori_n1372_), .B(ori_ori_n1183_), .Y(ori_ori_n2345_));
  NA4        o2296(.A(ori_ori_n2345_), .B(ori_ori_n2344_), .C(ori_ori_n2343_), .D(ori_ori_n2341_), .Y(ori_ori_n2346_));
  AOI210     o2297(.A0(ori_ori_n2333_), .A1(x7), .B0(ori_ori_n2346_), .Y(ori_ori_n2347_));
  NA3        o2298(.A(ori_ori_n2347_), .B(ori_ori_n2327_), .C(ori_ori_n2307_), .Y(ori34));
  NA2        o2299(.A(ori_ori_n431_), .B(x4), .Y(ori_ori_n2349_));
  NO2        o2300(.A(ori_ori_n1970_), .B(ori_ori_n863_), .Y(ori_ori_n2350_));
  AOI210     o2301(.A0(ori_ori_n2350_), .A1(ori_ori_n2349_), .B0(ori_ori_n317_), .Y(ori_ori_n2351_));
  NA2        o2302(.A(ori_ori_n283_), .B(ori_ori_n119_), .Y(ori_ori_n2352_));
  NO2        o2303(.A(ori_ori_n982_), .B(ori_ori_n2352_), .Y(ori_ori_n2353_));
  AOI210     o2304(.A0(ori_ori_n2051_), .A1(ori_ori_n543_), .B0(ori_ori_n135_), .Y(ori_ori_n2354_));
  NA2        o2305(.A(ori_ori_n1970_), .B(x0), .Y(ori_ori_n2355_));
  OAI210     o2306(.A0(ori_ori_n1847_), .A1(ori_ori_n986_), .B0(ori_ori_n2355_), .Y(ori_ori_n2356_));
  NO4        o2307(.A(ori_ori_n2356_), .B(ori_ori_n2354_), .C(ori_ori_n2353_), .D(ori_ori_n2351_), .Y(ori_ori_n2357_));
  NO2        o2308(.A(ori_ori_n2357_), .B(ori_ori_n476_), .Y(ori_ori_n2358_));
  NA2        o2309(.A(ori_ori_n738_), .B(x8), .Y(ori_ori_n2359_));
  AO210      o2310(.A0(ori_ori_n2359_), .A1(ori_ori_n486_), .B0(ori_ori_n664_), .Y(ori_ori_n2360_));
  NA2        o2311(.A(ori_ori_n674_), .B(ori_ori_n631_), .Y(ori_ori_n2361_));
  AOI210     o2312(.A0(ori_ori_n2361_), .A1(ori_ori_n2360_), .B0(ori_ori_n261_), .Y(ori_ori_n2362_));
  OAI210     o2313(.A0(ori_ori_n118_), .A1(ori_ori_n1062_), .B0(ori_ori_n1484_), .Y(ori_ori_n2363_));
  OAI210     o2314(.A0(ori_ori_n1625_), .A1(ori_ori_n58_), .B0(ori_ori_n2363_), .Y(ori_ori_n2364_));
  NA3        o2315(.A(ori_ori_n2364_), .B(ori_ori_n337_), .C(x8), .Y(ori_ori_n2365_));
  NO3        o2316(.A(ori_ori_n1003_), .B(ori_ori_n710_), .C(ori_ori_n455_), .Y(ori_ori_n2366_));
  AOI210     o2317(.A0(ori_ori_n1607_), .A1(ori_ori_n325_), .B0(ori_ori_n2366_), .Y(ori_ori_n2367_));
  NA2        o2318(.A(ori_ori_n668_), .B(ori_ori_n317_), .Y(ori_ori_n2368_));
  NA2        o2319(.A(ori_ori_n129_), .B(x0), .Y(ori_ori_n2369_));
  NAi31      o2320(.An(ori_ori_n2369_), .B(ori_ori_n2368_), .C(ori_ori_n804_), .Y(ori_ori_n2370_));
  NA3        o2321(.A(ori_ori_n1620_), .B(ori_ori_n1414_), .C(ori_ori_n50_), .Y(ori_ori_n2371_));
  NA4        o2322(.A(ori_ori_n2371_), .B(ori_ori_n2370_), .C(ori_ori_n2367_), .D(ori_ori_n2365_), .Y(ori_ori_n2372_));
  NA2        o2323(.A(ori_ori_n1121_), .B(ori_ori_n754_), .Y(ori_ori_n2373_));
  NA3        o2324(.A(ori_ori_n1161_), .B(ori_ori_n162_), .C(ori_ori_n1105_), .Y(ori_ori_n2374_));
  AOI210     o2325(.A0(ori_ori_n2374_), .A1(ori_ori_n2373_), .B0(ori_ori_n764_), .Y(ori_ori_n2375_));
  AOI210     o2326(.A0(ori_ori_n1793_), .A1(ori_ori_n125_), .B0(ori_ori_n2375_), .Y(ori_ori_n2376_));
  AOI210     o2327(.A0(ori_ori_n557_), .A1(ori_ori_n821_), .B0(ori_ori_n250_), .Y(ori_ori_n2377_));
  OAI220     o2328(.A0(ori_ori_n2377_), .A1(ori_ori_n59_), .B0(ori_ori_n1132_), .B1(ori_ori_n55_), .Y(ori_ori_n2378_));
  NA3        o2329(.A(ori_ori_n2378_), .B(ori_ori_n738_), .C(ori_ori_n56_), .Y(ori_ori_n2379_));
  OAI210     o2330(.A0(ori_ori_n2376_), .A1(ori_ori_n136_), .B0(ori_ori_n2379_), .Y(ori_ori_n2380_));
  NO4        o2331(.A(ori_ori_n2380_), .B(ori_ori_n2372_), .C(ori_ori_n2362_), .D(ori_ori_n2358_), .Y(ori_ori_n2381_));
  NO2        o2332(.A(ori_ori_n307_), .B(ori_ori_n963_), .Y(ori_ori_n2382_));
  NO3        o2333(.A(ori_ori_n2382_), .B(ori_ori_n443_), .C(ori_ori_n325_), .Y(ori_ori_n2383_));
  NA2        o2334(.A(ori_ori_n789_), .B(ori_ori_n155_), .Y(ori_ori_n2384_));
  NO3        o2335(.A(ori_ori_n2243_), .B(ori_ori_n300_), .C(ori_ori_n1105_), .Y(ori_ori_n2385_));
  OAI220     o2336(.A0(ori_ori_n2385_), .A1(ori_ori_n1577_), .B0(ori_ori_n2384_), .B1(ori_ori_n1187_), .Y(ori_ori_n2386_));
  OAI210     o2337(.A0(ori_ori_n2386_), .A1(ori_ori_n2383_), .B0(x2), .Y(ori_ori_n2387_));
  OAI210     o2338(.A0(ori_ori_n873_), .A1(ori_ori_n368_), .B0(ori_ori_n2387_), .Y(ori_ori_n2388_));
  NA2        o2339(.A(ori_ori_n310_), .B(x4), .Y(ori_ori_n2389_));
  OAI220     o2340(.A0(ori_ori_n750_), .A1(ori_ori_n55_), .B0(ori_ori_n276_), .B1(ori_ori_n103_), .Y(ori_ori_n2390_));
  NO4        o2341(.A(ori_ori_n447_), .B(ori_ori_n77_), .C(x7), .D(x3), .Y(ori_ori_n2391_));
  NO2        o2342(.A(ori_ori_n1121_), .B(ori_ori_n284_), .Y(ori_ori_n2392_));
  NO4        o2343(.A(ori_ori_n2392_), .B(ori_ori_n2391_), .C(ori_ori_n2390_), .D(ori_ori_n2389_), .Y(ori_ori_n2393_));
  NA2        o2344(.A(ori_ori_n1258_), .B(ori_ori_n1060_), .Y(ori_ori_n2394_));
  NA3        o2345(.A(ori_ori_n1411_), .B(ori_ori_n253_), .C(x7), .Y(ori_ori_n2395_));
  NA2        o2346(.A(ori_ori_n2395_), .B(ori_ori_n2394_), .Y(ori_ori_n2396_));
  OAI210     o2347(.A0(ori_ori_n2396_), .A1(ori_ori_n2393_), .B0(ori_ori_n159_), .Y(ori_ori_n2397_));
  NA3        o2348(.A(ori_ori_n868_), .B(ori_ori_n87_), .C(x0), .Y(ori_ori_n2398_));
  NA4        o2349(.A(ori_ori_n2398_), .B(ori_ori_n1165_), .C(ori_ori_n293_), .D(ori_ori_n588_), .Y(ori_ori_n2399_));
  NA2        o2350(.A(ori_ori_n1169_), .B(ori_ori_n679_), .Y(ori_ori_n2400_));
  OAI210     o2351(.A0(ori_ori_n2400_), .A1(ori_ori_n262_), .B0(ori_ori_n2179_), .Y(ori_ori_n2401_));
  AOI220     o2352(.A0(ori_ori_n2401_), .A1(x7), .B0(ori_ori_n1025_), .B1(ori_ori_n665_), .Y(ori_ori_n2402_));
  OAI210     o2353(.A0(ori_ori_n2064_), .A1(ori_ori_n258_), .B0(ori_ori_n742_), .Y(ori_ori_n2403_));
  AOI220     o2354(.A0(ori_ori_n408_), .A1(x8), .B0(ori_ori_n90_), .B1(x2), .Y(ori_ori_n2404_));
  AOI210     o2355(.A0(ori_ori_n266_), .A1(ori_ori_n53_), .B0(ori_ori_n656_), .Y(ori_ori_n2405_));
  OAI220     o2356(.A0(ori_ori_n2405_), .A1(ori_ori_n93_), .B0(ori_ori_n2404_), .B1(ori_ori_n1358_), .Y(ori_ori_n2406_));
  AOI220     o2357(.A0(ori_ori_n2406_), .A1(ori_ori_n1336_), .B0(ori_ori_n2403_), .B1(ori_ori_n1534_), .Y(ori_ori_n2407_));
  NA4        o2358(.A(ori_ori_n2407_), .B(ori_ori_n2402_), .C(ori_ori_n2399_), .D(ori_ori_n2397_), .Y(ori_ori_n2408_));
  AOI210     o2359(.A0(ori_ori_n2388_), .A1(ori_ori_n821_), .B0(ori_ori_n2408_), .Y(ori_ori_n2409_));
  OAI210     o2360(.A0(ori_ori_n2381_), .A1(x2), .B0(ori_ori_n2409_), .Y(ori35));
  NA2        o2361(.A(ori_ori_n505_), .B(ori_ori_n173_), .Y(ori_ori_n2411_));
  AOI220     o2362(.A0(ori_ori_n639_), .A1(ori_ori_n55_), .B0(ori_ori_n779_), .B1(ori_ori_n1238_), .Y(ori_ori_n2412_));
  AOI210     o2363(.A0(ori_ori_n2412_), .A1(ori_ori_n2411_), .B0(ori_ori_n71_), .Y(ori_ori_n2413_));
  NO3        o2364(.A(ori_ori_n513_), .B(ori_ori_n466_), .C(ori_ori_n336_), .Y(ori_ori_n2414_));
  OAI210     o2365(.A0(ori_ori_n2414_), .A1(ori_ori_n2413_), .B0(x2), .Y(ori_ori_n2415_));
  AOI210     o2366(.A0(ori_ori_n211_), .A1(x0), .B0(ori_ori_n270_), .Y(ori_ori_n2416_));
  OAI220     o2367(.A0(ori_ori_n2416_), .A1(ori_ori_n670_), .B0(ori_ori_n193_), .B1(x4), .Y(ori_ori_n2417_));
  NA2        o2368(.A(ori_ori_n2417_), .B(ori_ori_n133_), .Y(ori_ori_n2418_));
  NA3        o2369(.A(ori_ori_n408_), .B(x8), .C(ori_ori_n71_), .Y(ori_ori_n2419_));
  AOI210     o2370(.A0(ori_ori_n2419_), .A1(ori_ori_n1741_), .B0(ori_ori_n689_), .Y(ori_ori_n2420_));
  OAI210     o2371(.A0(ori_ori_n2334_), .A1(x6), .B0(ori_ori_n753_), .Y(ori_ori_n2421_));
  NO2        o2372(.A(ori_ori_n2421_), .B(ori_ori_n2420_), .Y(ori_ori_n2422_));
  NA3        o2373(.A(ori_ori_n2422_), .B(ori_ori_n2418_), .C(ori_ori_n2415_), .Y(ori_ori_n2423_));
  NAi21      o2374(.An(ori_ori_n1706_), .B(ori_ori_n1315_), .Y(ori_ori_n2424_));
  NA2        o2375(.A(ori_ori_n209_), .B(ori_ori_n575_), .Y(ori_ori_n2425_));
  NO2        o2376(.A(ori_ori_n431_), .B(ori_ori_n424_), .Y(ori_ori_n2426_));
  AOI220     o2377(.A0(ori_ori_n2426_), .A1(ori_ori_n2425_), .B0(ori_ori_n2424_), .B1(ori_ori_n56_), .Y(ori_ori_n2427_));
  NA2        o2378(.A(ori_ori_n768_), .B(ori_ori_n702_), .Y(ori_ori_n2428_));
  NO3        o2379(.A(ori_ori_n684_), .B(ori_ori_n55_), .C(x6), .Y(ori_ori_n2429_));
  OAI210     o2380(.A0(ori_ori_n2429_), .A1(ori_ori_n713_), .B0(ori_ori_n214_), .Y(ori_ori_n2430_));
  NA2        o2381(.A(ori_ori_n1344_), .B(ori_ori_n63_), .Y(ori_ori_n2431_));
  NA2        o2382(.A(x6), .B(ori_ori_n471_), .Y(ori_ori_n2432_));
  NA3        o2383(.A(ori_ori_n2432_), .B(ori_ori_n2431_), .C(ori_ori_n2430_), .Y(ori_ori_n2433_));
  NA3        o2384(.A(ori_ori_n1289_), .B(ori_ori_n756_), .C(x3), .Y(ori_ori_n2434_));
  NO3        o2385(.A(ori_ori_n2434_), .B(ori_ori_n686_), .C(ori_ori_n202_), .Y(ori_ori_n2435_));
  AOI210     o2386(.A0(ori_ori_n2433_), .A1(ori_ori_n50_), .B0(ori_ori_n2435_), .Y(ori_ori_n2436_));
  OAI210     o2387(.A0(ori_ori_n2428_), .A1(ori_ori_n2427_), .B0(ori_ori_n2436_), .Y(ori_ori_n2437_));
  AOI210     o2388(.A0(ori_ori_n2423_), .A1(ori_ori_n57_), .B0(ori_ori_n2437_), .Y(ori_ori_n2438_));
  NA2        o2389(.A(ori_ori_n972_), .B(ori_ori_n63_), .Y(ori_ori_n2439_));
  NO3        o2390(.A(ori_ori_n1084_), .B(ori_ori_n565_), .C(ori_ori_n119_), .Y(ori_ori_n2440_));
  OAI210     o2391(.A0(ori_ori_n152_), .A1(ori_ori_n67_), .B0(ori_ori_n2440_), .Y(ori_ori_n2441_));
  AOI210     o2392(.A0(ori_ori_n2441_), .A1(ori_ori_n2439_), .B0(ori_ori_n50_), .Y(ori_ori_n2442_));
  NA4        o2393(.A(ori_ori_n466_), .B(ori_ori_n226_), .C(ori_ori_n879_), .D(ori_ori_n100_), .Y(ori_ori_n2443_));
  OAI210     o2394(.A0(ori_ori_n972_), .A1(ori_ori_n251_), .B0(ori_ori_n757_), .Y(ori_ori_n2444_));
  OAI210     o2395(.A0(ori_ori_n251_), .A1(ori_ori_n587_), .B0(ori_ori_n2176_), .Y(ori_ori_n2445_));
  NA3        o2396(.A(ori_ori_n2445_), .B(ori_ori_n2444_), .C(ori_ori_n2443_), .Y(ori_ori_n2446_));
  OAI210     o2397(.A0(ori_ori_n2446_), .A1(ori_ori_n2442_), .B0(ori_ori_n59_), .Y(ori_ori_n2447_));
  AOI210     o2398(.A0(ori_ori_n868_), .A1(ori_ori_n534_), .B0(ori_ori_n1922_), .Y(ori_ori_n2448_));
  AOI210     o2399(.A0(ori_ori_n565_), .A1(ori_ori_n609_), .B0(ori_ori_n2448_), .Y(ori_ori_n2449_));
  NO4        o2400(.A(ori_ori_n964_), .B(ori_ori_n565_), .C(ori_ori_n360_), .D(ori_ori_n406_), .Y(ori_ori_n2450_));
  XN2        o2401(.A(x4), .B(x3), .Y(ori_ori_n2451_));
  NO3        o2402(.A(ori_ori_n2451_), .B(ori_ori_n669_), .C(ori_ori_n306_), .Y(ori_ori_n2452_));
  NO3        o2403(.A(ori_ori_n2452_), .B(ori_ori_n2450_), .C(ori_ori_n1480_), .Y(ori_ori_n2453_));
  OAI210     o2404(.A0(ori_ori_n2449_), .A1(x3), .B0(ori_ori_n2453_), .Y(ori_ori_n2454_));
  NO3        o2405(.A(ori_ori_n750_), .B(ori_ori_n870_), .C(ori_ori_n271_), .Y(ori_ori_n2455_));
  OAI210     o2406(.A0(ori_ori_n2455_), .A1(ori_ori_n1480_), .B0(ori_ori_n50_), .Y(ori_ori_n2456_));
  NA3        o2407(.A(ori_ori_n1092_), .B(ori_ori_n819_), .C(ori_ori_n250_), .Y(ori_ori_n2457_));
  NA2        o2408(.A(ori_ori_n2457_), .B(ori_ori_n2456_), .Y(ori_ori_n2458_));
  AOI210     o2409(.A0(ori_ori_n2454_), .A1(ori_ori_n590_), .B0(ori_ori_n2458_), .Y(ori_ori_n2459_));
  AOI210     o2410(.A0(ori_ori_n1450_), .A1(ori_ori_n646_), .B0(ori_ori_n686_), .Y(ori_ori_n2460_));
  NO2        o2411(.A(ori_ori_n879_), .B(ori_ori_n56_), .Y(ori_ori_n2461_));
  OAI210     o2412(.A0(ori_ori_n1973_), .A1(ori_ori_n609_), .B0(ori_ori_n2267_), .Y(ori_ori_n2462_));
  OAI210     o2413(.A0(ori_ori_n2359_), .A1(ori_ori_n2461_), .B0(ori_ori_n2462_), .Y(ori_ori_n2463_));
  OAI210     o2414(.A0(ori_ori_n2463_), .A1(ori_ori_n2460_), .B0(ori_ori_n90_), .Y(ori_ori_n2464_));
  NO2        o2415(.A(ori_ori_n861_), .B(ori_ori_n666_), .Y(ori_ori_n2465_));
  NO2        o2416(.A(ori_ori_n284_), .B(x6), .Y(ori_ori_n2466_));
  OAI210     o2417(.A0(ori_ori_n2465_), .A1(ori_ori_n1801_), .B0(ori_ori_n2466_), .Y(ori_ori_n2467_));
  NA4        o2418(.A(ori_ori_n2467_), .B(ori_ori_n2464_), .C(ori_ori_n2459_), .D(ori_ori_n2447_), .Y(ori_ori_n2468_));
  NA4        o2419(.A(ori_ori_n617_), .B(ori_ori_n689_), .C(ori_ori_n430_), .D(x6), .Y(ori_ori_n2469_));
  AOI210     o2420(.A0(ori_ori_n2469_), .A1(ori_ori_n425_), .B0(x1), .Y(ori_ori_n2470_));
  NO2        o2421(.A(ori_ori_n736_), .B(ori_ori_n686_), .Y(ori_ori_n2471_));
  OAI210     o2422(.A0(ori_ori_n466_), .A1(ori_ori_n163_), .B0(ori_ori_n801_), .Y(ori_ori_n2472_));
  AOI210     o2423(.A0(ori_ori_n2472_), .A1(ori_ori_n1030_), .B0(ori_ori_n53_), .Y(ori_ori_n2473_));
  NO3        o2424(.A(ori_ori_n2473_), .B(ori_ori_n2471_), .C(ori_ori_n2470_), .Y(ori_ori_n2474_));
  NA3        o2425(.A(ori_ori_n1452_), .B(ori_ori_n1290_), .C(ori_ori_n825_), .Y(ori_ori_n2475_));
  AOI220     o2426(.A0(ori_ori_n1962_), .A1(ori_ori_n133_), .B0(ori_ori_n417_), .B1(ori_ori_n122_), .Y(ori_ori_n2476_));
  AOI210     o2427(.A0(ori_ori_n2476_), .A1(ori_ori_n2475_), .B0(ori_ori_n1527_), .Y(ori_ori_n2477_));
  NO2        o2428(.A(ori_ori_n639_), .B(x3), .Y(ori_ori_n2478_));
  NO3        o2429(.A(ori_ori_n697_), .B(ori_ori_n1625_), .C(x2), .Y(ori_ori_n2479_));
  AOI220     o2430(.A0(ori_ori_n2479_), .A1(ori_ori_n2478_), .B0(ori_ori_n1936_), .B1(ori_ori_n775_), .Y(ori_ori_n2480_));
  NA3        o2431(.A(x6), .B(x4), .C(x0), .Y(ori_ori_n2481_));
  OAI220     o2432(.A0(ori_ori_n2481_), .A1(ori_ori_n192_), .B0(ori_ori_n684_), .B1(ori_ori_n530_), .Y(ori_ori_n2482_));
  OAI220     o2433(.A0(ori_ori_n1325_), .A1(x8), .B0(ori_ori_n372_), .B1(ori_ori_n350_), .Y(ori_ori_n2483_));
  AOI220     o2434(.A0(ori_ori_n2483_), .A1(ori_ori_n417_), .B0(ori_ori_n2482_), .B1(ori_ori_n925_), .Y(ori_ori_n2484_));
  OAI210     o2435(.A0(ori_ori_n2480_), .A1(ori_ori_n1178_), .B0(ori_ori_n2484_), .Y(ori_ori_n2485_));
  NO2        o2436(.A(ori_ori_n2485_), .B(ori_ori_n2477_), .Y(ori_ori_n2486_));
  OAI210     o2437(.A0(ori_ori_n2474_), .A1(ori_ori_n310_), .B0(ori_ori_n2486_), .Y(ori_ori_n2487_));
  AOI210     o2438(.A0(ori_ori_n2468_), .A1(x5), .B0(ori_ori_n2487_), .Y(ori_ori_n2488_));
  OAI210     o2439(.A0(ori_ori_n2438_), .A1(x5), .B0(ori_ori_n2488_), .Y(ori36));
  NO2        o2440(.A(ori_ori_n870_), .B(ori_ori_n299_), .Y(ori_ori_n2490_));
  NO3        o2441(.A(ori_ori_n118_), .B(ori_ori_n1062_), .C(ori_ori_n55_), .Y(ori_ori_n2491_));
  NO3        o2442(.A(ori_ori_n2491_), .B(ori_ori_n1992_), .C(ori_ori_n1084_), .Y(ori_ori_n2492_));
  OAI210     o2443(.A0(ori_ori_n2492_), .A1(ori_ori_n2490_), .B0(ori_ori_n106_), .Y(ori_ori_n2493_));
  OR4        o2444(.A(ori_ori_n965_), .B(ori_ori_n812_), .C(ori_ori_n375_), .D(ori_ori_n493_), .Y(ori_ori_n2494_));
  INV        o2445(.A(ori_ori_n1015_), .Y(ori_ori_n2495_));
  OAI210     o2446(.A0(ori_ori_n2229_), .A1(ori_ori_n2495_), .B0(ori_ori_n276_), .Y(ori_ori_n2496_));
  NA3        o2447(.A(ori_ori_n445_), .B(ori_ori_n223_), .C(ori_ori_n117_), .Y(ori_ori_n2497_));
  NA4        o2448(.A(ori_ori_n2497_), .B(ori_ori_n2496_), .C(ori_ori_n2494_), .D(ori_ori_n2493_), .Y(ori_ori_n2498_));
  NO2        o2449(.A(ori_ori_n1004_), .B(x8), .Y(ori_ori_n2499_));
  NO3        o2450(.A(ori_ori_n2499_), .B(ori_ori_n1000_), .C(ori_ori_n539_), .Y(ori_ori_n2500_));
  AOI220     o2451(.A0(ori_ori_n300_), .A1(x1), .B0(ori_ori_n132_), .B1(x6), .Y(ori_ori_n2501_));
  AOI210     o2452(.A0(ori_ori_n1105_), .A1(x6), .B0(ori_ori_n421_), .Y(ori_ori_n2502_));
  OAI220     o2453(.A0(ori_ori_n2502_), .A1(ori_ori_n359_), .B0(ori_ori_n2501_), .B1(ori_ori_n467_), .Y(ori_ori_n2503_));
  OAI210     o2454(.A0(ori_ori_n2503_), .A1(ori_ori_n2500_), .B0(ori_ori_n466_), .Y(ori_ori_n2504_));
  NA2        o2455(.A(ori_ori_n674_), .B(ori_ori_n493_), .Y(ori_ori_n2505_));
  AOI210     o2456(.A0(ori_ori_n2505_), .A1(ori_ori_n653_), .B0(ori_ori_n262_), .Y(ori_ori_n2506_));
  NO3        o2457(.A(ori_ori_n1893_), .B(ori_ori_n1624_), .C(ori_ori_n272_), .Y(ori_ori_n2507_));
  NO2        o2458(.A(ori_ori_n2439_), .B(ori_ori_n225_), .Y(ori_ori_n2508_));
  NO4        o2459(.A(ori_ori_n2508_), .B(ori_ori_n2507_), .C(ori_ori_n2506_), .D(ori_ori_n419_), .Y(ori_ori_n2509_));
  OAI210     o2460(.A0(ori_ori_n641_), .A1(ori_ori_n811_), .B0(ori_ori_n990_), .Y(ori_ori_n2510_));
  OAI220     o2461(.A0(ori_ori_n1670_), .A1(ori_ori_n1665_), .B0(ori_ori_n990_), .B1(ori_ori_n1105_), .Y(ori_ori_n2511_));
  AOI220     o2462(.A0(ori_ori_n2511_), .A1(ori_ori_n116_), .B0(ori_ori_n2510_), .B1(ori_ori_n631_), .Y(ori_ori_n2512_));
  NA3        o2463(.A(ori_ori_n2512_), .B(ori_ori_n2509_), .C(ori_ori_n2504_), .Y(ori_ori_n2513_));
  AOI210     o2464(.A0(ori_ori_n2498_), .A1(ori_ori_n337_), .B0(ori_ori_n2513_), .Y(ori_ori_n2514_));
  OAI210     o2465(.A0(ori_ori_n595_), .A1(ori_ori_n518_), .B0(ori_ori_n163_), .Y(ori_ori_n2515_));
  OAI210     o2466(.A0(ori_ori_n2007_), .A1(ori_ori_n70_), .B0(ori_ori_n2515_), .Y(ori_ori_n2516_));
  OAI210     o2467(.A0(ori_ori_n496_), .A1(ori_ori_n234_), .B0(ori_ori_n251_), .Y(ori_ori_n2517_));
  NO2        o2468(.A(ori_ori_n2016_), .B(ori_ori_n169_), .Y(ori_ori_n2518_));
  NA2        o2469(.A(ori_ori_n1225_), .B(ori_ori_n55_), .Y(ori_ori_n2519_));
  OAI210     o2470(.A0(ori_ori_n2519_), .A1(ori_ori_n2518_), .B0(ori_ori_n2517_), .Y(ori_ori_n2520_));
  OAI210     o2471(.A0(ori_ori_n2520_), .A1(ori_ori_n2516_), .B0(ori_ori_n904_), .Y(ori_ori_n2521_));
  AOI210     o2472(.A0(ori_ori_n103_), .A1(ori_ori_n106_), .B0(ori_ori_n339_), .Y(ori_ori_n2522_));
  NA2        o2473(.A(ori_ori_n674_), .B(ori_ori_n1625_), .Y(ori_ori_n2523_));
  OAI220     o2474(.A0(ori_ori_n2523_), .A1(ori_ori_n2522_), .B0(ori_ori_n753_), .B1(ori_ori_n1272_), .Y(ori_ori_n2524_));
  NO2        o2475(.A(ori_ori_n1414_), .B(ori_ori_n581_), .Y(ori_ori_n2525_));
  NO3        o2476(.A(ori_ori_n2525_), .B(ori_ori_n1809_), .C(ori_ori_n697_), .Y(ori_ori_n2526_));
  NOi31      o2477(.An(ori_ori_n2028_), .B(ori_ori_n2323_), .C(ori_ori_n763_), .Y(ori_ori_n2527_));
  NO3        o2478(.A(ori_ori_n2527_), .B(ori_ori_n2526_), .C(ori_ori_n2524_), .Y(ori_ori_n2528_));
  AOI210     o2479(.A0(ori_ori_n2528_), .A1(ori_ori_n2521_), .B0(x7), .Y(ori_ori_n2529_));
  NA2        o2480(.A(ori_ori_n132_), .B(ori_ori_n63_), .Y(ori_ori_n2530_));
  AOI210     o2481(.A0(ori_ori_n590_), .A1(ori_ori_n626_), .B0(ori_ori_n1203_), .Y(ori_ori_n2531_));
  NA4        o2482(.A(ori_ori_n2531_), .B(ori_ori_n2530_), .C(ori_ori_n1003_), .D(ori_ori_n897_), .Y(ori_ori_n2532_));
  NA2        o2483(.A(ori_ori_n2532_), .B(ori_ori_n505_), .Y(ori_ori_n2533_));
  AOI220     o2484(.A0(ori_ori_n1765_), .A1(ori_ori_n254_), .B0(ori_ori_n1060_), .B1(ori_ori_n122_), .Y(ori_ori_n2534_));
  NO2        o2485(.A(ori_ori_n2534_), .B(ori_ori_n445_), .Y(ori_ori_n2535_));
  NO2        o2486(.A(ori_ori_n406_), .B(ori_ori_n223_), .Y(ori_ori_n2536_));
  NO3        o2487(.A(ori_ori_n2536_), .B(ori_ori_n1294_), .C(ori_ori_n59_), .Y(ori_ori_n2537_));
  AOI210     o2488(.A0(ori_ori_n1242_), .A1(ori_ori_n407_), .B0(x6), .Y(ori_ori_n2538_));
  NA3        o2489(.A(ori_ori_n1697_), .B(ori_ori_n276_), .C(ori_ori_n266_), .Y(ori_ori_n2539_));
  NA2        o2490(.A(ori_ori_n2539_), .B(ori_ori_n1651_), .Y(ori_ori_n2540_));
  NO4        o2491(.A(ori_ori_n2540_), .B(ori_ori_n2538_), .C(ori_ori_n2537_), .D(ori_ori_n2535_), .Y(ori_ori_n2541_));
  AOI210     o2492(.A0(ori_ori_n2541_), .A1(ori_ori_n2533_), .B0(ori_ori_n455_), .Y(ori_ori_n2542_));
  NO3        o2493(.A(ori_ori_n2451_), .B(ori_ori_n910_), .C(ori_ori_n504_), .Y(ori_ori_n2543_));
  AOI210     o2494(.A0(ori_ori_n1292_), .A1(ori_ori_n265_), .B0(ori_ori_n2543_), .Y(ori_ori_n2544_));
  OAI210     o2495(.A0(ori_ori_n877_), .A1(ori_ori_n271_), .B0(ori_ori_n396_), .Y(ori_ori_n2545_));
  NA2        o2496(.A(ori_ori_n1225_), .B(ori_ori_n168_), .Y(ori_ori_n2546_));
  NO2        o2497(.A(ori_ori_n616_), .B(ori_ori_n106_), .Y(ori_ori_n2547_));
  AO210      o2498(.A0(ori_ori_n2547_), .A1(ori_ori_n2546_), .B0(ori_ori_n1780_), .Y(ori_ori_n2548_));
  NO2        o2499(.A(ori_ori_n462_), .B(ori_ori_n418_), .Y(ori_ori_n2549_));
  AOI220     o2500(.A0(ori_ori_n2549_), .A1(ori_ori_n2548_), .B0(ori_ori_n2545_), .B1(ori_ori_n291_), .Y(ori_ori_n2550_));
  OAI210     o2501(.A0(ori_ori_n2544_), .A1(x1), .B0(ori_ori_n2550_), .Y(ori_ori_n2551_));
  NO3        o2502(.A(ori_ori_n2551_), .B(ori_ori_n2542_), .C(ori_ori_n2529_), .Y(ori_ori_n2552_));
  OAI210     o2503(.A0(ori_ori_n2514_), .A1(ori_ori_n57_), .B0(ori_ori_n2552_), .Y(ori37));
  NA3        o2504(.A(ori_ori_n1081_), .B(ori_ori_n135_), .C(x3), .Y(ori_ori_n2554_));
  NA3        o2505(.A(ori_ori_n789_), .B(ori_ori_n155_), .C(ori_ori_n50_), .Y(ori_ori_n2555_));
  AOI210     o2506(.A0(ori_ori_n2555_), .A1(ori_ori_n2554_), .B0(ori_ori_n690_), .Y(ori_ori_n2556_));
  NO3        o2507(.A(ori_ori_n1081_), .B(ori_ori_n375_), .C(ori_ori_n512_), .Y(ori_ori_n2557_));
  OAI210     o2508(.A0(ori_ori_n2557_), .A1(ori_ori_n2556_), .B0(ori_ori_n56_), .Y(ori_ori_n2558_));
  NA2        o2509(.A(ori_ori_n604_), .B(ori_ori_n754_), .Y(ori_ori_n2559_));
  AOI210     o2510(.A0(ori_ori_n2559_), .A1(ori_ori_n1061_), .B0(x3), .Y(ori_ori_n2560_));
  AOI220     o2511(.A0(ori_ori_n604_), .A1(ori_ori_n754_), .B0(ori_ori_n466_), .B1(ori_ori_n1060_), .Y(ori_ori_n2561_));
  NO2        o2512(.A(ori_ori_n669_), .B(ori_ori_n176_), .Y(ori_ori_n2562_));
  OAI220     o2513(.A0(ori_ori_n2562_), .A1(ori_ori_n846_), .B0(ori_ori_n2561_), .B1(ori_ori_n106_), .Y(ori_ori_n2563_));
  OAI210     o2514(.A0(ori_ori_n2563_), .A1(ori_ori_n2560_), .B0(ori_ori_n71_), .Y(ori_ori_n2564_));
  NA2        o2515(.A(ori_ori_n1205_), .B(ori_ori_n1084_), .Y(ori_ori_n2565_));
  OAI210     o2516(.A0(ori_ori_n1227_), .A1(ori_ori_n186_), .B0(ori_ori_n456_), .Y(ori_ori_n2566_));
  NA4        o2517(.A(ori_ori_n2566_), .B(ori_ori_n2565_), .C(ori_ori_n2564_), .D(ori_ori_n2558_), .Y(ori_ori_n2567_));
  NA2        o2518(.A(ori_ori_n424_), .B(ori_ori_n132_), .Y(ori_ori_n2568_));
  NO2        o2519(.A(ori_ori_n1728_), .B(ori_ori_n105_), .Y(ori_ori_n2569_));
  AOI210     o2520(.A0(ori_ori_n1994_), .A1(ori_ori_n871_), .B0(ori_ori_n2569_), .Y(ori_ori_n2570_));
  OAI220     o2521(.A0(ori_ori_n2570_), .A1(ori_ori_n51_), .B0(ori_ori_n1626_), .B1(ori_ori_n2568_), .Y(ori_ori_n2571_));
  AOI210     o2522(.A0(ori_ori_n2567_), .A1(ori_ori_n68_), .B0(ori_ori_n2571_), .Y(ori_ori_n2572_));
  OAI210     o2523(.A0(ori_ori_n266_), .A1(ori_ori_n1109_), .B0(ori_ori_n487_), .Y(ori_ori_n2573_));
  NA3        o2524(.A(ori_ori_n2573_), .B(ori_ori_n262_), .C(ori_ori_n1062_), .Y(ori_ori_n2574_));
  OAI210     o2525(.A0(ori_ori_n226_), .A1(ori_ori_n214_), .B0(ori_ori_n1741_), .Y(ori_ori_n2575_));
  NA2        o2526(.A(ori_ori_n345_), .B(ori_ori_n270_), .Y(ori_ori_n2576_));
  NA3        o2527(.A(ori_ori_n402_), .B(ori_ori_n825_), .C(ori_ori_n106_), .Y(ori_ori_n2577_));
  NO2        o2528(.A(ori_ori_n531_), .B(ori_ori_n56_), .Y(ori_ori_n2578_));
  NA3        o2529(.A(ori_ori_n2578_), .B(ori_ori_n2577_), .C(ori_ori_n2576_), .Y(ori_ori_n2579_));
  AOI210     o2530(.A0(ori_ori_n2575_), .A1(ori_ori_n512_), .B0(ori_ori_n2579_), .Y(ori_ori_n2580_));
  NO2        o2531(.A(ori_ori_n1196_), .B(ori_ori_n271_), .Y(ori_ori_n2581_));
  OAI210     o2532(.A0(ori_ori_n291_), .A1(ori_ori_n260_), .B0(ori_ori_n2581_), .Y(ori_ori_n2582_));
  OAI210     o2533(.A0(ori_ori_n671_), .A1(ori_ori_n133_), .B0(x3), .Y(ori_ori_n2583_));
  AOI210     o2534(.A0(ori_ori_n671_), .A1(ori_ori_n364_), .B0(ori_ori_n2583_), .Y(ori_ori_n2584_));
  AOI210     o2535(.A0(ori_ori_n1625_), .A1(ori_ori_n50_), .B0(ori_ori_n345_), .Y(ori_ori_n2585_));
  OAI210     o2536(.A0(ori_ori_n2585_), .A1(ori_ori_n401_), .B0(ori_ori_n56_), .Y(ori_ori_n2586_));
  NO2        o2537(.A(ori_ori_n2586_), .B(ori_ori_n2584_), .Y(ori_ori_n2587_));
  AOI220     o2538(.A0(ori_ori_n2587_), .A1(ori_ori_n2582_), .B0(ori_ori_n2580_), .B1(ori_ori_n2574_), .Y(ori_ori_n2588_));
  NA2        o2539(.A(ori_ori_n2588_), .B(ori_ori_n98_), .Y(ori_ori_n2589_));
  NA2        o2540(.A(ori_ori_n697_), .B(ori_ori_n1210_), .Y(ori_ori_n2590_));
  NOi21      o2541(.An(ori_ori_n1378_), .B(ori_ori_n107_), .Y(ori_ori_n2591_));
  AOI210     o2542(.A0(ori_ori_n2591_), .A1(ori_ori_n2590_), .B0(ori_ori_n434_), .Y(ori_ori_n2592_));
  NO2        o2543(.A(ori_ori_n2240_), .B(ori_ori_n55_), .Y(ori_ori_n2593_));
  OAI210     o2544(.A0(ori_ori_n2593_), .A1(ori_ori_n2592_), .B0(ori_ori_n1838_), .Y(ori_ori_n2594_));
  NA2        o2545(.A(ori_ori_n173_), .B(ori_ori_n104_), .Y(ori_ori_n2595_));
  NA2        o2546(.A(ori_ori_n689_), .B(x6), .Y(ori_ori_n2596_));
  AOI210     o2547(.A0(ori_ori_n2596_), .A1(ori_ori_n486_), .B0(ori_ori_n2595_), .Y(ori_ori_n2597_));
  AOI210     o2548(.A0(ori_ori_n352_), .A1(ori_ori_n135_), .B0(ori_ori_n136_), .Y(ori_ori_n2598_));
  OAI210     o2549(.A0(ori_ori_n2598_), .A1(ori_ori_n2597_), .B0(ori_ori_n345_), .Y(ori_ori_n2599_));
  AOI210     o2550(.A0(ori_ori_n617_), .A1(ori_ori_n434_), .B0(ori_ori_n1304_), .Y(ori_ori_n2600_));
  NO3        o2551(.A(ori_ori_n2600_), .B(ori_ori_n262_), .C(ori_ori_n63_), .Y(ori_ori_n2601_));
  OAI220     o2552(.A0(ori_ori_n2359_), .A1(ori_ori_n484_), .B0(ori_ori_n2110_), .B1(ori_ori_n385_), .Y(ori_ori_n2602_));
  OAI210     o2553(.A0(ori_ori_n2602_), .A1(ori_ori_n2601_), .B0(ori_ori_n53_), .Y(ori_ori_n2603_));
  NO4        o2554(.A(ori_ori_n2369_), .B(ori_ori_n943_), .C(ori_ori_n435_), .D(ori_ori_n217_), .Y(ori_ori_n2604_));
  NO4        o2555(.A(ori_ori_n738_), .B(ori_ori_n605_), .C(ori_ori_n443_), .D(ori_ori_n1070_), .Y(ori_ori_n2605_));
  NO3        o2556(.A(ori_ori_n2605_), .B(ori_ori_n2604_), .C(ori_ori_n1076_), .Y(ori_ori_n2606_));
  NA4        o2557(.A(ori_ori_n2606_), .B(ori_ori_n2603_), .C(ori_ori_n2599_), .D(ori_ori_n2594_), .Y(ori_ori_n2607_));
  NO3        o2558(.A(ori_ori_n246_), .B(ori_ori_n351_), .C(ori_ori_n84_), .Y(ori_ori_n2608_));
  NO2        o2559(.A(ori_ori_n274_), .B(ori_ori_n779_), .Y(ori_ori_n2609_));
  NO3        o2560(.A(ori_ori_n2609_), .B(ori_ori_n1225_), .C(ori_ori_n1244_), .Y(ori_ori_n2610_));
  OAI220     o2561(.A0(ori_ori_n2610_), .A1(ori_ori_n2608_), .B0(ori_ori_n466_), .B1(ori_ori_n85_), .Y(ori_ori_n2611_));
  OR2        o2562(.A(ori_ori_n949_), .B(ori_ori_n756_), .Y(ori_ori_n2612_));
  NA2        o2563(.A(ori_ori_n1238_), .B(ori_ori_n55_), .Y(ori_ori_n2613_));
  NOi21      o2564(.An(ori_ori_n2613_), .B(ori_ori_n386_), .Y(ori_ori_n2614_));
  AOI210     o2565(.A0(ori_ori_n2614_), .A1(ori_ori_n2612_), .B0(x1), .Y(ori_ori_n2615_));
  NA2        o2566(.A(ori_ori_n261_), .B(ori_ori_n84_), .Y(ori_ori_n2616_));
  AOI210     o2567(.A0(ori_ori_n1577_), .A1(ori_ori_n401_), .B0(ori_ori_n2616_), .Y(ori_ori_n2617_));
  NA2        o2568(.A(ori_ori_n1121_), .B(ori_ori_n62_), .Y(ori_ori_n2618_));
  NA2        o2569(.A(ori_ori_n1169_), .B(ori_ori_n169_), .Y(ori_ori_n2619_));
  OAI210     o2570(.A0(ori_ori_n2618_), .A1(ori_ori_n309_), .B0(ori_ori_n2619_), .Y(ori_ori_n2620_));
  NO3        o2571(.A(ori_ori_n2620_), .B(ori_ori_n2617_), .C(ori_ori_n2615_), .Y(ori_ori_n2621_));
  OAI210     o2572(.A0(ori_ori_n2621_), .A1(x6), .B0(ori_ori_n2611_), .Y(ori_ori_n2622_));
  AOI220     o2573(.A0(ori_ori_n2622_), .A1(ori_ori_n1484_), .B0(ori_ori_n2607_), .B1(ori_ori_n57_), .Y(ori_ori_n2623_));
  NA3        o2574(.A(ori_ori_n2623_), .B(ori_ori_n2589_), .C(ori_ori_n2572_), .Y(ori38));
  NO2        o2575(.A(ori_ori_n182_), .B(ori_ori_n984_), .Y(ori_ori_n2625_));
  AOI210     o2576(.A0(ori_ori_n1242_), .A1(ori_ori_n580_), .B0(ori_ori_n1102_), .Y(ori_ori_n2626_));
  AOI210     o2577(.A0(ori_ori_n2613_), .A1(ori_ori_n1868_), .B0(ori_ori_n225_), .Y(ori_ori_n2627_));
  NO3        o2578(.A(ori_ori_n1314_), .B(ori_ori_n317_), .C(x8), .Y(ori_ori_n2628_));
  NO4        o2579(.A(ori_ori_n2628_), .B(ori_ori_n2627_), .C(ori_ori_n2626_), .D(ori_ori_n2625_), .Y(ori_ori_n2629_));
  NO2        o2580(.A(ori_ori_n2629_), .B(x6), .Y(ori_ori_n2630_));
  NA4        o2581(.A(ori_ori_n377_), .B(ori_ori_n253_), .C(ori_ori_n185_), .D(x8), .Y(ori_ori_n2631_));
  NA2        o2582(.A(ori_ori_n400_), .B(ori_ori_n104_), .Y(ori_ori_n2632_));
  AOI210     o2583(.A0(ori_ori_n2632_), .A1(ori_ori_n2631_), .B0(ori_ori_n136_), .Y(ori_ori_n2633_));
  AOI210     o2584(.A0(ori_ori_n435_), .A1(ori_ori_n405_), .B0(ori_ori_n1751_), .Y(ori_ori_n2634_));
  NO2        o2585(.A(ori_ori_n819_), .B(ori_ori_n90_), .Y(ori_ori_n2635_));
  OAI210     o2586(.A0(ori_ori_n1034_), .A1(ori_ori_n143_), .B0(ori_ori_n358_), .Y(ori_ori_n2636_));
  OAI220     o2587(.A0(ori_ori_n2636_), .A1(ori_ori_n2635_), .B0(ori_ori_n2634_), .B1(ori_ori_n185_), .Y(ori_ori_n2637_));
  OAI210     o2588(.A0(ori_ori_n2637_), .A1(ori_ori_n2633_), .B0(x6), .Y(ori_ori_n2638_));
  NO2        o2589(.A(ori_ori_n243_), .B(ori_ori_n779_), .Y(ori_ori_n2639_));
  NO3        o2590(.A(ori_ori_n2639_), .B(ori_ori_n1706_), .C(ori_ori_n253_), .Y(ori_ori_n2640_));
  NO3        o2591(.A(x3), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n2641_));
  OAI210     o2592(.A0(ori_ori_n524_), .A1(x2), .B0(ori_ori_n2641_), .Y(ori_ori_n2642_));
  NA3        o2593(.A(ori_ori_n434_), .B(ori_ori_n424_), .C(ori_ori_n290_), .Y(ori_ori_n2643_));
  NA2        o2594(.A(ori_ori_n2643_), .B(ori_ori_n2642_), .Y(ori_ori_n2644_));
  OAI210     o2595(.A0(ori_ori_n2644_), .A1(ori_ori_n2640_), .B0(ori_ori_n821_), .Y(ori_ori_n2645_));
  NO2        o2596(.A(ori_ori_n605_), .B(ori_ori_n272_), .Y(ori_ori_n2646_));
  AN3        o2597(.A(ori_ori_n826_), .B(ori_ori_n789_), .C(x0), .Y(ori_ori_n2647_));
  OAI210     o2598(.A0(ori_ori_n2647_), .A1(ori_ori_n2646_), .B0(ori_ori_n326_), .Y(ori_ori_n2648_));
  OAI220     o2599(.A0(ori_ori_n605_), .A1(ori_ori_n272_), .B0(ori_ori_n825_), .B1(ori_ori_n91_), .Y(ori_ori_n2649_));
  OAI210     o2600(.A0(ori_ori_n689_), .A1(x0), .B0(ori_ori_n51_), .Y(ori_ori_n2650_));
  AOI210     o2601(.A0(ori_ori_n586_), .A1(x4), .B0(ori_ori_n224_), .Y(ori_ori_n2651_));
  AOI220     o2602(.A0(ori_ori_n2651_), .A1(ori_ori_n2650_), .B0(ori_ori_n2649_), .B1(ori_ori_n402_), .Y(ori_ori_n2652_));
  NA4        o2603(.A(ori_ori_n2652_), .B(ori_ori_n2648_), .C(ori_ori_n2645_), .D(ori_ori_n2638_), .Y(ori_ori_n2653_));
  OAI210     o2604(.A0(ori_ori_n2653_), .A1(ori_ori_n2630_), .B0(x7), .Y(ori_ori_n2654_));
  AOI210     o2605(.A0(ori_ori_n373_), .A1(x1), .B0(ori_ori_n1250_), .Y(ori_ori_n2655_));
  NO2        o2606(.A(ori_ori_n2655_), .B(ori_ori_n51_), .Y(ori_ori_n2656_));
  AOI210     o2607(.A0(ori_ori_n90_), .A1(ori_ori_n71_), .B0(ori_ori_n2267_), .Y(ori_ori_n2657_));
  NA2        o2608(.A(ori_ori_n385_), .B(x3), .Y(ori_ori_n2658_));
  NO2        o2609(.A(ori_ori_n1771_), .B(ori_ori_n531_), .Y(ori_ori_n2659_));
  OAI210     o2610(.A0(ori_ori_n2658_), .A1(ori_ori_n2657_), .B0(ori_ori_n2659_), .Y(ori_ori_n2660_));
  OAI210     o2611(.A0(ori_ori_n2660_), .A1(ori_ori_n2656_), .B0(x4), .Y(ori_ori_n2661_));
  INV        o2612(.A(ori_ori_n460_), .Y(ori_ori_n2662_));
  NO3        o2613(.A(ori_ori_n2662_), .B(ori_ori_n401_), .C(ori_ori_n116_), .Y(ori_ori_n2663_));
  AOI210     o2614(.A0(ori_ori_n1070_), .A1(ori_ori_n237_), .B0(ori_ori_n394_), .Y(ori_ori_n2664_));
  AO210      o2615(.A0(ori_ori_n1319_), .A1(x6), .B0(ori_ori_n2664_), .Y(ori_ori_n2665_));
  NO2        o2616(.A(ori_ori_n1435_), .B(ori_ori_n133_), .Y(ori_ori_n2666_));
  NA2        o2617(.A(ori_ori_n1970_), .B(ori_ori_n320_), .Y(ori_ori_n2667_));
  OAI220     o2618(.A0(ori_ori_n2667_), .A1(ori_ori_n1089_), .B0(ori_ori_n2666_), .B1(ori_ori_n1852_), .Y(ori_ori_n2668_));
  NO3        o2619(.A(ori_ori_n2668_), .B(ori_ori_n2665_), .C(ori_ori_n2663_), .Y(ori_ori_n2669_));
  AOI210     o2620(.A0(ori_ori_n2669_), .A1(ori_ori_n2661_), .B0(ori_ori_n104_), .Y(ori_ori_n2670_));
  NA3        o2621(.A(ori_ori_n1962_), .B(ori_ori_n605_), .C(ori_ori_n159_), .Y(ori_ori_n2671_));
  AOI210     o2622(.A0(ori_ori_n2671_), .A1(ori_ori_n1446_), .B0(ori_ori_n226_), .Y(ori_ori_n2672_));
  AOI210     o2623(.A0(ori_ori_n505_), .A1(ori_ori_n493_), .B0(ori_ori_n685_), .Y(ori_ori_n2673_));
  OAI220     o2624(.A0(ori_ori_n2673_), .A1(ori_ori_n467_), .B0(ori_ori_n193_), .B1(ori_ori_n115_), .Y(ori_ori_n2674_));
  OAI210     o2625(.A0(ori_ori_n2674_), .A1(ori_ori_n2672_), .B0(x0), .Y(ori_ori_n2675_));
  NA3        o2626(.A(ori_ori_n405_), .B(ori_ori_n825_), .C(ori_ori_n272_), .Y(ori_ori_n2676_));
  AOI210     o2627(.A0(ori_ori_n2676_), .A1(ori_ori_n721_), .B0(ori_ori_n2224_), .Y(ori_ori_n2677_));
  NA2        o2628(.A(ori_ori_n1141_), .B(ori_ori_n963_), .Y(ori_ori_n2678_));
  NA4        o2629(.A(ori_ori_n684_), .B(ori_ori_n605_), .C(ori_ori_n173_), .D(x3), .Y(ori_ori_n2679_));
  AOI210     o2630(.A0(ori_ori_n2679_), .A1(ori_ori_n2678_), .B0(ori_ori_n499_), .Y(ori_ori_n2680_));
  NO4        o2631(.A(ori_ori_n1428_), .B(ori_ori_n520_), .C(ori_ori_n1244_), .D(ori_ori_n779_), .Y(ori_ori_n2681_));
  OAI220     o2632(.A0(ori_ori_n1799_), .A1(ori_ori_n2311_), .B0(ori_ori_n224_), .B1(ori_ori_n145_), .Y(ori_ori_n2682_));
  NO4        o2633(.A(ori_ori_n2682_), .B(ori_ori_n2681_), .C(ori_ori_n2680_), .D(ori_ori_n2677_), .Y(ori_ori_n2683_));
  NA2        o2634(.A(ori_ori_n2683_), .B(ori_ori_n2675_), .Y(ori_ori_n2684_));
  OAI210     o2635(.A0(ori_ori_n2684_), .A1(ori_ori_n2670_), .B0(ori_ori_n57_), .Y(ori_ori_n2685_));
  AOI210     o2636(.A0(ori_ori_n1839_), .A1(ori_ori_n272_), .B0(ori_ori_n686_), .Y(ori_ori_n2686_));
  OAI210     o2637(.A0(ori_ori_n1778_), .A1(ori_ori_n209_), .B0(ori_ori_n495_), .Y(ori_ori_n2687_));
  OAI210     o2638(.A0(ori_ori_n2687_), .A1(ori_ori_n2686_), .B0(ori_ori_n633_), .Y(ori_ori_n2688_));
  OAI220     o2639(.A0(ori_ori_n1783_), .A1(ori_ori_n272_), .B0(ori_ori_n252_), .B1(ori_ori_n100_), .Y(ori_ori_n2689_));
  NA2        o2640(.A(ori_ori_n1887_), .B(ori_ori_n353_), .Y(ori_ori_n2690_));
  OAI220     o2641(.A0(ori_ori_n2690_), .A1(ori_ori_n641_), .B0(ori_ori_n696_), .B1(ori_ori_n145_), .Y(ori_ori_n2691_));
  AOI210     o2642(.A0(ori_ori_n2689_), .A1(ori_ori_n1004_), .B0(ori_ori_n2691_), .Y(ori_ori_n2692_));
  NA4        o2643(.A(ori_ori_n2692_), .B(ori_ori_n2688_), .C(ori_ori_n2685_), .D(ori_ori_n2654_), .Y(ori39));
  INV        o2644(.A(ori_ori_n81_), .Y(ori_ori_n2696_));
  INV        m0000(.A(x3), .Y(mai_mai_n50_));
  NA2        m0001(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n51_));
  NA2        m0002(.A(x7), .B(x0), .Y(mai_mai_n52_));
  INV        m0003(.A(x1), .Y(mai_mai_n53_));
  NA2        m0004(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  INV        m0005(.A(x8), .Y(mai_mai_n55_));
  INV        m0006(.A(x4), .Y(mai_mai_n56_));
  INV        m0007(.A(x7), .Y(mai_mai_n57_));
  NA2        m0008(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0009(.A(x0), .Y(mai_mai_n59_));
  NA2        m0010(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n60_));
  NA4        m0011(.A(mai_mai_n60_), .B(mai_mai_n58_), .C(mai_mai_n55_), .D(x6), .Y(mai_mai_n61_));
  NA2        m0012(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n62_));
  NO2        m0013(.A(mai_mai_n55_), .B(x6), .Y(mai_mai_n63_));
  NA2        m0014(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n64_));
  NA3        m0015(.A(mai_mai_n64_), .B(mai_mai_n63_), .C(mai_mai_n62_), .Y(mai_mai_n65_));
  AOI210     m0016(.A0(mai_mai_n65_), .A1(mai_mai_n61_), .B0(mai_mai_n54_), .Y(mai_mai_n66_));
  NO2        m0017(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n67_));
  NO2        m0018(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n68_));
  NO2        m0019(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NAi21      m0020(.An(x5), .B(x1), .Y(mai_mai_n70_));
  INV        m0021(.A(x6), .Y(mai_mai_n71_));
  NA2        m0022(.A(mai_mai_n71_), .B(x4), .Y(mai_mai_n72_));
  NO3        m0023(.A(mai_mai_n72_), .B(mai_mai_n70_), .C(mai_mai_n69_), .Y(mai_mai_n73_));
  OAI210     m0024(.A0(mai_mai_n73_), .A1(mai_mai_n66_), .B0(mai_mai_n52_), .Y(mai_mai_n74_));
  NA2        m0025(.A(x7), .B(x4), .Y(mai_mai_n75_));
  NO2        m0026(.A(mai_mai_n75_), .B(x1), .Y(mai_mai_n76_));
  NO2        m0027(.A(mai_mai_n71_), .B(x5), .Y(mai_mai_n77_));
  NO2        m0028(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n78_));
  NA3        m0029(.A(mai_mai_n78_), .B(mai_mai_n77_), .C(mai_mai_n76_), .Y(mai_mai_n79_));
  AOI210     m0030(.A0(mai_mai_n79_), .A1(mai_mai_n74_), .B0(mai_mai_n51_), .Y(mai_mai_n80_));
  NA2        m0031(.A(x5), .B(x3), .Y(mai_mai_n81_));
  NO2        m0032(.A(x6), .B(x0), .Y(mai_mai_n82_));
  NO2        m0033(.A(mai_mai_n82_), .B(x4), .Y(mai_mai_n83_));
  NO2        m0034(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m0035(.A(mai_mai_n71_), .B(mai_mai_n59_), .Y(mai_mai_n85_));
  NO2        m0036(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n86_));
  NA2        m0037(.A(x8), .B(x1), .Y(mai_mai_n87_));
  NO2        m0038(.A(mai_mai_n87_), .B(x7), .Y(mai_mai_n88_));
  INV        m0039(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OR3        m0040(.A(mai_mai_n89_), .B(mai_mai_n86_), .C(mai_mai_n83_), .Y(mai_mai_n90_));
  NO3        m0041(.A(x8), .B(mai_mai_n57_), .C(x6), .Y(mai_mai_n91_));
  NO2        m0042(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n92_));
  NO2        m0043(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n93_));
  NA3        m0044(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n94_));
  AOI210     m0045(.A0(mai_mai_n94_), .A1(mai_mai_n90_), .B0(mai_mai_n81_), .Y(mai_mai_n95_));
  XO2        m0046(.A(x7), .B(x1), .Y(mai_mai_n96_));
  INV        m0047(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NO2        m0048(.A(mai_mai_n97_), .B(x6), .Y(mai_mai_n98_));
  NO2        m0049(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n99_));
  NA2        m0050(.A(mai_mai_n99_), .B(mai_mai_n55_), .Y(mai_mai_n100_));
  NO2        m0051(.A(x6), .B(x5), .Y(mai_mai_n101_));
  NO2        m0052(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n102_));
  NO2        m0053(.A(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  NA2        m0054(.A(x6), .B(x1), .Y(mai_mai_n104_));
  NA2        m0055(.A(mai_mai_n104_), .B(mai_mai_n84_), .Y(mai_mai_n105_));
  NO4        m0056(.A(mai_mai_n105_), .B(mai_mai_n103_), .C(mai_mai_n100_), .D(mai_mai_n98_), .Y(mai_mai_n106_));
  NA2        m0057(.A(x3), .B(x0), .Y(mai_mai_n107_));
  INV        m0058(.A(x5), .Y(mai_mai_n108_));
  NA2        m0059(.A(mai_mai_n71_), .B(mai_mai_n108_), .Y(mai_mai_n109_));
  INV        m0060(.A(x2), .Y(mai_mai_n110_));
  NO2        m0061(.A(mai_mai_n56_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  NA2        m0062(.A(mai_mai_n57_), .B(mai_mai_n108_), .Y(mai_mai_n112_));
  NA3        m0063(.A(mai_mai_n112_), .B(mai_mai_n111_), .C(mai_mai_n109_), .Y(mai_mai_n113_));
  NO3        m0064(.A(mai_mai_n113_), .B(mai_mai_n107_), .C(mai_mai_n53_), .Y(mai_mai_n114_));
  NO4        m0065(.A(mai_mai_n114_), .B(mai_mai_n106_), .C(mai_mai_n95_), .D(mai_mai_n80_), .Y(mai00));
  NO2        m0066(.A(x7), .B(x6), .Y(mai_mai_n116_));
  INV        m0067(.A(mai_mai_n116_), .Y(mai_mai_n117_));
  NO2        m0068(.A(mai_mai_n55_), .B(mai_mai_n53_), .Y(mai_mai_n118_));
  NA2        m0069(.A(mai_mai_n118_), .B(mai_mai_n56_), .Y(mai_mai_n119_));
  NO2        m0070(.A(mai_mai_n119_), .B(mai_mai_n117_), .Y(mai_mai_n120_));
  XN2        m0071(.A(x6), .B(x1), .Y(mai_mai_n121_));
  INV        m0072(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  NO2        m0073(.A(x6), .B(x4), .Y(mai_mai_n123_));
  NA2        m0074(.A(x6), .B(x4), .Y(mai_mai_n124_));
  NAi21      m0075(.An(mai_mai_n123_), .B(mai_mai_n124_), .Y(mai_mai_n125_));
  XN2        m0076(.A(x7), .B(x6), .Y(mai_mai_n126_));
  NO4        m0077(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n122_), .D(x8), .Y(mai_mai_n127_));
  NO2        m0078(.A(x3), .B(mai_mai_n110_), .Y(mai_mai_n128_));
  NA2        m0079(.A(mai_mai_n128_), .B(mai_mai_n108_), .Y(mai_mai_n129_));
  NO2        m0080(.A(mai_mai_n129_), .B(mai_mai_n59_), .Y(mai_mai_n130_));
  OAI210     m0081(.A0(mai_mai_n127_), .A1(mai_mai_n120_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NA2        m0082(.A(x3), .B(mai_mai_n110_), .Y(mai_mai_n132_));
  NO2        m0083(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n133_));
  NA2        m0084(.A(mai_mai_n133_), .B(mai_mai_n56_), .Y(mai_mai_n134_));
  NA2        m0085(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n135_));
  NA2        m0086(.A(mai_mai_n135_), .B(x2), .Y(mai_mai_n136_));
  NA2        m0087(.A(x8), .B(x3), .Y(mai_mai_n137_));
  NA2        m0088(.A(mai_mai_n137_), .B(mai_mai_n75_), .Y(mai_mai_n138_));
  OAI220     m0089(.A0(mai_mai_n138_), .A1(mai_mai_n136_), .B0(mai_mai_n134_), .B1(mai_mai_n132_), .Y(mai_mai_n139_));
  NO2        m0090(.A(x5), .B(x0), .Y(mai_mai_n140_));
  NO2        m0091(.A(x6), .B(x1), .Y(mai_mai_n141_));
  NA3        m0092(.A(mai_mai_n141_), .B(mai_mai_n140_), .C(mai_mai_n139_), .Y(mai_mai_n142_));
  NA2        m0093(.A(x8), .B(mai_mai_n108_), .Y(mai_mai_n143_));
  NA2        m0094(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n144_));
  NAi21      m0095(.An(x7), .B(x2), .Y(mai_mai_n145_));
  NO2        m0096(.A(mai_mai_n145_), .B(x0), .Y(mai_mai_n146_));
  XO2        m0097(.A(x8), .B(x7), .Y(mai_mai_n147_));
  NA2        m0098(.A(mai_mai_n147_), .B(mai_mai_n110_), .Y(mai_mai_n148_));
  NA2        m0099(.A(x6), .B(x5), .Y(mai_mai_n149_));
  NO2        m0100(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n150_));
  NO2        m0101(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n151_));
  NA2        m0102(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  NO3        m0103(.A(mai_mai_n152_), .B(mai_mai_n149_), .C(mai_mai_n148_), .Y(mai_mai_n153_));
  INV        m0104(.A(mai_mai_n153_), .Y(mai_mai_n154_));
  NA3        m0105(.A(mai_mai_n154_), .B(mai_mai_n142_), .C(mai_mai_n131_), .Y(mai01));
  NA2        m0106(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n156_));
  NO2        m0107(.A(x2), .B(x1), .Y(mai_mai_n157_));
  NA2        m0108(.A(x2), .B(x1), .Y(mai_mai_n158_));
  NOi21      m0109(.An(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NA2        m0110(.A(mai_mai_n108_), .B(mai_mai_n53_), .Y(mai_mai_n160_));
  NO2        m0111(.A(mai_mai_n160_), .B(x8), .Y(mai_mai_n161_));
  NAi21      m0112(.An(x8), .B(x1), .Y(mai_mai_n162_));
  NO2        m0113(.A(mai_mai_n162_), .B(x3), .Y(mai_mai_n163_));
  OAI210     m0114(.A0(mai_mai_n163_), .A1(mai_mai_n161_), .B0(mai_mai_n159_), .Y(mai_mai_n164_));
  NO2        m0115(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n165_));
  NO2        m0116(.A(mai_mai_n110_), .B(x1), .Y(mai_mai_n166_));
  NA2        m0117(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  AOI210     m0118(.A0(mai_mai_n167_), .A1(mai_mai_n164_), .B0(mai_mai_n156_), .Y(mai_mai_n168_));
  NAi21      m0119(.An(x7), .B(x0), .Y(mai_mai_n169_));
  NO2        m0120(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n170_));
  NO2        m0121(.A(mai_mai_n81_), .B(x1), .Y(mai_mai_n171_));
  NA2        m0122(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NA2        m0123(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n173_));
  NO2        m0124(.A(mai_mai_n173_), .B(mai_mai_n162_), .Y(mai_mai_n174_));
  NA2        m0125(.A(x8), .B(x5), .Y(mai_mai_n175_));
  NO2        m0126(.A(mai_mai_n175_), .B(mai_mai_n51_), .Y(mai_mai_n176_));
  NO3        m0127(.A(x3), .B(mai_mai_n110_), .C(mai_mai_n53_), .Y(mai_mai_n177_));
  NO3        m0128(.A(mai_mai_n177_), .B(mai_mai_n176_), .C(mai_mai_n174_), .Y(mai_mai_n178_));
  AOI210     m0129(.A0(mai_mai_n178_), .A1(mai_mai_n172_), .B0(mai_mai_n169_), .Y(mai_mai_n179_));
  NO2        m0130(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n180_));
  NO2        m0131(.A(mai_mai_n55_), .B(x0), .Y(mai_mai_n181_));
  NA3        m0132(.A(mai_mai_n108_), .B(mai_mai_n110_), .C(x1), .Y(mai_mai_n182_));
  NO2        m0133(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  NO2        m0134(.A(mai_mai_n87_), .B(mai_mai_n50_), .Y(mai_mai_n184_));
  NA2        m0135(.A(mai_mai_n108_), .B(x0), .Y(mai_mai_n185_));
  NO2        m0136(.A(mai_mai_n185_), .B(x2), .Y(mai_mai_n186_));
  AOI220     m0137(.A0(mai_mai_n186_), .A1(mai_mai_n184_), .B0(mai_mai_n183_), .B1(mai_mai_n180_), .Y(mai_mai_n187_));
  NA2        m0138(.A(x7), .B(mai_mai_n110_), .Y(mai_mai_n188_));
  NA2        m0139(.A(mai_mai_n165_), .B(x8), .Y(mai_mai_n189_));
  NA4        m0140(.A(x5), .B(x3), .C(x1), .D(x0), .Y(mai_mai_n190_));
  AO210      m0141(.A0(mai_mai_n190_), .A1(mai_mai_n189_), .B0(mai_mai_n188_), .Y(mai_mai_n191_));
  NO2        m0142(.A(mai_mai_n158_), .B(mai_mai_n50_), .Y(mai_mai_n192_));
  NAi21      m0143(.An(x1), .B(x2), .Y(mai_mai_n193_));
  NO2        m0144(.A(mai_mai_n173_), .B(mai_mai_n193_), .Y(mai_mai_n194_));
  NA2        m0145(.A(x8), .B(x7), .Y(mai_mai_n195_));
  NO2        m0146(.A(mai_mai_n195_), .B(x0), .Y(mai_mai_n196_));
  OAI210     m0147(.A0(mai_mai_n194_), .A1(mai_mai_n192_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  NA3        m0148(.A(mai_mai_n197_), .B(mai_mai_n191_), .C(mai_mai_n187_), .Y(mai_mai_n198_));
  NO3        m0149(.A(mai_mai_n198_), .B(mai_mai_n179_), .C(mai_mai_n168_), .Y(mai_mai_n199_));
  NA2        m0150(.A(x3), .B(x1), .Y(mai_mai_n200_));
  NA2        m0151(.A(mai_mai_n50_), .B(mai_mai_n110_), .Y(mai_mai_n201_));
  NO2        m0152(.A(mai_mai_n201_), .B(mai_mai_n70_), .Y(mai_mai_n202_));
  OAI210     m0153(.A0(mai_mai_n202_), .A1(mai_mai_n194_), .B0(mai_mai_n67_), .Y(mai_mai_n203_));
  NA2        m0154(.A(mai_mai_n133_), .B(mai_mai_n110_), .Y(mai_mai_n204_));
  OAI210     m0155(.A0(mai_mai_n204_), .A1(mai_mai_n200_), .B0(mai_mai_n203_), .Y(mai_mai_n205_));
  XO2        m0156(.A(x5), .B(x3), .Y(mai_mai_n206_));
  NA2        m0157(.A(mai_mai_n206_), .B(x8), .Y(mai_mai_n207_));
  NA2        m0158(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n208_));
  NA2        m0159(.A(mai_mai_n208_), .B(mai_mai_n137_), .Y(mai_mai_n209_));
  NA2        m0160(.A(x7), .B(mai_mai_n71_), .Y(mai_mai_n210_));
  NO2        m0161(.A(mai_mai_n193_), .B(mai_mai_n210_), .Y(mai_mai_n211_));
  OA210      m0162(.A0(mai_mai_n209_), .A1(mai_mai_n206_), .B0(mai_mai_n211_), .Y(mai_mai_n212_));
  AOI220     m0163(.A0(mai_mai_n212_), .A1(mai_mai_n207_), .B0(mai_mai_n205_), .B1(x0), .Y(mai_mai_n213_));
  OAI210     m0164(.A0(mai_mai_n199_), .A1(mai_mai_n71_), .B0(mai_mai_n213_), .Y(mai_mai_n214_));
  NO2        m0165(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n215_));
  NA4        m0166(.A(mai_mai_n55_), .B(x5), .C(x3), .D(x2), .Y(mai_mai_n216_));
  NA2        m0167(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n217_));
  NA2        m0168(.A(mai_mai_n217_), .B(x2), .Y(mai_mai_n218_));
  NA2        m0169(.A(mai_mai_n55_), .B(x3), .Y(mai_mai_n219_));
  NA4        m0170(.A(mai_mai_n219_), .B(mai_mai_n218_), .C(mai_mai_n206_), .D(mai_mai_n82_), .Y(mai_mai_n220_));
  AOI210     m0171(.A0(mai_mai_n220_), .A1(mai_mai_n216_), .B0(mai_mai_n53_), .Y(mai_mai_n221_));
  NO2        m0172(.A(mai_mai_n110_), .B(mai_mai_n59_), .Y(mai_mai_n222_));
  NA2        m0173(.A(x5), .B(x1), .Y(mai_mai_n223_));
  NO2        m0174(.A(mai_mai_n223_), .B(x6), .Y(mai_mai_n224_));
  NO2        m0175(.A(x3), .B(x1), .Y(mai_mai_n225_));
  AOI210     m0176(.A0(mai_mai_n225_), .A1(mai_mai_n77_), .B0(mai_mai_n224_), .Y(mai_mai_n226_));
  NO2        m0177(.A(mai_mai_n81_), .B(mai_mai_n55_), .Y(mai_mai_n227_));
  NO2        m0178(.A(mai_mai_n104_), .B(mai_mai_n50_), .Y(mai_mai_n228_));
  NO2        m0179(.A(mai_mai_n228_), .B(mai_mai_n227_), .Y(mai_mai_n229_));
  OAI210     m0180(.A0(mai_mai_n226_), .A1(x8), .B0(mai_mai_n229_), .Y(mai_mai_n230_));
  NO2        m0181(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n231_));
  NA2        m0182(.A(mai_mai_n231_), .B(mai_mai_n71_), .Y(mai_mai_n232_));
  NAi21      m0183(.An(x2), .B(x5), .Y(mai_mai_n233_));
  NA2        m0184(.A(x8), .B(x6), .Y(mai_mai_n234_));
  OAI210     m0185(.A0(mai_mai_n234_), .A1(mai_mai_n233_), .B0(mai_mai_n232_), .Y(mai_mai_n235_));
  NA2        m0186(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n236_));
  NO2        m0187(.A(mai_mai_n236_), .B(mai_mai_n59_), .Y(mai_mai_n237_));
  AO220      m0188(.A0(mai_mai_n237_), .A1(mai_mai_n235_), .B0(mai_mai_n230_), .B1(mai_mai_n222_), .Y(mai_mai_n238_));
  OAI210     m0189(.A0(mai_mai_n238_), .A1(mai_mai_n221_), .B0(mai_mai_n215_), .Y(mai_mai_n239_));
  NA2        m0190(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n240_));
  NO2        m0191(.A(mai_mai_n240_), .B(x7), .Y(mai_mai_n241_));
  NO2        m0192(.A(mai_mai_n108_), .B(mai_mai_n53_), .Y(mai_mai_n242_));
  NA2        m0193(.A(mai_mai_n242_), .B(mai_mai_n110_), .Y(mai_mai_n243_));
  AOI210     m0194(.A0(mai_mai_n243_), .A1(mai_mai_n167_), .B0(mai_mai_n59_), .Y(mai_mai_n244_));
  NA2        m0195(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n245_));
  NO2        m0196(.A(mai_mai_n182_), .B(mai_mai_n245_), .Y(mai_mai_n246_));
  OA210      m0197(.A0(mai_mai_n246_), .A1(mai_mai_n244_), .B0(x8), .Y(mai_mai_n247_));
  NO2        m0198(.A(x1), .B(x0), .Y(mai_mai_n248_));
  NA2        m0199(.A(mai_mai_n248_), .B(mai_mai_n110_), .Y(mai_mai_n249_));
  NA2        m0200(.A(mai_mai_n108_), .B(mai_mai_n50_), .Y(mai_mai_n250_));
  XN2        m0201(.A(x3), .B(x2), .Y(mai_mai_n251_));
  NA2        m0202(.A(mai_mai_n251_), .B(mai_mai_n159_), .Y(mai_mai_n252_));
  NO2        m0203(.A(mai_mai_n108_), .B(x0), .Y(mai_mai_n253_));
  NA2        m0204(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n254_));
  NA2        m0205(.A(mai_mai_n254_), .B(mai_mai_n253_), .Y(mai_mai_n255_));
  OAI220     m0206(.A0(mai_mai_n255_), .A1(mai_mai_n252_), .B0(mai_mai_n250_), .B1(mai_mai_n249_), .Y(mai_mai_n256_));
  OAI210     m0207(.A0(mai_mai_n256_), .A1(mai_mai_n247_), .B0(mai_mai_n241_), .Y(mai_mai_n257_));
  NO2        m0208(.A(x7), .B(x1), .Y(mai_mai_n258_));
  NOi21      m0209(.An(x8), .B(x3), .Y(mai_mai_n259_));
  NA2        m0210(.A(mai_mai_n259_), .B(mai_mai_n59_), .Y(mai_mai_n260_));
  NA2        m0211(.A(x5), .B(x0), .Y(mai_mai_n261_));
  NAi21      m0212(.An(mai_mai_n140_), .B(mai_mai_n261_), .Y(mai_mai_n262_));
  NA2        m0213(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n263_));
  OAI210     m0214(.A0(mai_mai_n263_), .A1(mai_mai_n262_), .B0(mai_mai_n260_), .Y(mai_mai_n264_));
  NA3        m0215(.A(mai_mai_n264_), .B(mai_mai_n143_), .C(mai_mai_n258_), .Y(mai_mai_n265_));
  NA2        m0216(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n266_));
  NO2        m0217(.A(mai_mai_n266_), .B(x5), .Y(mai_mai_n267_));
  NO2        m0218(.A(mai_mai_n151_), .B(mai_mai_n71_), .Y(mai_mai_n268_));
  NA2        m0219(.A(x1), .B(x0), .Y(mai_mai_n269_));
  NA2        m0220(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n270_));
  NA2        m0221(.A(mai_mai_n265_), .B(mai_mai_n190_), .Y(mai_mai_n271_));
  NO2        m0222(.A(mai_mai_n108_), .B(x3), .Y(mai_mai_n272_));
  NO2        m0223(.A(mai_mai_n110_), .B(x0), .Y(mai_mai_n273_));
  NA2        m0224(.A(mai_mai_n273_), .B(mai_mai_n272_), .Y(mai_mai_n274_));
  NO2        m0225(.A(mai_mai_n55_), .B(x7), .Y(mai_mai_n275_));
  NA2        m0226(.A(mai_mai_n275_), .B(mai_mai_n141_), .Y(mai_mai_n276_));
  NO3        m0227(.A(x8), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n277_));
  NAi21      m0228(.An(x8), .B(x0), .Y(mai_mai_n278_));
  NAi21      m0229(.An(x1), .B(x3), .Y(mai_mai_n279_));
  NO2        m0230(.A(mai_mai_n279_), .B(mai_mai_n278_), .Y(mai_mai_n280_));
  NO2        m0231(.A(x2), .B(mai_mai_n53_), .Y(mai_mai_n281_));
  AOI210     m0232(.A0(mai_mai_n281_), .A1(mai_mai_n277_), .B0(mai_mai_n280_), .Y(mai_mai_n282_));
  NOi21      m0233(.An(x5), .B(x6), .Y(mai_mai_n283_));
  NO2        m0234(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n284_));
  NA2        m0235(.A(mai_mai_n284_), .B(mai_mai_n283_), .Y(mai_mai_n285_));
  OAI220     m0236(.A0(mai_mai_n285_), .A1(mai_mai_n282_), .B0(mai_mai_n276_), .B1(mai_mai_n274_), .Y(mai_mai_n286_));
  AOI210     m0237(.A0(mai_mai_n271_), .A1(mai_mai_n111_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  NA3        m0238(.A(mai_mai_n287_), .B(mai_mai_n257_), .C(mai_mai_n239_), .Y(mai_mai_n288_));
  AOI210     m0239(.A0(mai_mai_n214_), .A1(mai_mai_n56_), .B0(mai_mai_n288_), .Y(mai02));
  NO2        m0240(.A(x8), .B(mai_mai_n108_), .Y(mai_mai_n290_));
  XN2        m0241(.A(x7), .B(x3), .Y(mai_mai_n291_));
  INV        m0242(.A(mai_mai_n291_), .Y(mai_mai_n292_));
  NO2        m0243(.A(x2), .B(x0), .Y(mai_mai_n293_));
  NA2        m0244(.A(mai_mai_n293_), .B(mai_mai_n71_), .Y(mai_mai_n294_));
  NO2        m0245(.A(mai_mai_n57_), .B(x1), .Y(mai_mai_n295_));
  NO3        m0246(.A(mai_mai_n295_), .B(mai_mai_n294_), .C(mai_mai_n292_), .Y(mai_mai_n296_));
  NA2        m0247(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n297_));
  NO2        m0248(.A(mai_mai_n279_), .B(x6), .Y(mai_mai_n298_));
  XO2        m0249(.A(x7), .B(x0), .Y(mai_mai_n299_));
  NO2        m0250(.A(mai_mai_n299_), .B(mai_mai_n293_), .Y(mai_mai_n300_));
  NA2        m0251(.A(mai_mai_n300_), .B(mai_mai_n298_), .Y(mai_mai_n301_));
  AN2        m0252(.A(x7), .B(x2), .Y(mai_mai_n302_));
  NA2        m0253(.A(mai_mai_n302_), .B(mai_mai_n50_), .Y(mai_mai_n303_));
  OAI210     m0254(.A0(mai_mai_n303_), .A1(mai_mai_n297_), .B0(mai_mai_n301_), .Y(mai_mai_n304_));
  OAI210     m0255(.A0(mai_mai_n304_), .A1(mai_mai_n296_), .B0(mai_mai_n290_), .Y(mai_mai_n305_));
  NAi21      m0256(.An(x8), .B(x6), .Y(mai_mai_n306_));
  NO2        m0257(.A(mai_mai_n108_), .B(mai_mai_n59_), .Y(mai_mai_n307_));
  NA2        m0258(.A(x7), .B(x3), .Y(mai_mai_n308_));
  NO2        m0259(.A(mai_mai_n308_), .B(x2), .Y(mai_mai_n309_));
  NA2        m0260(.A(x2), .B(x0), .Y(mai_mai_n310_));
  NA2        m0261(.A(mai_mai_n110_), .B(mai_mai_n59_), .Y(mai_mai_n311_));
  NA2        m0262(.A(mai_mai_n311_), .B(mai_mai_n310_), .Y(mai_mai_n312_));
  NAi21      m0263(.An(x7), .B(x1), .Y(mai_mai_n313_));
  NO2        m0264(.A(mai_mai_n313_), .B(x3), .Y(mai_mai_n314_));
  AOI220     m0265(.A0(mai_mai_n314_), .A1(mai_mai_n312_), .B0(mai_mai_n309_), .B1(mai_mai_n307_), .Y(mai_mai_n315_));
  NA2        m0266(.A(mai_mai_n281_), .B(mai_mai_n50_), .Y(mai_mai_n316_));
  NA3        m0267(.A(x7), .B(mai_mai_n108_), .C(x0), .Y(mai_mai_n317_));
  NA2        m0268(.A(mai_mai_n273_), .B(mai_mai_n53_), .Y(mai_mai_n318_));
  NA2        m0269(.A(mai_mai_n165_), .B(mai_mai_n57_), .Y(mai_mai_n319_));
  OA220      m0270(.A0(mai_mai_n319_), .A1(mai_mai_n318_), .B0(mai_mai_n317_), .B1(mai_mai_n316_), .Y(mai_mai_n320_));
  AOI210     m0271(.A0(mai_mai_n320_), .A1(mai_mai_n315_), .B0(mai_mai_n306_), .Y(mai_mai_n321_));
  INV        m0272(.A(mai_mai_n299_), .Y(mai_mai_n322_));
  NO2        m0273(.A(x7), .B(mai_mai_n71_), .Y(mai_mai_n323_));
  NA2        m0274(.A(mai_mai_n108_), .B(x3), .Y(mai_mai_n324_));
  NO2        m0275(.A(mai_mai_n324_), .B(mai_mai_n323_), .Y(mai_mai_n325_));
  NA2        m0276(.A(mai_mai_n325_), .B(mai_mai_n322_), .Y(mai_mai_n326_));
  NA2        m0277(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n327_));
  NO2        m0278(.A(mai_mai_n327_), .B(x7), .Y(mai_mai_n328_));
  NA2        m0279(.A(mai_mai_n328_), .B(mai_mai_n283_), .Y(mai_mai_n329_));
  NA2        m0280(.A(mai_mai_n170_), .B(x1), .Y(mai_mai_n330_));
  AOI210     m0281(.A0(mai_mai_n329_), .A1(mai_mai_n326_), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  NO2        m0282(.A(mai_mai_n57_), .B(mai_mai_n50_), .Y(mai_mai_n332_));
  NO2        m0283(.A(mai_mai_n55_), .B(mai_mai_n110_), .Y(mai_mai_n333_));
  NA3        m0284(.A(mai_mai_n333_), .B(mai_mai_n332_), .C(mai_mai_n59_), .Y(mai_mai_n334_));
  NO2        m0285(.A(mai_mai_n160_), .B(x6), .Y(mai_mai_n335_));
  NO2        m0286(.A(mai_mai_n104_), .B(mai_mai_n108_), .Y(mai_mai_n336_));
  NA2        m0287(.A(mai_mai_n57_), .B(mai_mai_n110_), .Y(mai_mai_n337_));
  NO2        m0288(.A(mai_mai_n337_), .B(mai_mai_n270_), .Y(mai_mai_n338_));
  OAI210     m0289(.A0(mai_mai_n336_), .A1(mai_mai_n335_), .B0(mai_mai_n338_), .Y(mai_mai_n339_));
  OAI210     m0290(.A0(mai_mai_n334_), .A1(mai_mai_n104_), .B0(mai_mai_n339_), .Y(mai_mai_n340_));
  NO3        m0291(.A(mai_mai_n340_), .B(mai_mai_n331_), .C(mai_mai_n321_), .Y(mai_mai_n341_));
  AOI210     m0292(.A0(mai_mai_n341_), .A1(mai_mai_n305_), .B0(x4), .Y(mai_mai_n342_));
  NA2        m0293(.A(x8), .B(mai_mai_n71_), .Y(mai_mai_n343_));
  NO2        m0294(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n344_));
  NA3        m0295(.A(mai_mai_n344_), .B(mai_mai_n108_), .C(mai_mai_n53_), .Y(mai_mai_n345_));
  NO2        m0296(.A(x3), .B(x0), .Y(mai_mai_n346_));
  NAi21      m0297(.An(mai_mai_n346_), .B(mai_mai_n107_), .Y(mai_mai_n347_));
  NA2        m0298(.A(x5), .B(x2), .Y(mai_mai_n348_));
  NO2        m0299(.A(mai_mai_n348_), .B(mai_mai_n225_), .Y(mai_mai_n349_));
  AOI210     m0300(.A0(mai_mai_n349_), .A1(mai_mai_n347_), .B0(mai_mai_n246_), .Y(mai_mai_n350_));
  AO210      m0301(.A0(mai_mai_n350_), .A1(mai_mai_n345_), .B0(mai_mai_n343_), .Y(mai_mai_n351_));
  NO2        m0302(.A(mai_mai_n110_), .B(mai_mai_n53_), .Y(mai_mai_n352_));
  NA2        m0303(.A(mai_mai_n352_), .B(x3), .Y(mai_mai_n353_));
  NO2        m0304(.A(mai_mai_n55_), .B(x1), .Y(mai_mai_n354_));
  NA2        m0305(.A(mai_mai_n354_), .B(mai_mai_n110_), .Y(mai_mai_n355_));
  OAI210     m0306(.A0(mai_mai_n355_), .A1(mai_mai_n173_), .B0(mai_mai_n353_), .Y(mai_mai_n356_));
  NAi32      m0307(.An(x3), .Bn(x0), .C(x2), .Y(mai_mai_n357_));
  NO2        m0308(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n358_));
  NAi21      m0309(.An(x6), .B(x5), .Y(mai_mai_n359_));
  NO2        m0310(.A(x2), .B(mai_mai_n59_), .Y(mai_mai_n360_));
  NO4        m0311(.A(mai_mai_n360_), .B(mai_mai_n359_), .C(mai_mai_n162_), .D(mai_mai_n358_), .Y(mai_mai_n361_));
  AOI220     m0312(.A0(mai_mai_n361_), .A1(mai_mai_n357_), .B0(mai_mai_n356_), .B1(mai_mai_n85_), .Y(mai_mai_n362_));
  AOI210     m0313(.A0(mai_mai_n362_), .A1(mai_mai_n351_), .B0(mai_mai_n75_), .Y(mai_mai_n363_));
  NA2        m0314(.A(mai_mai_n354_), .B(mai_mai_n56_), .Y(mai_mai_n364_));
  NO2        m0315(.A(mai_mai_n108_), .B(mai_mai_n50_), .Y(mai_mai_n365_));
  NO2        m0316(.A(mai_mai_n293_), .B(mai_mai_n222_), .Y(mai_mai_n366_));
  XO2        m0317(.A(x7), .B(x2), .Y(mai_mai_n367_));
  INV        m0318(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  XO2        m0319(.A(x6), .B(x2), .Y(mai_mai_n369_));
  NA4        m0320(.A(mai_mai_n369_), .B(mai_mai_n368_), .C(mai_mai_n366_), .D(mai_mai_n365_), .Y(mai_mai_n370_));
  NAi21      m0321(.An(x0), .B(x6), .Y(mai_mai_n371_));
  AOI210     m0322(.A0(mai_mai_n371_), .A1(mai_mai_n145_), .B0(mai_mai_n273_), .Y(mai_mai_n372_));
  XN2        m0323(.A(x7), .B(x5), .Y(mai_mai_n373_));
  NA2        m0324(.A(mai_mai_n373_), .B(mai_mai_n71_), .Y(mai_mai_n374_));
  NA2        m0325(.A(x7), .B(x5), .Y(mai_mai_n375_));
  AOI210     m0326(.A0(mai_mai_n375_), .A1(x6), .B0(mai_mai_n357_), .Y(mai_mai_n376_));
  AOI220     m0327(.A0(mai_mai_n376_), .A1(mai_mai_n374_), .B0(mai_mai_n372_), .B1(mai_mai_n325_), .Y(mai_mai_n377_));
  AOI210     m0328(.A0(mai_mai_n377_), .A1(mai_mai_n370_), .B0(mai_mai_n364_), .Y(mai_mai_n378_));
  NO2        m0329(.A(x8), .B(x6), .Y(mai_mai_n379_));
  NAi21      m0330(.An(mai_mai_n379_), .B(mai_mai_n234_), .Y(mai_mai_n380_));
  NA2        m0331(.A(mai_mai_n108_), .B(x2), .Y(mai_mai_n381_));
  NO2        m0332(.A(mai_mai_n381_), .B(mai_mai_n64_), .Y(mai_mai_n382_));
  NA2        m0333(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n383_));
  NA2        m0334(.A(x4), .B(x2), .Y(mai_mai_n384_));
  NO2        m0335(.A(mai_mai_n384_), .B(mai_mai_n108_), .Y(mai_mai_n385_));
  NAi21      m0336(.An(x1), .B(x6), .Y(mai_mai_n386_));
  NA2        m0337(.A(mai_mai_n346_), .B(mai_mai_n275_), .Y(mai_mai_n387_));
  OAI220     m0338(.A0(mai_mai_n387_), .A1(mai_mai_n386_), .B0(mai_mai_n107_), .B1(mai_mai_n53_), .Y(mai_mai_n388_));
  NA2        m0339(.A(x8), .B(x2), .Y(mai_mai_n389_));
  NO2        m0340(.A(mai_mai_n389_), .B(mai_mai_n50_), .Y(mai_mai_n390_));
  INV        m0341(.A(mai_mai_n224_), .Y(mai_mai_n391_));
  NO2        m0342(.A(mai_mai_n391_), .B(mai_mai_n52_), .Y(mai_mai_n392_));
  AOI220     m0343(.A0(mai_mai_n392_), .A1(mai_mai_n390_), .B0(mai_mai_n388_), .B1(mai_mai_n385_), .Y(mai_mai_n393_));
  INV        m0344(.A(mai_mai_n393_), .Y(mai_mai_n394_));
  NO4        m0345(.A(mai_mai_n394_), .B(mai_mai_n378_), .C(mai_mai_n363_), .D(mai_mai_n342_), .Y(mai03));
  NAi21      m0346(.An(x2), .B(x0), .Y(mai_mai_n396_));
  NO3        m0347(.A(x8), .B(x6), .C(x4), .Y(mai_mai_n397_));
  INV        m0348(.A(mai_mai_n397_), .Y(mai_mai_n398_));
  NO2        m0349(.A(mai_mai_n398_), .B(mai_mai_n396_), .Y(mai_mai_n399_));
  NA2        m0350(.A(mai_mai_n111_), .B(mai_mai_n59_), .Y(mai_mai_n400_));
  NO2        m0351(.A(mai_mai_n400_), .B(mai_mai_n55_), .Y(mai_mai_n401_));
  OAI210     m0352(.A0(mai_mai_n401_), .A1(mai_mai_n399_), .B0(mai_mai_n165_), .Y(mai_mai_n402_));
  NA2        m0353(.A(x3), .B(x2), .Y(mai_mai_n403_));
  NO2        m0354(.A(mai_mai_n162_), .B(x0), .Y(mai_mai_n404_));
  NA2        m0355(.A(x8), .B(x0), .Y(mai_mai_n405_));
  NO2        m0356(.A(mai_mai_n405_), .B(x6), .Y(mai_mai_n406_));
  AOI210     m0357(.A0(mai_mai_n406_), .A1(x5), .B0(mai_mai_n404_), .Y(mai_mai_n407_));
  NO2        m0358(.A(mai_mai_n407_), .B(mai_mai_n403_), .Y(mai_mai_n408_));
  NO2        m0359(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n409_));
  NO2        m0360(.A(x3), .B(x2), .Y(mai_mai_n410_));
  NA2        m0361(.A(mai_mai_n410_), .B(mai_mai_n409_), .Y(mai_mai_n411_));
  NO2        m0362(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n412_));
  NA2        m0363(.A(mai_mai_n412_), .B(x5), .Y(mai_mai_n413_));
  AOI210     m0364(.A0(mai_mai_n413_), .A1(mai_mai_n411_), .B0(mai_mai_n306_), .Y(mai_mai_n414_));
  NA2        m0365(.A(mai_mai_n260_), .B(mai_mai_n175_), .Y(mai_mai_n415_));
  NO2        m0366(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n416_));
  NO2        m0367(.A(mai_mai_n71_), .B(x0), .Y(mai_mai_n417_));
  NO4        m0368(.A(mai_mai_n417_), .B(mai_mai_n416_), .C(x2), .D(mai_mai_n53_), .Y(mai_mai_n418_));
  AO210      m0369(.A0(mai_mai_n418_), .A1(mai_mai_n415_), .B0(mai_mai_n414_), .Y(mai_mai_n419_));
  OAI210     m0370(.A0(mai_mai_n419_), .A1(mai_mai_n408_), .B0(x4), .Y(mai_mai_n420_));
  NO2        m0371(.A(x4), .B(mai_mai_n53_), .Y(mai_mai_n421_));
  NA2        m0372(.A(mai_mai_n421_), .B(mai_mai_n59_), .Y(mai_mai_n422_));
  NO3        m0373(.A(mai_mai_n422_), .B(mai_mai_n234_), .C(x5), .Y(mai_mai_n423_));
  NA2        m0374(.A(x7), .B(mai_mai_n108_), .Y(mai_mai_n424_));
  NO3        m0375(.A(x5), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n425_));
  INV        m0376(.A(mai_mai_n425_), .Y(mai_mai_n426_));
  NO2        m0377(.A(x6), .B(mai_mai_n56_), .Y(mai_mai_n427_));
  NO2        m0378(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n428_));
  NA2        m0379(.A(mai_mai_n428_), .B(mai_mai_n427_), .Y(mai_mai_n429_));
  OAI210     m0380(.A0(mai_mai_n429_), .A1(mai_mai_n426_), .B0(mai_mai_n424_), .Y(mai_mai_n430_));
  AOI210     m0381(.A0(mai_mai_n423_), .A1(x2), .B0(mai_mai_n430_), .Y(mai_mai_n431_));
  AOI220     m0382(.A0(mai_mai_n431_), .A1(mai_mai_n420_), .B0(mai_mai_n402_), .B1(x7), .Y(mai_mai_n432_));
  NA2        m0383(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n433_));
  NO2        m0384(.A(mai_mai_n259_), .B(mai_mai_n110_), .Y(mai_mai_n434_));
  NO2        m0385(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n435_));
  NO3        m0386(.A(mai_mai_n435_), .B(mai_mai_n434_), .C(mai_mai_n149_), .Y(mai_mai_n436_));
  AOI210     m0387(.A0(mai_mai_n209_), .A1(mai_mai_n101_), .B0(mai_mai_n436_), .Y(mai_mai_n437_));
  NO2        m0388(.A(x5), .B(x2), .Y(mai_mai_n438_));
  NO2        m0389(.A(x8), .B(x3), .Y(mai_mai_n439_));
  NA2        m0390(.A(mai_mai_n439_), .B(mai_mai_n438_), .Y(mai_mai_n440_));
  NO2        m0391(.A(mai_mai_n440_), .B(x6), .Y(mai_mai_n441_));
  NA2        m0392(.A(mai_mai_n208_), .B(x2), .Y(mai_mai_n442_));
  NO3        m0393(.A(mai_mai_n439_), .B(mai_mai_n347_), .C(mai_mai_n359_), .Y(mai_mai_n443_));
  AOI210     m0394(.A0(mai_mai_n443_), .A1(mai_mai_n442_), .B0(mai_mai_n441_), .Y(mai_mai_n444_));
  OAI210     m0395(.A0(mai_mai_n437_), .A1(mai_mai_n293_), .B0(mai_mai_n444_), .Y(mai_mai_n445_));
  NA2        m0396(.A(mai_mai_n445_), .B(x4), .Y(mai_mai_n446_));
  NA2        m0397(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n447_));
  NO2        m0398(.A(mai_mai_n447_), .B(x5), .Y(mai_mai_n448_));
  NAi21      m0399(.An(x4), .B(x6), .Y(mai_mai_n449_));
  NO2        m0400(.A(mai_mai_n449_), .B(mai_mai_n51_), .Y(mai_mai_n450_));
  NO2        m0401(.A(mai_mai_n55_), .B(mai_mai_n71_), .Y(mai_mai_n451_));
  NO2        m0402(.A(mai_mai_n50_), .B(mai_mai_n110_), .Y(mai_mai_n452_));
  NO2        m0403(.A(mai_mai_n234_), .B(x0), .Y(mai_mai_n453_));
  NO2        m0404(.A(mai_mai_n359_), .B(x8), .Y(mai_mai_n454_));
  OAI210     m0405(.A0(mai_mai_n454_), .A1(mai_mai_n453_), .B0(mai_mai_n452_), .Y(mai_mai_n455_));
  OAI210     m0406(.A0(mai_mai_n411_), .A1(mai_mai_n451_), .B0(mai_mai_n455_), .Y(mai_mai_n456_));
  AOI220     m0407(.A0(mai_mai_n456_), .A1(mai_mai_n56_), .B0(mai_mai_n450_), .B1(mai_mai_n448_), .Y(mai_mai_n457_));
  AOI210     m0408(.A0(mai_mai_n457_), .A1(mai_mai_n446_), .B0(mai_mai_n433_), .Y(mai_mai_n458_));
  NA2        m0409(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n459_));
  NO2        m0410(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n460_));
  NA2        m0411(.A(mai_mai_n358_), .B(mai_mai_n59_), .Y(mai_mai_n461_));
  OAI220     m0412(.A0(mai_mai_n461_), .A1(mai_mai_n55_), .B0(mai_mai_n201_), .B1(mai_mai_n278_), .Y(mai_mai_n462_));
  NA2        m0413(.A(mai_mai_n462_), .B(mai_mai_n460_), .Y(mai_mai_n463_));
  NO3        m0414(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n464_));
  NA2        m0415(.A(mai_mai_n435_), .B(x5), .Y(mai_mai_n465_));
  NO2        m0416(.A(x8), .B(x5), .Y(mai_mai_n466_));
  NAi21      m0417(.An(mai_mai_n466_), .B(mai_mai_n175_), .Y(mai_mai_n467_));
  OAI210     m0418(.A0(mai_mai_n467_), .A1(mai_mai_n311_), .B0(mai_mai_n465_), .Y(mai_mai_n468_));
  NA2        m0419(.A(mai_mai_n366_), .B(mai_mai_n77_), .Y(mai_mai_n469_));
  NOi21      m0420(.An(x3), .B(x4), .Y(mai_mai_n470_));
  NA2        m0421(.A(mai_mai_n55_), .B(mai_mai_n110_), .Y(mai_mai_n471_));
  NA2        m0422(.A(mai_mai_n471_), .B(mai_mai_n470_), .Y(mai_mai_n472_));
  NO2        m0423(.A(mai_mai_n51_), .B(x6), .Y(mai_mai_n473_));
  NO2        m0424(.A(mai_mai_n149_), .B(mai_mai_n55_), .Y(mai_mai_n474_));
  NO3        m0425(.A(mai_mai_n56_), .B(x2), .C(x0), .Y(mai_mai_n475_));
  AOI220     m0426(.A0(mai_mai_n475_), .A1(mai_mai_n474_), .B0(mai_mai_n473_), .B1(mai_mai_n448_), .Y(mai_mai_n476_));
  OAI210     m0427(.A0(mai_mai_n472_), .A1(mai_mai_n469_), .B0(mai_mai_n476_), .Y(mai_mai_n477_));
  AOI210     m0428(.A0(mai_mai_n468_), .A1(mai_mai_n464_), .B0(mai_mai_n477_), .Y(mai_mai_n478_));
  AOI210     m0429(.A0(mai_mai_n478_), .A1(mai_mai_n463_), .B0(mai_mai_n459_), .Y(mai_mai_n479_));
  NA2        m0430(.A(x7), .B(x1), .Y(mai_mai_n480_));
  NO3        m0431(.A(x5), .B(x4), .C(x2), .Y(mai_mai_n481_));
  AN2        m0432(.A(mai_mai_n481_), .B(mai_mai_n379_), .Y(mai_mai_n482_));
  NO2        m0433(.A(mai_mai_n482_), .B(mai_mai_n385_), .Y(mai_mai_n483_));
  OAI210     m0434(.A0(mai_mai_n379_), .A1(mai_mai_n84_), .B0(mai_mai_n346_), .Y(mai_mai_n484_));
  NO2        m0435(.A(mai_mai_n484_), .B(mai_mai_n483_), .Y(mai_mai_n485_));
  NO2        m0436(.A(x4), .B(mai_mai_n110_), .Y(mai_mai_n486_));
  NA2        m0437(.A(mai_mai_n486_), .B(x6), .Y(mai_mai_n487_));
  NA3        m0438(.A(mai_mai_n108_), .B(x4), .C(mai_mai_n110_), .Y(mai_mai_n488_));
  AOI210     m0439(.A0(mai_mai_n488_), .A1(mai_mai_n487_), .B0(mai_mai_n100_), .Y(mai_mai_n489_));
  NA2        m0440(.A(mai_mai_n470_), .B(mai_mai_n71_), .Y(mai_mai_n490_));
  NA2        m0441(.A(mai_mai_n170_), .B(mai_mai_n59_), .Y(mai_mai_n491_));
  NO2        m0442(.A(mai_mai_n491_), .B(mai_mai_n490_), .Y(mai_mai_n492_));
  NA2        m0443(.A(mai_mai_n452_), .B(x4), .Y(mai_mai_n493_));
  NO3        m0444(.A(mai_mai_n493_), .B(mai_mai_n379_), .C(mai_mai_n417_), .Y(mai_mai_n494_));
  NO4        m0445(.A(mai_mai_n494_), .B(mai_mai_n492_), .C(mai_mai_n489_), .D(mai_mai_n485_), .Y(mai_mai_n495_));
  NA2        m0446(.A(x5), .B(x4), .Y(mai_mai_n496_));
  NO2        m0447(.A(mai_mai_n71_), .B(mai_mai_n53_), .Y(mai_mai_n497_));
  NO3        m0448(.A(x8), .B(x3), .C(x2), .Y(mai_mai_n498_));
  NA3        m0449(.A(mai_mai_n498_), .B(mai_mai_n497_), .C(mai_mai_n59_), .Y(mai_mai_n499_));
  NO3        m0450(.A(x6), .B(x5), .C(x2), .Y(mai_mai_n500_));
  NO2        m0451(.A(mai_mai_n499_), .B(mai_mai_n496_), .Y(mai_mai_n501_));
  NA2        m0452(.A(mai_mai_n71_), .B(x2), .Y(mai_mai_n502_));
  NO3        m0453(.A(x4), .B(x3), .C(mai_mai_n59_), .Y(mai_mai_n503_));
  NA2        m0454(.A(mai_mai_n503_), .B(mai_mai_n231_), .Y(mai_mai_n504_));
  NO3        m0455(.A(mai_mai_n504_), .B(mai_mai_n502_), .C(mai_mai_n96_), .Y(mai_mai_n505_));
  XO2        m0456(.A(x4), .B(x0), .Y(mai_mai_n506_));
  NA2        m0457(.A(mai_mai_n270_), .B(x5), .Y(mai_mai_n507_));
  NO2        m0458(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n508_));
  NO2        m0459(.A(mai_mai_n508_), .B(mai_mai_n63_), .Y(mai_mai_n509_));
  NO4        m0460(.A(mai_mai_n509_), .B(mai_mai_n507_), .C(mai_mai_n506_), .D(mai_mai_n158_), .Y(mai_mai_n510_));
  NO3        m0461(.A(mai_mai_n510_), .B(mai_mai_n505_), .C(mai_mai_n501_), .Y(mai_mai_n511_));
  OAI210     m0462(.A0(mai_mai_n495_), .A1(mai_mai_n480_), .B0(mai_mai_n511_), .Y(mai_mai_n512_));
  NO4        m0463(.A(mai_mai_n512_), .B(mai_mai_n479_), .C(mai_mai_n458_), .D(mai_mai_n432_), .Y(mai04));
  NO2        m0464(.A(x7), .B(x2), .Y(mai_mai_n514_));
  NO2        m0465(.A(x3), .B(mai_mai_n53_), .Y(mai_mai_n515_));
  NO2        m0466(.A(mai_mai_n515_), .B(mai_mai_n151_), .Y(mai_mai_n516_));
  XN2        m0467(.A(x8), .B(x1), .Y(mai_mai_n517_));
  NO2        m0468(.A(mai_mai_n517_), .B(mai_mai_n149_), .Y(mai_mai_n518_));
  NA2        m0469(.A(mai_mai_n518_), .B(mai_mai_n516_), .Y(mai_mai_n519_));
  NA2        m0470(.A(x6), .B(x3), .Y(mai_mai_n520_));
  NO2        m0471(.A(mai_mai_n520_), .B(x5), .Y(mai_mai_n521_));
  NA2        m0472(.A(mai_mai_n71_), .B(x1), .Y(mai_mai_n522_));
  NO2        m0473(.A(mai_mai_n466_), .B(mai_mai_n259_), .Y(mai_mai_n523_));
  NO3        m0474(.A(mai_mai_n523_), .B(mai_mai_n439_), .C(mai_mai_n522_), .Y(mai_mai_n524_));
  AOI210     m0475(.A0(mai_mai_n521_), .A1(mai_mai_n354_), .B0(mai_mai_n524_), .Y(mai_mai_n525_));
  AOI210     m0476(.A0(mai_mai_n525_), .A1(mai_mai_n519_), .B0(x0), .Y(mai_mai_n526_));
  NOi21      m0477(.An(mai_mai_n175_), .B(mai_mai_n466_), .Y(mai_mai_n527_));
  NA2        m0478(.A(mai_mai_n109_), .B(x1), .Y(mai_mai_n528_));
  NO3        m0479(.A(mai_mai_n528_), .B(mai_mai_n527_), .C(mai_mai_n327_), .Y(mai_mai_n529_));
  OAI210     m0480(.A0(mai_mai_n529_), .A1(mai_mai_n526_), .B0(mai_mai_n514_), .Y(mai_mai_n530_));
  NA2        m0481(.A(mai_mai_n137_), .B(mai_mai_n245_), .Y(mai_mai_n531_));
  OR4        m0482(.A(mai_mai_n531_), .B(mai_mai_n380_), .C(mai_mai_n82_), .D(mai_mai_n54_), .Y(mai_mai_n532_));
  OR2        m0483(.A(x6), .B(x0), .Y(mai_mai_n533_));
  NO3        m0484(.A(mai_mai_n533_), .B(x3), .C(x1), .Y(mai_mai_n534_));
  AOI220     m0485(.A0(mai_mai_n534_), .A1(mai_mai_n108_), .B0(mai_mai_n283_), .B1(mai_mai_n277_), .Y(mai_mai_n535_));
  AOI210     m0486(.A0(mai_mai_n535_), .A1(mai_mai_n532_), .B0(mai_mai_n188_), .Y(mai_mai_n536_));
  NA2        m0487(.A(x7), .B(x2), .Y(mai_mai_n537_));
  INV        m0488(.A(mai_mai_n137_), .Y(mai_mai_n538_));
  OAI210     m0489(.A0(mai_mai_n174_), .A1(mai_mai_n538_), .B0(mai_mai_n82_), .Y(mai_mai_n539_));
  NO2        m0490(.A(mai_mai_n324_), .B(mai_mai_n55_), .Y(mai_mai_n540_));
  NO3        m0491(.A(x3), .B(x1), .C(x0), .Y(mai_mai_n541_));
  OR2        m0492(.A(x6), .B(x1), .Y(mai_mai_n542_));
  NA2        m0493(.A(mai_mai_n542_), .B(x0), .Y(mai_mai_n543_));
  AOI220     m0494(.A0(mai_mai_n543_), .A1(mai_mai_n540_), .B0(mai_mai_n541_), .B1(mai_mai_n474_), .Y(mai_mai_n544_));
  AOI210     m0495(.A0(mai_mai_n544_), .A1(mai_mai_n539_), .B0(mai_mai_n537_), .Y(mai_mai_n545_));
  NA2        m0496(.A(mai_mai_n71_), .B(x0), .Y(mai_mai_n546_));
  NOi31      m0497(.An(mai_mai_n349_), .B(mai_mai_n546_), .C(mai_mai_n266_), .Y(mai_mai_n547_));
  NO4        m0498(.A(mai_mai_n547_), .B(mai_mai_n545_), .C(mai_mai_n536_), .D(mai_mai_n56_), .Y(mai_mai_n548_));
  NA2        m0499(.A(mai_mai_n548_), .B(mai_mai_n530_), .Y(mai_mai_n549_));
  NA3        m0500(.A(x8), .B(x7), .C(x0), .Y(mai_mai_n550_));
  INV        m0501(.A(mai_mai_n550_), .Y(mai_mai_n551_));
  AOI210     m0502(.A0(mai_mai_n275_), .A1(mai_mai_n99_), .B0(mai_mai_n551_), .Y(mai_mai_n552_));
  NO2        m0503(.A(mai_mai_n552_), .B(mai_mai_n158_), .Y(mai_mai_n553_));
  NA2        m0504(.A(mai_mai_n435_), .B(mai_mai_n57_), .Y(mai_mai_n554_));
  NO2        m0505(.A(x8), .B(x0), .Y(mai_mai_n555_));
  NA2        m0506(.A(mai_mai_n555_), .B(mai_mai_n368_), .Y(mai_mai_n556_));
  AOI210     m0507(.A0(mai_mai_n556_), .A1(mai_mai_n554_), .B0(mai_mai_n279_), .Y(mai_mai_n557_));
  OAI210     m0508(.A0(mai_mai_n557_), .A1(mai_mai_n553_), .B0(mai_mai_n283_), .Y(mai_mai_n558_));
  NO2        m0509(.A(mai_mai_n71_), .B(mai_mai_n110_), .Y(mai_mai_n559_));
  NO2        m0510(.A(mai_mai_n375_), .B(x8), .Y(mai_mai_n560_));
  NO2        m0511(.A(mai_mai_n560_), .B(mai_mai_n267_), .Y(mai_mai_n561_));
  NO3        m0512(.A(mai_mai_n561_), .B(mai_mai_n383_), .C(mai_mai_n272_), .Y(mai_mai_n562_));
  NO2        m0513(.A(mai_mai_n292_), .B(x8), .Y(mai_mai_n563_));
  OAI210     m0514(.A0(mai_mai_n466_), .A1(mai_mai_n332_), .B0(mai_mai_n248_), .Y(mai_mai_n564_));
  NA2        m0515(.A(mai_mai_n354_), .B(mai_mai_n180_), .Y(mai_mai_n565_));
  OAI220     m0516(.A0(mai_mai_n565_), .A1(mai_mai_n59_), .B0(mai_mai_n564_), .B1(mai_mai_n563_), .Y(mai_mai_n566_));
  OAI210     m0517(.A0(mai_mai_n566_), .A1(mai_mai_n562_), .B0(mai_mai_n559_), .Y(mai_mai_n567_));
  NO2        m0518(.A(x8), .B(x2), .Y(mai_mai_n568_));
  NO2        m0519(.A(mai_mai_n225_), .B(mai_mai_n57_), .Y(mai_mai_n569_));
  NA3        m0520(.A(mai_mai_n569_), .B(mai_mai_n568_), .C(mai_mai_n347_), .Y(mai_mai_n570_));
  NO2        m0521(.A(mai_mai_n249_), .B(mai_mai_n137_), .Y(mai_mai_n571_));
  AOI210     m0522(.A0(mai_mai_n328_), .A1(mai_mai_n166_), .B0(mai_mai_n571_), .Y(mai_mai_n572_));
  AOI210     m0523(.A0(mai_mai_n572_), .A1(mai_mai_n570_), .B0(mai_mai_n109_), .Y(mai_mai_n573_));
  NA2        m0524(.A(mai_mai_n344_), .B(x2), .Y(mai_mai_n574_));
  NO2        m0525(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n575_));
  NA2        m0526(.A(mai_mai_n575_), .B(mai_mai_n63_), .Y(mai_mai_n576_));
  AOI210     m0527(.A0(mai_mai_n574_), .A1(mai_mai_n461_), .B0(mai_mai_n576_), .Y(mai_mai_n577_));
  NA2        m0528(.A(mai_mai_n110_), .B(mai_mai_n53_), .Y(mai_mai_n578_));
  NO2        m0529(.A(mai_mai_n578_), .B(x8), .Y(mai_mai_n579_));
  NA2        m0530(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n580_));
  NO2        m0531(.A(mai_mai_n185_), .B(mai_mai_n580_), .Y(mai_mai_n581_));
  AN2        m0532(.A(mai_mai_n581_), .B(mai_mai_n579_), .Y(mai_mai_n582_));
  NA2        m0533(.A(mai_mai_n409_), .B(mai_mai_n151_), .Y(mai_mai_n583_));
  NO2        m0534(.A(mai_mai_n71_), .B(x2), .Y(mai_mai_n584_));
  NA2        m0535(.A(mai_mai_n584_), .B(mai_mai_n275_), .Y(mai_mai_n585_));
  OAI210     m0536(.A0(mai_mai_n585_), .A1(mai_mai_n583_), .B0(mai_mai_n56_), .Y(mai_mai_n586_));
  NO4        m0537(.A(mai_mai_n586_), .B(mai_mai_n582_), .C(mai_mai_n577_), .D(mai_mai_n573_), .Y(mai_mai_n587_));
  NA3        m0538(.A(mai_mai_n587_), .B(mai_mai_n567_), .C(mai_mai_n558_), .Y(mai_mai_n588_));
  NA2        m0539(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n589_));
  NOi21      m0540(.An(x2), .B(x7), .Y(mai_mai_n590_));
  NO2        m0541(.A(x6), .B(x3), .Y(mai_mai_n591_));
  NA2        m0542(.A(mai_mai_n591_), .B(mai_mai_n590_), .Y(mai_mai_n592_));
  NO2        m0543(.A(x6), .B(mai_mai_n59_), .Y(mai_mai_n593_));
  NO3        m0544(.A(mai_mai_n57_), .B(x2), .C(x1), .Y(mai_mai_n594_));
  NO3        m0545(.A(mai_mai_n57_), .B(x2), .C(x0), .Y(mai_mai_n595_));
  AOI220     m0546(.A0(mai_mai_n595_), .A1(mai_mai_n228_), .B0(mai_mai_n594_), .B1(mai_mai_n593_), .Y(mai_mai_n596_));
  OAI210     m0547(.A0(mai_mai_n592_), .A1(mai_mai_n589_), .B0(mai_mai_n596_), .Y(mai_mai_n597_));
  NO2        m0548(.A(mai_mai_n101_), .B(mai_mai_n53_), .Y(mai_mai_n598_));
  NA2        m0549(.A(mai_mai_n223_), .B(mai_mai_n57_), .Y(mai_mai_n599_));
  OAI210     m0550(.A0(mai_mai_n598_), .A1(mai_mai_n454_), .B0(mai_mai_n599_), .Y(mai_mai_n600_));
  NO3        m0551(.A(mai_mai_n600_), .B(mai_mai_n493_), .C(mai_mai_n59_), .Y(mai_mai_n601_));
  AO210      m0552(.A0(mai_mai_n597_), .A1(mai_mai_n466_), .B0(mai_mai_n601_), .Y(mai_mai_n602_));
  AOI210     m0553(.A0(mai_mai_n588_), .A1(mai_mai_n549_), .B0(mai_mai_n602_), .Y(mai05));
  AOI210     m0554(.A0(mai_mai_n165_), .A1(mai_mai_n55_), .B0(mai_mai_n508_), .Y(mai_mai_n604_));
  OR2        m0555(.A(mai_mai_n604_), .B(mai_mai_n57_), .Y(mai_mai_n605_));
  NO2        m0556(.A(x7), .B(mai_mai_n108_), .Y(mai_mai_n606_));
  NO2        m0557(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n607_));
  NA2        m0558(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n608_));
  NO2        m0559(.A(mai_mai_n608_), .B(mai_mai_n580_), .Y(mai_mai_n609_));
  AOI210     m0560(.A0(mai_mai_n607_), .A1(mai_mai_n606_), .B0(mai_mai_n609_), .Y(mai_mai_n610_));
  AOI210     m0561(.A0(mai_mai_n610_), .A1(mai_mai_n605_), .B0(mai_mai_n110_), .Y(mai_mai_n611_));
  NO2        m0562(.A(x7), .B(x4), .Y(mai_mai_n612_));
  NO2        m0563(.A(mai_mai_n64_), .B(mai_mai_n55_), .Y(mai_mai_n613_));
  NO2        m0564(.A(mai_mai_n201_), .B(x5), .Y(mai_mai_n614_));
  NA2        m0565(.A(mai_mai_n108_), .B(mai_mai_n110_), .Y(mai_mai_n615_));
  NO2        m0566(.A(mai_mai_n615_), .B(mai_mai_n219_), .Y(mai_mai_n616_));
  AO220      m0567(.A0(mai_mai_n616_), .A1(mai_mai_n612_), .B0(mai_mai_n614_), .B1(mai_mai_n613_), .Y(mai_mai_n617_));
  OAI210     m0568(.A0(mai_mai_n617_), .A1(mai_mai_n611_), .B0(mai_mai_n497_), .Y(mai_mai_n618_));
  NO2        m0569(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n619_));
  NA2        m0570(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n620_));
  NO2        m0571(.A(mai_mai_n108_), .B(mai_mai_n110_), .Y(mai_mai_n621_));
  NA2        m0572(.A(mai_mai_n621_), .B(x7), .Y(mai_mai_n622_));
  NA2        m0573(.A(mai_mai_n438_), .B(mai_mai_n258_), .Y(mai_mai_n623_));
  AOI210     m0574(.A0(mai_mai_n623_), .A1(mai_mai_n622_), .B0(mai_mai_n620_), .Y(mai_mai_n624_));
  NA2        m0575(.A(mai_mai_n108_), .B(x4), .Y(mai_mai_n625_));
  XO2        m0576(.A(x7), .B(x5), .Y(mai_mai_n626_));
  NO2        m0577(.A(mai_mai_n626_), .B(mai_mai_n53_), .Y(mai_mai_n627_));
  NA3        m0578(.A(mai_mai_n627_), .B(mai_mai_n625_), .C(mai_mai_n333_), .Y(mai_mai_n628_));
  NO2        m0579(.A(mai_mai_n108_), .B(x2), .Y(mai_mai_n629_));
  NO2        m0580(.A(mai_mai_n75_), .B(mai_mai_n55_), .Y(mai_mai_n630_));
  NA2        m0581(.A(mai_mai_n630_), .B(mai_mai_n629_), .Y(mai_mai_n631_));
  NA2        m0582(.A(mai_mai_n631_), .B(mai_mai_n628_), .Y(mai_mai_n632_));
  OAI210     m0583(.A0(mai_mai_n632_), .A1(mai_mai_n624_), .B0(mai_mai_n619_), .Y(mai_mai_n633_));
  NO2        m0584(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n634_));
  NO2        m0585(.A(mai_mai_n195_), .B(x4), .Y(mai_mai_n635_));
  NO2        m0586(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n636_));
  XO2        m0587(.A(x5), .B(x2), .Y(mai_mai_n637_));
  NO3        m0588(.A(x8), .B(x7), .C(mai_mai_n110_), .Y(mai_mai_n638_));
  AN2        m0589(.A(mai_mai_n637_), .B(mai_mai_n635_), .Y(mai_mai_n639_));
  NA3        m0590(.A(mai_mai_n639_), .B(mai_mai_n634_), .C(mai_mai_n53_), .Y(mai_mai_n640_));
  NA2        m0591(.A(mai_mai_n272_), .B(mai_mai_n590_), .Y(mai_mai_n641_));
  NOi21      m0592(.An(x4), .B(x1), .Y(mai_mai_n642_));
  NA2        m0593(.A(mai_mai_n642_), .B(mai_mai_n63_), .Y(mai_mai_n643_));
  NA2        m0594(.A(x4), .B(x1), .Y(mai_mai_n644_));
  NO2        m0595(.A(mai_mai_n644_), .B(mai_mai_n50_), .Y(mai_mai_n645_));
  AOI210     m0596(.A0(mai_mai_n645_), .A1(mai_mai_n621_), .B0(mai_mai_n59_), .Y(mai_mai_n646_));
  OA210      m0597(.A0(mai_mai_n643_), .A1(mai_mai_n641_), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  NA4        m0598(.A(mai_mai_n647_), .B(mai_mai_n640_), .C(mai_mai_n633_), .D(mai_mai_n618_), .Y(mai_mai_n648_));
  NA2        m0599(.A(mai_mai_n634_), .B(mai_mai_n56_), .Y(mai_mai_n649_));
  NA2        m0600(.A(mai_mai_n568_), .B(mai_mai_n606_), .Y(mai_mai_n650_));
  NO2        m0601(.A(mai_mai_n650_), .B(mai_mai_n649_), .Y(mai_mai_n651_));
  NA2        m0602(.A(mai_mai_n275_), .B(mai_mai_n123_), .Y(mai_mai_n652_));
  OAI210     m0603(.A0(mai_mai_n652_), .A1(mai_mai_n167_), .B0(mai_mai_n59_), .Y(mai_mai_n653_));
  NA2        m0604(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n654_));
  AOI210     m0605(.A0(mai_mai_n654_), .A1(x3), .B0(mai_mai_n91_), .Y(mai_mai_n655_));
  NA2        m0606(.A(mai_mai_n636_), .B(mai_mai_n157_), .Y(mai_mai_n656_));
  NO3        m0607(.A(mai_mai_n656_), .B(mai_mai_n655_), .C(mai_mai_n428_), .Y(mai_mai_n657_));
  NA2        m0608(.A(mai_mai_n284_), .B(mai_mai_n71_), .Y(mai_mai_n658_));
  NO2        m0609(.A(mai_mai_n389_), .B(x3), .Y(mai_mai_n659_));
  NA2        m0610(.A(mai_mai_n659_), .B(mai_mai_n242_), .Y(mai_mai_n660_));
  NO2        m0611(.A(mai_mai_n428_), .B(mai_mai_n635_), .Y(mai_mai_n661_));
  NO2        m0612(.A(mai_mai_n470_), .B(mai_mai_n108_), .Y(mai_mai_n662_));
  NO2        m0613(.A(mai_mai_n578_), .B(x6), .Y(mai_mai_n663_));
  NA2        m0614(.A(mai_mai_n663_), .B(mai_mai_n662_), .Y(mai_mai_n664_));
  OAI220     m0615(.A0(mai_mai_n664_), .A1(mai_mai_n661_), .B0(mai_mai_n660_), .B1(mai_mai_n658_), .Y(mai_mai_n665_));
  NO4        m0616(.A(mai_mai_n665_), .B(mai_mai_n657_), .C(mai_mai_n653_), .D(mai_mai_n651_), .Y(mai_mai_n666_));
  NA2        m0617(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n667_));
  NO2        m0618(.A(mai_mai_n667_), .B(x1), .Y(mai_mai_n668_));
  NA2        m0619(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n669_));
  NO2        m0620(.A(mai_mai_n669_), .B(mai_mai_n132_), .Y(mai_mai_n670_));
  NA2        m0621(.A(x8), .B(x4), .Y(mai_mai_n671_));
  NO2        m0622(.A(x8), .B(x4), .Y(mai_mai_n672_));
  NAi21      m0623(.An(mai_mai_n672_), .B(mai_mai_n671_), .Y(mai_mai_n673_));
  NAi21      m0624(.An(mai_mai_n568_), .B(mai_mai_n389_), .Y(mai_mai_n674_));
  NO4        m0625(.A(mai_mai_n674_), .B(mai_mai_n673_), .C(mai_mai_n428_), .D(mai_mai_n71_), .Y(mai_mai_n675_));
  OAI210     m0626(.A0(mai_mai_n675_), .A1(mai_mai_n670_), .B0(mai_mai_n668_), .Y(mai_mai_n676_));
  NO3        m0627(.A(x8), .B(mai_mai_n108_), .C(x4), .Y(mai_mai_n677_));
  INV        m0628(.A(mai_mai_n677_), .Y(mai_mai_n678_));
  NO2        m0629(.A(mai_mai_n678_), .B(mai_mai_n110_), .Y(mai_mai_n679_));
  NO2        m0630(.A(x5), .B(x4), .Y(mai_mai_n680_));
  NA3        m0631(.A(mai_mai_n680_), .B(mai_mai_n63_), .C(mai_mai_n110_), .Y(mai_mai_n681_));
  NO2        m0632(.A(x6), .B(mai_mai_n110_), .Y(mai_mai_n682_));
  NA2        m0633(.A(mai_mai_n669_), .B(mai_mai_n682_), .Y(mai_mai_n683_));
  OAI210     m0634(.A0(mai_mai_n683_), .A1(mai_mai_n527_), .B0(mai_mai_n681_), .Y(mai_mai_n684_));
  OAI210     m0635(.A0(mai_mai_n684_), .A1(mai_mai_n679_), .B0(mai_mai_n314_), .Y(mai_mai_n685_));
  NA3        m0636(.A(mai_mai_n685_), .B(mai_mai_n676_), .C(mai_mai_n666_), .Y(mai_mai_n686_));
  OR2        m0637(.A(x4), .B(x1), .Y(mai_mai_n687_));
  NO2        m0638(.A(mai_mai_n687_), .B(x3), .Y(mai_mai_n688_));
  NA2        m0639(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n689_));
  NO3        m0640(.A(mai_mai_n373_), .B(mai_mai_n689_), .C(x6), .Y(mai_mai_n690_));
  AOI220     m0641(.A0(mai_mai_n690_), .A1(mai_mai_n688_), .B0(mai_mai_n686_), .B1(mai_mai_n648_), .Y(mai06));
  NA2        m0642(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n692_));
  NA2        m0643(.A(x6), .B(mai_mai_n110_), .Y(mai_mai_n693_));
  NA2        m0644(.A(mai_mai_n693_), .B(mai_mai_n55_), .Y(mai_mai_n694_));
  NA2        m0645(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n695_));
  NO2        m0646(.A(mai_mai_n695_), .B(mai_mai_n118_), .Y(mai_mai_n696_));
  NA3        m0647(.A(mai_mai_n696_), .B(mai_mai_n694_), .C(mai_mai_n502_), .Y(mai_mai_n697_));
  NO2        m0648(.A(mai_mai_n389_), .B(x0), .Y(mai_mai_n698_));
  NA2        m0649(.A(mai_mai_n343_), .B(x2), .Y(mai_mai_n699_));
  NOi21      m0650(.An(x6), .B(x8), .Y(mai_mai_n700_));
  NO2        m0651(.A(mai_mai_n700_), .B(x2), .Y(mai_mai_n701_));
  NO3        m0652(.A(mai_mai_n701_), .B(mai_mai_n70_), .C(mai_mai_n59_), .Y(mai_mai_n702_));
  AOI220     m0653(.A0(mai_mai_n702_), .A1(mai_mai_n699_), .B0(mai_mai_n698_), .B1(mai_mai_n335_), .Y(mai_mai_n703_));
  AOI210     m0654(.A0(mai_mai_n703_), .A1(mai_mai_n697_), .B0(mai_mai_n692_), .Y(mai_mai_n704_));
  NA2        m0655(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n705_));
  NA2        m0656(.A(mai_mai_n371_), .B(mai_mai_n359_), .Y(mai_mai_n706_));
  NO2        m0657(.A(mai_mai_n71_), .B(mai_mai_n108_), .Y(mai_mai_n707_));
  NO2        m0658(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n708_));
  NO4        m0659(.A(mai_mai_n708_), .B(mai_mai_n689_), .C(mai_mai_n707_), .D(mai_mai_n497_), .Y(mai_mai_n709_));
  AOI220     m0660(.A0(mai_mai_n709_), .A1(mai_mai_n706_), .B0(mai_mai_n425_), .B1(mai_mai_n63_), .Y(mai_mai_n710_));
  NO2        m0661(.A(mai_mai_n710_), .B(mai_mai_n705_), .Y(mai_mai_n711_));
  NO2        m0662(.A(mai_mai_n54_), .B(x0), .Y(mai_mai_n712_));
  NA2        m0663(.A(x4), .B(x3), .Y(mai_mai_n713_));
  OAI210     m0664(.A0(mai_mai_n713_), .A1(x8), .B0(mai_mai_n520_), .Y(mai_mai_n714_));
  NA2        m0665(.A(mai_mai_n714_), .B(mai_mai_n712_), .Y(mai_mai_n715_));
  NO2        m0666(.A(mai_mai_n104_), .B(mai_mai_n56_), .Y(mai_mai_n716_));
  NA3        m0667(.A(mai_mai_n716_), .B(mai_mai_n259_), .C(mai_mai_n409_), .Y(mai_mai_n717_));
  AOI210     m0668(.A0(mai_mai_n717_), .A1(mai_mai_n715_), .B0(x2), .Y(mai_mai_n718_));
  INV        m0669(.A(mai_mai_n385_), .Y(mai_mai_n719_));
  NO2        m0670(.A(mai_mai_n412_), .B(x8), .Y(mai_mai_n720_));
  NO2        m0671(.A(mai_mai_n260_), .B(mai_mai_n522_), .Y(mai_mai_n721_));
  AOI210     m0672(.A0(mai_mai_n720_), .A1(mai_mai_n268_), .B0(mai_mai_n721_), .Y(mai_mai_n722_));
  NO2        m0673(.A(x5), .B(x3), .Y(mai_mai_n723_));
  NA3        m0674(.A(mai_mai_n555_), .B(mai_mai_n723_), .C(x1), .Y(mai_mai_n724_));
  OR2        m0675(.A(mai_mai_n724_), .B(mai_mai_n502_), .Y(mai_mai_n725_));
  OAI210     m0676(.A0(mai_mai_n722_), .A1(mai_mai_n719_), .B0(mai_mai_n725_), .Y(mai_mai_n726_));
  OR4        m0677(.A(mai_mai_n726_), .B(mai_mai_n718_), .C(mai_mai_n711_), .D(mai_mai_n704_), .Y(mai_mai_n727_));
  NA2        m0678(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n728_));
  NO2        m0679(.A(mai_mai_n621_), .B(mai_mai_n59_), .Y(mai_mai_n729_));
  NA2        m0680(.A(mai_mai_n729_), .B(mai_mai_n634_), .Y(mai_mai_n730_));
  NO2        m0681(.A(mai_mai_n173_), .B(x6), .Y(mai_mai_n731_));
  NA2        m0682(.A(mai_mai_n731_), .B(mai_mai_n293_), .Y(mai_mai_n732_));
  AOI210     m0683(.A0(mai_mai_n732_), .A1(mai_mai_n730_), .B0(mai_mai_n728_), .Y(mai_mai_n733_));
  AN2        m0684(.A(mai_mai_n475_), .B(mai_mai_n325_), .Y(mai_mai_n734_));
  OAI210     m0685(.A0(mai_mai_n734_), .A1(mai_mai_n733_), .B0(mai_mai_n354_), .Y(mai_mai_n735_));
  NO2        m0686(.A(mai_mai_n310_), .B(mai_mai_n108_), .Y(mai_mai_n736_));
  NO2        m0687(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n737_));
  NA2        m0688(.A(mai_mai_n737_), .B(mai_mai_n71_), .Y(mai_mai_n738_));
  NO2        m0689(.A(mai_mai_n738_), .B(mai_mai_n254_), .Y(mai_mai_n739_));
  NO2        m0690(.A(mai_mai_n71_), .B(x3), .Y(mai_mai_n740_));
  NA3        m0691(.A(mai_mai_n740_), .B(mai_mai_n575_), .C(mai_mai_n56_), .Y(mai_mai_n741_));
  NO2        m0692(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n742_));
  NA2        m0693(.A(mai_mai_n184_), .B(mai_mai_n742_), .Y(mai_mai_n743_));
  NA3        m0694(.A(mai_mai_n607_), .B(mai_mai_n332_), .C(mai_mai_n71_), .Y(mai_mai_n744_));
  NA3        m0695(.A(mai_mai_n744_), .B(mai_mai_n743_), .C(mai_mai_n741_), .Y(mai_mai_n745_));
  OR3        m0696(.A(mai_mai_n745_), .B(mai_mai_n739_), .C(mai_mai_n645_), .Y(mai_mai_n746_));
  NA2        m0697(.A(mai_mai_n746_), .B(mai_mai_n736_), .Y(mai_mai_n747_));
  NA2        m0698(.A(mai_mai_n712_), .B(mai_mai_n634_), .Y(mai_mai_n748_));
  NA4        m0699(.A(mai_mai_n269_), .B(mai_mai_n591_), .C(mai_mai_n223_), .D(mai_mai_n261_), .Y(mai_mai_n749_));
  NA2        m0700(.A(mai_mai_n486_), .B(mai_mai_n67_), .Y(mai_mai_n750_));
  AOI210     m0701(.A0(mai_mai_n749_), .A1(mai_mai_n748_), .B0(mai_mai_n750_), .Y(mai_mai_n751_));
  NA2        m0702(.A(x7), .B(x6), .Y(mai_mai_n752_));
  NA3        m0703(.A(x2), .B(x1), .C(x0), .Y(mai_mai_n753_));
  NO3        m0704(.A(mai_mai_n753_), .B(mai_mai_n752_), .C(mai_mai_n604_), .Y(mai_mai_n754_));
  NA2        m0705(.A(mai_mai_n498_), .B(mai_mai_n150_), .Y(mai_mai_n755_));
  NO2        m0706(.A(x5), .B(x1), .Y(mai_mai_n756_));
  NA2        m0707(.A(mai_mai_n756_), .B(mai_mai_n742_), .Y(mai_mai_n757_));
  NA2        m0708(.A(x4), .B(x0), .Y(mai_mai_n758_));
  NO3        m0709(.A(mai_mai_n57_), .B(x6), .C(x2), .Y(mai_mai_n759_));
  NA2        m0710(.A(mai_mai_n759_), .B(mai_mai_n227_), .Y(mai_mai_n760_));
  OAI220     m0711(.A0(mai_mai_n760_), .A1(mai_mai_n758_), .B0(mai_mai_n757_), .B1(mai_mai_n755_), .Y(mai_mai_n761_));
  NO3        m0712(.A(mai_mai_n761_), .B(mai_mai_n754_), .C(mai_mai_n751_), .Y(mai_mai_n762_));
  NA3        m0713(.A(mai_mai_n762_), .B(mai_mai_n747_), .C(mai_mai_n735_), .Y(mai_mai_n763_));
  AOI210     m0714(.A0(mai_mai_n727_), .A1(mai_mai_n57_), .B0(mai_mai_n763_), .Y(mai07));
  NA2        m0715(.A(mai_mai_n108_), .B(mai_mai_n59_), .Y(mai_mai_n765_));
  NOi21      m0716(.An(mai_mai_n752_), .B(mai_mai_n116_), .Y(mai_mai_n766_));
  NO3        m0717(.A(mai_mai_n57_), .B(x5), .C(x1), .Y(mai_mai_n767_));
  NA2        m0718(.A(mai_mai_n767_), .B(mai_mai_n379_), .Y(mai_mai_n768_));
  NO2        m0719(.A(mai_mai_n57_), .B(mai_mai_n71_), .Y(mai_mai_n769_));
  NO2        m0720(.A(mai_mai_n156_), .B(mai_mai_n109_), .Y(mai_mai_n770_));
  AOI210     m0721(.A0(mai_mai_n769_), .A1(mai_mai_n92_), .B0(mai_mai_n770_), .Y(mai_mai_n771_));
  OAI220     m0722(.A0(mai_mai_n771_), .A1(mai_mai_n137_), .B0(mai_mai_n768_), .B1(mai_mai_n327_), .Y(mai_mai_n772_));
  NA2        m0723(.A(mai_mai_n772_), .B(x2), .Y(mai_mai_n773_));
  NAi21      m0724(.An(mai_mai_n157_), .B(mai_mai_n158_), .Y(mai_mai_n774_));
  NA3        m0725(.A(mai_mai_n774_), .B(mai_mai_n91_), .C(x3), .Y(mai_mai_n775_));
  NO3        m0726(.A(mai_mai_n55_), .B(x3), .C(x1), .Y(mai_mai_n776_));
  NO2        m0727(.A(mai_mai_n515_), .B(x2), .Y(mai_mai_n777_));
  AOI210     m0728(.A0(mai_mai_n777_), .A1(mai_mai_n517_), .B0(mai_mai_n776_), .Y(mai_mai_n778_));
  OAI210     m0729(.A0(mai_mai_n778_), .A1(mai_mai_n654_), .B0(mai_mai_n775_), .Y(mai_mai_n779_));
  NO2        m0730(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n780_));
  NA2        m0731(.A(mai_mai_n780_), .B(mai_mai_n59_), .Y(mai_mai_n781_));
  NA2        m0732(.A(mai_mai_n360_), .B(mai_mai_n354_), .Y(mai_mai_n782_));
  NO2        m0733(.A(x7), .B(x3), .Y(mai_mai_n783_));
  NA2        m0734(.A(mai_mai_n783_), .B(mai_mai_n101_), .Y(mai_mai_n784_));
  AOI210     m0735(.A0(mai_mai_n782_), .A1(mai_mai_n781_), .B0(mai_mai_n784_), .Y(mai_mai_n785_));
  AOI210     m0736(.A0(mai_mai_n779_), .A1(mai_mai_n253_), .B0(mai_mai_n785_), .Y(mai_mai_n786_));
  AOI210     m0737(.A0(mai_mai_n786_), .A1(mai_mai_n773_), .B0(x4), .Y(mai_mai_n787_));
  NO2        m0738(.A(mai_mai_n600_), .B(mai_mai_n110_), .Y(mai_mai_n788_));
  XO2        m0739(.A(x5), .B(x1), .Y(mai_mai_n789_));
  NO4        m0740(.A(mai_mai_n789_), .B(mai_mai_n166_), .C(mai_mai_n210_), .D(mai_mai_n55_), .Y(mai_mai_n790_));
  OAI210     m0741(.A0(mai_mai_n790_), .A1(mai_mai_n788_), .B0(mai_mai_n416_), .Y(mai_mai_n791_));
  NO3        m0742(.A(mai_mai_n50_), .B(x2), .C(x0), .Y(mai_mai_n792_));
  NO2        m0743(.A(mai_mai_n313_), .B(mai_mai_n108_), .Y(mai_mai_n793_));
  NA2        m0744(.A(x6), .B(x0), .Y(mai_mai_n794_));
  NO2        m0745(.A(mai_mai_n689_), .B(mai_mai_n794_), .Y(mai_mai_n795_));
  NO2        m0746(.A(mai_mai_n789_), .B(mai_mai_n700_), .Y(mai_mai_n796_));
  OAI210     m0747(.A0(mai_mai_n756_), .A1(mai_mai_n63_), .B0(mai_mai_n57_), .Y(mai_mai_n797_));
  OAI210     m0748(.A0(mai_mai_n797_), .A1(mai_mai_n796_), .B0(mai_mai_n768_), .Y(mai_mai_n798_));
  AOI220     m0749(.A0(mai_mai_n798_), .A1(mai_mai_n792_), .B0(mai_mai_n795_), .B1(mai_mai_n793_), .Y(mai_mai_n799_));
  AOI210     m0750(.A0(mai_mai_n799_), .A1(mai_mai_n791_), .B0(mai_mai_n56_), .Y(mai_mai_n800_));
  NOi21      m0751(.An(mai_mai_n234_), .B(mai_mai_n379_), .Y(mai_mai_n801_));
  NO3        m0752(.A(mai_mai_n801_), .B(mai_mai_n243_), .C(mai_mai_n67_), .Y(mai_mai_n802_));
  NO2        m0753(.A(mai_mai_n193_), .B(mai_mai_n71_), .Y(mai_mai_n803_));
  NO2        m0754(.A(mai_mai_n313_), .B(x6), .Y(mai_mai_n804_));
  AO220      m0755(.A0(mai_mai_n804_), .A1(mai_mai_n333_), .B0(mai_mai_n803_), .B1(mai_mai_n560_), .Y(mai_mai_n805_));
  OAI210     m0756(.A0(mai_mai_n805_), .A1(mai_mai_n802_), .B0(mai_mai_n59_), .Y(mai_mai_n806_));
  NA2        m0757(.A(mai_mai_n92_), .B(mai_mai_n71_), .Y(mai_mai_n807_));
  NO2        m0758(.A(mai_mai_n807_), .B(mai_mai_n650_), .Y(mai_mai_n808_));
  NAi21      m0759(.An(x8), .B(x7), .Y(mai_mai_n809_));
  NA2        m0760(.A(mai_mai_n801_), .B(mai_mai_n809_), .Y(mai_mai_n810_));
  NA2        m0761(.A(mai_mai_n409_), .B(mai_mai_n110_), .Y(mai_mai_n811_));
  NO2        m0762(.A(mai_mai_n700_), .B(x1), .Y(mai_mai_n812_));
  NO3        m0763(.A(mai_mai_n812_), .B(mai_mai_n811_), .C(mai_mai_n575_), .Y(mai_mai_n813_));
  AOI210     m0764(.A0(mai_mai_n813_), .A1(mai_mai_n810_), .B0(mai_mai_n808_), .Y(mai_mai_n814_));
  AOI210     m0765(.A0(mai_mai_n814_), .A1(mai_mai_n806_), .B0(mai_mai_n144_), .Y(mai_mai_n815_));
  NO2        m0766(.A(x8), .B(x7), .Y(mai_mai_n816_));
  NO2        m0767(.A(mai_mai_n816_), .B(x3), .Y(mai_mai_n817_));
  NA3        m0768(.A(mai_mai_n817_), .B(mai_mai_n368_), .C(x1), .Y(mai_mai_n818_));
  NO2        m0769(.A(x8), .B(mai_mai_n110_), .Y(mai_mai_n819_));
  AOI220     m0770(.A0(mai_mai_n332_), .A1(mai_mai_n354_), .B0(mai_mai_n819_), .B1(mai_mai_n258_), .Y(mai_mai_n820_));
  NO2        m0771(.A(mai_mai_n71_), .B(x4), .Y(mai_mai_n821_));
  NA2        m0772(.A(mai_mai_n821_), .B(mai_mai_n307_), .Y(mai_mai_n822_));
  AOI210     m0773(.A0(mai_mai_n820_), .A1(mai_mai_n818_), .B0(mai_mai_n822_), .Y(mai_mai_n823_));
  NO4        m0774(.A(mai_mai_n823_), .B(mai_mai_n815_), .C(mai_mai_n800_), .D(mai_mai_n787_), .Y(mai08));
  NA2        m0775(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n825_));
  XN2        m0776(.A(x5), .B(x4), .Y(mai_mai_n826_));
  INV        m0777(.A(mai_mai_n826_), .Y(mai_mai_n827_));
  AOI220     m0778(.A0(mai_mai_n827_), .A1(mai_mai_n360_), .B0(mai_mai_n140_), .B1(mai_mai_n56_), .Y(mai_mai_n828_));
  NO2        m0779(.A(mai_mai_n245_), .B(mai_mai_n108_), .Y(mai_mai_n829_));
  AOI210     m0780(.A0(mai_mai_n829_), .A1(mai_mai_n281_), .B0(mai_mai_n194_), .Y(mai_mai_n830_));
  OAI220     m0781(.A0(mai_mai_n830_), .A1(x4), .B0(mai_mai_n828_), .B1(mai_mai_n825_), .Y(mai_mai_n831_));
  NA2        m0782(.A(mai_mai_n831_), .B(mai_mai_n275_), .Y(mai_mai_n832_));
  AOI210     m0783(.A0(mai_mai_n274_), .A1(mai_mai_n811_), .B0(mai_mai_n620_), .Y(mai_mai_n833_));
  NA2        m0784(.A(mai_mai_n615_), .B(mai_mai_n173_), .Y(mai_mai_n834_));
  OAI220     m0785(.A0(mai_mai_n834_), .A1(mai_mai_n669_), .B0(mai_mai_n488_), .B1(mai_mai_n50_), .Y(mai_mai_n835_));
  AO210      m0786(.A0(mai_mai_n835_), .A1(mai_mai_n347_), .B0(mai_mai_n833_), .Y(mai_mai_n836_));
  NA2        m0787(.A(mai_mai_n281_), .B(mai_mai_n150_), .Y(mai_mai_n837_));
  NA2        m0788(.A(mai_mai_n144_), .B(x7), .Y(mai_mai_n838_));
  OR3        m0789(.A(mai_mai_n753_), .B(mai_mai_n470_), .C(mai_mai_n723_), .Y(mai_mai_n839_));
  OAI220     m0790(.A0(mai_mai_n839_), .A1(mai_mai_n838_), .B0(mai_mai_n837_), .B1(mai_mai_n207_), .Y(mai_mai_n840_));
  AOI210     m0791(.A0(mai_mai_n836_), .A1(mai_mai_n295_), .B0(mai_mai_n840_), .Y(mai_mai_n841_));
  AOI210     m0792(.A0(mai_mai_n841_), .A1(mai_mai_n832_), .B0(mai_mai_n71_), .Y(mai_mai_n842_));
  NO2        m0793(.A(mai_mai_n816_), .B(mai_mai_n110_), .Y(mai_mai_n843_));
  NA2        m0794(.A(mai_mai_n843_), .B(mai_mai_n195_), .Y(mai_mai_n844_));
  OAI210     m0795(.A0(mai_mai_n412_), .A1(mai_mai_n307_), .B0(mai_mai_n347_), .Y(mai_mai_n845_));
  NA2        m0796(.A(mai_mai_n438_), .B(mai_mai_n236_), .Y(mai_mai_n846_));
  NA2        m0797(.A(mai_mai_n720_), .B(mai_mai_n107_), .Y(mai_mai_n847_));
  OAI220     m0798(.A0(mai_mai_n847_), .A1(mai_mai_n846_), .B0(mai_mai_n845_), .B1(mai_mai_n844_), .Y(mai_mai_n848_));
  NA2        m0799(.A(mai_mai_n848_), .B(mai_mai_n291_), .Y(mai_mai_n849_));
  NA2        m0800(.A(mai_mai_n337_), .B(mai_mai_n53_), .Y(mai_mai_n850_));
  NO3        m0801(.A(mai_mai_n412_), .B(mai_mai_n137_), .C(mai_mai_n68_), .Y(mai_mai_n851_));
  NO2        m0802(.A(mai_mai_n708_), .B(mai_mai_n248_), .Y(mai_mai_n852_));
  NO3        m0803(.A(mai_mai_n569_), .B(mai_mai_n471_), .C(mai_mai_n99_), .Y(mai_mai_n853_));
  AO220      m0804(.A0(mai_mai_n853_), .A1(mai_mai_n852_), .B0(mai_mai_n851_), .B1(mai_mai_n850_), .Y(mai_mai_n854_));
  NA2        m0805(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n855_));
  NO3        m0806(.A(mai_mai_n316_), .B(mai_mai_n855_), .C(mai_mai_n290_), .Y(mai_mai_n856_));
  AOI210     m0807(.A0(mai_mai_n854_), .A1(x5), .B0(mai_mai_n856_), .Y(mai_mai_n857_));
  AOI210     m0808(.A0(mai_mai_n857_), .A1(mai_mai_n849_), .B0(mai_mai_n72_), .Y(mai_mai_n858_));
  NO2        m0809(.A(mai_mai_n70_), .B(x3), .Y(mai_mai_n859_));
  OAI210     m0810(.A0(mai_mai_n859_), .A1(mai_mai_n267_), .B0(mai_mai_n148_), .Y(mai_mai_n860_));
  MUX2       m0811(.S(x3), .A(mai_mai_n166_), .B(mai_mai_n774_), .Y(mai_mai_n861_));
  NA2        m0812(.A(mai_mai_n861_), .B(mai_mai_n560_), .Y(mai_mai_n862_));
  NO3        m0813(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n863_));
  INV        m0814(.A(mai_mai_n863_), .Y(mai_mai_n864_));
  AOI210     m0815(.A0(mai_mai_n862_), .A1(mai_mai_n860_), .B0(mai_mai_n864_), .Y(mai_mai_n865_));
  NO3        m0816(.A(x5), .B(x3), .C(mai_mai_n110_), .Y(mai_mai_n866_));
  AOI220     m0817(.A0(mai_mai_n827_), .A1(mai_mai_n312_), .B0(mai_mai_n866_), .B1(mai_mai_n59_), .Y(mai_mai_n867_));
  OR2        m0818(.A(x8), .B(x1), .Y(mai_mai_n868_));
  NO3        m0819(.A(mai_mai_n868_), .B(mai_mai_n867_), .C(mai_mai_n737_), .Y(mai_mai_n869_));
  NAi21      m0820(.An(x4), .B(x1), .Y(mai_mai_n870_));
  NO2        m0821(.A(mai_mai_n870_), .B(x0), .Y(mai_mai_n871_));
  NA2        m0822(.A(mai_mai_n614_), .B(mai_mai_n871_), .Y(mai_mai_n872_));
  NA3        m0823(.A(mai_mai_n55_), .B(x1), .C(x0), .Y(mai_mai_n873_));
  OAI210     m0824(.A0(mai_mai_n873_), .A1(mai_mai_n719_), .B0(mai_mai_n872_), .Y(mai_mai_n874_));
  OAI210     m0825(.A0(mai_mai_n874_), .A1(mai_mai_n869_), .B0(mai_mai_n323_), .Y(mai_mai_n875_));
  AO210      m0826(.A0(mai_mai_n293_), .A1(mai_mai_n267_), .B0(mai_mai_n736_), .Y(mai_mai_n876_));
  NA2        m0827(.A(mai_mai_n108_), .B(mai_mai_n56_), .Y(mai_mai_n877_));
  NO2        m0828(.A(mai_mai_n877_), .B(mai_mai_n263_), .Y(mai_mai_n878_));
  NO2        m0829(.A(mai_mai_n57_), .B(x2), .Y(mai_mai_n879_));
  NO4        m0830(.A(mai_mai_n333_), .B(mai_mai_n879_), .C(mai_mai_n816_), .D(mai_mai_n297_), .Y(mai_mai_n880_));
  AOI220     m0831(.A0(mai_mai_n880_), .A1(mai_mai_n878_), .B0(mai_mai_n876_), .B1(mai_mai_n645_), .Y(mai_mai_n881_));
  NA2        m0832(.A(mai_mai_n881_), .B(mai_mai_n875_), .Y(mai_mai_n882_));
  NO4        m0833(.A(mai_mai_n882_), .B(mai_mai_n865_), .C(mai_mai_n858_), .D(mai_mai_n842_), .Y(mai09));
  NO3        m0834(.A(mai_mai_n789_), .B(mai_mai_n121_), .C(mai_mai_n96_), .Y(mai_mai_n884_));
  AOI220     m0835(.A0(mai_mai_n302_), .A1(mai_mai_n70_), .B0(mai_mai_n590_), .B1(mai_mai_n542_), .Y(mai_mai_n885_));
  OAI210     m0836(.A0(mai_mai_n884_), .A1(x2), .B0(mai_mai_n885_), .Y(mai_mai_n886_));
  AOI210     m0837(.A0(mai_mai_n886_), .A1(mai_mai_n757_), .B0(mai_mai_n447_), .Y(mai_mai_n887_));
  NO2        m0838(.A(mai_mai_n589_), .B(mai_mai_n266_), .Y(mai_mai_n888_));
  NO2        m0839(.A(mai_mai_n756_), .B(mai_mai_n343_), .Y(mai_mai_n889_));
  NO3        m0840(.A(mai_mai_n606_), .B(mai_mai_n102_), .C(mai_mai_n110_), .Y(mai_mai_n890_));
  AO220      m0841(.A0(mai_mai_n890_), .A1(mai_mai_n889_), .B0(mai_mai_n888_), .B1(mai_mai_n621_), .Y(mai_mai_n891_));
  OAI210     m0842(.A0(mai_mai_n891_), .A1(mai_mai_n887_), .B0(x4), .Y(mai_mai_n892_));
  OAI220     m0843(.A0(mai_mai_n371_), .A1(mai_mai_n145_), .B0(mai_mai_n396_), .B1(mai_mai_n283_), .Y(mai_mai_n893_));
  NO2        m0844(.A(mai_mai_n193_), .B(mai_mai_n108_), .Y(mai_mai_n894_));
  AOI220     m0845(.A0(mai_mai_n894_), .A1(mai_mai_n126_), .B0(mai_mai_n893_), .B1(mai_mai_n627_), .Y(mai_mai_n895_));
  NO2        m0846(.A(mai_mai_n789_), .B(mai_mai_n96_), .Y(mai_mai_n896_));
  NAi21      m0847(.An(x0), .B(x2), .Y(mai_mai_n897_));
  NO2        m0848(.A(mai_mai_n306_), .B(mai_mai_n897_), .Y(mai_mai_n898_));
  OAI210     m0849(.A0(mai_mai_n480_), .A1(mai_mai_n278_), .B0(mai_mai_n193_), .Y(mai_mai_n899_));
  AOI210     m0850(.A0(mai_mai_n169_), .A1(mai_mai_n809_), .B0(mai_mai_n359_), .Y(mai_mai_n900_));
  AOI220     m0851(.A0(mai_mai_n900_), .A1(mai_mai_n899_), .B0(mai_mai_n898_), .B1(mai_mai_n896_), .Y(mai_mai_n901_));
  OAI210     m0852(.A0(mai_mai_n895_), .A1(mai_mai_n55_), .B0(mai_mai_n901_), .Y(mai_mai_n902_));
  NA2        m0853(.A(mai_mai_n902_), .B(mai_mai_n56_), .Y(mai_mai_n903_));
  NO2        m0854(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n904_));
  INV        m0855(.A(mai_mai_n126_), .Y(mai_mai_n905_));
  NA2        m0856(.A(mai_mai_n756_), .B(mai_mai_n55_), .Y(mai_mai_n906_));
  AOI210     m0857(.A0(x6), .A1(x1), .B0(x5), .Y(mai_mai_n907_));
  OAI210     m0858(.A0(mai_mai_n907_), .A1(mai_mai_n336_), .B0(x2), .Y(mai_mai_n908_));
  AOI210     m0859(.A0(mai_mai_n908_), .A1(mai_mai_n906_), .B0(mai_mai_n905_), .Y(mai_mai_n909_));
  NA2        m0860(.A(mai_mai_n559_), .B(mai_mai_n55_), .Y(mai_mai_n910_));
  NO4        m0861(.A(mai_mai_n57_), .B(x6), .C(x5), .D(x1), .Y(mai_mai_n911_));
  NO2        m0862(.A(mai_mai_n233_), .B(mai_mai_n386_), .Y(mai_mai_n912_));
  NO2        m0863(.A(mai_mai_n313_), .B(mai_mai_n149_), .Y(mai_mai_n913_));
  NO3        m0864(.A(mai_mai_n913_), .B(mai_mai_n912_), .C(mai_mai_n911_), .Y(mai_mai_n914_));
  OAI220     m0865(.A0(mai_mai_n914_), .A1(mai_mai_n55_), .B0(mai_mai_n910_), .B1(mai_mai_n459_), .Y(mai_mai_n915_));
  OAI210     m0866(.A0(mai_mai_n915_), .A1(mai_mai_n909_), .B0(mai_mai_n904_), .Y(mai_mai_n916_));
  NO2        m0867(.A(mai_mai_n405_), .B(mai_mai_n108_), .Y(mai_mai_n917_));
  NO2        m0868(.A(mai_mai_n337_), .B(mai_mai_n497_), .Y(mai_mai_n918_));
  AOI220     m0869(.A0(mai_mai_n918_), .A1(mai_mai_n917_), .B0(mai_mai_n211_), .B1(mai_mai_n231_), .Y(mai_mai_n919_));
  NA4        m0870(.A(mai_mai_n919_), .B(mai_mai_n916_), .C(mai_mai_n903_), .D(mai_mai_n892_), .Y(mai_mai_n920_));
  NA2        m0871(.A(mai_mai_n920_), .B(mai_mai_n50_), .Y(mai_mai_n921_));
  NO2        m0872(.A(mai_mai_n381_), .B(mai_mai_n162_), .Y(mai_mai_n922_));
  NA2        m0873(.A(mai_mai_n242_), .B(mai_mai_n590_), .Y(mai_mai_n923_));
  NO2        m0874(.A(mai_mai_n433_), .B(mai_mai_n819_), .Y(mai_mai_n924_));
  OAI210     m0875(.A0(mai_mai_n924_), .A1(mai_mai_n922_), .B0(x0), .Y(mai_mai_n925_));
  NO3        m0876(.A(x8), .B(x7), .C(x2), .Y(mai_mai_n926_));
  NO3        m0877(.A(mai_mai_n57_), .B(x5), .C(x2), .Y(mai_mai_n927_));
  OAI210     m0878(.A0(mai_mai_n927_), .A1(mai_mai_n926_), .B0(mai_mai_n517_), .Y(mai_mai_n928_));
  AOI210     m0879(.A0(mai_mai_n928_), .A1(mai_mai_n925_), .B0(x4), .Y(mai_mai_n929_));
  NO2        m0880(.A(mai_mai_n426_), .B(mai_mai_n148_), .Y(mai_mai_n930_));
  NO2        m0881(.A(mai_mai_n52_), .B(x2), .Y(mai_mai_n931_));
  NO2        m0882(.A(mai_mai_n108_), .B(mai_mai_n56_), .Y(mai_mai_n932_));
  NA2        m0883(.A(mai_mai_n932_), .B(x8), .Y(mai_mai_n933_));
  OAI210     m0884(.A0(mai_mai_n930_), .A1(mai_mai_n929_), .B0(mai_mai_n619_), .Y(mai_mai_n934_));
  NO2        m0885(.A(mai_mai_n262_), .B(mai_mai_n119_), .Y(mai_mai_n935_));
  OAI210     m0886(.A0(x4), .A1(x2), .B0(x0), .Y(mai_mai_n936_));
  NA3        m0887(.A(mai_mai_n608_), .B(mai_mai_n620_), .C(mai_mai_n348_), .Y(mai_mai_n937_));
  OAI210     m0888(.A0(mai_mai_n936_), .A1(mai_mai_n290_), .B0(mai_mai_n53_), .Y(mai_mai_n938_));
  AOI210     m0889(.A0(mai_mai_n937_), .A1(mai_mai_n936_), .B0(mai_mai_n938_), .Y(mai_mai_n939_));
  OAI210     m0890(.A0(mai_mai_n939_), .A1(mai_mai_n935_), .B0(mai_mai_n332_), .Y(mai_mai_n940_));
  AOI220     m0891(.A0(mai_mai_n671_), .A1(mai_mai_n352_), .B0(mai_mai_n354_), .B1(mai_mai_n93_), .Y(mai_mai_n941_));
  NA2        m0892(.A(mai_mai_n93_), .B(x5), .Y(mai_mai_n942_));
  OAI220     m0893(.A0(mai_mai_n942_), .A1(mai_mai_n868_), .B0(mai_mai_n941_), .B1(mai_mai_n324_), .Y(mai_mai_n943_));
  NA2        m0894(.A(mai_mai_n943_), .B(mai_mai_n68_), .Y(mai_mai_n944_));
  NA2        m0895(.A(mai_mai_n409_), .B(mai_mai_n774_), .Y(mai_mai_n945_));
  NA2        m0896(.A(mai_mai_n253_), .B(mai_mai_n166_), .Y(mai_mai_n946_));
  AO210      m0897(.A0(mai_mai_n946_), .A1(mai_mai_n945_), .B0(mai_mai_n134_), .Y(mai_mai_n947_));
  NO2        m0898(.A(mai_mai_n439_), .B(x2), .Y(mai_mai_n948_));
  NO2        m0899(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n949_));
  NA2        m0900(.A(mai_mai_n949_), .B(x5), .Y(mai_mai_n950_));
  NO2        m0901(.A(mai_mai_n950_), .B(mai_mai_n60_), .Y(mai_mai_n951_));
  AOI220     m0902(.A0(mai_mai_n951_), .A1(mai_mai_n948_), .B0(mai_mai_n672_), .B1(mai_mai_n246_), .Y(mai_mai_n952_));
  NA4        m0903(.A(mai_mai_n952_), .B(mai_mai_n947_), .C(mai_mai_n944_), .D(mai_mai_n940_), .Y(mai_mai_n953_));
  NO4        m0904(.A(mai_mai_n937_), .B(mai_mai_n636_), .C(mai_mai_n459_), .D(mai_mai_n50_), .Y(mai_mai_n954_));
  AOI220     m0905(.A0(mai_mai_n607_), .A1(mai_mai_n606_), .B0(mai_mai_n284_), .B1(x5), .Y(mai_mai_n955_));
  NO2        m0906(.A(mai_mai_n680_), .B(mai_mai_n193_), .Y(mai_mai_n956_));
  NA3        m0907(.A(mai_mai_n956_), .B(mai_mai_n673_), .C(x7), .Y(mai_mai_n957_));
  OAI210     m0908(.A0(mai_mai_n955_), .A1(mai_mai_n353_), .B0(mai_mai_n957_), .Y(mai_mai_n958_));
  OAI210     m0909(.A0(mai_mai_n958_), .A1(mai_mai_n954_), .B0(mai_mai_n82_), .Y(mai_mai_n959_));
  NA2        m0910(.A(mai_mai_n780_), .B(x2), .Y(mai_mai_n960_));
  NO2        m0911(.A(mai_mai_n960_), .B(mai_mai_n58_), .Y(mai_mai_n961_));
  NO2        m0912(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n962_));
  NAi21      m0913(.An(x1), .B(x4), .Y(mai_mai_n963_));
  NA2        m0914(.A(mai_mai_n963_), .B(mai_mai_n870_), .Y(mai_mai_n964_));
  NO3        m0915(.A(mai_mai_n964_), .B(mai_mai_n204_), .C(mai_mai_n962_), .Y(mai_mai_n965_));
  OAI210     m0916(.A0(mai_mai_n965_), .A1(mai_mai_n961_), .B0(mai_mai_n416_), .Y(mai_mai_n966_));
  NA3        m0917(.A(mai_mai_n399_), .B(mai_mai_n756_), .C(mai_mai_n57_), .Y(mai_mai_n967_));
  NA3        m0918(.A(mai_mai_n967_), .B(mai_mai_n966_), .C(mai_mai_n959_), .Y(mai_mai_n968_));
  AOI210     m0919(.A0(mai_mai_n953_), .A1(x6), .B0(mai_mai_n968_), .Y(mai_mai_n969_));
  NA3        m0920(.A(mai_mai_n969_), .B(mai_mai_n934_), .C(mai_mai_n921_), .Y(mai10));
  NO2        m0921(.A(x4), .B(x1), .Y(mai_mai_n971_));
  NO2        m0922(.A(mai_mai_n971_), .B(mai_mai_n150_), .Y(mai_mai_n972_));
  NA3        m0923(.A(x5), .B(x4), .C(x0), .Y(mai_mai_n973_));
  OAI220     m0924(.A0(mai_mai_n973_), .A1(mai_mai_n279_), .B0(mai_mai_n708_), .B1(mai_mai_n250_), .Y(mai_mai_n974_));
  NA2        m0925(.A(mai_mai_n974_), .B(mai_mai_n972_), .Y(mai_mai_n975_));
  NO3        m0926(.A(mai_mai_n360_), .B(mai_mai_n324_), .C(mai_mai_n92_), .Y(mai_mai_n976_));
  NA3        m0927(.A(mai_mai_n976_), .B(mai_mai_n384_), .C(mai_mai_n62_), .Y(mai_mai_n977_));
  AOI210     m0928(.A0(mai_mai_n977_), .A1(mai_mai_n975_), .B0(mai_mai_n306_), .Y(mai_mai_n978_));
  NOi21      m0929(.An(mai_mai_n261_), .B(mai_mai_n140_), .Y(mai_mai_n979_));
  AOI210     m0930(.A0(mai_mai_n503_), .A1(mai_mai_n621_), .B0(mai_mai_n333_), .Y(mai_mai_n980_));
  NO2        m0931(.A(mai_mai_n904_), .B(mai_mai_n346_), .Y(mai_mai_n981_));
  NOi31      m0932(.An(mai_mai_n981_), .B(mai_mai_n980_), .C(mai_mai_n979_), .Y(mai_mai_n982_));
  NA2        m0933(.A(x4), .B(mai_mai_n110_), .Y(mai_mai_n983_));
  NO2        m0934(.A(mai_mai_n327_), .B(mai_mai_n983_), .Y(mai_mai_n984_));
  NA2        m0935(.A(mai_mai_n99_), .B(x5), .Y(mai_mai_n985_));
  NO3        m0936(.A(mai_mai_n985_), .B(mai_mai_n111_), .C(mai_mai_n55_), .Y(mai_mai_n986_));
  NO3        m0937(.A(mai_mai_n986_), .B(mai_mai_n984_), .C(mai_mai_n982_), .Y(mai_mai_n987_));
  NA2        m0938(.A(mai_mai_n962_), .B(mai_mai_n50_), .Y(mai_mai_n988_));
  NA2        m0939(.A(mai_mai_n607_), .B(mai_mai_n273_), .Y(mai_mai_n989_));
  NO2        m0940(.A(mai_mai_n989_), .B(mai_mai_n988_), .Y(mai_mai_n990_));
  OAI220     m0941(.A0(mai_mai_n933_), .A1(mai_mai_n107_), .B0(mai_mai_n877_), .B1(mai_mai_n447_), .Y(mai_mai_n991_));
  AOI210     m0942(.A0(mai_mai_n991_), .A1(mai_mai_n281_), .B0(mai_mai_n990_), .Y(mai_mai_n992_));
  OAI210     m0943(.A0(mai_mai_n987_), .A1(mai_mai_n386_), .B0(mai_mai_n992_), .Y(mai_mai_n993_));
  OAI210     m0944(.A0(mai_mai_n993_), .A1(mai_mai_n978_), .B0(x7), .Y(mai_mai_n994_));
  NA2        m0945(.A(mai_mai_n55_), .B(mai_mai_n71_), .Y(mai_mai_n995_));
  AOI210     m0946(.A0(mai_mai_n447_), .A1(mai_mai_n359_), .B0(mai_mai_n983_), .Y(mai_mai_n996_));
  NO3        m0947(.A(mai_mai_n449_), .B(mai_mai_n897_), .C(x5), .Y(mai_mai_n997_));
  OAI210     m0948(.A0(mai_mai_n997_), .A1(mai_mai_n996_), .B0(mai_mai_n995_), .Y(mai_mai_n998_));
  NO2        m0949(.A(mai_mai_n360_), .B(mai_mai_n143_), .Y(mai_mai_n999_));
  NA2        m0950(.A(mai_mai_n999_), .B(mai_mai_n427_), .Y(mai_mai_n1000_));
  AOI210     m0951(.A0(mai_mai_n1000_), .A1(mai_mai_n998_), .B0(x3), .Y(mai_mai_n1001_));
  NA2        m0952(.A(mai_mai_n700_), .B(mai_mai_n253_), .Y(mai_mai_n1002_));
  NO2        m0953(.A(x5), .B(mai_mai_n110_), .Y(mai_mai_n1003_));
  OAI210     m0954(.A0(mai_mai_n1003_), .A1(mai_mai_n240_), .B0(mai_mai_n942_), .Y(mai_mai_n1004_));
  NA3        m0955(.A(mai_mai_n466_), .B(mai_mai_n132_), .C(mai_mai_n427_), .Y(mai_mai_n1005_));
  OAI210     m0956(.A0(mai_mai_n449_), .A1(mai_mai_n216_), .B0(mai_mai_n1005_), .Y(mai_mai_n1006_));
  AOI210     m0957(.A0(mai_mai_n1004_), .A1(mai_mai_n259_), .B0(mai_mai_n1006_), .Y(mai_mai_n1007_));
  OAI220     m0958(.A0(mai_mai_n1007_), .A1(mai_mai_n59_), .B0(mai_mai_n1002_), .B1(mai_mai_n713_), .Y(mai_mai_n1008_));
  OAI210     m0959(.A0(mai_mai_n1008_), .A1(mai_mai_n1001_), .B0(mai_mai_n949_), .Y(mai_mai_n1009_));
  NO2        m0960(.A(x4), .B(x3), .Y(mai_mai_n1010_));
  NO3        m0961(.A(mai_mai_n1010_), .B(mai_mai_n347_), .C(mai_mai_n87_), .Y(mai_mai_n1011_));
  OAI210     m0962(.A0(mai_mai_n1011_), .A1(mai_mai_n280_), .B0(mai_mai_n438_), .Y(mai_mai_n1012_));
  AOI210     m0963(.A0(mai_mai_n400_), .A1(mai_mai_n129_), .B0(mai_mai_n254_), .Y(mai_mai_n1013_));
  NA2        m0964(.A(mai_mai_n971_), .B(mai_mai_n55_), .Y(mai_mai_n1014_));
  NO2        m0965(.A(mai_mai_n1014_), .B(mai_mai_n985_), .Y(mai_mai_n1015_));
  NO2        m0966(.A(mai_mai_n527_), .B(mai_mai_n365_), .Y(mai_mai_n1016_));
  NO3        m0967(.A(x4), .B(mai_mai_n110_), .C(mai_mai_n59_), .Y(mai_mai_n1017_));
  NO2        m0968(.A(mai_mai_n439_), .B(x1), .Y(mai_mai_n1018_));
  NOi31      m0969(.An(mai_mai_n1017_), .B(mai_mai_n1018_), .C(mai_mai_n1016_), .Y(mai_mai_n1019_));
  NA2        m0970(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n1020_));
  NO4        m0971(.A(mai_mai_n972_), .B(mai_mai_n516_), .C(mai_mai_n1020_), .D(x2), .Y(mai_mai_n1021_));
  NO4        m0972(.A(mai_mai_n1021_), .B(mai_mai_n1019_), .C(mai_mai_n1015_), .D(mai_mai_n1013_), .Y(mai_mai_n1022_));
  AOI210     m0973(.A0(mai_mai_n1022_), .A1(mai_mai_n1012_), .B0(mai_mai_n210_), .Y(mai_mai_n1023_));
  NO2        m0974(.A(mai_mai_n669_), .B(mai_mai_n502_), .Y(mai_mai_n1024_));
  NO2        m0975(.A(x6), .B(x2), .Y(mai_mai_n1025_));
  NO3        m0976(.A(mai_mai_n1025_), .B(mai_mai_n700_), .C(mai_mai_n60_), .Y(mai_mai_n1026_));
  OAI210     m0977(.A0(mai_mai_n1026_), .A1(mai_mai_n1024_), .B0(mai_mai_n272_), .Y(mai_mai_n1027_));
  NO2        m0978(.A(mai_mai_n877_), .B(mai_mai_n447_), .Y(mai_mai_n1028_));
  NA3        m0979(.A(x4), .B(x3), .C(mai_mai_n110_), .Y(mai_mai_n1029_));
  NO3        m0980(.A(mai_mai_n1029_), .B(mai_mai_n706_), .C(mai_mai_n466_), .Y(mai_mai_n1030_));
  AOI210     m0981(.A0(mai_mai_n1028_), .A1(mai_mai_n473_), .B0(mai_mai_n1030_), .Y(mai_mai_n1031_));
  AOI210     m0982(.A0(mai_mai_n1031_), .A1(mai_mai_n1027_), .B0(mai_mai_n459_), .Y(mai_mai_n1032_));
  NO2        m0983(.A(mai_mai_n55_), .B(mai_mai_n56_), .Y(mai_mai_n1033_));
  OAI220     m0984(.A0(mai_mai_n827_), .A1(mai_mai_n461_), .B0(mai_mai_n758_), .B1(mai_mai_n129_), .Y(mai_mai_n1034_));
  NOi21      m0985(.An(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n1035_));
  NO3        m0986(.A(mai_mai_n348_), .B(mai_mai_n327_), .C(mai_mai_n1035_), .Y(mai_mai_n1036_));
  AOI220     m0987(.A0(mai_mai_n1036_), .A1(mai_mai_n258_), .B0(mai_mai_n1034_), .B1(mai_mai_n116_), .Y(mai_mai_n1037_));
  NO2        m0988(.A(mai_mai_n1037_), .B(mai_mai_n1033_), .Y(mai_mai_n1038_));
  NA2        m0989(.A(mai_mai_n520_), .B(mai_mai_n263_), .Y(mai_mai_n1039_));
  NO2        m0990(.A(mai_mai_n488_), .B(mai_mai_n589_), .Y(mai_mai_n1040_));
  NA3        m0991(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n55_), .Y(mai_mai_n1041_));
  NO2        m0992(.A(mai_mai_n185_), .B(mai_mai_n110_), .Y(mai_mai_n1042_));
  NA3        m0993(.A(mai_mai_n1042_), .B(mai_mai_n184_), .C(mai_mai_n123_), .Y(mai_mai_n1043_));
  NA2        m0994(.A(mai_mai_n1043_), .B(mai_mai_n1041_), .Y(mai_mai_n1044_));
  NO4        m0995(.A(mai_mai_n1044_), .B(mai_mai_n1038_), .C(mai_mai_n1032_), .D(mai_mai_n1023_), .Y(mai_mai_n1045_));
  NA3        m0996(.A(mai_mai_n1045_), .B(mai_mai_n1009_), .C(mai_mai_n994_), .Y(mai11));
  NA2        m0997(.A(mai_mai_n380_), .B(mai_mai_n92_), .Y(mai_mai_n1047_));
  INV        m0998(.A(mai_mai_n898_), .Y(mai_mai_n1048_));
  OAI220     m0999(.A0(mai_mai_n1048_), .A1(mai_mai_n53_), .B0(mai_mai_n1047_), .B1(mai_mai_n369_), .Y(mai_mai_n1049_));
  NO2        m1000(.A(mai_mai_n774_), .B(x5), .Y(mai_mai_n1050_));
  NO2        m1001(.A(mai_mai_n170_), .B(mai_mai_n533_), .Y(mai_mai_n1051_));
  AOI220     m1002(.A0(mai_mai_n1051_), .A1(mai_mai_n1050_), .B0(mai_mai_n1049_), .B1(x5), .Y(mai_mai_n1052_));
  OAI220     m1003(.A0(mai_mai_n979_), .A1(mai_mai_n219_), .B0(mai_mai_n217_), .B1(mai_mai_n185_), .Y(mai_mai_n1053_));
  NO2        m1004(.A(mai_mai_n344_), .B(mai_mai_n428_), .Y(mai_mai_n1054_));
  AOI220     m1005(.A0(mai_mai_n1054_), .A1(mai_mai_n183_), .B0(mai_mai_n1053_), .B1(mai_mai_n166_), .Y(mai_mai_n1055_));
  NO2        m1006(.A(mai_mai_n1055_), .B(mai_mai_n449_), .Y(mai_mai_n1056_));
  NO2        m1007(.A(mai_mai_n254_), .B(x2), .Y(mai_mai_n1057_));
  OAI210     m1008(.A0(mai_mai_n922_), .A1(mai_mai_n1057_), .B0(mai_mai_n417_), .Y(mai_mai_n1058_));
  NO2        m1009(.A(mai_mai_n55_), .B(mai_mai_n108_), .Y(mai_mai_n1059_));
  NA2        m1010(.A(mai_mai_n281_), .B(mai_mai_n1059_), .Y(mai_mai_n1060_));
  NO2        m1011(.A(mai_mai_n71_), .B(x1), .Y(mai_mai_n1061_));
  NA2        m1012(.A(mai_mai_n1061_), .B(mai_mai_n78_), .Y(mai_mai_n1062_));
  OR2        m1013(.A(mai_mai_n1062_), .B(mai_mai_n615_), .Y(mai_mai_n1063_));
  AOI210     m1014(.A0(mai_mai_n1063_), .A1(mai_mai_n1058_), .B0(mai_mai_n713_), .Y(mai_mai_n1064_));
  NO2        m1015(.A(mai_mai_n307_), .B(mai_mai_n53_), .Y(mai_mai_n1065_));
  NO2        m1016(.A(mai_mai_n438_), .B(x3), .Y(mai_mai_n1066_));
  NA3        m1017(.A(mai_mai_n1066_), .B(mai_mai_n1065_), .C(mai_mai_n897_), .Y(mai_mai_n1067_));
  AOI210     m1018(.A0(mai_mai_n1067_), .A1(mai_mai_n946_), .B0(mai_mai_n398_), .Y(mai_mai_n1068_));
  NA2        m1019(.A(mai_mai_n110_), .B(x1), .Y(mai_mai_n1069_));
  NO2        m1020(.A(mai_mai_n621_), .B(mai_mai_n222_), .Y(mai_mai_n1070_));
  NA4        m1021(.A(mai_mai_n1070_), .B(mai_mai_n889_), .C(mai_mai_n470_), .D(mai_mai_n1069_), .Y(mai_mai_n1071_));
  NA3        m1022(.A(x6), .B(x5), .C(mai_mai_n110_), .Y(mai_mai_n1072_));
  NO2        m1023(.A(mai_mai_n1072_), .B(mai_mai_n279_), .Y(mai_mai_n1073_));
  NO2        m1024(.A(mai_mai_n449_), .B(x0), .Y(mai_mai_n1074_));
  NOi31      m1025(.An(mai_mai_n1074_), .B(mai_mai_n175_), .C(mai_mai_n51_), .Y(mai_mai_n1075_));
  AOI210     m1026(.A0(mai_mai_n1073_), .A1(mai_mai_n181_), .B0(mai_mai_n1075_), .Y(mai_mai_n1076_));
  NA2        m1027(.A(mai_mai_n1076_), .B(mai_mai_n1071_), .Y(mai_mai_n1077_));
  NO4        m1028(.A(mai_mai_n1077_), .B(mai_mai_n1068_), .C(mai_mai_n1064_), .D(mai_mai_n1056_), .Y(mai_mai_n1078_));
  OAI210     m1029(.A0(mai_mai_n1052_), .A1(mai_mai_n144_), .B0(mai_mai_n1078_), .Y(mai_mai_n1079_));
  NA2        m1030(.A(mai_mai_n868_), .B(mai_mai_n87_), .Y(mai_mai_n1080_));
  NO3        m1031(.A(mai_mai_n467_), .B(mai_mai_n780_), .C(mai_mai_n124_), .Y(mai_mai_n1081_));
  AOI210     m1032(.A0(mai_mai_n1080_), .A1(mai_mai_n101_), .B0(mai_mai_n1081_), .Y(mai_mai_n1082_));
  NO2        m1033(.A(x8), .B(x1), .Y(mai_mai_n1083_));
  NO3        m1034(.A(mai_mai_n1083_), .B(mai_mai_n692_), .C(mai_mai_n451_), .Y(mai_mai_n1084_));
  OAI210     m1035(.A0(mai_mai_n77_), .A1(mai_mai_n53_), .B0(mai_mai_n1084_), .Y(mai_mai_n1085_));
  OAI210     m1036(.A0(mai_mai_n1082_), .A1(x3), .B0(mai_mai_n1085_), .Y(mai_mai_n1086_));
  NO2        m1037(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n1087_));
  OAI210     m1038(.A0(mai_mai_n1087_), .A1(x2), .B0(mai_mai_n236_), .Y(mai_mai_n1088_));
  NO2        m1039(.A(mai_mai_n608_), .B(mai_mai_n234_), .Y(mai_mai_n1089_));
  NA2        m1040(.A(mai_mai_n1089_), .B(mai_mai_n1088_), .Y(mai_mai_n1090_));
  NO2        m1041(.A(mai_mai_n520_), .B(x4), .Y(mai_mai_n1091_));
  NO3        m1042(.A(mai_mai_n55_), .B(x6), .C(x1), .Y(mai_mai_n1092_));
  NOi21      m1043(.An(mai_mai_n1092_), .B(mai_mai_n488_), .Y(mai_mai_n1093_));
  AOI210     m1044(.A0(mai_mai_n1091_), .A1(mai_mai_n579_), .B0(mai_mai_n1093_), .Y(mai_mai_n1094_));
  NA2        m1045(.A(mai_mai_n1094_), .B(mai_mai_n1090_), .Y(mai_mai_n1095_));
  AOI210     m1046(.A0(mai_mai_n1086_), .A1(x2), .B0(mai_mai_n1095_), .Y(mai_mai_n1096_));
  NO2        m1047(.A(mai_mai_n234_), .B(x2), .Y(mai_mai_n1097_));
  NA2        m1048(.A(mai_mai_n1097_), .B(mai_mai_n1010_), .Y(mai_mai_n1098_));
  NOi21      m1049(.An(mai_mai_n389_), .B(mai_mai_n568_), .Y(mai_mai_n1099_));
  NO3        m1050(.A(mai_mai_n1099_), .B(mai_mai_n607_), .C(mai_mai_n327_), .Y(mai_mai_n1100_));
  NA2        m1051(.A(x8), .B(mai_mai_n110_), .Y(mai_mai_n1101_));
  OAI220     m1052(.A0(mai_mai_n713_), .A1(mai_mai_n1101_), .B0(mai_mai_n327_), .B1(mai_mai_n384_), .Y(mai_mai_n1102_));
  OAI210     m1053(.A0(mai_mai_n1102_), .A1(mai_mai_n1100_), .B0(mai_mai_n71_), .Y(mai_mai_n1103_));
  NO2        m1054(.A(mai_mai_n108_), .B(x1), .Y(mai_mai_n1104_));
  NA2        m1055(.A(mai_mai_n1104_), .B(x7), .Y(mai_mai_n1105_));
  AOI210     m1056(.A0(mai_mai_n1103_), .A1(mai_mai_n1098_), .B0(mai_mai_n1105_), .Y(mai_mai_n1106_));
  NA2        m1057(.A(mai_mai_n84_), .B(mai_mai_n71_), .Y(mai_mai_n1107_));
  INV        m1058(.A(mai_mai_n251_), .Y(mai_mai_n1108_));
  NA2        m1059(.A(mai_mai_n1108_), .B(mai_mai_n150_), .Y(mai_mai_n1109_));
  OAI220     m1060(.A0(mai_mai_n1109_), .A1(mai_mai_n369_), .B0(mai_mai_n1107_), .B1(mai_mai_n327_), .Y(mai_mai_n1110_));
  NO2        m1061(.A(mai_mai_n160_), .B(mai_mai_n55_), .Y(mai_mai_n1111_));
  AOI210     m1062(.A0(mai_mai_n1111_), .A1(mai_mai_n1110_), .B0(mai_mai_n1106_), .Y(mai_mai_n1112_));
  OAI210     m1063(.A0(mai_mai_n1096_), .A1(mai_mai_n855_), .B0(mai_mai_n1112_), .Y(mai_mai_n1113_));
  AO210      m1064(.A0(mai_mai_n1079_), .A1(mai_mai_n57_), .B0(mai_mai_n1113_), .Y(mai12));
  NA2        m1065(.A(mai_mai_n888_), .B(mai_mai_n250_), .Y(mai_mai_n1115_));
  NO2        m1066(.A(mai_mai_n625_), .B(x7), .Y(mai_mai_n1116_));
  NA2        m1067(.A(mai_mai_n1116_), .B(mai_mai_n280_), .Y(mai_mai_n1117_));
  NA2        m1068(.A(mai_mai_n705_), .B(mai_mai_n877_), .Y(mai_mai_n1118_));
  AOI210     m1069(.A0(mai_mai_n1117_), .A1(mai_mai_n1115_), .B0(mai_mai_n1118_), .Y(mai_mai_n1119_));
  NOi21      m1070(.An(mai_mai_n405_), .B(mai_mai_n555_), .Y(mai_mai_n1120_));
  NO2        m1071(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n1121_));
  NO2        m1072(.A(mai_mai_n608_), .B(mai_mai_n1121_), .Y(mai_mai_n1122_));
  NO3        m1073(.A(mai_mai_n870_), .B(mai_mai_n112_), .C(mai_mai_n99_), .Y(mai_mai_n1123_));
  AOI210     m1074(.A0(mai_mai_n1122_), .A1(mai_mai_n1018_), .B0(mai_mai_n1123_), .Y(mai_mai_n1124_));
  NA2        m1075(.A(mai_mai_n1059_), .B(mai_mai_n56_), .Y(mai_mai_n1125_));
  OAI220     m1076(.A0(mai_mai_n1125_), .A1(mai_mai_n580_), .B0(mai_mai_n1124_), .B1(mai_mai_n1120_), .Y(mai_mai_n1126_));
  OAI210     m1077(.A0(mai_mai_n1126_), .A1(mai_mai_n1119_), .B0(mai_mai_n584_), .Y(mai_mai_n1127_));
  NA2        m1078(.A(mai_mai_n87_), .B(x5), .Y(mai_mai_n1128_));
  OAI210     m1079(.A0(mai_mai_n1128_), .A1(mai_mai_n327_), .B0(mai_mai_n724_), .Y(mai_mai_n1129_));
  INV        m1080(.A(mai_mai_n1129_), .Y(mai_mai_n1130_));
  NA2        m1081(.A(mai_mai_n606_), .B(mai_mai_n53_), .Y(mai_mai_n1131_));
  NA2        m1082(.A(mai_mai_n290_), .B(mai_mai_n50_), .Y(mai_mai_n1132_));
  OAI220     m1083(.A0(mai_mai_n1132_), .A1(mai_mai_n313_), .B0(mai_mai_n1131_), .B1(mai_mai_n137_), .Y(mai_mai_n1133_));
  NO2        m1084(.A(mai_mai_n1080_), .B(mai_mai_n515_), .Y(mai_mai_n1134_));
  NO4        m1085(.A(mai_mai_n242_), .B(mai_mai_n272_), .C(mai_mai_n60_), .D(mai_mai_n57_), .Y(mai_mai_n1135_));
  AOI220     m1086(.A0(mai_mai_n1135_), .A1(mai_mai_n1134_), .B0(mai_mai_n1133_), .B1(mai_mai_n56_), .Y(mai_mai_n1136_));
  OAI210     m1087(.A0(mai_mai_n1130_), .A1(mai_mai_n64_), .B0(mai_mai_n1136_), .Y(mai_mai_n1137_));
  NO2        m1088(.A(mai_mai_n57_), .B(x0), .Y(mai_mai_n1138_));
  NO2        m1089(.A(mai_mai_n669_), .B(mai_mai_n324_), .Y(mai_mai_n1139_));
  NO2        m1090(.A(mai_mai_n758_), .B(x3), .Y(mai_mai_n1140_));
  NO2        m1091(.A(mai_mai_n667_), .B(x8), .Y(mai_mai_n1141_));
  AOI220     m1092(.A0(mai_mai_n1141_), .A1(mai_mai_n1140_), .B0(mai_mai_n1139_), .B1(mai_mai_n1138_), .Y(mai_mai_n1142_));
  AOI210     m1093(.A0(mai_mai_n692_), .A1(mai_mai_n250_), .B0(x7), .Y(mai_mai_n1143_));
  NO3        m1094(.A(mai_mai_n1143_), .B(mai_mai_n609_), .C(x8), .Y(mai_mai_n1144_));
  NA4        m1095(.A(mai_mai_n671_), .B(mai_mai_n663_), .C(mai_mai_n207_), .D(x0), .Y(mai_mai_n1145_));
  OAI220     m1096(.A0(mai_mai_n1145_), .A1(mai_mai_n1144_), .B0(mai_mai_n1142_), .B1(mai_mai_n578_), .Y(mai_mai_n1146_));
  AOI210     m1097(.A0(mai_mai_n1137_), .A1(mai_mai_n1025_), .B0(mai_mai_n1146_), .Y(mai_mai_n1147_));
  NO2        m1098(.A(mai_mai_n250_), .B(mai_mai_n55_), .Y(mai_mai_n1148_));
  NO2        m1099(.A(mai_mai_n258_), .B(x8), .Y(mai_mai_n1149_));
  NOi32      m1100(.An(mai_mai_n1149_), .Bn(mai_mai_n206_), .C(mai_mai_n569_), .Y(mai_mai_n1150_));
  INV        m1101(.A(mai_mai_n60_), .Y(mai_mai_n1151_));
  OAI210     m1102(.A0(mai_mai_n1150_), .A1(mai_mai_n1148_), .B0(mai_mai_n1151_), .Y(mai_mai_n1152_));
  NO2        m1103(.A(mai_mai_n949_), .B(mai_mai_n100_), .Y(mai_mai_n1153_));
  NO2        m1104(.A(mai_mai_n169_), .B(mai_mai_n53_), .Y(mai_mai_n1154_));
  AOI210     m1105(.A0(mai_mai_n344_), .A1(x8), .B0(mai_mai_n1154_), .Y(mai_mai_n1155_));
  AOI210     m1106(.A0(mai_mai_n219_), .A1(mai_mai_n96_), .B0(mai_mai_n1155_), .Y(mai_mai_n1156_));
  OAI210     m1107(.A0(mai_mai_n1156_), .A1(mai_mai_n1153_), .B0(mai_mai_n680_), .Y(mai_mai_n1157_));
  NO2        m1108(.A(x7), .B(x0), .Y(mai_mai_n1158_));
  NO3        m1109(.A(mai_mai_n160_), .B(mai_mai_n1158_), .C(mai_mai_n147_), .Y(mai_mai_n1159_));
  XN2        m1110(.A(x8), .B(x7), .Y(mai_mai_n1160_));
  NO3        m1111(.A(mai_mai_n1083_), .B(mai_mai_n261_), .C(mai_mai_n1160_), .Y(mai_mai_n1161_));
  OAI210     m1112(.A0(mai_mai_n1161_), .A1(mai_mai_n1159_), .B0(mai_mai_n737_), .Y(mai_mai_n1162_));
  NO2        m1113(.A(mai_mai_n270_), .B(mai_mai_n266_), .Y(mai_mai_n1163_));
  NO2        m1114(.A(mai_mai_n108_), .B(x4), .Y(mai_mai_n1164_));
  OAI210     m1115(.A0(mai_mai_n1163_), .A1(mai_mai_n280_), .B0(mai_mai_n1164_), .Y(mai_mai_n1165_));
  NA4        m1116(.A(mai_mai_n1165_), .B(mai_mai_n1162_), .C(mai_mai_n1157_), .D(mai_mai_n1152_), .Y(mai_mai_n1166_));
  NA2        m1117(.A(mai_mai_n1166_), .B(mai_mai_n559_), .Y(mai_mai_n1167_));
  NO2        m1118(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n1168_));
  NA2        m1119(.A(mai_mai_n1168_), .B(mai_mai_n165_), .Y(mai_mai_n1169_));
  NO2        m1120(.A(mai_mai_n673_), .B(mai_mai_n261_), .Y(mai_mai_n1170_));
  OAI210     m1121(.A0(mai_mai_n1170_), .A1(mai_mai_n1028_), .B0(mai_mai_n50_), .Y(mai_mai_n1171_));
  AOI210     m1122(.A0(mai_mai_n1171_), .A1(mai_mai_n1169_), .B0(mai_mai_n433_), .Y(mai_mai_n1172_));
  OAI220     m1123(.A0(mai_mai_n292_), .A1(mai_mai_n278_), .B0(mai_mai_n266_), .B1(mai_mai_n245_), .Y(mai_mai_n1173_));
  NA3        m1124(.A(mai_mai_n1173_), .B(mai_mai_n680_), .C(x1), .Y(mai_mai_n1174_));
  OAI210     m1125(.A0(x8), .A1(x0), .B0(x4), .Y(mai_mai_n1175_));
  NO2        m1126(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n1176_));
  NO2        m1127(.A(mai_mai_n68_), .B(mai_mai_n1176_), .Y(mai_mai_n1177_));
  NOi21      m1128(.An(mai_mai_n1175_), .B(mai_mai_n1177_), .Y(mai_mai_n1178_));
  NO2        m1129(.A(mai_mai_n671_), .B(mai_mai_n327_), .Y(mai_mai_n1179_));
  NO2        m1130(.A(mai_mai_n783_), .B(mai_mai_n223_), .Y(mai_mai_n1180_));
  OAI210     m1131(.A0(mai_mai_n1179_), .A1(mai_mai_n1178_), .B0(mai_mai_n1180_), .Y(mai_mai_n1181_));
  NO2        m1132(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n1182_));
  NO2        m1133(.A(mai_mai_n608_), .B(mai_mai_n447_), .Y(mai_mai_n1183_));
  OAI210     m1134(.A0(mai_mai_n1183_), .A1(mai_mai_n1182_), .B0(mai_mai_n258_), .Y(mai_mai_n1184_));
  NO2        m1135(.A(mai_mai_n825_), .B(mai_mai_n424_), .Y(mai_mai_n1185_));
  NA2        m1136(.A(mai_mai_n332_), .B(mai_mai_n59_), .Y(mai_mai_n1186_));
  NO2        m1137(.A(mai_mai_n1125_), .B(mai_mai_n1186_), .Y(mai_mai_n1187_));
  AOI210     m1138(.A0(mai_mai_n1185_), .A1(mai_mai_n181_), .B0(mai_mai_n1187_), .Y(mai_mai_n1188_));
  NA4        m1139(.A(mai_mai_n1188_), .B(mai_mai_n1184_), .C(mai_mai_n1181_), .D(mai_mai_n1174_), .Y(mai_mai_n1189_));
  OAI210     m1140(.A0(mai_mai_n1189_), .A1(mai_mai_n1172_), .B0(mai_mai_n682_), .Y(mai_mai_n1190_));
  NA4        m1141(.A(mai_mai_n1190_), .B(mai_mai_n1167_), .C(mai_mai_n1147_), .D(mai_mai_n1127_), .Y(mai13));
  NO2        m1142(.A(mai_mai_n466_), .B(mai_mai_n354_), .Y(mai_mai_n1192_));
  NOi41      m1143(.An(mai_mai_n1192_), .B(mai_mai_n680_), .C(mai_mai_n294_), .D(mai_mai_n242_), .Y(mai_mai_n1193_));
  NO2        m1144(.A(mai_mai_n870_), .B(mai_mai_n185_), .Y(mai_mai_n1194_));
  NO2        m1145(.A(mai_mai_n159_), .B(mai_mai_n71_), .Y(mai_mai_n1195_));
  XN2        m1146(.A(x4), .B(x0), .Y(mai_mai_n1196_));
  NO3        m1147(.A(mai_mai_n1196_), .B(mai_mai_n111_), .C(mai_mai_n424_), .Y(mai_mai_n1197_));
  AO220      m1148(.A0(mai_mai_n1197_), .A1(mai_mai_n1195_), .B0(mai_mai_n1194_), .B1(mai_mai_n333_), .Y(mai_mai_n1198_));
  OAI210     m1149(.A0(mai_mai_n1198_), .A1(mai_mai_n1193_), .B0(x3), .Y(mai_mai_n1199_));
  NO2        m1150(.A(mai_mai_n870_), .B(x6), .Y(mai_mai_n1200_));
  NO2        m1151(.A(mai_mai_n1132_), .B(mai_mai_n396_), .Y(mai_mai_n1201_));
  NO3        m1152(.A(x8), .B(x5), .C(mai_mai_n110_), .Y(mai_mai_n1202_));
  NA2        m1153(.A(mai_mai_n1202_), .B(mai_mai_n645_), .Y(mai_mai_n1203_));
  NO2        m1154(.A(mai_mai_n608_), .B(mai_mai_n201_), .Y(mai_mai_n1204_));
  NA2        m1155(.A(mai_mai_n1204_), .B(mai_mai_n1092_), .Y(mai_mai_n1205_));
  NA2        m1156(.A(mai_mai_n451_), .B(mai_mai_n53_), .Y(mai_mai_n1206_));
  NO2        m1157(.A(mai_mai_n1206_), .B(mai_mai_n942_), .Y(mai_mai_n1207_));
  NA2        m1158(.A(mai_mai_n1125_), .B(mai_mai_n471_), .Y(mai_mai_n1208_));
  NA2        m1159(.A(mai_mai_n56_), .B(mai_mai_n110_), .Y(mai_mai_n1209_));
  NA2        m1160(.A(mai_mai_n1209_), .B(x1), .Y(mai_mai_n1210_));
  NO2        m1161(.A(mai_mai_n1210_), .B(mai_mai_n263_), .Y(mai_mai_n1211_));
  NO2        m1162(.A(mai_mai_n324_), .B(x6), .Y(mai_mai_n1212_));
  OAI210     m1163(.A0(mai_mai_n254_), .A1(mai_mai_n983_), .B0(mai_mai_n960_), .Y(mai_mai_n1213_));
  AOI220     m1164(.A0(mai_mai_n1213_), .A1(mai_mai_n1212_), .B0(mai_mai_n1211_), .B1(mai_mai_n1208_), .Y(mai_mai_n1214_));
  NAi41      m1165(.An(mai_mai_n1207_), .B(mai_mai_n1214_), .C(mai_mai_n1205_), .D(mai_mai_n1203_), .Y(mai_mai_n1215_));
  AOI220     m1166(.A0(mai_mai_n1215_), .A1(mai_mai_n68_), .B0(mai_mai_n1201_), .B1(mai_mai_n1200_), .Y(mai_mai_n1216_));
  NA2        m1167(.A(mai_mai_n71_), .B(x3), .Y(mai_mai_n1217_));
  NA2        m1168(.A(mai_mai_n1217_), .B(mai_mai_n906_), .Y(mai_mai_n1218_));
  OAI220     m1169(.A0(mai_mai_n306_), .A1(mai_mai_n825_), .B0(mai_mai_n87_), .B1(mai_mai_n77_), .Y(mai_mai_n1219_));
  AOI210     m1170(.A0(mai_mai_n1128_), .A1(mai_mai_n619_), .B0(mai_mai_n983_), .Y(mai_mai_n1220_));
  OA210      m1171(.A0(mai_mai_n1219_), .A1(mai_mai_n1218_), .B0(mai_mai_n1220_), .Y(mai_mai_n1221_));
  NA2        m1172(.A(mai_mai_n621_), .B(mai_mai_n55_), .Y(mai_mai_n1222_));
  NA2        m1173(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n1223_));
  NA2        m1174(.A(mai_mai_n1223_), .B(mai_mai_n542_), .Y(mai_mai_n1224_));
  NO2        m1175(.A(mai_mai_n162_), .B(mai_mai_n132_), .Y(mai_mai_n1225_));
  AOI210     m1176(.A0(mai_mai_n1224_), .A1(mai_mai_n434_), .B0(mai_mai_n1225_), .Y(mai_mai_n1226_));
  NO2        m1177(.A(mai_mai_n1226_), .B(mai_mai_n877_), .Y(mai_mai_n1227_));
  OAI210     m1178(.A0(mai_mai_n1227_), .A1(mai_mai_n1221_), .B0(mai_mai_n1158_), .Y(mai_mai_n1228_));
  NAi21      m1179(.An(mai_mai_n84_), .B(mai_mai_n384_), .Y(mai_mai_n1229_));
  NO2        m1180(.A(mai_mai_n1229_), .B(mai_mai_n71_), .Y(mai_mai_n1230_));
  AOI210     m1181(.A0(mai_mai_n165_), .A1(x4), .B0(mai_mai_n177_), .Y(mai_mai_n1231_));
  NO2        m1182(.A(mai_mai_n1231_), .B(x0), .Y(mai_mai_n1232_));
  NO2        m1183(.A(mai_mai_n173_), .B(mai_mai_n297_), .Y(mai_mai_n1233_));
  OAI210     m1184(.A0(mai_mai_n1233_), .A1(mai_mai_n1232_), .B0(mai_mai_n1230_), .Y(mai_mai_n1234_));
  NA3        m1185(.A(mai_mai_n1164_), .B(mai_mai_n192_), .C(mai_mai_n71_), .Y(mai_mai_n1235_));
  NO2        m1186(.A(x4), .B(x0), .Y(mai_mai_n1236_));
  NO3        m1187(.A(mai_mai_n1003_), .B(mai_mai_n251_), .C(mai_mai_n542_), .Y(mai_mai_n1237_));
  OAI210     m1188(.A0(mai_mai_n1237_), .A1(mai_mai_n202_), .B0(mai_mai_n1236_), .Y(mai_mai_n1238_));
  NA3        m1189(.A(mai_mai_n1238_), .B(mai_mai_n1235_), .C(mai_mai_n1234_), .Y(mai_mai_n1239_));
  NA2        m1190(.A(mai_mai_n253_), .B(mai_mai_n737_), .Y(mai_mai_n1240_));
  NO2        m1191(.A(mai_mai_n1240_), .B(mai_mai_n522_), .Y(mai_mai_n1241_));
  NA2        m1192(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n1242_));
  NO3        m1193(.A(mai_mai_n1242_), .B(mai_mai_n497_), .C(mai_mai_n81_), .Y(mai_mai_n1243_));
  OAI210     m1194(.A0(mai_mai_n1243_), .A1(mai_mai_n1241_), .B0(x2), .Y(mai_mai_n1244_));
  NO2        m1195(.A(mai_mai_n327_), .B(mai_mai_n384_), .Y(mai_mai_n1245_));
  NO2        m1196(.A(mai_mai_n692_), .B(x0), .Y(mai_mai_n1246_));
  OAI210     m1197(.A0(mai_mai_n1246_), .A1(mai_mai_n1245_), .B0(mai_mai_n336_), .Y(mai_mai_n1247_));
  NO2        m1198(.A(mai_mai_n794_), .B(x1), .Y(mai_mai_n1248_));
  AOI220     m1199(.A0(mai_mai_n1248_), .A1(mai_mai_n614_), .B0(mai_mai_n481_), .B1(mai_mai_n298_), .Y(mai_mai_n1249_));
  NA2        m1200(.A(mai_mai_n502_), .B(mai_mai_n50_), .Y(mai_mai_n1250_));
  AOI220     m1201(.A0(mai_mai_n1250_), .A1(mai_mai_n1194_), .B0(mai_mai_n984_), .B1(mai_mai_n101_), .Y(mai_mai_n1251_));
  NA4        m1202(.A(mai_mai_n1251_), .B(mai_mai_n1249_), .C(mai_mai_n1247_), .D(mai_mai_n1244_), .Y(mai_mai_n1252_));
  AOI220     m1203(.A0(mai_mai_n1252_), .A1(mai_mai_n133_), .B0(mai_mai_n1239_), .B1(mai_mai_n67_), .Y(mai_mai_n1253_));
  NA4        m1204(.A(mai_mai_n1253_), .B(mai_mai_n1228_), .C(mai_mai_n1216_), .D(mai_mai_n1199_), .Y(mai14));
  NO2        m1205(.A(mai_mai_n375_), .B(mai_mai_n71_), .Y(mai_mai_n1255_));
  NO3        m1206(.A(x7), .B(x6), .C(x0), .Y(mai_mai_n1256_));
  OAI210     m1207(.A0(mai_mai_n1256_), .A1(mai_mai_n1255_), .B0(x8), .Y(mai_mai_n1257_));
  NA2        m1208(.A(mai_mai_n1141_), .B(mai_mai_n85_), .Y(mai_mai_n1258_));
  AOI210     m1209(.A0(mai_mai_n1258_), .A1(mai_mai_n1257_), .B0(mai_mai_n158_), .Y(mai_mai_n1259_));
  AOI220     m1210(.A0(mai_mai_n379_), .A1(mai_mai_n855_), .B0(mai_mai_n451_), .B1(mai_mai_n424_), .Y(mai_mai_n1260_));
  NA2        m1211(.A(mai_mai_n281_), .B(mai_mai_n979_), .Y(mai_mai_n1261_));
  OAI220     m1212(.A0(mai_mai_n1261_), .A1(mai_mai_n1260_), .B0(mai_mai_n469_), .B1(mai_mai_n809_), .Y(mai_mai_n1262_));
  OA210      m1213(.A0(mai_mai_n1262_), .A1(mai_mai_n1259_), .B0(x4), .Y(mai_mai_n1263_));
  NO2        m1214(.A(mai_mai_n143_), .B(mai_mai_n612_), .Y(mai_mai_n1264_));
  NA2        m1215(.A(x6), .B(x2), .Y(mai_mai_n1265_));
  NO2        m1216(.A(mai_mai_n630_), .B(mai_mai_n1265_), .Y(mai_mai_n1266_));
  OA210      m1217(.A0(mai_mai_n1264_), .A1(mai_mai_n215_), .B0(mai_mai_n1266_), .Y(mai_mai_n1267_));
  NO4        m1218(.A(mai_mai_n608_), .B(mai_mai_n380_), .C(mai_mai_n302_), .D(mai_mai_n116_), .Y(mai_mai_n1268_));
  OAI210     m1219(.A0(mai_mai_n1268_), .A1(mai_mai_n1267_), .B0(mai_mai_n59_), .Y(mai_mai_n1269_));
  NA2        m1220(.A(x6), .B(mai_mai_n108_), .Y(mai_mai_n1270_));
  NO2        m1221(.A(mai_mai_n669_), .B(mai_mai_n1270_), .Y(mai_mai_n1271_));
  NA2        m1222(.A(mai_mai_n1271_), .B(mai_mai_n931_), .Y(mai_mai_n1272_));
  AOI210     m1223(.A0(mai_mai_n1141_), .A1(mai_mai_n1017_), .B0(x1), .Y(mai_mai_n1273_));
  NO2        m1224(.A(mai_mai_n537_), .B(x5), .Y(mai_mai_n1274_));
  NA3        m1225(.A(mai_mai_n1274_), .B(mai_mai_n123_), .C(x0), .Y(mai_mai_n1275_));
  NA4        m1226(.A(mai_mai_n699_), .B(mai_mai_n932_), .C(mai_mai_n306_), .D(mai_mai_n68_), .Y(mai_mai_n1276_));
  AN4        m1227(.A(mai_mai_n1276_), .B(mai_mai_n1275_), .C(mai_mai_n1273_), .D(mai_mai_n1272_), .Y(mai_mai_n1277_));
  NO2        m1228(.A(mai_mai_n706_), .B(mai_mai_n1101_), .Y(mai_mai_n1278_));
  NO2        m1229(.A(mai_mai_n77_), .B(mai_mai_n58_), .Y(mai_mai_n1279_));
  OAI210     m1230(.A0(mai_mai_n1278_), .A1(mai_mai_n448_), .B0(mai_mai_n1279_), .Y(mai_mai_n1280_));
  AO210      m1231(.A0(mai_mai_n1255_), .A1(mai_mai_n1017_), .B0(mai_mai_n53_), .Y(mai_mai_n1281_));
  AOI210     m1232(.A0(mai_mai_n770_), .A1(mai_mai_n819_), .B0(mai_mai_n1281_), .Y(mai_mai_n1282_));
  AOI220     m1233(.A0(mai_mai_n1282_), .A1(mai_mai_n1280_), .B0(mai_mai_n1277_), .B1(mai_mai_n1269_), .Y(mai_mai_n1283_));
  NO2        m1234(.A(mai_mai_n681_), .B(mai_mai_n169_), .Y(mai_mai_n1284_));
  NO3        m1235(.A(mai_mai_n1284_), .B(mai_mai_n1283_), .C(mai_mai_n1263_), .Y(mai_mai_n1285_));
  NO2        m1236(.A(mai_mai_n324_), .B(x2), .Y(mai_mai_n1286_));
  XN2        m1237(.A(x4), .B(x1), .Y(mai_mai_n1287_));
  NO2        m1238(.A(mai_mai_n1287_), .B(mai_mai_n306_), .Y(mai_mai_n1288_));
  NOi21      m1239(.An(mai_mai_n1288_), .B(mai_mai_n412_), .Y(mai_mai_n1289_));
  NO2        m1240(.A(mai_mai_n343_), .B(mai_mai_n60_), .Y(mai_mai_n1290_));
  OAI210     m1241(.A0(mai_mai_n1290_), .A1(mai_mai_n1289_), .B0(mai_mai_n1286_), .Y(mai_mai_n1291_));
  NA2        m1242(.A(mai_mai_n693_), .B(mai_mai_n56_), .Y(mai_mai_n1292_));
  OAI220     m1243(.A0(mai_mai_n1292_), .A1(mai_mai_n159_), .B0(mai_mai_n193_), .B1(mai_mai_n71_), .Y(mai_mai_n1293_));
  NO2        m1244(.A(mai_mai_n219_), .B(mai_mai_n261_), .Y(mai_mai_n1294_));
  NA2        m1245(.A(mai_mai_n253_), .B(mai_mai_n358_), .Y(mai_mai_n1295_));
  NA2        m1246(.A(mai_mai_n644_), .B(mai_mai_n1035_), .Y(mai_mai_n1296_));
  NO2        m1247(.A(mai_mai_n1296_), .B(mai_mai_n1295_), .Y(mai_mai_n1297_));
  AOI210     m1248(.A0(mai_mai_n1294_), .A1(mai_mai_n1293_), .B0(mai_mai_n1297_), .Y(mai_mai_n1298_));
  AOI210     m1249(.A0(mai_mai_n1298_), .A1(mai_mai_n1291_), .B0(x7), .Y(mai_mai_n1299_));
  NO2        m1250(.A(mai_mai_n496_), .B(x6), .Y(mai_mai_n1300_));
  AOI210     m1251(.A0(mai_mai_n821_), .A1(mai_mai_n962_), .B0(mai_mai_n1300_), .Y(mai_mai_n1301_));
  OAI220     m1252(.A0(mai_mai_n1301_), .A1(mai_mai_n55_), .B0(mai_mai_n496_), .B1(mai_mai_n104_), .Y(mai_mai_n1302_));
  NA2        m1253(.A(mai_mai_n1302_), .B(mai_mai_n360_), .Y(mai_mai_n1303_));
  NA3        m1254(.A(mai_mai_n615_), .B(mai_mai_n1069_), .C(mai_mai_n70_), .Y(mai_mai_n1304_));
  NO4        m1255(.A(mai_mai_n1304_), .B(mai_mai_n1242_), .C(mai_mai_n121_), .D(mai_mai_n55_), .Y(mai_mai_n1305_));
  NO3        m1256(.A(mai_mai_n1062_), .B(mai_mai_n827_), .C(mai_mai_n486_), .Y(mai_mai_n1306_));
  NO3        m1257(.A(mai_mai_n758_), .B(mai_mai_n502_), .C(mai_mai_n54_), .Y(mai_mai_n1307_));
  NO4        m1258(.A(mai_mai_n1307_), .B(mai_mai_n1306_), .C(mai_mai_n1305_), .D(mai_mai_n1040_), .Y(mai_mai_n1308_));
  AOI210     m1259(.A0(mai_mai_n1308_), .A1(mai_mai_n1303_), .B0(mai_mai_n308_), .Y(mai_mai_n1309_));
  NA2        m1260(.A(mai_mai_n904_), .B(mai_mai_n53_), .Y(mai_mai_n1310_));
  OAI210     m1261(.A0(mai_mai_n248_), .A1(mai_mai_n118_), .B0(x2), .Y(mai_mai_n1311_));
  NA2        m1262(.A(mai_mai_n371_), .B(mai_mai_n56_), .Y(mai_mai_n1312_));
  OA220      m1263(.A0(mai_mai_n1312_), .A1(mai_mai_n1311_), .B0(mai_mai_n1310_), .B1(mai_mai_n379_), .Y(mai_mai_n1313_));
  NA3        m1264(.A(mai_mai_n1040_), .B(mai_mai_n742_), .C(mai_mai_n55_), .Y(mai_mai_n1314_));
  NA2        m1265(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n1315_));
  NO2        m1266(.A(mai_mai_n1315_), .B(mai_mai_n200_), .Y(mai_mai_n1316_));
  NA4        m1267(.A(mai_mai_n1316_), .B(mai_mai_n371_), .C(mai_mai_n261_), .D(mai_mai_n67_), .Y(mai_mai_n1317_));
  NA3        m1268(.A(mai_mai_n1248_), .B(mai_mai_n621_), .C(mai_mai_n635_), .Y(mai_mai_n1318_));
  AN3        m1269(.A(mai_mai_n1318_), .B(mai_mai_n1317_), .C(mai_mai_n1314_), .Y(mai_mai_n1319_));
  OAI210     m1270(.A0(mai_mai_n1313_), .A1(mai_mai_n319_), .B0(mai_mai_n1319_), .Y(mai_mai_n1320_));
  NO3        m1271(.A(mai_mai_n1320_), .B(mai_mai_n1309_), .C(mai_mai_n1299_), .Y(mai_mai_n1321_));
  OAI210     m1272(.A0(mai_mai_n1285_), .A1(x3), .B0(mai_mai_n1321_), .Y(mai15));
  NA2        m1273(.A(mai_mai_n590_), .B(mai_mai_n59_), .Y(mai_mai_n1323_));
  NAi41      m1274(.An(x2), .B(x7), .C(x6), .D(x0), .Y(mai_mai_n1324_));
  AOI210     m1275(.A0(mai_mai_n1324_), .A1(mai_mai_n1323_), .B0(mai_mai_n53_), .Y(mai_mai_n1325_));
  NA3        m1276(.A(mai_mai_n57_), .B(x6), .C(mai_mai_n110_), .Y(mai_mai_n1326_));
  NO2        m1277(.A(mai_mai_n1326_), .B(mai_mai_n297_), .Y(mai_mai_n1327_));
  OAI210     m1278(.A0(mai_mai_n1327_), .A1(mai_mai_n1325_), .B0(mai_mai_n1164_), .Y(mai_mai_n1328_));
  NA2        m1279(.A(mai_mai_n112_), .B(mai_mai_n110_), .Y(mai_mai_n1329_));
  NA4        m1280(.A(mai_mai_n1329_), .B(mai_mai_n642_), .C(mai_mai_n312_), .D(x6), .Y(mai_mai_n1330_));
  AOI210     m1281(.A0(mai_mai_n736_), .A1(mai_mai_n76_), .B0(x3), .Y(mai_mai_n1331_));
  NA3        m1282(.A(mai_mai_n1331_), .B(mai_mai_n1330_), .C(mai_mai_n1328_), .Y(mai_mai_n1332_));
  AOI210     m1283(.A0(mai_mai_n1074_), .A1(mai_mai_n594_), .B0(mai_mai_n50_), .Y(mai_mai_n1333_));
  NO2        m1284(.A(mai_mai_n297_), .B(mai_mai_n110_), .Y(mai_mai_n1334_));
  NO2        m1285(.A(mai_mai_n240_), .B(x5), .Y(mai_mai_n1335_));
  NA2        m1286(.A(mai_mai_n1335_), .B(mai_mai_n1334_), .Y(mai_mai_n1336_));
  NA3        m1287(.A(mai_mai_n1248_), .B(mai_mai_n629_), .C(mai_mai_n1176_), .Y(mai_mai_n1337_));
  NA4        m1288(.A(mai_mai_n1337_), .B(mai_mai_n1336_), .C(mai_mai_n1333_), .D(mai_mai_n1275_), .Y(mai_mai_n1338_));
  NA2        m1289(.A(mai_mai_n337_), .B(mai_mai_n346_), .Y(mai_mai_n1339_));
  AOI210     m1290(.A0(mai_mai_n1210_), .A1(mai_mai_n58_), .B0(mai_mai_n1339_), .Y(mai_mai_n1340_));
  NA4        m1291(.A(mai_mai_n1210_), .B(mai_mai_n705_), .C(mai_mai_n1138_), .D(mai_mai_n384_), .Y(mai_mai_n1341_));
  NA2        m1292(.A(mai_mai_n594_), .B(mai_mai_n470_), .Y(mai_mai_n1342_));
  NO2        m1293(.A(mai_mai_n758_), .B(mai_mai_n53_), .Y(mai_mai_n1343_));
  NO2        m1294(.A(mai_mai_n783_), .B(mai_mai_n302_), .Y(mai_mai_n1344_));
  NA2        m1295(.A(mai_mai_n1344_), .B(mai_mai_n1343_), .Y(mai_mai_n1345_));
  NA3        m1296(.A(mai_mai_n1345_), .B(mai_mai_n1342_), .C(mai_mai_n1341_), .Y(mai_mai_n1346_));
  OAI210     m1297(.A0(mai_mai_n1346_), .A1(mai_mai_n1340_), .B0(mai_mai_n77_), .Y(mai_mai_n1347_));
  NA2        m1298(.A(mai_mai_n373_), .B(mai_mai_n708_), .Y(mai_mai_n1348_));
  NA2        m1299(.A(mai_mai_n575_), .B(mai_mai_n56_), .Y(mai_mai_n1349_));
  NA3        m1300(.A(mai_mai_n1349_), .B(mai_mai_n346_), .C(mai_mai_n112_), .Y(mai_mai_n1350_));
  AOI210     m1301(.A0(mai_mai_n1350_), .A1(mai_mai_n1348_), .B0(mai_mai_n502_), .Y(mai_mai_n1351_));
  NO3        m1302(.A(mai_mai_n807_), .B(mai_mai_n626_), .C(mai_mai_n201_), .Y(mai_mai_n1352_));
  OAI210     m1303(.A0(mai_mai_n1352_), .A1(mai_mai_n1351_), .B0(mai_mai_n496_), .Y(mai_mai_n1353_));
  NO2        m1304(.A(mai_mai_n877_), .B(mai_mai_n50_), .Y(mai_mai_n1354_));
  NO2        m1305(.A(mai_mai_n250_), .B(mai_mai_n64_), .Y(mai_mai_n1355_));
  OA210      m1306(.A0(mai_mai_n1355_), .A1(mai_mai_n1354_), .B0(mai_mai_n412_), .Y(mai_mai_n1356_));
  NA2        m1307(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n1357_));
  AOI210     m1308(.A0(mai_mai_n985_), .A1(mai_mai_n1357_), .B0(mai_mai_n687_), .Y(mai_mai_n1358_));
  OAI210     m1309(.A0(mai_mai_n1358_), .A1(mai_mai_n1356_), .B0(mai_mai_n1025_), .Y(mai_mai_n1359_));
  NA2        m1310(.A(mai_mai_n1316_), .B(mai_mai_n68_), .Y(mai_mai_n1360_));
  NO2        m1311(.A(mai_mai_n1265_), .B(x0), .Y(mai_mai_n1361_));
  AOI210     m1312(.A0(mai_mai_n1361_), .A1(mai_mai_n609_), .B0(x8), .Y(mai_mai_n1362_));
  NO2        m1313(.A(mai_mai_n433_), .B(mai_mai_n81_), .Y(mai_mai_n1363_));
  NO2        m1314(.A(mai_mai_n936_), .B(mai_mai_n71_), .Y(mai_mai_n1364_));
  NA2        m1315(.A(mai_mai_n1364_), .B(mai_mai_n1363_), .Y(mai_mai_n1365_));
  NO2        m1316(.A(mai_mai_n983_), .B(x6), .Y(mai_mai_n1366_));
  NA4        m1317(.A(mai_mai_n1366_), .B(mai_mai_n599_), .C(mai_mai_n160_), .D(mai_mai_n416_), .Y(mai_mai_n1367_));
  AN4        m1318(.A(mai_mai_n1367_), .B(mai_mai_n1365_), .C(mai_mai_n1362_), .D(mai_mai_n1360_), .Y(mai_mai_n1368_));
  NA4        m1319(.A(mai_mai_n1368_), .B(mai_mai_n1359_), .C(mai_mai_n1353_), .D(mai_mai_n1347_), .Y(mai_mai_n1369_));
  NA2        m1320(.A(mai_mai_n166_), .B(mai_mai_n742_), .Y(mai_mai_n1370_));
  NO2        m1321(.A(mai_mai_n654_), .B(x2), .Y(mai_mai_n1371_));
  OAI210     m1322(.A0(mai_mai_n68_), .A1(mai_mai_n53_), .B0(mai_mai_n145_), .Y(mai_mai_n1372_));
  OAI210     m1323(.A0(mai_mai_n1371_), .A1(mai_mai_n85_), .B0(mai_mai_n1372_), .Y(mai_mai_n1373_));
  AOI210     m1324(.A0(mai_mai_n1373_), .A1(mai_mai_n1370_), .B0(mai_mai_n324_), .Y(mai_mai_n1374_));
  NO3        m1325(.A(mai_mai_n1326_), .B(mai_mai_n269_), .C(mai_mai_n250_), .Y(mai_mai_n1375_));
  NA3        m1326(.A(mai_mai_n57_), .B(x1), .C(x0), .Y(mai_mai_n1376_));
  NA3        m1327(.A(mai_mai_n71_), .B(x5), .C(x2), .Y(mai_mai_n1377_));
  NA4        m1328(.A(x7), .B(x3), .C(mai_mai_n53_), .D(x0), .Y(mai_mai_n1378_));
  OAI220     m1329(.A0(mai_mai_n1378_), .A1(x6), .B0(mai_mai_n1377_), .B1(mai_mai_n1376_), .Y(mai_mai_n1379_));
  NO2        m1330(.A(mai_mai_n1379_), .B(mai_mai_n1375_), .Y(mai_mai_n1380_));
  NAi21      m1331(.An(mai_mai_n116_), .B(mai_mai_n752_), .Y(mai_mai_n1381_));
  NA4        m1332(.A(mai_mai_n1381_), .B(mai_mai_n322_), .C(mai_mai_n292_), .D(mai_mai_n629_), .Y(mai_mai_n1382_));
  OAI220     m1333(.A0(mai_mai_n327_), .A1(x7), .B0(mai_mai_n132_), .B1(mai_mai_n71_), .Y(mai_mai_n1383_));
  NA3        m1334(.A(mai_mai_n1383_), .B(mai_mai_n794_), .C(mai_mai_n1104_), .Y(mai_mai_n1384_));
  NA2        m1335(.A(mai_mai_n82_), .B(mai_mai_n50_), .Y(mai_mai_n1385_));
  AO210      m1336(.A0(mai_mai_n1385_), .A1(mai_mai_n317_), .B0(mai_mai_n158_), .Y(mai_mai_n1386_));
  NA4        m1337(.A(mai_mai_n1386_), .B(mai_mai_n1384_), .C(mai_mai_n1382_), .D(mai_mai_n1380_), .Y(mai_mai_n1387_));
  OAI210     m1338(.A0(mai_mai_n1387_), .A1(mai_mai_n1374_), .B0(mai_mai_n56_), .Y(mai_mai_n1388_));
  AOI210     m1339(.A0(mai_mai_n695_), .A1(x4), .B0(mai_mai_n962_), .Y(mai_mai_n1389_));
  OAI220     m1340(.A0(mai_mai_n1389_), .A1(mai_mai_n303_), .B0(mai_mai_n1029_), .B1(mai_mai_n950_), .Y(mai_mai_n1390_));
  NA2        m1341(.A(mai_mai_n838_), .B(mai_mai_n409_), .Y(mai_mai_n1391_));
  OAI210     m1342(.A0(mai_mai_n1363_), .A1(mai_mai_n1355_), .B0(mai_mai_n293_), .Y(mai_mai_n1392_));
  OAI210     m1343(.A0(mai_mai_n1391_), .A1(mai_mai_n850_), .B0(mai_mai_n1392_), .Y(mai_mai_n1393_));
  OAI210     m1344(.A0(mai_mai_n1393_), .A1(mai_mai_n1390_), .B0(x6), .Y(mai_mai_n1394_));
  NO2        m1345(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n1395_));
  NO2        m1346(.A(x7), .B(x5), .Y(mai_mai_n1396_));
  AOI220     m1347(.A0(mai_mai_n859_), .A1(mai_mai_n1395_), .B0(mai_mai_n541_), .B1(mai_mai_n1396_), .Y(mai_mai_n1397_));
  NA2        m1348(.A(mai_mai_n767_), .B(mai_mai_n293_), .Y(mai_mai_n1398_));
  NA3        m1349(.A(mai_mai_n621_), .B(mai_mai_n295_), .C(mai_mai_n245_), .Y(mai_mai_n1399_));
  NA3        m1350(.A(mai_mai_n1399_), .B(mai_mai_n1398_), .C(mai_mai_n1397_), .Y(mai_mai_n1400_));
  NA2        m1351(.A(mai_mai_n1400_), .B(mai_mai_n427_), .Y(mai_mai_n1401_));
  AOI210     m1352(.A0(mai_mai_n382_), .A1(mai_mai_n344_), .B0(mai_mai_n55_), .Y(mai_mai_n1402_));
  NA4        m1353(.A(mai_mai_n1402_), .B(mai_mai_n1401_), .C(mai_mai_n1394_), .D(mai_mai_n1388_), .Y(mai_mai_n1403_));
  AO220      m1354(.A0(mai_mai_n1403_), .A1(mai_mai_n1369_), .B0(mai_mai_n1338_), .B1(mai_mai_n1332_), .Y(mai16));
  NO2        m1355(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n1405_));
  NA2        m1356(.A(mai_mai_n668_), .B(mai_mai_n538_), .Y(mai_mai_n1406_));
  NA3        m1357(.A(mai_mai_n234_), .B(mai_mai_n434_), .C(mai_mai_n962_), .Y(mai_mai_n1407_));
  NA2        m1358(.A(mai_mai_n135_), .B(mai_mai_n210_), .Y(mai_mai_n1408_));
  AOI210     m1359(.A0(mai_mai_n1407_), .A1(mai_mai_n1406_), .B0(mai_mai_n1408_), .Y(mai_mai_n1409_));
  NO3        m1360(.A(x8), .B(x6), .C(mai_mai_n50_), .Y(mai_mai_n1410_));
  NO2        m1361(.A(mai_mai_n740_), .B(mai_mai_n188_), .Y(mai_mai_n1411_));
  OAI210     m1362(.A0(mai_mai_n1410_), .A1(mai_mai_n242_), .B0(mai_mai_n1411_), .Y(mai_mai_n1412_));
  NO2        m1363(.A(mai_mai_n162_), .B(x5), .Y(mai_mai_n1413_));
  NA2        m1364(.A(mai_mai_n1413_), .B(mai_mai_n1371_), .Y(mai_mai_n1414_));
  NA3        m1365(.A(mai_mai_n584_), .B(mai_mai_n540_), .C(mai_mai_n480_), .Y(mai_mai_n1415_));
  NA3        m1366(.A(mai_mai_n1415_), .B(mai_mai_n1414_), .C(mai_mai_n1412_), .Y(mai_mai_n1416_));
  OAI210     m1367(.A0(mai_mai_n1416_), .A1(mai_mai_n1409_), .B0(mai_mai_n1405_), .Y(mai_mai_n1417_));
  NO2        m1368(.A(mai_mai_n324_), .B(x7), .Y(mai_mai_n1418_));
  NA2        m1369(.A(mai_mai_n1418_), .B(x0), .Y(mai_mai_n1419_));
  NO2        m1370(.A(mai_mai_n1419_), .B(mai_mai_n643_), .Y(mai_mai_n1420_));
  NA2        m1371(.A(mai_mai_n1083_), .B(mai_mai_n201_), .Y(mai_mai_n1421_));
  NA2        m1372(.A(mai_mai_n55_), .B(mai_mai_n108_), .Y(mai_mai_n1422_));
  NA2        m1373(.A(mai_mai_n1422_), .B(mai_mai_n689_), .Y(mai_mai_n1423_));
  NA2        m1374(.A(mai_mai_n381_), .B(mai_mai_n1087_), .Y(mai_mai_n1424_));
  OA220      m1375(.A0(mai_mai_n1424_), .A1(mai_mai_n1423_), .B0(mai_mai_n1421_), .B1(mai_mai_n637_), .Y(mai_mai_n1425_));
  NO2        m1376(.A(mai_mai_n1425_), .B(mai_mai_n658_), .Y(mai_mai_n1426_));
  INV        m1377(.A(mai_mai_n1025_), .Y(mai_mai_n1427_));
  NO2        m1378(.A(mai_mai_n1427_), .B(mai_mai_n62_), .Y(mai_mai_n1428_));
  AOI220     m1379(.A0(mai_mai_n1428_), .A1(mai_mai_n272_), .B0(mai_mai_n1271_), .B1(mai_mai_n128_), .Y(mai_mai_n1429_));
  AOI220     m1380(.A0(mai_mai_n642_), .A1(mai_mai_n367_), .B0(mai_mai_n629_), .B1(mai_mai_n88_), .Y(mai_mai_n1430_));
  NA3        m1381(.A(mai_mai_n467_), .B(mai_mai_n591_), .C(mai_mai_n195_), .Y(mai_mai_n1431_));
  OAI220     m1382(.A0(mai_mai_n1431_), .A1(mai_mai_n1430_), .B0(mai_mai_n1429_), .B1(mai_mai_n313_), .Y(mai_mai_n1432_));
  NO3        m1383(.A(mai_mai_n1432_), .B(mai_mai_n1426_), .C(mai_mai_n1420_), .Y(mai_mai_n1433_));
  NO3        m1384(.A(x6), .B(x4), .C(x3), .Y(mai_mai_n1434_));
  NA2        m1385(.A(mai_mai_n1434_), .B(mai_mai_n537_), .Y(mai_mai_n1435_));
  NA4        m1386(.A(mai_mai_n713_), .B(mai_mai_n188_), .C(mai_mai_n58_), .D(x6), .Y(mai_mai_n1436_));
  AOI210     m1387(.A0(mai_mai_n1436_), .A1(mai_mai_n1435_), .B0(mai_mai_n54_), .Y(mai_mai_n1437_));
  NO2        m1388(.A(mai_mai_n728_), .B(x3), .Y(mai_mai_n1438_));
  NO3        m1389(.A(mai_mai_n502_), .B(mai_mai_n223_), .C(mai_mai_n75_), .Y(mai_mai_n1439_));
  NO2        m1390(.A(mai_mai_n767_), .B(mai_mai_n514_), .Y(mai_mai_n1440_));
  NO3        m1391(.A(mai_mai_n1440_), .B(mai_mai_n263_), .C(mai_mai_n157_), .Y(mai_mai_n1441_));
  NO3        m1392(.A(mai_mai_n1441_), .B(mai_mai_n1439_), .C(mai_mai_n1437_), .Y(mai_mai_n1442_));
  NA2        m1393(.A(mai_mai_n410_), .B(mai_mai_n962_), .Y(mai_mai_n1443_));
  NA4        m1394(.A(mai_mai_n486_), .B(mai_mai_n375_), .C(mai_mai_n225_), .D(x6), .Y(mai_mai_n1444_));
  OAI210     m1395(.A0(mai_mai_n728_), .A1(mai_mai_n1443_), .B0(mai_mai_n1444_), .Y(mai_mai_n1445_));
  NA2        m1396(.A(mai_mai_n913_), .B(mai_mai_n1315_), .Y(mai_mai_n1446_));
  NA2        m1397(.A(mai_mai_n737_), .B(x7), .Y(mai_mai_n1447_));
  OAI210     m1398(.A0(mai_mai_n1447_), .A1(mai_mai_n391_), .B0(mai_mai_n1446_), .Y(mai_mai_n1448_));
  NA2        m1399(.A(mai_mai_n279_), .B(x2), .Y(mai_mai_n1449_));
  NO3        m1400(.A(mai_mai_n1449_), .B(mai_mai_n599_), .C(mai_mai_n72_), .Y(mai_mai_n1450_));
  OA210      m1401(.A0(mai_mai_n1270_), .A1(mai_mai_n58_), .B0(mai_mai_n784_), .Y(mai_mai_n1451_));
  AOI210     m1402(.A0(mai_mai_n584_), .A1(mai_mai_n50_), .B0(mai_mai_n594_), .Y(mai_mai_n1452_));
  OAI210     m1403(.A0(mai_mai_n932_), .A1(mai_mai_n949_), .B0(mai_mai_n386_), .Y(mai_mai_n1453_));
  OAI220     m1404(.A0(mai_mai_n1453_), .A1(mai_mai_n1452_), .B0(mai_mai_n1451_), .B1(mai_mai_n193_), .Y(mai_mai_n1454_));
  NO4        m1405(.A(mai_mai_n1454_), .B(mai_mai_n1450_), .C(mai_mai_n1448_), .D(mai_mai_n1445_), .Y(mai_mai_n1455_));
  OA220      m1406(.A0(mai_mai_n1455_), .A1(mai_mai_n447_), .B0(mai_mai_n1442_), .B1(mai_mai_n208_), .Y(mai_mai_n1456_));
  NO2        m1407(.A(mai_mai_n927_), .B(mai_mai_n55_), .Y(mai_mai_n1457_));
  NA2        m1408(.A(mai_mai_n421_), .B(mai_mai_n809_), .Y(mai_mai_n1458_));
  NO2        m1409(.A(mai_mai_n1458_), .B(mai_mai_n1457_), .Y(mai_mai_n1459_));
  NO3        m1410(.A(mai_mai_n963_), .B(mai_mai_n337_), .C(x8), .Y(mai_mai_n1460_));
  OAI210     m1411(.A0(mai_mai_n1460_), .A1(mai_mai_n1459_), .B0(x6), .Y(mai_mai_n1461_));
  NO2        m1412(.A(mai_mai_n1099_), .B(mai_mai_n1061_), .Y(mai_mai_n1462_));
  NA2        m1413(.A(mai_mai_n193_), .B(x7), .Y(mai_mai_n1463_));
  OAI220     m1414(.A0(mai_mai_n1463_), .A1(mai_mai_n1462_), .B0(mai_mai_n769_), .B1(mai_mai_n87_), .Y(mai_mai_n1464_));
  NA2        m1415(.A(mai_mai_n1464_), .B(mai_mai_n932_), .Y(mai_mai_n1465_));
  NA2        m1416(.A(mai_mai_n879_), .B(mai_mai_n71_), .Y(mai_mai_n1466_));
  OAI210     m1417(.A0(mai_mai_n1466_), .A1(mai_mai_n160_), .B0(mai_mai_n1014_), .Y(mai_mai_n1467_));
  AOI210     m1418(.A0(mai_mai_n502_), .A1(mai_mai_n57_), .B0(mai_mai_n637_), .Y(mai_mai_n1468_));
  NA3        m1419(.A(mai_mai_n231_), .B(mai_mai_n76_), .C(mai_mai_n71_), .Y(mai_mai_n1469_));
  OAI210     m1420(.A0(mai_mai_n923_), .A1(mai_mai_n234_), .B0(mai_mai_n1469_), .Y(mai_mai_n1470_));
  AOI210     m1421(.A0(mai_mai_n1468_), .A1(mai_mai_n1467_), .B0(mai_mai_n1470_), .Y(mai_mai_n1471_));
  NA3        m1422(.A(mai_mai_n1471_), .B(mai_mai_n1465_), .C(mai_mai_n1461_), .Y(mai_mai_n1472_));
  NO2        m1423(.A(mai_mai_n644_), .B(x6), .Y(mai_mai_n1473_));
  OAI210     m1424(.A0(mai_mai_n386_), .A1(mai_mai_n84_), .B0(mai_mai_n384_), .Y(mai_mai_n1474_));
  OA210      m1425(.A0(mai_mai_n1474_), .A1(mai_mai_n1473_), .B0(mai_mai_n133_), .Y(mai_mai_n1475_));
  NO3        m1426(.A(mai_mai_n449_), .B(mai_mai_n389_), .C(x7), .Y(mai_mai_n1476_));
  NO3        m1427(.A(mai_mai_n162_), .B(mai_mai_n75_), .C(x2), .Y(mai_mai_n1477_));
  NO3        m1428(.A(mai_mai_n1477_), .B(mai_mai_n1476_), .C(mai_mai_n1475_), .Y(mai_mai_n1478_));
  NO2        m1429(.A(mai_mai_n234_), .B(x1), .Y(mai_mai_n1479_));
  OAI210     m1430(.A0(mai_mai_n1479_), .A1(mai_mai_n454_), .B0(mai_mai_n514_), .Y(mai_mai_n1480_));
  NO2        m1431(.A(mai_mai_n57_), .B(mai_mai_n108_), .Y(mai_mai_n1481_));
  NA2        m1432(.A(mai_mai_n1092_), .B(mai_mai_n1481_), .Y(mai_mai_n1482_));
  AOI210     m1433(.A0(mai_mai_n1482_), .A1(mai_mai_n1480_), .B0(mai_mai_n56_), .Y(mai_mai_n1483_));
  AOI220     m1434(.A0(mai_mai_n769_), .A1(mai_mai_n780_), .B0(mai_mai_n517_), .B1(mai_mai_n283_), .Y(mai_mai_n1484_));
  NO2        m1435(.A(mai_mai_n1484_), .B(mai_mai_n1315_), .Y(mai_mai_n1485_));
  NO3        m1436(.A(mai_mai_n537_), .B(mai_mai_n175_), .C(mai_mai_n1061_), .Y(mai_mai_n1486_));
  NA2        m1437(.A(mai_mai_n949_), .B(x4), .Y(mai_mai_n1487_));
  OAI220     m1438(.A0(mai_mai_n1487_), .A1(mai_mai_n694_), .B0(mai_mai_n652_), .B1(mai_mai_n615_), .Y(mai_mai_n1488_));
  NO4        m1439(.A(mai_mai_n1488_), .B(mai_mai_n1486_), .C(mai_mai_n1485_), .D(mai_mai_n1483_), .Y(mai_mai_n1489_));
  OAI210     m1440(.A0(mai_mai_n1478_), .A1(x5), .B0(mai_mai_n1489_), .Y(mai_mai_n1490_));
  AOI220     m1441(.A0(mai_mai_n1490_), .A1(mai_mai_n99_), .B0(mai_mai_n1472_), .B1(mai_mai_n344_), .Y(mai_mai_n1491_));
  NA4        m1442(.A(mai_mai_n1491_), .B(mai_mai_n1456_), .C(mai_mai_n1433_), .D(mai_mai_n1417_), .Y(mai17));
  NO4        m1443(.A(mai_mai_n606_), .B(mai_mai_n707_), .C(mai_mai_n102_), .D(mai_mai_n101_), .Y(mai_mai_n1493_));
  NO2        m1444(.A(mai_mai_n126_), .B(mai_mai_n1176_), .Y(mai_mai_n1494_));
  AOI220     m1445(.A0(mai_mai_n1494_), .A1(mai_mai_n723_), .B0(mai_mai_n1493_), .B1(mai_mai_n508_), .Y(mai_mai_n1495_));
  NA2        m1446(.A(mai_mai_n166_), .B(mai_mai_n78_), .Y(mai_mai_n1496_));
  NOi21      m1447(.An(mai_mai_n384_), .B(mai_mai_n84_), .Y(mai_mai_n1497_));
  OAI210     m1448(.A0(mai_mai_n629_), .A1(mai_mai_n55_), .B0(mai_mai_n1497_), .Y(mai_mai_n1498_));
  NA2        m1449(.A(mai_mai_n1229_), .B(mai_mai_n1020_), .Y(mai_mai_n1499_));
  NA4        m1450(.A(mai_mai_n1499_), .B(mai_mai_n1498_), .C(mai_mai_n740_), .D(mai_mai_n57_), .Y(mai_mai_n1500_));
  OAI210     m1451(.A0(mai_mai_n713_), .A1(x8), .B0(mai_mai_n1315_), .Y(mai_mai_n1501_));
  NA3        m1452(.A(mai_mai_n1501_), .B(mai_mai_n1255_), .C(mai_mai_n403_), .Y(mai_mai_n1502_));
  NA3        m1453(.A(mai_mai_n397_), .B(mai_mai_n272_), .C(mai_mai_n590_), .Y(mai_mai_n1503_));
  OA210      m1454(.A0(mai_mai_n1326_), .A1(mai_mai_n1169_), .B0(mai_mai_n760_), .Y(mai_mai_n1504_));
  NA4        m1455(.A(mai_mai_n1504_), .B(mai_mai_n1503_), .C(mai_mai_n1502_), .D(mai_mai_n1500_), .Y(mai_mai_n1505_));
  NA3        m1456(.A(mai_mai_n165_), .B(mai_mai_n635_), .C(mai_mai_n1061_), .Y(mai_mai_n1506_));
  AOI210     m1457(.A0(mai_mai_n1089_), .A1(mai_mai_n309_), .B0(mai_mai_n59_), .Y(mai_mai_n1507_));
  NA2        m1458(.A(mai_mai_n1507_), .B(mai_mai_n1506_), .Y(mai_mai_n1508_));
  AOI210     m1459(.A0(mai_mai_n1505_), .A1(x1), .B0(mai_mai_n1508_), .Y(mai_mai_n1509_));
  NO2        m1460(.A(mai_mai_n988_), .B(mai_mai_n502_), .Y(mai_mai_n1510_));
  OAI210     m1461(.A0(mai_mai_n1510_), .A1(mai_mai_n1073_), .B0(mai_mai_n612_), .Y(mai_mai_n1511_));
  NO3        m1462(.A(mai_mai_n637_), .B(mai_mai_n559_), .C(mai_mai_n528_), .Y(mai_mai_n1512_));
  OAI210     m1463(.A0(mai_mai_n1512_), .A1(mai_mai_n912_), .B0(mai_mai_n1438_), .Y(mai_mai_n1513_));
  AOI210     m1464(.A0(mai_mai_n1513_), .A1(mai_mai_n1511_), .B0(x8), .Y(mai_mai_n1514_));
  NA3        m1465(.A(mai_mai_n637_), .B(mai_mai_n275_), .C(mai_mai_n123_), .Y(mai_mai_n1515_));
  NO2        m1466(.A(mai_mai_n145_), .B(mai_mai_n144_), .Y(mai_mai_n1516_));
  NO3        m1467(.A(mai_mai_n907_), .B(mai_mai_n780_), .C(mai_mai_n707_), .Y(mai_mai_n1517_));
  AOI210     m1468(.A0(mai_mai_n1517_), .A1(mai_mai_n1516_), .B0(x0), .Y(mai_mai_n1518_));
  OAI210     m1469(.A0(mai_mai_n1515_), .A1(mai_mai_n252_), .B0(mai_mai_n1518_), .Y(mai_mai_n1519_));
  NO2        m1470(.A(mai_mai_n1519_), .B(mai_mai_n1514_), .Y(mai_mai_n1520_));
  OAI220     m1471(.A0(mai_mai_n1520_), .A1(mai_mai_n1509_), .B0(mai_mai_n1496_), .B1(mai_mai_n1495_), .Y(mai18));
  AOI210     m1472(.A0(x8), .A1(x0), .B0(x5), .Y(mai_mai_n1522_));
  NOi31      m1473(.An(mai_mai_n309_), .B(mai_mai_n1522_), .C(mai_mai_n1059_), .Y(mai_mai_n1523_));
  NA2        m1474(.A(mai_mai_n606_), .B(mai_mai_n59_), .Y(mai_mai_n1524_));
  AOI210     m1475(.A0(mai_mai_n1421_), .A1(mai_mai_n355_), .B0(mai_mai_n1524_), .Y(mai_mai_n1525_));
  NO2        m1476(.A(mai_mai_n622_), .B(mai_mai_n781_), .Y(mai_mai_n1526_));
  NO4        m1477(.A(mai_mai_n259_), .B(mai_mai_n819_), .C(mai_mai_n156_), .D(mai_mai_n70_), .Y(mai_mai_n1527_));
  NO4        m1478(.A(mai_mai_n1527_), .B(mai_mai_n1526_), .C(mai_mai_n1525_), .D(mai_mai_n1523_), .Y(mai_mai_n1528_));
  NA3        m1479(.A(mai_mai_n523_), .B(mai_mai_n219_), .C(x0), .Y(mai_mai_n1529_));
  NAi21      m1480(.An(mai_mai_n390_), .B(mai_mai_n1529_), .Y(mai_mai_n1530_));
  NO2        m1481(.A(mai_mai_n897_), .B(x5), .Y(mai_mai_n1531_));
  AOI210     m1482(.A0(mai_mai_n1154_), .A1(x5), .B0(mai_mai_n1531_), .Y(mai_mai_n1532_));
  OA220      m1483(.A0(mai_mai_n523_), .A1(mai_mai_n337_), .B0(mai_mai_n403_), .B1(x5), .Y(mai_mai_n1533_));
  OAI220     m1484(.A0(mai_mai_n1533_), .A1(mai_mai_n297_), .B0(mai_mai_n1532_), .B1(mai_mai_n217_), .Y(mai_mai_n1534_));
  AOI210     m1485(.A0(mai_mai_n1530_), .A1(mai_mai_n295_), .B0(mai_mai_n1534_), .Y(mai_mai_n1535_));
  AOI210     m1486(.A0(mai_mai_n1535_), .A1(mai_mai_n1528_), .B0(x6), .Y(mai_mai_n1536_));
  NA3        m1487(.A(mai_mai_n527_), .B(mai_mai_n424_), .C(x2), .Y(mai_mai_n1537_));
  NA3        m1488(.A(mai_mai_n1059_), .B(mai_mai_n51_), .C(mai_mai_n57_), .Y(mai_mai_n1538_));
  AOI210     m1489(.A0(mai_mai_n1538_), .A1(mai_mai_n1537_), .B0(mai_mai_n794_), .Y(mai_mai_n1539_));
  AOI210     m1490(.A0(mai_mai_n428_), .A1(mai_mai_n140_), .B0(mai_mai_n792_), .Y(mai_mai_n1540_));
  NA2        m1491(.A(mai_mai_n272_), .B(x6), .Y(mai_mai_n1541_));
  OAI210     m1492(.A0(mai_mai_n181_), .A1(mai_mai_n110_), .B0(mai_mai_n1160_), .Y(mai_mai_n1542_));
  OAI220     m1493(.A0(mai_mai_n1542_), .A1(mai_mai_n1541_), .B0(mai_mai_n1540_), .B1(mai_mai_n752_), .Y(mai_mai_n1543_));
  OAI210     m1494(.A0(mai_mai_n1543_), .A1(mai_mai_n1539_), .B0(mai_mai_n53_), .Y(mai_mai_n1544_));
  NO2        m1495(.A(mai_mai_n693_), .B(mai_mai_n266_), .Y(mai_mai_n1545_));
  NO2        m1496(.A(mai_mai_n269_), .B(x3), .Y(mai_mai_n1546_));
  NO3        m1497(.A(mai_mai_n438_), .B(mai_mai_n606_), .C(mai_mai_n843_), .Y(mai_mai_n1547_));
  OAI210     m1498(.A0(mai_mai_n1547_), .A1(mai_mai_n1545_), .B0(mai_mai_n1546_), .Y(mai_mai_n1548_));
  AOI210     m1499(.A0(mai_mai_n1163_), .A1(mai_mai_n621_), .B0(x4), .Y(mai_mai_n1549_));
  OAI210     m1500(.A0(mai_mai_n559_), .A1(mai_mai_n606_), .B0(mai_mai_n59_), .Y(mai_mai_n1550_));
  OAI210     m1501(.A0(mai_mai_n629_), .A1(mai_mai_n654_), .B0(mai_mai_n1550_), .Y(mai_mai_n1551_));
  AO220      m1502(.A0(mai_mai_n1274_), .A1(mai_mai_n740_), .B0(mai_mai_n560_), .B1(mai_mai_n360_), .Y(mai_mai_n1552_));
  AOI220     m1503(.A0(mai_mai_n1552_), .A1(x1), .B0(mai_mai_n1551_), .B1(mai_mai_n163_), .Y(mai_mai_n1553_));
  NA4        m1504(.A(mai_mai_n1553_), .B(mai_mai_n1549_), .C(mai_mai_n1548_), .D(mai_mai_n1544_), .Y(mai_mai_n1554_));
  NO3        m1505(.A(mai_mai_n1080_), .B(mai_mai_n133_), .C(mai_mai_n132_), .Y(mai_mai_n1555_));
  OAI210     m1506(.A0(mai_mai_n1555_), .A1(mai_mai_n659_), .B0(mai_mai_n108_), .Y(mai_mai_n1556_));
  AOI210     m1507(.A0(mai_mai_n1556_), .A1(mai_mai_n565_), .B0(mai_mai_n794_), .Y(mai_mai_n1557_));
  NA3        m1508(.A(mai_mai_n1222_), .B(mai_mai_n193_), .C(mai_mai_n143_), .Y(mai_mai_n1558_));
  NA3        m1509(.A(mai_mai_n1083_), .B(mai_mai_n783_), .C(mai_mai_n348_), .Y(mai_mai_n1559_));
  NA2        m1510(.A(mai_mai_n173_), .B(mai_mai_n780_), .Y(mai_mai_n1560_));
  OAI210     m1511(.A0(mai_mai_n1560_), .A1(mai_mai_n1329_), .B0(mai_mai_n1559_), .Y(mai_mai_n1561_));
  AOI210     m1512(.A0(mai_mai_n1558_), .A1(mai_mai_n180_), .B0(mai_mai_n1561_), .Y(mai_mai_n1562_));
  OAI210     m1513(.A0(mai_mai_n1562_), .A1(mai_mai_n546_), .B0(x4), .Y(mai_mai_n1563_));
  OAI220     m1514(.A0(mai_mai_n1563_), .A1(mai_mai_n1557_), .B0(mai_mai_n1554_), .B1(mai_mai_n1536_), .Y(mai_mai_n1564_));
  NO2        m1515(.A(mai_mai_n148_), .B(mai_mai_n124_), .Y(mai_mai_n1565_));
  NO2        m1516(.A(mai_mai_n193_), .B(mai_mai_n809_), .Y(mai_mai_n1566_));
  AOI210     m1517(.A0(mai_mai_n607_), .A1(mai_mai_n514_), .B0(mai_mai_n1566_), .Y(mai_mai_n1567_));
  NO2        m1518(.A(mai_mai_n1567_), .B(x6), .Y(mai_mai_n1568_));
  NO2        m1519(.A(mai_mai_n389_), .B(mai_mai_n258_), .Y(mai_mai_n1569_));
  NO2        m1520(.A(mai_mai_n133_), .B(mai_mai_n742_), .Y(mai_mai_n1570_));
  NO2        m1521(.A(mai_mai_n963_), .B(mai_mai_n590_), .Y(mai_mai_n1571_));
  AO220      m1522(.A0(mai_mai_n1571_), .A1(mai_mai_n1570_), .B0(mai_mai_n1569_), .B1(mai_mai_n126_), .Y(mai_mai_n1572_));
  NO3        m1523(.A(mai_mai_n1572_), .B(mai_mai_n1568_), .C(mai_mai_n1565_), .Y(mai_mai_n1573_));
  NA2        m1524(.A(mai_mai_n1080_), .B(x3), .Y(mai_mai_n1574_));
  NA2        m1525(.A(mai_mai_n1366_), .B(mai_mai_n135_), .Y(mai_mai_n1575_));
  OAI220     m1526(.A0(mai_mai_n1575_), .A1(mai_mai_n1574_), .B0(mai_mai_n1573_), .B1(x3), .Y(mai_mai_n1576_));
  NO3        m1527(.A(mai_mai_n1010_), .B(mai_mai_n693_), .C(mai_mai_n332_), .Y(mai_mai_n1577_));
  AO210      m1528(.A0(mai_mai_n1039_), .A1(mai_mai_n302_), .B0(mai_mai_n1577_), .Y(mai_mai_n1578_));
  AOI220     m1529(.A0(mai_mai_n1578_), .A1(x8), .B0(mai_mai_n1366_), .B1(mai_mai_n439_), .Y(mai_mai_n1579_));
  NA2        m1530(.A(mai_mai_n756_), .B(mai_mai_n323_), .Y(mai_mai_n1580_));
  NO4        m1531(.A(mai_mai_n373_), .B(mai_mai_n206_), .C(mai_mai_n343_), .D(x2), .Y(mai_mai_n1581_));
  NA2        m1532(.A(mai_mai_n1422_), .B(mai_mai_n110_), .Y(mai_mai_n1582_));
  NO3        m1533(.A(mai_mai_n1223_), .B(mai_mai_n1003_), .C(mai_mai_n1160_), .Y(mai_mai_n1583_));
  AOI210     m1534(.A0(mai_mai_n1583_), .A1(mai_mai_n1582_), .B0(mai_mai_n1581_), .Y(mai_mai_n1584_));
  OA220      m1535(.A0(mai_mai_n1584_), .A1(mai_mai_n963_), .B0(mai_mai_n1580_), .B1(mai_mai_n574_), .Y(mai_mai_n1585_));
  OAI210     m1536(.A0(mai_mai_n1579_), .A1(mai_mai_n413_), .B0(mai_mai_n1585_), .Y(mai_mai_n1586_));
  AOI210     m1537(.A0(mai_mai_n1576_), .A1(mai_mai_n140_), .B0(mai_mai_n1586_), .Y(mai_mai_n1587_));
  NA2        m1538(.A(mai_mai_n1587_), .B(mai_mai_n1564_), .Y(mai19));
  NO2        m1539(.A(mai_mai_n1466_), .B(mai_mai_n262_), .Y(mai_mai_n1589_));
  NA2        m1540(.A(mai_mai_n654_), .B(x3), .Y(mai_mai_n1590_));
  OAI210     m1541(.A0(mai_mai_n156_), .A1(mai_mai_n109_), .B0(mai_mai_n81_), .Y(mai_mai_n1591_));
  NA3        m1542(.A(mai_mai_n1591_), .B(mai_mai_n1590_), .C(mai_mai_n245_), .Y(mai_mai_n1592_));
  NO2        m1543(.A(mai_mai_n1324_), .B(mai_mai_n173_), .Y(mai_mai_n1593_));
  AOI210     m1544(.A0(mai_mai_n1493_), .A1(mai_mai_n358_), .B0(mai_mai_n1593_), .Y(mai_mai_n1594_));
  AOI210     m1545(.A0(mai_mai_n1594_), .A1(mai_mai_n1592_), .B0(mai_mai_n56_), .Y(mai_mai_n1595_));
  NO2        m1546(.A(mai_mai_n868_), .B(mai_mai_n1236_), .Y(mai_mai_n1596_));
  OAI210     m1547(.A0(mai_mai_n1595_), .A1(mai_mai_n1589_), .B0(mai_mai_n1596_), .Y(mai_mai_n1597_));
  NOi21      m1548(.An(mai_mai_n616_), .B(mai_mai_n658_), .Y(mai_mai_n1598_));
  AOI210     m1549(.A0(mai_mai_n358_), .A1(x6), .B0(mai_mai_n123_), .Y(mai_mai_n1599_));
  NO3        m1550(.A(mai_mai_n1599_), .B(mai_mai_n765_), .C(mai_mai_n128_), .Y(mai_mai_n1600_));
  NA2        m1551(.A(mai_mai_n1217_), .B(mai_mai_n124_), .Y(mai_mai_n1601_));
  NO4        m1552(.A(mai_mai_n1601_), .B(mai_mai_n1010_), .C(mai_mai_n897_), .D(mai_mai_n77_), .Y(mai_mai_n1602_));
  NO3        m1553(.A(mai_mai_n1602_), .B(mai_mai_n1600_), .C(mai_mai_n1036_), .Y(mai_mai_n1603_));
  NO2        m1554(.A(mai_mai_n546_), .B(mai_mai_n625_), .Y(mai_mai_n1604_));
  NA2        m1555(.A(mai_mai_n1270_), .B(mai_mai_n50_), .Y(mai_mai_n1605_));
  NO3        m1556(.A(mai_mai_n521_), .B(mai_mai_n311_), .C(mai_mai_n64_), .Y(mai_mai_n1606_));
  AOI220     m1557(.A0(mai_mai_n1606_), .A1(mai_mai_n1605_), .B0(mai_mai_n1604_), .B1(mai_mai_n783_), .Y(mai_mai_n1607_));
  OAI210     m1558(.A0(mai_mai_n1603_), .A1(mai_mai_n57_), .B0(mai_mai_n1607_), .Y(mai_mai_n1608_));
  AOI210     m1559(.A0(mai_mai_n1608_), .A1(mai_mai_n780_), .B0(mai_mai_n1598_), .Y(mai_mai_n1609_));
  AOI210     m1560(.A0(mai_mai_n829_), .A1(mai_mai_n742_), .B0(mai_mai_n770_), .Y(mai_mai_n1610_));
  NO2        m1561(.A(mai_mai_n1610_), .B(x4), .Y(mai_mai_n1611_));
  NA3        m1562(.A(mai_mai_n740_), .B(mai_mai_n261_), .C(x7), .Y(mai_mai_n1612_));
  AOI220     m1563(.A0(mai_mai_n1418_), .A1(mai_mai_n794_), .B0(mai_mai_n707_), .B1(mai_mai_n1176_), .Y(mai_mai_n1613_));
  AOI210     m1564(.A0(mai_mai_n1613_), .A1(mai_mai_n1612_), .B0(mai_mai_n506_), .Y(mai_mai_n1614_));
  OAI210     m1565(.A0(mai_mai_n1614_), .A1(mai_mai_n1611_), .B0(mai_mai_n819_), .Y(mai_mai_n1615_));
  NO2        m1566(.A(mai_mai_n752_), .B(mai_mai_n327_), .Y(mai_mai_n1616_));
  NO2        m1567(.A(mai_mai_n156_), .B(mai_mai_n1035_), .Y(mai_mai_n1617_));
  AOI220     m1568(.A0(mai_mai_n1617_), .A1(mai_mai_n1286_), .B0(mai_mai_n1616_), .B1(mai_mai_n481_), .Y(mai_mai_n1618_));
  AO210      m1569(.A0(mai_mai_n1618_), .A1(mai_mai_n1615_), .B0(x1), .Y(mai_mai_n1619_));
  NA3        m1570(.A(mai_mai_n637_), .B(mai_mai_n1061_), .C(mai_mai_n1209_), .Y(mai_mai_n1620_));
  NA2        m1571(.A(mai_mai_n149_), .B(mai_mai_n111_), .Y(mai_mai_n1621_));
  NOi21      m1572(.An(x1), .B(x6), .Y(mai_mai_n1622_));
  NA2        m1573(.A(mai_mai_n1622_), .B(mai_mai_n84_), .Y(mai_mai_n1623_));
  NA3        m1574(.A(mai_mai_n1623_), .B(mai_mai_n1621_), .C(mai_mai_n1620_), .Y(mai_mai_n1624_));
  AOI220     m1575(.A0(mai_mai_n1624_), .A1(x3), .B0(mai_mai_n1224_), .B1(mai_mai_n385_), .Y(mai_mai_n1625_));
  NA3        m1576(.A(mai_mai_n1229_), .B(mai_mai_n804_), .C(mai_mai_n608_), .Y(mai_mai_n1626_));
  AOI220     m1577(.A0(mai_mai_n1274_), .A1(mai_mai_n123_), .B0(mai_mai_n927_), .B1(mai_mai_n821_), .Y(mai_mai_n1627_));
  AOI210     m1578(.A0(mai_mai_n1627_), .A1(mai_mai_n1626_), .B0(mai_mai_n327_), .Y(mai_mai_n1628_));
  NA2        m1579(.A(mai_mai_n949_), .B(mai_mai_n50_), .Y(mai_mai_n1629_));
  NA3        m1580(.A(mai_mai_n1217_), .B(mai_mai_n386_), .C(mai_mai_n110_), .Y(mai_mai_n1630_));
  AOI210     m1581(.A0(mai_mai_n1630_), .A1(mai_mai_n1629_), .B0(mai_mai_n973_), .Y(mai_mai_n1631_));
  NO3        m1582(.A(mai_mai_n623_), .B(mai_mai_n520_), .C(mai_mai_n1242_), .Y(mai_mai_n1632_));
  NO3        m1583(.A(mai_mai_n1632_), .B(mai_mai_n1631_), .C(mai_mai_n1628_), .Y(mai_mai_n1633_));
  OAI210     m1584(.A0(mai_mai_n1625_), .A1(mai_mai_n855_), .B0(mai_mai_n1633_), .Y(mai_mai_n1634_));
  NO2        m1585(.A(mai_mai_n559_), .B(mai_mai_n68_), .Y(mai_mai_n1635_));
  OAI220     m1586(.A0(mai_mai_n1635_), .A1(mai_mai_n1590_), .B0(mai_mai_n310_), .B1(mai_mai_n905_), .Y(mai_mai_n1636_));
  AOI220     m1587(.A0(mai_mai_n1636_), .A1(mai_mai_n56_), .B0(mai_mai_n1371_), .B1(mai_mai_n737_), .Y(mai_mai_n1637_));
  NO2        m1588(.A(mai_mai_n54_), .B(mai_mai_n71_), .Y(mai_mai_n1638_));
  AO220      m1589(.A0(mai_mai_n1638_), .A1(mai_mai_n1010_), .B0(mai_mai_n821_), .B1(mai_mai_n962_), .Y(mai_mai_n1639_));
  NA2        m1590(.A(mai_mai_n1200_), .B(mai_mai_n365_), .Y(mai_mai_n1640_));
  NO2        m1591(.A(mai_mai_n1003_), .B(mai_mai_n1622_), .Y(mai_mai_n1641_));
  NA2        m1592(.A(mai_mai_n502_), .B(mai_mai_n737_), .Y(mai_mai_n1642_));
  OAI210     m1593(.A0(mai_mai_n1642_), .A1(mai_mai_n1641_), .B0(mai_mai_n1640_), .Y(mai_mai_n1643_));
  AOI210     m1594(.A0(mai_mai_n1639_), .A1(x2), .B0(mai_mai_n1643_), .Y(mai_mai_n1644_));
  OAI220     m1595(.A0(mai_mai_n1644_), .A1(mai_mai_n156_), .B0(mai_mai_n1637_), .B1(mai_mai_n54_), .Y(mai_mai_n1645_));
  OAI210     m1596(.A0(mai_mai_n1645_), .A1(mai_mai_n1634_), .B0(x8), .Y(mai_mai_n1646_));
  NA4        m1597(.A(mai_mai_n1646_), .B(mai_mai_n1619_), .C(mai_mai_n1609_), .D(mai_mai_n1597_), .Y(mai20));
  NA2        m1598(.A(mai_mai_n481_), .B(mai_mai_n417_), .Y(mai_mai_n1648_));
  NO2        m1599(.A(mai_mai_n1648_), .B(mai_mai_n87_), .Y(mai_mai_n1649_));
  AOI210     m1600(.A0(mai_mai_n1065_), .A1(mai_mai_n62_), .B0(mai_mai_n1604_), .Y(mai_mai_n1650_));
  AOI210     m1601(.A0(mai_mai_n997_), .A1(mai_mai_n354_), .B0(mai_mai_n1207_), .Y(mai_mai_n1651_));
  OAI210     m1602(.A0(mai_mai_n1650_), .A1(mai_mai_n689_), .B0(mai_mai_n1651_), .Y(mai_mai_n1652_));
  OAI210     m1603(.A0(mai_mai_n1652_), .A1(mai_mai_n1649_), .B0(mai_mai_n1121_), .Y(mai_mai_n1653_));
  NAi21      m1604(.An(mai_mai_n555_), .B(mai_mai_n405_), .Y(mai_mai_n1654_));
  NA3        m1605(.A(mai_mai_n1654_), .B(mai_mai_n995_), .C(mai_mai_n962_), .Y(mai_mai_n1655_));
  NA3        m1606(.A(mai_mai_n1120_), .B(mai_mai_n283_), .C(mai_mai_n589_), .Y(mai_mai_n1656_));
  AOI210     m1607(.A0(mai_mai_n1656_), .A1(mai_mai_n1655_), .B0(mai_mai_n1315_), .Y(mai_mai_n1657_));
  NO2        m1608(.A(mai_mai_n756_), .B(mai_mai_n983_), .Y(mai_mai_n1658_));
  NOi31      m1609(.An(mai_mai_n1658_), .B(mai_mai_n1192_), .C(mai_mai_n533_), .Y(mai_mai_n1659_));
  OAI210     m1610(.A0(mai_mai_n1659_), .A1(mai_mai_n1657_), .B0(mai_mai_n332_), .Y(mai_mai_n1660_));
  NO4        m1611(.A(mai_mai_n550_), .B(mai_mai_n240_), .C(x5), .D(x2), .Y(mai_mai_n1661_));
  NA2        m1612(.A(mai_mai_n323_), .B(mai_mai_n93_), .Y(mai_mai_n1662_));
  NA2        m1613(.A(mai_mai_n333_), .B(mai_mai_n108_), .Y(mai_mai_n1663_));
  NA2        m1614(.A(mai_mai_n427_), .B(mai_mai_n52_), .Y(mai_mai_n1664_));
  OAI220     m1615(.A0(mai_mai_n1664_), .A1(mai_mai_n1663_), .B0(mai_mai_n1662_), .B1(mai_mai_n278_), .Y(mai_mai_n1665_));
  OAI210     m1616(.A0(mai_mai_n1665_), .A1(mai_mai_n1661_), .B0(mai_mai_n225_), .Y(mai_mai_n1666_));
  NO2        m1617(.A(mai_mai_n673_), .B(mai_mai_n612_), .Y(mai_mai_n1667_));
  NA2        m1618(.A(mai_mai_n963_), .B(mai_mai_n50_), .Y(mai_mai_n1668_));
  NO3        m1619(.A(mai_mai_n1668_), .B(mai_mai_n371_), .C(mai_mai_n233_), .Y(mai_mai_n1669_));
  NA4        m1620(.A(mai_mai_n344_), .B(mai_mai_n242_), .C(mai_mai_n809_), .D(mai_mai_n64_), .Y(mai_mai_n1670_));
  OAI220     m1621(.A0(mai_mai_n1670_), .A1(mai_mai_n683_), .B0(mai_mai_n1487_), .B1(mai_mai_n1048_), .Y(mai_mai_n1671_));
  AOI210     m1622(.A0(mai_mai_n1669_), .A1(mai_mai_n1667_), .B0(mai_mai_n1671_), .Y(mai_mai_n1672_));
  NA4        m1623(.A(mai_mai_n1672_), .B(mai_mai_n1666_), .C(mai_mai_n1660_), .D(mai_mai_n1653_), .Y(mai21));
  OAI210     m1624(.A0(mai_mai_n410_), .A1(mai_mai_n54_), .B0(x7), .Y(mai_mai_n1674_));
  OAI220     m1625(.A0(mai_mai_n1674_), .A1(mai_mai_n1304_), .B0(mai_mai_n1066_), .B1(mai_mai_n96_), .Y(mai_mai_n1675_));
  NA2        m1626(.A(mai_mai_n1675_), .B(mai_mai_n78_), .Y(mai_mai_n1676_));
  NA2        m1627(.A(mai_mai_n295_), .B(mai_mai_n866_), .Y(mai_mai_n1677_));
  AOI220     m1628(.A0(mai_mai_n1677_), .A1(mai_mai_n313_), .B0(mai_mai_n574_), .B1(mai_mai_n465_), .Y(mai_mai_n1678_));
  NA2        m1629(.A(mai_mai_n949_), .B(mai_mai_n277_), .Y(mai_mai_n1679_));
  NA2        m1630(.A(mai_mai_n541_), .B(mai_mai_n466_), .Y(mai_mai_n1680_));
  NA4        m1631(.A(mai_mai_n1680_), .B(mai_mai_n1679_), .C(mai_mai_n1398_), .D(mai_mai_n56_), .Y(mai_mai_n1681_));
  NO2        m1632(.A(mai_mai_n783_), .B(mai_mai_n438_), .Y(mai_mai_n1682_));
  NO3        m1633(.A(mai_mai_n1682_), .B(mai_mai_n729_), .C(mai_mai_n254_), .Y(mai_mai_n1683_));
  NOi31      m1634(.An(mai_mai_n196_), .B(mai_mai_n637_), .C(mai_mai_n1104_), .Y(mai_mai_n1684_));
  NO4        m1635(.A(mai_mai_n1684_), .B(mai_mai_n1683_), .C(mai_mai_n1681_), .D(mai_mai_n1678_), .Y(mai_mai_n1685_));
  NO3        m1636(.A(mai_mai_n438_), .B(mai_mai_n281_), .C(mai_mai_n52_), .Y(mai_mai_n1686_));
  OA210      m1637(.A0(mai_mai_n1686_), .A1(mai_mai_n894_), .B0(x3), .Y(mai_mai_n1687_));
  OAI210     m1638(.A0(mai_mai_n793_), .A1(mai_mai_n594_), .B0(mai_mai_n346_), .Y(mai_mai_n1688_));
  NO2        m1639(.A(mai_mai_n70_), .B(x2), .Y(mai_mai_n1689_));
  OAI210     m1640(.A0(mai_mai_n180_), .A1(x0), .B0(mai_mai_n1689_), .Y(mai_mai_n1690_));
  NA2        m1641(.A(mai_mai_n146_), .B(mai_mai_n108_), .Y(mai_mai_n1691_));
  NA3        m1642(.A(mai_mai_n1691_), .B(mai_mai_n1690_), .C(mai_mai_n1688_), .Y(mai_mai_n1692_));
  OAI210     m1643(.A0(mai_mai_n1692_), .A1(mai_mai_n1687_), .B0(x8), .Y(mai_mai_n1693_));
  NO3        m1644(.A(mai_mai_n781_), .B(mai_mai_n626_), .C(mai_mai_n590_), .Y(mai_mai_n1694_));
  NA2        m1645(.A(mai_mai_n55_), .B(mai_mai_n50_), .Y(mai_mai_n1695_));
  MUX2       m1646(.S(mai_mai_n606_), .A(mai_mai_n1695_), .B(mai_mai_n107_), .Y(mai_mai_n1696_));
  AOI210     m1647(.A0(mai_mai_n1376_), .A1(mai_mai_n243_), .B0(mai_mai_n1696_), .Y(mai_mai_n1697_));
  OAI210     m1648(.A0(mai_mai_n650_), .A1(mai_mai_n589_), .B0(x4), .Y(mai_mai_n1698_));
  NO3        m1649(.A(mai_mai_n1698_), .B(mai_mai_n1697_), .C(mai_mai_n1694_), .Y(mai_mai_n1699_));
  AO220      m1650(.A0(mai_mai_n1699_), .A1(mai_mai_n1693_), .B0(mai_mai_n1685_), .B1(mai_mai_n1676_), .Y(mai_mai_n1700_));
  AO220      m1651(.A0(mai_mai_n638_), .A1(mai_mai_n327_), .B0(mai_mai_n595_), .B1(x8), .Y(mai_mai_n1701_));
  NO2        m1652(.A(mai_mai_n868_), .B(x0), .Y(mai_mai_n1702_));
  NO3        m1653(.A(mai_mai_n1702_), .B(mai_mai_n551_), .C(mai_mai_n88_), .Y(mai_mai_n1703_));
  NO2        m1654(.A(mai_mai_n162_), .B(x2), .Y(mai_mai_n1704_));
  NO3        m1655(.A(mai_mai_n383_), .B(mai_mai_n259_), .C(mai_mai_n188_), .Y(mai_mai_n1705_));
  AOI210     m1656(.A0(mai_mai_n1704_), .A1(mai_mai_n68_), .B0(mai_mai_n1705_), .Y(mai_mai_n1706_));
  OAI210     m1657(.A0(mai_mai_n1703_), .A1(mai_mai_n403_), .B0(mai_mai_n1706_), .Y(mai_mai_n1707_));
  AOI220     m1658(.A0(mai_mai_n1707_), .A1(x5), .B0(mai_mai_n1701_), .B1(mai_mai_n756_), .Y(mai_mai_n1708_));
  AOI210     m1659(.A0(mai_mai_n1708_), .A1(mai_mai_n1700_), .B0(mai_mai_n71_), .Y(mai_mai_n1709_));
  NO2        m1660(.A(mai_mai_n917_), .B(mai_mai_n171_), .Y(mai_mai_n1710_));
  NOi41      m1661(.An(mai_mai_n1449_), .B(mai_mai_n1522_), .C(mai_mai_n1175_), .D(mai_mai_n859_), .Y(mai_mai_n1711_));
  NA2        m1662(.A(mai_mai_n1711_), .B(mai_mai_n1710_), .Y(mai_mai_n1712_));
  NO2        m1663(.A(mai_mai_n78_), .B(x4), .Y(mai_mai_n1713_));
  OAI210     m1664(.A0(mai_mai_n293_), .A1(mai_mai_n160_), .B0(mai_mai_n1713_), .Y(mai_mai_n1714_));
  OAI210     m1665(.A0(mai_mai_n412_), .A1(mai_mai_n428_), .B0(mai_mai_n233_), .Y(mai_mai_n1715_));
  NO2        m1666(.A(mai_mai_n261_), .B(mai_mai_n50_), .Y(mai_mai_n1716_));
  NO2        m1667(.A(mai_mai_n1716_), .B(mai_mai_n57_), .Y(mai_mai_n1717_));
  NA2        m1668(.A(mai_mai_n1717_), .B(mai_mai_n1715_), .Y(mai_mai_n1718_));
  AOI210     m1669(.A0(mai_mai_n1714_), .A1(mai_mai_n1712_), .B0(mai_mai_n1718_), .Y(mai_mai_n1719_));
  NA2        m1670(.A(mai_mai_n767_), .B(mai_mai_n555_), .Y(mai_mai_n1720_));
  AO210      m1671(.A0(mai_mai_n1720_), .A1(mai_mai_n973_), .B0(mai_mai_n50_), .Y(mai_mai_n1721_));
  NO2        m1672(.A(mai_mai_n1654_), .B(mai_mai_n1236_), .Y(mai_mai_n1722_));
  AOI220     m1673(.A0(mai_mai_n1722_), .A1(mai_mai_n1185_), .B0(mai_mai_n1343_), .B1(mai_mai_n1059_), .Y(mai_mai_n1723_));
  AOI210     m1674(.A0(mai_mai_n1723_), .A1(mai_mai_n1721_), .B0(mai_mai_n110_), .Y(mai_mai_n1724_));
  NA2        m1675(.A(mai_mai_n302_), .B(mai_mai_n108_), .Y(mai_mai_n1725_));
  NA2        m1676(.A(mai_mai_n904_), .B(mai_mai_n55_), .Y(mai_mai_n1726_));
  NO2        m1677(.A(mai_mai_n1726_), .B(mai_mai_n1725_), .Y(mai_mai_n1727_));
  NO2        m1678(.A(mai_mai_n678_), .B(mai_mai_n1069_), .Y(mai_mai_n1728_));
  NO4        m1679(.A(mai_mai_n1728_), .B(mai_mai_n1727_), .C(mai_mai_n1724_), .D(mai_mai_n1719_), .Y(mai_mai_n1729_));
  NO2        m1680(.A(mai_mai_n1729_), .B(x6), .Y(mai_mai_n1730_));
  AOI210     m1681(.A0(mai_mai_n615_), .A1(mai_mai_n1069_), .B0(mai_mai_n1522_), .Y(mai_mai_n1731_));
  OAI210     m1682(.A0(mai_mai_n1731_), .A1(mai_mai_n696_), .B0(mai_mai_n56_), .Y(mai_mai_n1732_));
  NO2        m1683(.A(mai_mai_n758_), .B(mai_mai_n54_), .Y(mai_mai_n1733_));
  NO4        m1684(.A(mai_mai_n971_), .B(mai_mai_n281_), .C(mai_mai_n780_), .D(mai_mai_n765_), .Y(mai_mai_n1734_));
  NO2        m1685(.A(mai_mai_n873_), .B(x5), .Y(mai_mai_n1735_));
  NO4        m1686(.A(mai_mai_n1735_), .B(mai_mai_n1734_), .C(mai_mai_n1733_), .D(mai_mai_n956_), .Y(mai_mai_n1736_));
  AOI210     m1687(.A0(mai_mai_n1736_), .A1(mai_mai_n1732_), .B0(mai_mai_n50_), .Y(mai_mai_n1737_));
  NA2        m1688(.A(mai_mai_n162_), .B(mai_mai_n108_), .Y(mai_mai_n1738_));
  OA220      m1689(.A0(mai_mai_n1738_), .A1(mai_mai_n442_), .B0(mai_mai_n471_), .B1(mai_mai_n756_), .Y(mai_mai_n1739_));
  NA3        m1690(.A(mai_mai_n55_), .B(x2), .C(x0), .Y(mai_mai_n1740_));
  AOI220     m1691(.A0(mai_mai_n1740_), .A1(mai_mai_n173_), .B0(mai_mai_n873_), .B1(mai_mai_n158_), .Y(mai_mai_n1741_));
  NO2        m1692(.A(mai_mai_n689_), .B(mai_mai_n261_), .Y(mai_mai_n1742_));
  NO3        m1693(.A(mai_mai_n249_), .B(mai_mai_n231_), .C(mai_mai_n365_), .Y(mai_mai_n1743_));
  NO3        m1694(.A(mai_mai_n1743_), .B(mai_mai_n1742_), .C(mai_mai_n1741_), .Y(mai_mai_n1744_));
  OAI220     m1695(.A0(mai_mai_n1744_), .A1(mai_mai_n56_), .B0(mai_mai_n1739_), .B1(mai_mai_n705_), .Y(mai_mai_n1745_));
  OAI210     m1696(.A0(mai_mai_n1745_), .A1(mai_mai_n1737_), .B0(mai_mai_n116_), .Y(mai_mai_n1746_));
  NO2        m1697(.A(mai_mai_n620_), .B(mai_mai_n308_), .Y(mai_mai_n1747_));
  AOI210     m1698(.A0(mai_mai_n613_), .A1(x5), .B0(mai_mai_n1747_), .Y(mai_mai_n1748_));
  NO2        m1699(.A(mai_mai_n1748_), .B(mai_mai_n110_), .Y(mai_mai_n1749_));
  NA2        m1700(.A(mai_mai_n713_), .B(mai_mai_n81_), .Y(mai_mai_n1750_));
  NA3        m1701(.A(mai_mai_n1750_), .B(mai_mai_n435_), .C(mai_mai_n57_), .Y(mai_mai_n1751_));
  OAI210     m1702(.A0(mai_mai_n1726_), .A1(mai_mai_n1725_), .B0(mai_mai_n1751_), .Y(mai_mai_n1752_));
  OAI210     m1703(.A0(mai_mai_n1752_), .A1(mai_mai_n1749_), .B0(x1), .Y(mai_mai_n1753_));
  NO4        m1704(.A(mai_mai_n421_), .B(mai_mai_n78_), .C(mai_mai_n150_), .D(x3), .Y(mai_mai_n1754_));
  NO2        m1705(.A(mai_mai_n333_), .B(mai_mai_n112_), .Y(mai_mai_n1755_));
  OAI210     m1706(.A0(mai_mai_n1754_), .A1(mai_mai_n1316_), .B0(mai_mai_n1755_), .Y(mai_mai_n1756_));
  NO2        m1707(.A(mai_mai_n60_), .B(mai_mai_n108_), .Y(mai_mai_n1757_));
  NO4        m1708(.A(mai_mai_n1725_), .B(mai_mai_n971_), .C(mai_mai_n673_), .D(mai_mai_n50_), .Y(mai_mai_n1758_));
  AOI210     m1709(.A0(mai_mai_n1757_), .A1(mai_mai_n1566_), .B0(mai_mai_n1758_), .Y(mai_mai_n1759_));
  NA4        m1710(.A(mai_mai_n1759_), .B(mai_mai_n1756_), .C(mai_mai_n1753_), .D(mai_mai_n1746_), .Y(mai_mai_n1760_));
  NO3        m1711(.A(mai_mai_n1760_), .B(mai_mai_n1730_), .C(mai_mai_n1709_), .Y(mai22));
  AOI210     m1712(.A0(mai_mai_n527_), .A1(mai_mai_n71_), .B0(mai_mai_n474_), .Y(mai_mai_n1762_));
  NO3        m1713(.A(mai_mai_n1212_), .B(mai_mai_n559_), .C(mai_mai_n707_), .Y(mai_mai_n1763_));
  AOI210     m1714(.A0(x5), .A1(x2), .B0(x8), .Y(mai_mai_n1764_));
  NA2        m1715(.A(mai_mai_n1764_), .B(mai_mai_n59_), .Y(mai_mai_n1765_));
  OAI220     m1716(.A0(mai_mai_n1765_), .A1(mai_mai_n1763_), .B0(mai_mai_n1762_), .B1(mai_mai_n403_), .Y(mai_mai_n1766_));
  NA2        m1717(.A(mai_mai_n589_), .B(mai_mai_n87_), .Y(mai_mai_n1767_));
  NA2        m1718(.A(mai_mai_n278_), .B(mai_mai_n77_), .Y(mai_mai_n1768_));
  OA220      m1719(.A0(mai_mai_n1768_), .A1(mai_mai_n1767_), .B0(mai_mai_n852_), .B1(mai_mai_n1020_), .Y(mai_mai_n1769_));
  NO4        m1720(.A(mai_mai_n389_), .B(mai_mai_n223_), .C(mai_mai_n71_), .D(x3), .Y(mai_mai_n1770_));
  NO3        m1721(.A(mai_mai_n1265_), .B(mai_mai_n87_), .C(x0), .Y(mai_mai_n1771_));
  OAI210     m1722(.A0(mai_mai_n403_), .A1(mai_mai_n208_), .B0(x4), .Y(mai_mai_n1772_));
  NO2        m1723(.A(mai_mai_n1772_), .B(mai_mai_n1770_), .Y(mai_mai_n1773_));
  OAI210     m1724(.A0(mai_mai_n1769_), .A1(mai_mai_n201_), .B0(mai_mai_n1773_), .Y(mai_mai_n1774_));
  AOI210     m1725(.A0(mai_mai_n1766_), .A1(mai_mai_n53_), .B0(mai_mai_n1774_), .Y(mai_mai_n1775_));
  NA2        m1726(.A(mai_mai_n306_), .B(mai_mai_n311_), .Y(mai_mai_n1776_));
  NA3        m1727(.A(mai_mai_n1776_), .B(mai_mai_n225_), .C(mai_mai_n310_), .Y(mai_mai_n1777_));
  NA2        m1728(.A(mai_mai_n584_), .B(mai_mai_n248_), .Y(mai_mai_n1778_));
  NO3        m1729(.A(mai_mai_n502_), .B(mai_mai_n269_), .C(mai_mai_n217_), .Y(mai_mai_n1779_));
  NAi31      m1730(.An(mai_mai_n1779_), .B(mai_mai_n1778_), .C(mai_mai_n1777_), .Y(mai_mai_n1780_));
  NO2        m1731(.A(mai_mai_n471_), .B(mai_mai_n263_), .Y(mai_mai_n1781_));
  NO2        m1732(.A(mai_mai_n1265_), .B(x3), .Y(mai_mai_n1782_));
  AOI210     m1733(.A0(mai_mai_n1782_), .A1(mai_mai_n354_), .B0(mai_mai_n1781_), .Y(mai_mai_n1783_));
  OAI210     m1734(.A0(mai_mai_n1099_), .A1(mai_mai_n190_), .B0(mai_mai_n56_), .Y(mai_mai_n1784_));
  NA3        m1735(.A(mai_mai_n55_), .B(mai_mai_n71_), .C(x0), .Y(mai_mai_n1785_));
  OAI220     m1736(.A0(mai_mai_n1785_), .A1(mai_mai_n1069_), .B0(mai_mai_n371_), .B1(mai_mai_n216_), .Y(mai_mai_n1786_));
  NO2        m1737(.A(mai_mai_n1786_), .B(mai_mai_n1784_), .Y(mai_mai_n1787_));
  OAI210     m1738(.A0(mai_mai_n1783_), .A1(mai_mai_n261_), .B0(mai_mai_n1787_), .Y(mai_mai_n1788_));
  AOI210     m1739(.A0(mai_mai_n1780_), .A1(mai_mai_n108_), .B0(mai_mai_n1788_), .Y(mai_mai_n1789_));
  AOI210     m1740(.A0(mai_mai_n960_), .A1(mai_mai_n782_), .B0(mai_mai_n877_), .Y(mai_mai_n1790_));
  OAI210     m1741(.A0(mai_mai_n811_), .A1(mai_mai_n162_), .B0(mai_mai_n946_), .Y(mai_mai_n1791_));
  OAI210     m1742(.A0(mai_mai_n1791_), .A1(mai_mai_n1790_), .B0(mai_mai_n619_), .Y(mai_mai_n1792_));
  OA210      m1743(.A0(mai_mai_n1789_), .A1(mai_mai_n1775_), .B0(mai_mai_n1792_), .Y(mai_mai_n1793_));
  OAI210     m1744(.A0(mai_mai_n1194_), .A1(mai_mai_n712_), .B0(mai_mai_n700_), .Y(mai_mai_n1794_));
  NO2        m1745(.A(mai_mai_n359_), .B(x0), .Y(mai_mai_n1795_));
  NA3        m1746(.A(mai_mai_n1795_), .B(mai_mai_n354_), .C(mai_mai_n56_), .Y(mai_mai_n1796_));
  AOI210     m1747(.A0(mai_mai_n1796_), .A1(mai_mai_n1794_), .B0(mai_mai_n403_), .Y(mai_mai_n1797_));
  NO3        m1748(.A(mai_mai_n173_), .B(mai_mai_n162_), .C(mai_mai_n62_), .Y(mai_mai_n1798_));
  OAI210     m1749(.A0(mai_mai_n1798_), .A1(mai_mai_n423_), .B0(mai_mai_n110_), .Y(mai_mai_n1799_));
  NA2        m1750(.A(mai_mai_n143_), .B(mai_mai_n794_), .Y(mai_mai_n1800_));
  NA2        m1751(.A(mai_mai_n421_), .B(x3), .Y(mai_mai_n1801_));
  NAi31      m1752(.An(mai_mai_n1801_), .B(mai_mai_n1800_), .C(mai_mai_n1582_), .Y(mai_mai_n1802_));
  NO3        m1753(.A(mai_mai_n868_), .B(mai_mai_n470_), .C(mai_mai_n110_), .Y(mai_mai_n1803_));
  NO2        m1754(.A(mai_mai_n1101_), .B(mai_mai_n144_), .Y(mai_mai_n1804_));
  NO3        m1755(.A(mai_mai_n907_), .B(mai_mai_n417_), .C(mai_mai_n307_), .Y(mai_mai_n1805_));
  AOI220     m1756(.A0(mai_mai_n1805_), .A1(mai_mai_n1804_), .B0(mai_mai_n1803_), .B1(mai_mai_n1795_), .Y(mai_mai_n1806_));
  NA3        m1757(.A(mai_mai_n417_), .B(mai_mai_n93_), .C(mai_mai_n81_), .Y(mai_mai_n1807_));
  AOI210     m1758(.A0(mai_mai_n615_), .A1(mai_mai_n460_), .B0(mai_mai_n500_), .Y(mai_mai_n1808_));
  NA2        m1759(.A(mai_mai_n1196_), .B(x3), .Y(mai_mai_n1809_));
  OAI210     m1760(.A0(mai_mai_n1809_), .A1(mai_mai_n1808_), .B0(mai_mai_n1807_), .Y(mai_mai_n1810_));
  NA3        m1761(.A(mai_mai_n56_), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n1811_));
  NOi21      m1762(.An(mai_mai_n83_), .B(mai_mai_n740_), .Y(mai_mai_n1812_));
  NA3        m1763(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n1813_));
  NA3        m1764(.A(mai_mai_n1813_), .B(mai_mai_n1003_), .C(mai_mai_n270_), .Y(mai_mai_n1814_));
  OAI220     m1765(.A0(mai_mai_n1814_), .A1(mai_mai_n1812_), .B0(mai_mai_n1072_), .B1(mai_mai_n1811_), .Y(mai_mai_n1815_));
  AOI220     m1766(.A0(mai_mai_n1815_), .A1(mai_mai_n1083_), .B0(mai_mai_n1810_), .B1(mai_mai_n354_), .Y(mai_mai_n1816_));
  NA4        m1767(.A(mai_mai_n1816_), .B(mai_mai_n1806_), .C(mai_mai_n1802_), .D(mai_mai_n1799_), .Y(mai_mai_n1817_));
  AOI210     m1768(.A0(mai_mai_n1817_), .A1(x7), .B0(mai_mai_n1797_), .Y(mai_mai_n1818_));
  OAI210     m1769(.A0(mai_mai_n1793_), .A1(x7), .B0(mai_mai_n1818_), .Y(mai23));
  OR2        m1770(.A(mai_mai_n521_), .B(mai_mai_n225_), .Y(mai_mai_n1820_));
  AOI220     m1771(.A0(mai_mai_n1820_), .A1(mai_mai_n1658_), .B0(mai_mai_n621_), .B1(mai_mai_n298_), .Y(mai_mai_n1821_));
  NO3        m1772(.A(mai_mai_n852_), .B(mai_mai_n598_), .C(mai_mai_n493_), .Y(mai_mai_n1822_));
  NO3        m1773(.A(mai_mai_n964_), .B(mai_mai_n151_), .C(mai_mai_n117_), .Y(mai_mai_n1823_));
  AOI210     m1774(.A0(mai_mai_n1823_), .A1(mai_mai_n1042_), .B0(mai_mai_n1822_), .Y(mai_mai_n1824_));
  OAI210     m1775(.A0(mai_mai_n1821_), .A1(mai_mai_n156_), .B0(mai_mai_n1824_), .Y(mai_mai_n1825_));
  NA2        m1776(.A(mai_mai_n1825_), .B(mai_mai_n55_), .Y(mai_mai_n1826_));
  NO2        m1777(.A(mai_mai_n971_), .B(mai_mai_n519_), .Y(mai_mai_n1827_));
  AO220      m1778(.A0(mai_mai_n1300_), .A1(mai_mai_n184_), .B0(mai_mai_n1010_), .B1(mai_mai_n756_), .Y(mai_mai_n1828_));
  OAI210     m1779(.A0(mai_mai_n1828_), .A1(mai_mai_n1827_), .B0(mai_mai_n595_), .Y(mai_mai_n1829_));
  NA2        m1780(.A(mai_mai_n181_), .B(mai_mai_n171_), .Y(mai_mai_n1830_));
  NA2        m1781(.A(mai_mai_n409_), .B(mai_mai_n163_), .Y(mai_mai_n1831_));
  AOI210     m1782(.A0(mai_mai_n1831_), .A1(mai_mai_n1830_), .B0(mai_mai_n240_), .Y(mai_mai_n1832_));
  NA3        m1783(.A(mai_mai_n877_), .B(mai_mai_n428_), .C(mai_mai_n261_), .Y(mai_mai_n1833_));
  AOI210     m1784(.A0(mai_mai_n1833_), .A1(mai_mai_n504_), .B0(mai_mai_n386_), .Y(mai_mai_n1834_));
  OAI210     m1785(.A0(mai_mai_n1834_), .A1(mai_mai_n1832_), .B0(mai_mai_n302_), .Y(mai_mai_n1835_));
  NA3        m1786(.A(mai_mai_n57_), .B(x4), .C(x3), .Y(mai_mai_n1836_));
  NO3        m1787(.A(mai_mai_n1836_), .B(mai_mai_n753_), .C(mai_mai_n143_), .Y(mai_mai_n1837_));
  INV        m1788(.A(mai_mai_n1837_), .Y(mai_mai_n1838_));
  NA4        m1789(.A(mai_mai_n1838_), .B(mai_mai_n1835_), .C(mai_mai_n1829_), .D(mai_mai_n1826_), .Y(mai24));
  NO2        m1790(.A(mai_mai_n245_), .B(x1), .Y(mai_mai_n1840_));
  NA2        m1791(.A(mai_mai_n344_), .B(mai_mai_n497_), .Y(mai_mai_n1841_));
  NO3        m1792(.A(mai_mai_n546_), .B(mai_mai_n692_), .C(mai_mai_n158_), .Y(mai_mai_n1842_));
  AOI210     m1793(.A0(mai_mai_n1840_), .A1(mai_mai_n93_), .B0(mai_mai_n1842_), .Y(mai_mai_n1843_));
  NA2        m1794(.A(mai_mai_n102_), .B(x8), .Y(mai_mai_n1844_));
  NO3        m1795(.A(mai_mai_n1080_), .B(mai_mai_n1357_), .C(mai_mai_n1061_), .Y(mai_mai_n1845_));
  AOI210     m1796(.A0(mai_mai_n995_), .A1(mai_mai_n56_), .B0(mai_mai_n1473_), .Y(mai_mai_n1846_));
  AO220      m1797(.A0(mai_mai_n1846_), .A1(mai_mai_n1845_), .B0(mai_mai_n1288_), .B1(mai_mai_n332_), .Y(mai_mai_n1847_));
  NA2        m1798(.A(mai_mai_n460_), .B(x8), .Y(mai_mai_n1848_));
  NA2        m1799(.A(mai_mai_n674_), .B(mai_mai_n126_), .Y(mai_mai_n1849_));
  OAI220     m1800(.A0(mai_mai_n1849_), .A1(mai_mai_n1458_), .B0(mai_mai_n1848_), .B1(mai_mai_n850_), .Y(mai_mai_n1850_));
  AOI220     m1801(.A0(mai_mai_n1850_), .A1(mai_mai_n1716_), .B0(mai_mai_n1847_), .B1(mai_mai_n1042_), .Y(mai_mai_n1851_));
  OAI210     m1802(.A0(mai_mai_n1844_), .A1(mai_mai_n1843_), .B0(mai_mai_n1851_), .Y(mai25));
  NA2        m1803(.A(mai_mai_n333_), .B(mai_mai_n59_), .Y(mai_mai_n1853_));
  NO2        m1804(.A(mai_mai_n1853_), .B(mai_mai_n324_), .Y(mai_mai_n1854_));
  OAI210     m1805(.A0(mai_mai_n1854_), .A1(mai_mai_n1201_), .B0(mai_mai_n116_), .Y(mai_mai_n1855_));
  INV        m1806(.A(mai_mai_n1295_), .Y(mai_mai_n1856_));
  NO2        m1807(.A(mai_mai_n752_), .B(mai_mai_n55_), .Y(mai_mai_n1857_));
  AOI220     m1808(.A0(mai_mai_n1857_), .A1(mai_mai_n1856_), .B0(mai_mai_n1616_), .B1(mai_mai_n1202_), .Y(mai_mai_n1858_));
  AOI210     m1809(.A0(mai_mai_n1858_), .A1(mai_mai_n1855_), .B0(mai_mai_n687_), .Y(mai_mai_n1859_));
  NO3        m1810(.A(mai_mai_n1054_), .B(mai_mai_n145_), .C(mai_mai_n78_), .Y(mai_mai_n1860_));
  OAI210     m1811(.A0(mai_mai_n201_), .A1(mai_mai_n278_), .B0(mai_mai_n334_), .Y(mai_mai_n1861_));
  OAI210     m1812(.A0(mai_mai_n1861_), .A1(mai_mai_n1860_), .B0(mai_mai_n1200_), .Y(mai_mai_n1862_));
  NO2        m1813(.A(mai_mai_n1410_), .B(mai_mai_n453_), .Y(mai_mai_n1863_));
  NO3        m1814(.A(mai_mai_n1863_), .B(mai_mai_n537_), .C(mai_mai_n99_), .Y(mai_mai_n1864_));
  NA2        m1815(.A(mai_mai_n514_), .B(mai_mai_n55_), .Y(mai_mai_n1865_));
  NO2        m1816(.A(mai_mai_n1865_), .B(mai_mai_n245_), .Y(mai_mai_n1866_));
  OAI210     m1817(.A0(mai_mai_n1866_), .A1(mai_mai_n1864_), .B0(mai_mai_n642_), .Y(mai_mai_n1867_));
  NA2        m1818(.A(mai_mai_n1781_), .B(mai_mai_n1154_), .Y(mai_mai_n1868_));
  NA3        m1819(.A(mai_mai_n1868_), .B(mai_mai_n1867_), .C(mai_mai_n1862_), .Y(mai_mai_n1869_));
  AO210      m1820(.A0(mai_mai_n1869_), .A1(mai_mai_n108_), .B0(mai_mai_n1859_), .Y(mai26));
  NA2        m1821(.A(mai_mai_n780_), .B(mai_mai_n50_), .Y(mai_mai_n1871_));
  OAI220     m1822(.A0(mai_mai_n308_), .A1(mai_mai_n254_), .B0(mai_mai_n1871_), .B1(x7), .Y(mai_mai_n1872_));
  AOI220     m1823(.A0(mai_mai_n1872_), .A1(mai_mai_n93_), .B0(mai_mai_n1316_), .B1(mai_mai_n1160_), .Y(mai_mai_n1873_));
  NA2        m1824(.A(mai_mai_n630_), .B(mai_mai_n584_), .Y(mai_mai_n1874_));
  OAI210     m1825(.A0(mai_mai_n638_), .A1(mai_mai_n630_), .B0(mai_mai_n756_), .Y(mai_mai_n1875_));
  AOI210     m1826(.A0(mai_mai_n1874_), .A1(mai_mai_n1223_), .B0(mai_mai_n1875_), .Y(mai_mai_n1876_));
  NA2        m1827(.A(mai_mai_n1033_), .B(mai_mai_n590_), .Y(mai_mai_n1877_));
  NA2        m1828(.A(mai_mai_n1804_), .B(mai_mai_n1481_), .Y(mai_mai_n1878_));
  NO2        m1829(.A(mai_mai_n1101_), .B(mai_mai_n75_), .Y(mai_mai_n1879_));
  NA2        m1830(.A(mai_mai_n819_), .B(mai_mai_n180_), .Y(mai_mai_n1880_));
  NO2        m1831(.A(mai_mai_n1880_), .B(mai_mai_n542_), .Y(mai_mai_n1881_));
  AOI210     m1832(.A0(mai_mai_n1879_), .A1(mai_mai_n591_), .B0(mai_mai_n1881_), .Y(mai_mai_n1882_));
  OAI220     m1833(.A0(mai_mai_n1882_), .A1(mai_mai_n108_), .B0(mai_mai_n1878_), .B1(mai_mai_n53_), .Y(mai_mai_n1883_));
  NA2        m1834(.A(mai_mai_n607_), .B(mai_mai_n514_), .Y(mai_mai_n1884_));
  NO2        m1835(.A(mai_mai_n136_), .B(mai_mai_n133_), .Y(mai_mai_n1885_));
  NA2        m1836(.A(mai_mai_n1885_), .B(mai_mai_n123_), .Y(mai_mai_n1886_));
  NA2        m1837(.A(mai_mai_n756_), .B(x3), .Y(mai_mai_n1887_));
  AOI210     m1838(.A0(mai_mai_n1886_), .A1(mai_mai_n1884_), .B0(mai_mai_n1887_), .Y(mai_mai_n1888_));
  NO2        m1839(.A(mai_mai_n1020_), .B(x3), .Y(mai_mai_n1889_));
  AOI210     m1840(.A0(mai_mai_n451_), .A1(mai_mai_n108_), .B0(mai_mai_n1889_), .Y(mai_mai_n1890_));
  NA3        m1841(.A(mai_mai_n575_), .B(mai_mai_n51_), .C(mai_mai_n56_), .Y(mai_mai_n1891_));
  AOI210     m1842(.A0(mai_mai_n1667_), .A1(mai_mai_n1073_), .B0(x0), .Y(mai_mai_n1892_));
  OAI210     m1843(.A0(mai_mai_n1891_), .A1(mai_mai_n1890_), .B0(mai_mai_n1892_), .Y(mai_mai_n1893_));
  NO4        m1844(.A(mai_mai_n1893_), .B(mai_mai_n1888_), .C(mai_mai_n1883_), .D(mai_mai_n1876_), .Y(mai_mai_n1894_));
  AOI210     m1845(.A0(x8), .A1(x6), .B0(x5), .Y(mai_mai_n1895_));
  AO220      m1846(.A0(mai_mai_n1895_), .A1(mai_mai_n147_), .B0(mai_mai_n598_), .B1(mai_mai_n143_), .Y(mai_mai_n1896_));
  NA2        m1847(.A(mai_mai_n1896_), .B(mai_mai_n452_), .Y(mai_mai_n1897_));
  NO2        m1848(.A(mai_mai_n766_), .B(mai_mai_n147_), .Y(mai_mai_n1898_));
  NA3        m1849(.A(mai_mai_n1898_), .B(mai_mai_n1689_), .C(mai_mai_n137_), .Y(mai_mai_n1899_));
  NO2        m1850(.A(mai_mai_n403_), .B(mai_mai_n1396_), .Y(mai_mai_n1900_));
  OAI210     m1851(.A0(mai_mai_n1900_), .A1(mai_mai_n1363_), .B0(mai_mai_n451_), .Y(mai_mai_n1901_));
  NA3        m1852(.A(mai_mai_n1901_), .B(mai_mai_n1899_), .C(mai_mai_n1897_), .Y(mai_mai_n1902_));
  NO2        m1853(.A(mai_mai_n2696_), .B(mai_mai_n117_), .Y(mai_mai_n1903_));
  NA3        m1854(.A(mai_mai_n821_), .B(mai_mai_n1020_), .C(x7), .Y(mai_mai_n1904_));
  AOI210     m1855(.A0(mai_mai_n348_), .A1(mai_mai_n219_), .B0(mai_mai_n1904_), .Y(mai_mai_n1905_));
  OAI220     m1856(.A0(mai_mai_n910_), .A1(mai_mai_n308_), .B0(mai_mai_n650_), .B1(mai_mai_n692_), .Y(mai_mai_n1906_));
  NO3        m1857(.A(mai_mai_n1906_), .B(mai_mai_n1905_), .C(mai_mai_n1903_), .Y(mai_mai_n1907_));
  NA3        m1858(.A(mai_mai_n674_), .B(mai_mai_n195_), .C(mai_mai_n962_), .Y(mai_mai_n1908_));
  NA2        m1859(.A(mai_mai_n1908_), .B(mai_mai_n650_), .Y(mai_mai_n1909_));
  NA2        m1860(.A(mai_mai_n143_), .B(mai_mai_n135_), .Y(mai_mai_n1910_));
  OAI210     m1861(.A0(mai_mai_n1910_), .A1(mai_mai_n1444_), .B0(x0), .Y(mai_mai_n1911_));
  AOI210     m1862(.A0(mai_mai_n1909_), .A1(mai_mai_n1434_), .B0(mai_mai_n1911_), .Y(mai_mai_n1912_));
  OAI210     m1863(.A0(mai_mai_n1907_), .A1(mai_mai_n53_), .B0(mai_mai_n1912_), .Y(mai_mai_n1913_));
  AOI210     m1864(.A0(mai_mai_n1902_), .A1(x4), .B0(mai_mai_n1913_), .Y(mai_mai_n1914_));
  OA220      m1865(.A0(mai_mai_n1914_), .A1(mai_mai_n1894_), .B0(mai_mai_n1873_), .B1(mai_mai_n109_), .Y(mai27));
  NA2        m1866(.A(mai_mai_n1164_), .B(mai_mai_n451_), .Y(mai_mai_n1916_));
  NO2        m1867(.A(mai_mai_n1916_), .B(mai_mai_n303_), .Y(mai_mai_n1917_));
  NA2        m1868(.A(mai_mai_n927_), .B(mai_mai_n821_), .Y(mai_mai_n1918_));
  NA3        m1869(.A(mai_mai_n827_), .B(mai_mai_n368_), .C(mai_mai_n1035_), .Y(mai_mai_n1919_));
  AOI210     m1870(.A0(mai_mai_n1919_), .A1(mai_mai_n1918_), .B0(mai_mai_n219_), .Y(mai_mai_n1920_));
  OAI210     m1871(.A0(mai_mai_n1920_), .A1(mai_mai_n1917_), .B0(mai_mai_n708_), .Y(mai_mai_n1921_));
  XO2        m1872(.A(x8), .B(x4), .Y(mai_mai_n1922_));
  NO3        m1873(.A(mai_mai_n1922_), .B(mai_mai_n451_), .C(mai_mai_n173_), .Y(mai_mai_n1923_));
  OA210      m1874(.A0(mai_mai_n1923_), .A1(mai_mai_n1271_), .B0(mai_mai_n281_), .Y(mai_mai_n1924_));
  NO2        m1875(.A(mai_mai_n398_), .B(mai_mai_n167_), .Y(mai_mai_n1925_));
  OAI210     m1876(.A0(mai_mai_n1925_), .A1(mai_mai_n1924_), .B0(mai_mai_n1138_), .Y(mai_mai_n1926_));
  AOI210     m1877(.A0(mai_mai_n638_), .A1(mai_mai_n56_), .B0(mai_mai_n1879_), .Y(mai_mai_n1927_));
  OAI220     m1878(.A0(mai_mai_n1927_), .A1(mai_mai_n1270_), .B0(mai_mai_n1222_), .B1(mai_mai_n210_), .Y(mai_mai_n1928_));
  NO2        m1879(.A(mai_mai_n705_), .B(mai_mai_n145_), .Y(mai_mai_n1929_));
  NO2        m1880(.A(mai_mai_n1206_), .B(mai_mai_n261_), .Y(mai_mai_n1930_));
  AOI220     m1881(.A0(mai_mai_n1930_), .A1(mai_mai_n1929_), .B0(mai_mai_n1928_), .B1(mai_mai_n541_), .Y(mai_mai_n1931_));
  NA3        m1882(.A(mai_mai_n1931_), .B(mai_mai_n1926_), .C(mai_mai_n1921_), .Y(mai28));
  NO3        m1883(.A(mai_mai_n1922_), .B(mai_mai_n1405_), .C(mai_mai_n149_), .Y(mai_mai_n1933_));
  OAI210     m1884(.A0(mai_mai_n1933_), .A1(mai_mai_n1290_), .B0(mai_mai_n590_), .Y(mai_mai_n1934_));
  NA3        m1885(.A(mai_mai_n1202_), .B(mai_mai_n904_), .C(x7), .Y(mai_mai_n1935_));
  NA3        m1886(.A(mai_mai_n500_), .B(mai_mai_n78_), .C(mai_mai_n612_), .Y(mai_mai_n1936_));
  NA3        m1887(.A(mai_mai_n1936_), .B(mai_mai_n1935_), .C(mai_mai_n1934_), .Y(mai_mai_n1937_));
  NA2        m1888(.A(mai_mai_n1265_), .B(mai_mai_n449_), .Y(mai_mai_n1938_));
  NA3        m1889(.A(mai_mai_n1938_), .B(mai_mai_n1423_), .C(mai_mai_n416_), .Y(mai_mai_n1939_));
  NO2        m1890(.A(mai_mai_n311_), .B(x4), .Y(mai_mai_n1940_));
  AOI220     m1891(.A0(mai_mai_n1940_), .A1(mai_mai_n1889_), .B0(mai_mai_n1139_), .B1(mai_mai_n682_), .Y(mai_mai_n1941_));
  NA2        m1892(.A(mai_mai_n1941_), .B(mai_mai_n1939_), .Y(mai_mai_n1942_));
  NO2        m1893(.A(mai_mai_n1265_), .B(mai_mai_n1242_), .Y(mai_mai_n1943_));
  NO4        m1894(.A(x6), .B(mai_mai_n56_), .C(x2), .D(x0), .Y(mai_mai_n1944_));
  OAI210     m1895(.A0(mai_mai_n1944_), .A1(mai_mai_n1943_), .B0(mai_mai_n1059_), .Y(mai_mai_n1945_));
  NA2        m1896(.A(mai_mai_n1196_), .B(mai_mai_n108_), .Y(mai_mai_n1946_));
  NA2        m1897(.A(mai_mai_n1097_), .B(mai_mai_n107_), .Y(mai_mai_n1947_));
  OAI210     m1898(.A0(mai_mai_n1947_), .A1(mai_mai_n1946_), .B0(mai_mai_n1945_), .Y(mai_mai_n1948_));
  OAI210     m1899(.A0(mai_mai_n1948_), .A1(mai_mai_n1942_), .B0(x7), .Y(mai_mai_n1949_));
  NO2        m1900(.A(mai_mai_n389_), .B(x7), .Y(mai_mai_n1950_));
  NO3        m1901(.A(mai_mai_n403_), .B(mai_mai_n275_), .C(mai_mai_n124_), .Y(mai_mai_n1951_));
  OAI210     m1902(.A0(mai_mai_n877_), .A1(mai_mai_n263_), .B0(mai_mai_n81_), .Y(mai_mai_n1952_));
  OAI220     m1903(.A0(mai_mai_n1952_), .A1(mai_mai_n1951_), .B0(mai_mai_n1950_), .B1(mai_mai_n111_), .Y(mai_mai_n1953_));
  NA2        m1904(.A(mai_mai_n1813_), .B(mai_mai_n662_), .Y(mai_mai_n1954_));
  NO2        m1905(.A(mai_mai_n1865_), .B(mai_mai_n77_), .Y(mai_mai_n1955_));
  AOI220     m1906(.A0(mai_mai_n1955_), .A1(mai_mai_n1954_), .B0(mai_mai_n482_), .B1(mai_mai_n50_), .Y(mai_mai_n1956_));
  AOI210     m1907(.A0(mai_mai_n1956_), .A1(mai_mai_n1953_), .B0(mai_mai_n59_), .Y(mai_mai_n1957_));
  AOI220     m1908(.A0(mai_mai_n1410_), .A1(mai_mai_n680_), .B0(mai_mai_n415_), .B1(mai_mai_n460_), .Y(mai_mai_n1958_));
  OAI210     m1909(.A0(mai_mai_n1958_), .A1(mai_mai_n145_), .B0(x1), .Y(mai_mai_n1959_));
  NO2        m1910(.A(mai_mai_n1959_), .B(mai_mai_n1957_), .Y(mai_mai_n1960_));
  AOI210     m1911(.A0(mai_mai_n1601_), .A1(mai_mai_n403_), .B0(mai_mai_n672_), .Y(mai_mai_n1961_));
  NO2        m1912(.A(mai_mai_n403_), .B(x5), .Y(mai_mai_n1962_));
  NO2        m1913(.A(mai_mai_n1962_), .B(mai_mai_n231_), .Y(mai_mai_n1963_));
  NO2        m1914(.A(mai_mai_n1963_), .B(mai_mai_n1961_), .Y(mai_mai_n1964_));
  NOi21      m1915(.An(mai_mai_n713_), .B(mai_mai_n1010_), .Y(mai_mai_n1965_));
  NA3        m1916(.A(mai_mai_n1965_), .B(mai_mai_n1097_), .C(mai_mai_n877_), .Y(mai_mai_n1966_));
  OAI210     m1917(.A0(mai_mai_n1377_), .A1(mai_mai_n1695_), .B0(mai_mai_n1966_), .Y(mai_mai_n1967_));
  OAI210     m1918(.A0(mai_mai_n1967_), .A1(mai_mai_n1964_), .B0(mai_mai_n1138_), .Y(mai_mai_n1968_));
  OAI210     m1919(.A0(mai_mai_n449_), .A1(mai_mai_n51_), .B0(mai_mai_n1029_), .Y(mai_mai_n1969_));
  AOI220     m1920(.A0(mai_mai_n1969_), .A1(mai_mai_n466_), .B0(mai_mai_n449_), .B1(mai_mai_n390_), .Y(mai_mai_n1970_));
  NO2        m1921(.A(mai_mai_n1970_), .B(mai_mai_n156_), .Y(mai_mai_n1971_));
  NA2        m1922(.A(mai_mai_n165_), .B(mai_mai_n71_), .Y(mai_mai_n1972_));
  OAI210     m1923(.A0(mai_mai_n1877_), .A1(mai_mai_n1972_), .B0(mai_mai_n53_), .Y(mai_mai_n1973_));
  OAI220     m1924(.A0(mai_mai_n693_), .A1(mai_mai_n266_), .B0(mai_mai_n689_), .B1(x6), .Y(mai_mai_n1974_));
  NO2        m1925(.A(mai_mai_n306_), .B(x4), .Y(mai_mai_n1975_));
  AOI220     m1926(.A0(mai_mai_n1975_), .A1(mai_mai_n368_), .B0(mai_mai_n1974_), .B1(x4), .Y(mai_mai_n1976_));
  NO3        m1927(.A(mai_mai_n1976_), .B(mai_mai_n327_), .C(x5), .Y(mai_mai_n1977_));
  NO2        m1928(.A(mai_mai_n713_), .B(mai_mai_n57_), .Y(mai_mai_n1978_));
  OAI210     m1929(.A0(mai_mai_n1978_), .A1(mai_mai_n1929_), .B0(mai_mai_n451_), .Y(mai_mai_n1979_));
  AOI220     m1930(.A0(mai_mai_n670_), .A1(mai_mai_n742_), .B0(mai_mai_n498_), .B1(mai_mai_n241_), .Y(mai_mai_n1980_));
  AOI210     m1931(.A0(mai_mai_n1980_), .A1(mai_mai_n1979_), .B0(mai_mai_n261_), .Y(mai_mai_n1981_));
  NO4        m1932(.A(mai_mai_n1981_), .B(mai_mai_n1977_), .C(mai_mai_n1973_), .D(mai_mai_n1971_), .Y(mai_mai_n1982_));
  AOI220     m1933(.A0(mai_mai_n1982_), .A1(mai_mai_n1968_), .B0(mai_mai_n1960_), .B1(mai_mai_n1949_), .Y(mai_mai_n1983_));
  AOI210     m1934(.A0(mai_mai_n1937_), .A1(x3), .B0(mai_mai_n1983_), .Y(mai29));
  OAI210     m1935(.A0(mai_mai_n560_), .A1(mai_mai_n267_), .B0(mai_mai_n737_), .Y(mai_mai_n1985_));
  NA2        m1936(.A(mai_mai_n758_), .B(mai_mai_n1059_), .Y(mai_mai_n1986_));
  AO210      m1937(.A0(mai_mai_n1177_), .A1(mai_mai_n1186_), .B0(mai_mai_n1986_), .Y(mai_mai_n1987_));
  AOI210     m1938(.A0(mai_mai_n185_), .A1(mai_mai_n169_), .B0(mai_mai_n713_), .Y(mai_mai_n1988_));
  AOI210     m1939(.A0(mai_mai_n1438_), .A1(mai_mai_n78_), .B0(mai_mai_n1988_), .Y(mai_mai_n1989_));
  NA3        m1940(.A(mai_mai_n1989_), .B(mai_mai_n1987_), .C(mai_mai_n1985_), .Y(mai_mai_n1990_));
  NO3        m1941(.A(mai_mai_n672_), .B(mai_mai_n1160_), .C(mai_mai_n50_), .Y(mai_mai_n1991_));
  NO3        m1942(.A(mai_mai_n1991_), .B(mai_mai_n1264_), .C(mai_mai_n560_), .Y(mai_mai_n1992_));
  NO2        m1943(.A(mai_mai_n447_), .B(mai_mai_n58_), .Y(mai_mai_n1993_));
  AOI220     m1944(.A0(mai_mai_n1993_), .A1(mai_mai_n1223_), .B0(mai_mai_n677_), .B1(mai_mai_n1395_), .Y(mai_mai_n1994_));
  OAI210     m1945(.A0(mai_mai_n1992_), .A1(mai_mai_n546_), .B0(mai_mai_n1994_), .Y(mai_mai_n1995_));
  AOI210     m1946(.A0(mai_mai_n1990_), .A1(x6), .B0(mai_mai_n1995_), .Y(mai_mai_n1996_));
  OAI210     m1947(.A0(x8), .A1(x4), .B0(x5), .Y(mai_mai_n1997_));
  NA2        m1948(.A(mai_mai_n1997_), .B(mai_mai_n112_), .Y(mai_mai_n1998_));
  NA2        m1949(.A(mai_mai_n306_), .B(mai_mai_n149_), .Y(mai_mai_n1999_));
  NA4        m1950(.A(mai_mai_n1999_), .B(mai_mai_n1998_), .C(mai_mai_n671_), .D(mai_mai_n64_), .Y(mai_mai_n2000_));
  AOI210     m1951(.A0(mai_mai_n1335_), .A1(mai_mai_n275_), .B0(mai_mai_n1747_), .Y(mai_mai_n2001_));
  AOI210     m1952(.A0(mai_mai_n2001_), .A1(mai_mai_n2000_), .B0(mai_mai_n897_), .Y(mai_mai_n2002_));
  NA4        m1953(.A(mai_mai_n672_), .B(mai_mai_n311_), .C(mai_mai_n185_), .D(mai_mai_n169_), .Y(mai_mai_n2003_));
  NA3        m1954(.A(mai_mai_n636_), .B(mai_mai_n299_), .C(mai_mai_n809_), .Y(mai_mai_n2004_));
  AOI210     m1955(.A0(mai_mai_n2004_), .A1(mai_mai_n2003_), .B0(mai_mai_n1223_), .Y(mai_mai_n2005_));
  OAI210     m1956(.A0(mai_mai_n904_), .A1(x8), .B0(x7), .Y(mai_mai_n2006_));
  NO2        m1957(.A(mai_mai_n2006_), .B(mai_mai_n129_), .Y(mai_mai_n2007_));
  OA210      m1958(.A0(mai_mai_n877_), .A1(mai_mai_n278_), .B0(mai_mai_n1997_), .Y(mai_mai_n2008_));
  OAI220     m1959(.A0(mai_mai_n2008_), .A1(mai_mai_n592_), .B0(mai_mai_n1524_), .B1(mai_mai_n398_), .Y(mai_mai_n2009_));
  NO4        m1960(.A(mai_mai_n2009_), .B(mai_mai_n2007_), .C(mai_mai_n2005_), .D(mai_mai_n2002_), .Y(mai_mai_n2010_));
  OAI210     m1961(.A0(mai_mai_n1996_), .A1(x2), .B0(mai_mai_n2010_), .Y(mai_mai_n2011_));
  NA3        m1962(.A(x6), .B(mai_mai_n50_), .C(x2), .Y(mai_mai_n2012_));
  OAI210     m1963(.A0(mai_mai_n1242_), .A1(mai_mai_n358_), .B0(mai_mai_n2012_), .Y(mai_mai_n2013_));
  NO3        m1964(.A(mai_mai_n449_), .B(x3), .C(x0), .Y(mai_mai_n2014_));
  AO220      m1965(.A0(mai_mai_n2014_), .A1(x5), .B0(mai_mai_n1944_), .B1(mai_mai_n81_), .Y(mai_mai_n2015_));
  AOI210     m1966(.A0(mai_mai_n2013_), .A1(mai_mai_n348_), .B0(mai_mai_n2015_), .Y(mai_mai_n2016_));
  NO3        m1967(.A(mai_mai_n706_), .B(mai_mai_n369_), .C(mai_mai_n144_), .Y(mai_mai_n2017_));
  AOI210     m1968(.A0(mai_mai_n736_), .A1(mai_mai_n619_), .B0(mai_mai_n2017_), .Y(mai_mai_n2018_));
  OAI210     m1969(.A0(mai_mai_n2016_), .A1(x7), .B0(mai_mai_n2018_), .Y(mai_mai_n2019_));
  AOI210     m1970(.A0(mai_mai_n1107_), .A1(mai_mai_n403_), .B0(mai_mai_n1422_), .Y(mai_mai_n2020_));
  NO2        m1971(.A(mai_mai_n149_), .B(x2), .Y(mai_mai_n2021_));
  OA210      m1972(.A0(mai_mai_n2021_), .A1(mai_mai_n634_), .B0(mai_mai_n672_), .Y(mai_mai_n2022_));
  OAI210     m1973(.A0(mai_mai_n2022_), .A1(mai_mai_n2020_), .B0(mai_mai_n68_), .Y(mai_mai_n2023_));
  NO2        m1974(.A(mai_mai_n201_), .B(mai_mai_n85_), .Y(mai_mai_n2024_));
  OAI210     m1975(.A0(mai_mai_n2024_), .A1(mai_mai_n795_), .B0(mai_mai_n1116_), .Y(mai_mai_n2025_));
  NA3        m1976(.A(mai_mai_n1962_), .B(mai_mai_n234_), .C(mai_mai_n83_), .Y(mai_mai_n2026_));
  NA3        m1977(.A(mai_mai_n2026_), .B(mai_mai_n2025_), .C(mai_mai_n2023_), .Y(mai_mai_n2027_));
  AOI210     m1978(.A0(mai_mai_n2019_), .A1(x8), .B0(mai_mai_n2027_), .Y(mai_mai_n2028_));
  OAI210     m1979(.A0(mai_mai_n447_), .A1(mai_mai_n250_), .B0(mai_mai_n973_), .Y(mai_mai_n2029_));
  OAI210     m1980(.A0(mai_mai_n2029_), .A1(mai_mai_n1139_), .B0(mai_mai_n682_), .Y(mai_mai_n2030_));
  NO3        m1981(.A(mai_mai_n1033_), .B(mai_mai_n359_), .C(mai_mai_n150_), .Y(mai_mai_n2031_));
  NA3        m1982(.A(mai_mai_n2031_), .B(mai_mai_n1315_), .C(mai_mai_n50_), .Y(mai_mai_n2032_));
  NO2        m1983(.A(mai_mai_n137_), .B(mai_mai_n93_), .Y(mai_mai_n2033_));
  AOI220     m1984(.A0(mai_mai_n2033_), .A1(mai_mai_n593_), .B0(mai_mai_n1943_), .B1(mai_mai_n365_), .Y(mai_mai_n2034_));
  NOi31      m1985(.An(mai_mai_n1140_), .B(mai_mai_n1895_), .C(mai_mai_n629_), .Y(mai_mai_n2035_));
  NA2        m1986(.A(mai_mai_n175_), .B(x4), .Y(mai_mai_n2036_));
  NO3        m1987(.A(mai_mai_n1497_), .B(mai_mai_n245_), .C(mai_mai_n71_), .Y(mai_mai_n2037_));
  AOI210     m1988(.A0(mai_mai_n2037_), .A1(mai_mai_n2036_), .B0(mai_mai_n2035_), .Y(mai_mai_n2038_));
  NA4        m1989(.A(mai_mai_n2038_), .B(mai_mai_n2034_), .C(mai_mai_n2032_), .D(mai_mai_n2030_), .Y(mai_mai_n2039_));
  NO4        m1990(.A(mai_mai_n1242_), .B(mai_mai_n173_), .C(mai_mai_n55_), .D(mai_mai_n71_), .Y(mai_mai_n2040_));
  NO4        m1991(.A(mai_mai_n1217_), .B(mai_mai_n506_), .C(mai_mai_n1395_), .D(mai_mai_n108_), .Y(mai_mai_n2041_));
  OAI210     m1992(.A0(mai_mai_n2041_), .A1(mai_mai_n2040_), .B0(mai_mai_n110_), .Y(mai_mai_n2042_));
  AOI210     m1993(.A0(mai_mai_n310_), .A1(x4), .B0(mai_mai_n195_), .Y(mai_mai_n2043_));
  OAI210     m1994(.A0(mai_mai_n2043_), .A1(mai_mai_n1993_), .B0(mai_mai_n731_), .Y(mai_mai_n2044_));
  OR3        m1995(.A(mai_mai_n1768_), .B(mai_mai_n1447_), .C(mai_mai_n1099_), .Y(mai_mai_n2045_));
  NA2        m1996(.A(mai_mai_n1944_), .B(mai_mai_n816_), .Y(mai_mai_n2046_));
  OA220      m1997(.A0(mai_mai_n2046_), .A1(mai_mai_n250_), .B0(mai_mai_n585_), .B1(mai_mai_n1811_), .Y(mai_mai_n2047_));
  NA4        m1998(.A(mai_mai_n2047_), .B(mai_mai_n2045_), .C(mai_mai_n2044_), .D(mai_mai_n2042_), .Y(mai_mai_n2048_));
  AOI210     m1999(.A0(mai_mai_n2039_), .A1(mai_mai_n295_), .B0(mai_mai_n2048_), .Y(mai_mai_n2049_));
  OAI210     m2000(.A0(mai_mai_n2028_), .A1(x1), .B0(mai_mai_n2049_), .Y(mai_mai_n2050_));
  AO210      m2001(.A0(mai_mai_n2011_), .A1(x1), .B0(mai_mai_n2050_), .Y(mai30));
  NO3        m2002(.A(mai_mai_n1795_), .B(mai_mai_n581_), .C(mai_mai_n99_), .Y(mai_mai_n2052_));
  NO3        m2003(.A(mai_mai_n1158_), .B(mai_mai_n140_), .C(mai_mai_n386_), .Y(mai_mai_n2053_));
  AOI210     m2004(.A0(mai_mai_n731_), .A1(mai_mai_n258_), .B0(mai_mai_n2053_), .Y(mai_mai_n2054_));
  AOI210     m2005(.A0(mai_mai_n2054_), .A1(mai_mai_n2052_), .B0(mai_mai_n56_), .Y(mai_mai_n2055_));
  NA2        m2006(.A(mai_mai_n821_), .B(mai_mai_n346_), .Y(mai_mai_n2056_));
  NA2        m2007(.A(mai_mai_n2056_), .B(mai_mai_n1378_), .Y(mai_mai_n2057_));
  OAI210     m2008(.A0(mai_mai_n2057_), .A1(mai_mai_n2055_), .B0(mai_mai_n110_), .Y(mai_mai_n2058_));
  OAI210     m2009(.A0(mai_mai_n1010_), .A1(mai_mai_n575_), .B0(mai_mai_n682_), .Y(mai_mai_n2059_));
  AOI220     m2010(.A0(mai_mai_n452_), .A1(mai_mai_n949_), .B0(mai_mai_n332_), .B1(mai_mai_n460_), .Y(mai_mai_n2060_));
  AOI210     m2011(.A0(mai_mai_n2060_), .A1(mai_mai_n2059_), .B0(mai_mai_n261_), .Y(mai_mai_n2061_));
  NO3        m2012(.A(mai_mai_n284_), .B(mai_mai_n125_), .C(x0), .Y(mai_mai_n2062_));
  AOI210     m2013(.A0(mai_mai_n508_), .A1(x6), .B0(mai_mai_n2062_), .Y(mai_mai_n2063_));
  AOI220     m2014(.A0(mai_mai_n1154_), .A1(mai_mai_n427_), .B0(mai_mai_n769_), .B1(mai_mai_n92_), .Y(mai_mai_n2064_));
  OAI220     m2015(.A0(mai_mai_n2064_), .A1(mai_mai_n250_), .B0(mai_mai_n2063_), .B1(mai_mai_n54_), .Y(mai_mai_n2065_));
  NA3        m2016(.A(mai_mai_n328_), .B(mai_mai_n166_), .C(mai_mai_n71_), .Y(mai_mai_n2066_));
  AO210      m2017(.A0(mai_mai_n574_), .A1(mai_mai_n522_), .B0(x5), .Y(mai_mai_n2067_));
  AOI210     m2018(.A0(mai_mai_n2066_), .A1(mai_mai_n728_), .B0(mai_mai_n2067_), .Y(mai_mai_n2068_));
  AOI210     m2019(.A0(mai_mai_n1622_), .A1(mai_mai_n50_), .B0(mai_mai_n460_), .Y(mai_mai_n2069_));
  NA2        m2020(.A(mai_mai_n200_), .B(x2), .Y(mai_mai_n2070_));
  OA220      m2021(.A0(mai_mai_n2070_), .A1(mai_mai_n2069_), .B0(mai_mai_n279_), .B1(x6), .Y(mai_mai_n2071_));
  OAI210     m2022(.A0(x7), .A1(x6), .B0(x1), .Y(mai_mai_n2072_));
  NA3        m2023(.A(mai_mai_n57_), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n2073_));
  AOI220     m2024(.A0(mai_mai_n2073_), .A1(mai_mai_n1385_), .B0(mai_mai_n2072_), .B1(mai_mai_n1836_), .Y(mai_mai_n2074_));
  NO3        m2025(.A(mai_mai_n1381_), .B(mai_mai_n348_), .C(mai_mai_n1035_), .Y(mai_mai_n2075_));
  NO2        m2026(.A(mai_mai_n520_), .B(mai_mai_n870_), .Y(mai_mai_n2076_));
  NOi21      m2027(.An(mai_mai_n2076_), .B(mai_mai_n855_), .Y(mai_mai_n2077_));
  NO3        m2028(.A(mai_mai_n1315_), .B(mai_mai_n236_), .C(mai_mai_n654_), .Y(mai_mai_n2078_));
  NO4        m2029(.A(mai_mai_n2078_), .B(mai_mai_n2077_), .C(mai_mai_n2075_), .D(mai_mai_n2074_), .Y(mai_mai_n2079_));
  OAI210     m2030(.A0(mai_mai_n2071_), .A1(mai_mai_n765_), .B0(mai_mai_n2079_), .Y(mai_mai_n2080_));
  NO4        m2031(.A(mai_mai_n2080_), .B(mai_mai_n2068_), .C(mai_mai_n2065_), .D(mai_mai_n2061_), .Y(mai_mai_n2081_));
  AOI210     m2032(.A0(mai_mai_n2081_), .A1(mai_mai_n2058_), .B0(x8), .Y(mai_mai_n2082_));
  NO3        m2033(.A(mai_mai_n496_), .B(mai_mai_n792_), .C(mai_mai_n53_), .Y(mai_mai_n2083_));
  OAI220     m2034(.A0(mai_mai_n1811_), .A1(mai_mai_n348_), .B0(mai_mai_n488_), .B1(mai_mai_n589_), .Y(mai_mai_n2084_));
  OAI210     m2035(.A0(mai_mai_n2084_), .A1(mai_mai_n2083_), .B0(x6), .Y(mai_mai_n2085_));
  OAI210     m2036(.A0(mai_mai_n1050_), .A1(mai_mai_n541_), .B0(mai_mai_n821_), .Y(mai_mai_n2086_));
  OAI210     m2037(.A0(mai_mai_n1757_), .A1(mai_mai_n335_), .B0(mai_mai_n128_), .Y(mai_mai_n2087_));
  AOI210     m2038(.A0(mai_mai_n383_), .A1(mai_mai_n233_), .B0(mai_mai_n72_), .Y(mai_mai_n2088_));
  AOI210     m2039(.A0(mai_mai_n1010_), .A1(mai_mai_n756_), .B0(mai_mai_n2088_), .Y(mai_mai_n2089_));
  NA4        m2040(.A(mai_mai_n2089_), .B(mai_mai_n2087_), .C(mai_mai_n2086_), .D(mai_mai_n2085_), .Y(mai_mai_n2090_));
  NA2        m2041(.A(mai_mai_n1104_), .B(mai_mai_n59_), .Y(mai_mai_n2091_));
  AOI210     m2042(.A0(mai_mai_n932_), .A1(mai_mai_n497_), .B0(mai_mai_n688_), .Y(mai_mai_n2092_));
  OAI220     m2043(.A0(mai_mai_n2092_), .A1(mai_mai_n310_), .B0(mai_mai_n2091_), .B1(mai_mai_n487_), .Y(mai_mai_n2093_));
  AOI210     m2044(.A0(mai_mai_n2090_), .A1(x8), .B0(mai_mai_n2093_), .Y(mai_mai_n2094_));
  NO2        m2045(.A(mai_mai_n2094_), .B(mai_mai_n57_), .Y(mai_mai_n2095_));
  NA2        m2046(.A(mai_mai_n438_), .B(mai_mai_n855_), .Y(mai_mai_n2096_));
  NO2        m2047(.A(mai_mai_n931_), .B(mai_mai_n668_), .Y(mai_mai_n2097_));
  AOI210     m2048(.A0(mai_mai_n2097_), .A1(mai_mai_n2096_), .B0(mai_mai_n449_), .Y(mai_mai_n2098_));
  NO3        m2049(.A(mai_mai_n642_), .B(mai_mai_n412_), .C(mai_mai_n1158_), .Y(mai_mai_n2099_));
  NO3        m2050(.A(mai_mai_n2099_), .B(mai_mai_n1270_), .C(mai_mai_n1395_), .Y(mai_mai_n2100_));
  AOI210     m2051(.A0(mai_mai_n307_), .A1(x1), .B0(mai_mai_n150_), .Y(mai_mai_n2101_));
  NO2        m2052(.A(mai_mai_n313_), .B(x5), .Y(mai_mai_n2102_));
  NO2        m2053(.A(mai_mai_n2102_), .B(mai_mai_n863_), .Y(mai_mai_n2103_));
  OAI220     m2054(.A0(mai_mai_n2103_), .A1(mai_mai_n1070_), .B0(mai_mai_n2101_), .B1(mai_mai_n210_), .Y(mai_mai_n2104_));
  NO3        m2055(.A(mai_mai_n2104_), .B(mai_mai_n2100_), .C(mai_mai_n2098_), .Y(mai_mai_n2105_));
  NA2        m2056(.A(mai_mai_n971_), .B(mai_mai_n82_), .Y(mai_mai_n2106_));
  AO210      m2057(.A0(mai_mai_n2106_), .A1(mai_mai_n1623_), .B0(x3), .Y(mai_mai_n2107_));
  NO2        m2058(.A(mai_mai_n222_), .B(mai_mai_n56_), .Y(mai_mai_n2108_));
  OAI220     m2059(.A0(mai_mai_n383_), .A1(mai_mai_n1270_), .B0(mai_mai_n359_), .B1(mai_mai_n236_), .Y(mai_mai_n2109_));
  AOI220     m2060(.A0(mai_mai_n2109_), .A1(x2), .B0(mai_mai_n2108_), .B1(mai_mai_n1638_), .Y(mai_mai_n2110_));
  AOI210     m2061(.A0(mai_mai_n2110_), .A1(mai_mai_n2107_), .B0(mai_mai_n266_), .Y(mai_mai_n2111_));
  NO2        m2062(.A(mai_mai_n307_), .B(mai_mai_n124_), .Y(mai_mai_n2112_));
  NO3        m2063(.A(mai_mai_n826_), .B(mai_mai_n707_), .C(mai_mai_n169_), .Y(mai_mai_n2113_));
  OAI210     m2064(.A0(mai_mai_n2113_), .A1(mai_mai_n2112_), .B0(mai_mai_n157_), .Y(mai_mai_n2114_));
  NA3        m2065(.A(x5), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n2115_));
  AOI210     m2066(.A0(mai_mai_n2115_), .A1(mai_mai_n1323_), .B0(mai_mai_n542_), .Y(mai_mai_n2116_));
  AOI210     m2067(.A0(mai_mai_n1343_), .A1(x2), .B0(mai_mai_n2116_), .Y(mai_mai_n2117_));
  AOI210     m2068(.A0(mai_mai_n2117_), .A1(mai_mai_n2114_), .B0(mai_mai_n50_), .Y(mai_mai_n2118_));
  NA3        m2069(.A(mai_mai_n1494_), .B(mai_mai_n1149_), .C(mai_mai_n480_), .Y(mai_mai_n2119_));
  AOI210     m2070(.A0(mai_mai_n2119_), .A1(mai_mai_n2106_), .B0(mai_mai_n615_), .Y(mai_mai_n2120_));
  AOI210     m2071(.A0(mai_mai_n1035_), .A1(x1), .B0(mai_mai_n1335_), .Y(mai_mai_n2121_));
  OAI220     m2072(.A0(mai_mai_n311_), .A1(x4), .B0(mai_mai_n51_), .B1(x6), .Y(mai_mai_n2122_));
  NO2        m2073(.A(mai_mai_n123_), .B(mai_mai_n112_), .Y(mai_mai_n2123_));
  AOI220     m2074(.A0(mai_mai_n2123_), .A1(mai_mai_n2122_), .B0(mai_mai_n1179_), .B1(mai_mai_n629_), .Y(mai_mai_n2124_));
  OAI210     m2075(.A0(mai_mai_n2121_), .A1(mai_mai_n491_), .B0(mai_mai_n2124_), .Y(mai_mai_n2125_));
  NO4        m2076(.A(mai_mai_n2125_), .B(mai_mai_n2120_), .C(mai_mai_n2118_), .D(mai_mai_n2111_), .Y(mai_mai_n2126_));
  OAI210     m2077(.A0(mai_mai_n2105_), .A1(mai_mai_n137_), .B0(mai_mai_n2126_), .Y(mai_mai_n2127_));
  NO3        m2078(.A(mai_mai_n2127_), .B(mai_mai_n2095_), .C(mai_mai_n2082_), .Y(mai31));
  NA2        m2079(.A(mai_mai_n995_), .B(mai_mai_n360_), .Y(mai_mai_n2129_));
  NO2        m2080(.A(mai_mai_n453_), .B(mai_mai_n682_), .Y(mai_mai_n2130_));
  AOI210     m2081(.A0(mai_mai_n2130_), .A1(mai_mai_n2129_), .B0(mai_mai_n58_), .Y(mai_mai_n2131_));
  NO2        m2082(.A(mai_mai_n794_), .B(mai_mai_n56_), .Y(mai_mai_n2132_));
  AOI220     m2083(.A0(mai_mai_n2132_), .A1(x2), .B0(mai_mai_n91_), .B1(x0), .Y(mai_mai_n2133_));
  NA3        m2084(.A(mai_mai_n2133_), .B(mai_mai_n2046_), .C(mai_mai_n1874_), .Y(mai_mai_n2134_));
  OAI210     m2085(.A0(mai_mai_n2134_), .A1(mai_mai_n2131_), .B0(mai_mai_n53_), .Y(mai_mai_n2135_));
  NO2        m2086(.A(mai_mai_n435_), .B(mai_mai_n682_), .Y(mai_mai_n2136_));
  NO3        m2087(.A(mai_mai_n1975_), .B(mai_mai_n1944_), .C(mai_mai_n898_), .Y(mai_mai_n2137_));
  OA220      m2088(.A0(mai_mai_n2137_), .A1(mai_mai_n480_), .B0(mai_mai_n2136_), .B1(mai_mai_n1487_), .Y(mai_mai_n2138_));
  AOI210     m2089(.A0(mai_mai_n2138_), .A1(mai_mai_n2135_), .B0(mai_mai_n108_), .Y(mai_mai_n2139_));
  NO2        m2090(.A(mai_mai_n502_), .B(mai_mai_n75_), .Y(mai_mai_n2140_));
  NA2        m2091(.A(mai_mai_n449_), .B(mai_mai_n57_), .Y(mai_mai_n2141_));
  AOI210     m2092(.A0(mai_mai_n310_), .A1(mai_mai_n86_), .B0(mai_mai_n2141_), .Y(mai_mai_n2142_));
  OAI210     m2093(.A0(mai_mai_n2142_), .A1(mai_mai_n2140_), .B0(mai_mai_n780_), .Y(mai_mai_n2143_));
  NO4        m2094(.A(mai_mai_n1175_), .B(mai_mai_n369_), .C(mai_mai_n1622_), .D(mai_mai_n67_), .Y(mai_mai_n2144_));
  AOI210     m2095(.A0(mai_mai_n1662_), .A1(mai_mai_n1370_), .B0(mai_mai_n447_), .Y(mai_mai_n2145_));
  OAI220     m2096(.A0(mai_mai_n1324_), .A1(mai_mai_n963_), .B0(mai_mai_n782_), .B1(mai_mai_n117_), .Y(mai_mai_n2146_));
  NO3        m2097(.A(mai_mai_n2146_), .B(mai_mai_n2145_), .C(mai_mai_n2144_), .Y(mai_mai_n2147_));
  AOI210     m2098(.A0(mai_mai_n2147_), .A1(mai_mai_n2143_), .B0(x5), .Y(mai_mai_n2148_));
  AOI220     m2099(.A0(mai_mai_n451_), .A1(mai_mai_n629_), .B0(mai_mai_n575_), .B1(mai_mai_n63_), .Y(mai_mai_n2149_));
  AOI210     m2100(.A0(mai_mai_n2149_), .A1(mai_mai_n585_), .B0(mai_mai_n1242_), .Y(mai_mai_n2150_));
  AOI220     m2101(.A0(mai_mai_n972_), .A1(mai_mai_n742_), .B0(mai_mai_n1158_), .B1(mai_mai_n122_), .Y(mai_mai_n2151_));
  OAI220     m2102(.A0(mai_mai_n2151_), .A1(mai_mai_n389_), .B0(mai_mai_n487_), .B1(mai_mai_n781_), .Y(mai_mai_n2152_));
  NO4        m2103(.A(mai_mai_n2152_), .B(mai_mai_n2150_), .C(mai_mai_n2148_), .D(mai_mai_n2139_), .Y(mai_mai_n2153_));
  NA2        m2104(.A(mai_mai_n497_), .B(mai_mai_n59_), .Y(mai_mai_n2154_));
  AOI210     m2105(.A0(mai_mai_n546_), .A1(mai_mai_n2154_), .B0(mai_mai_n143_), .Y(mai_mai_n2155_));
  OAI210     m2106(.A0(mai_mai_n104_), .A1(mai_mai_n278_), .B0(mai_mai_n2091_), .Y(mai_mai_n2156_));
  OAI210     m2107(.A0(mai_mai_n2156_), .A1(mai_mai_n2155_), .B0(x7), .Y(mai_mai_n2157_));
  NO3        m2108(.A(mai_mai_n383_), .B(mai_mai_n55_), .C(x7), .Y(mai_mai_n2158_));
  OA210      m2109(.A0(mai_mai_n2158_), .A1(mai_mai_n1334_), .B0(mai_mai_n101_), .Y(mai_mai_n2159_));
  NA2        m2110(.A(mai_mai_n1101_), .B(mai_mai_n92_), .Y(mai_mai_n2160_));
  AOI210     m2111(.A0(mai_mai_n910_), .A1(mai_mai_n112_), .B0(mai_mai_n2160_), .Y(mai_mai_n2161_));
  NA2        m2112(.A(mai_mai_n1569_), .B(x6), .Y(mai_mai_n2162_));
  AOI210     m2113(.A0(mai_mai_n2162_), .A1(mai_mai_n294_), .B0(mai_mai_n108_), .Y(mai_mai_n2163_));
  NA2        m2114(.A(mai_mai_n1202_), .B(mai_mai_n323_), .Y(mai_mai_n2164_));
  AOI210     m2115(.A0(mai_mai_n2164_), .A1(mai_mai_n650_), .B0(mai_mai_n53_), .Y(mai_mai_n2165_));
  NO4        m2116(.A(mai_mai_n2165_), .B(mai_mai_n2163_), .C(mai_mai_n2161_), .D(mai_mai_n2159_), .Y(mai_mai_n2166_));
  AOI210     m2117(.A0(mai_mai_n2166_), .A1(mai_mai_n2157_), .B0(mai_mai_n692_), .Y(mai_mai_n2167_));
  NOi21      m2118(.An(mai_mai_n1785_), .B(mai_mai_n1074_), .Y(mai_mai_n2168_));
  OAI220     m2119(.A0(mai_mai_n2168_), .A1(mai_mai_n1946_), .B0(mai_mai_n933_), .B1(mai_mai_n2154_), .Y(mai_mai_n2169_));
  NA2        m2120(.A(mai_mai_n2169_), .B(x3), .Y(mai_mai_n2170_));
  AOI220     m2121(.A0(mai_mai_n1405_), .A1(x8), .B0(mai_mai_n60_), .B1(x1), .Y(mai_mai_n2171_));
  NO3        m2122(.A(mai_mai_n2171_), .B(mai_mai_n1128_), .C(x6), .Y(mai_mai_n2172_));
  AOI220     m2123(.A0(mai_mai_n619_), .A1(mai_mai_n412_), .B0(mai_mai_n497_), .B1(mai_mai_n78_), .Y(mai_mai_n2173_));
  NA2        m2124(.A(mai_mai_n118_), .B(mai_mai_n533_), .Y(mai_mai_n2174_));
  OAI220     m2125(.A0(mai_mai_n2174_), .A1(mai_mai_n1946_), .B0(mai_mai_n2173_), .B1(x4), .Y(mai_mai_n2175_));
  NO2        m2126(.A(mai_mai_n2175_), .B(mai_mai_n2172_), .Y(mai_mai_n2176_));
  AOI210     m2127(.A0(mai_mai_n2176_), .A1(mai_mai_n2170_), .B0(mai_mai_n188_), .Y(mai_mai_n2177_));
  NO4        m2128(.A(mai_mai_n620_), .B(mai_mai_n593_), .C(mai_mai_n708_), .D(mai_mai_n707_), .Y(mai_mai_n2178_));
  OAI210     m2129(.A0(mai_mai_n2178_), .A1(mai_mai_n1092_), .B0(x3), .Y(mai_mai_n2179_));
  NO4        m2130(.A(mai_mai_n812_), .B(mai_mai_n1242_), .C(mai_mai_n780_), .D(x5), .Y(mai_mai_n2180_));
  NO3        m2131(.A(x6), .B(mai_mai_n56_), .C(x1), .Y(mai_mai_n2181_));
  NA2        m2132(.A(mai_mai_n2181_), .B(mai_mai_n290_), .Y(mai_mai_n2182_));
  OAI210     m2133(.A0(mai_mai_n1916_), .A1(mai_mai_n383_), .B0(mai_mai_n2182_), .Y(mai_mai_n2183_));
  NA4        m2134(.A(mai_mai_n642_), .B(mai_mai_n181_), .C(x6), .D(mai_mai_n108_), .Y(mai_mai_n2184_));
  NO2        m2135(.A(mai_mai_n864_), .B(mai_mai_n254_), .Y(mai_mai_n2185_));
  NOi41      m2136(.An(mai_mai_n2184_), .B(mai_mai_n2185_), .C(mai_mai_n2183_), .D(mai_mai_n2180_), .Y(mai_mai_n2186_));
  AOI210     m2137(.A0(mai_mai_n2186_), .A1(mai_mai_n2179_), .B0(mai_mai_n537_), .Y(mai_mai_n2187_));
  OAI210     m2138(.A0(mai_mai_n619_), .A1(mai_mai_n474_), .B0(mai_mai_n949_), .Y(mai_mai_n2188_));
  NO3        m2139(.A(mai_mai_n379_), .B(mai_mai_n77_), .C(mai_mai_n53_), .Y(mai_mai_n2189_));
  NO3        m2140(.A(mai_mai_n466_), .B(mai_mai_n354_), .C(mai_mai_n50_), .Y(mai_mai_n2190_));
  OAI210     m2141(.A0(mai_mai_n2190_), .A1(mai_mai_n2189_), .B0(mai_mai_n1176_), .Y(mai_mai_n2191_));
  AOI210     m2142(.A0(mai_mai_n2191_), .A1(mai_mai_n2188_), .B0(mai_mai_n396_), .Y(mai_mai_n2192_));
  NO2        m2143(.A(mai_mai_n219_), .B(mai_mai_n542_), .Y(mai_mai_n2193_));
  OAI210     m2144(.A0(mai_mai_n140_), .A1(x2), .B0(mai_mai_n2193_), .Y(mai_mai_n2194_));
  NO2        m2145(.A(mai_mai_n2194_), .B(mai_mai_n64_), .Y(mai_mai_n2195_));
  NA2        m2146(.A(mai_mai_n123_), .B(mai_mai_n57_), .Y(mai_mai_n2196_));
  AOI220     m2147(.A0(mai_mai_n1601_), .A1(mai_mai_n917_), .B0(mai_mai_n277_), .B1(x4), .Y(mai_mai_n2197_));
  AOI220     m2148(.A0(mai_mai_n1654_), .A1(mai_mai_n621_), .B0(mai_mai_n729_), .B1(mai_mai_n780_), .Y(mai_mai_n2198_));
  OAI220     m2149(.A0(mai_mai_n2198_), .A1(mai_mai_n2196_), .B0(mai_mai_n2197_), .B1(mai_mai_n193_), .Y(mai_mai_n2199_));
  OR3        m2150(.A(mai_mai_n2199_), .B(mai_mai_n2195_), .C(mai_mai_n2192_), .Y(mai_mai_n2200_));
  NO4        m2151(.A(mai_mai_n2200_), .B(mai_mai_n2187_), .C(mai_mai_n2177_), .D(mai_mai_n2167_), .Y(mai_mai_n2201_));
  OAI210     m2152(.A0(mai_mai_n2153_), .A1(x3), .B0(mai_mai_n2201_), .Y(mai32));
  OAI210     m2153(.A0(mai_mai_n568_), .A1(mai_mai_n53_), .B0(mai_mai_n417_), .Y(mai_mai_n2203_));
  NA2        m2154(.A(mai_mai_n517_), .B(x2), .Y(mai_mai_n2204_));
  AOI210     m2155(.A0(mai_mai_n2204_), .A1(mai_mai_n2203_), .B0(mai_mai_n57_), .Y(mai_mai_n2205_));
  OAI210     m2156(.A0(mai_mai_n2205_), .A1(mai_mai_n795_), .B0(mai_mai_n56_), .Y(mai_mai_n2206_));
  OAI210     m2157(.A0(mai_mai_n1726_), .A1(mai_mai_n1466_), .B0(mai_mai_n1496_), .Y(mai_mai_n2207_));
  AOI210     m2158(.A0(mai_mai_n2132_), .A1(mai_mai_n281_), .B0(mai_mai_n2207_), .Y(mai_mai_n2208_));
  AOI210     m2159(.A0(mai_mai_n2208_), .A1(mai_mai_n2206_), .B0(mai_mai_n50_), .Y(mai_mai_n2209_));
  NA3        m2160(.A(mai_mai_n1570_), .B(mai_mai_n810_), .C(mai_mai_n293_), .Y(mai_mai_n2210_));
  NA2        m2161(.A(mai_mai_n753_), .B(mai_mai_n550_), .Y(mai_mai_n2211_));
  OAI220     m2162(.A0(mai_mai_n1069_), .A1(mai_mai_n234_), .B0(mai_mai_n689_), .B1(mai_mai_n210_), .Y(mai_mai_n2212_));
  NO3        m2163(.A(mai_mai_n380_), .B(mai_mai_n578_), .C(mai_mai_n816_), .Y(mai_mai_n2213_));
  NO3        m2164(.A(mai_mai_n1381_), .B(mai_mai_n589_), .C(mai_mai_n275_), .Y(mai_mai_n2214_));
  NO4        m2165(.A(mai_mai_n2214_), .B(mai_mai_n2213_), .C(mai_mai_n2212_), .D(mai_mai_n2211_), .Y(mai_mai_n2215_));
  AOI210     m2166(.A0(mai_mai_n2215_), .A1(mai_mai_n2210_), .B0(mai_mai_n144_), .Y(mai_mai_n2216_));
  OAI220     m2167(.A0(mai_mai_n405_), .A1(x7), .B0(mai_mai_n306_), .B1(mai_mai_n299_), .Y(mai_mai_n2217_));
  NA2        m2168(.A(mai_mai_n2217_), .B(mai_mai_n971_), .Y(mai_mai_n2218_));
  NO2        m2169(.A(mai_mai_n555_), .B(mai_mai_n870_), .Y(mai_mai_n2219_));
  AOI220     m2170(.A0(mai_mai_n2219_), .A1(mai_mai_n1898_), .B0(mai_mai_n534_), .B1(mai_mai_n133_), .Y(mai_mai_n2220_));
  AOI210     m2171(.A0(mai_mai_n2220_), .A1(mai_mai_n2218_), .B0(mai_mai_n110_), .Y(mai_mai_n2221_));
  NA3        m2172(.A(mai_mai_n1334_), .B(mai_mai_n1160_), .C(mai_mai_n117_), .Y(mai_mai_n2222_));
  NA2        m2173(.A(mai_mai_n1371_), .B(mai_mai_n708_), .Y(mai_mai_n2223_));
  AOI210     m2174(.A0(mai_mai_n2223_), .A1(mai_mai_n2222_), .B0(mai_mai_n56_), .Y(mai_mai_n2224_));
  NA2        m2175(.A(mai_mai_n971_), .B(mai_mai_n57_), .Y(mai_mai_n2225_));
  NOi21      m2176(.An(mai_mai_n2225_), .B(mai_mai_n133_), .Y(mai_mai_n2226_));
  NA2        m2177(.A(mai_mai_n1025_), .B(mai_mai_n254_), .Y(mai_mai_n2227_));
  NO3        m2178(.A(mai_mai_n2227_), .B(mai_mai_n2226_), .C(mai_mai_n59_), .Y(mai_mai_n2228_));
  OR4        m2179(.A(mai_mai_n2228_), .B(mai_mai_n2224_), .C(mai_mai_n2221_), .D(mai_mai_n2216_), .Y(mai_mai_n2229_));
  OAI210     m2180(.A0(mai_mai_n2229_), .A1(mai_mai_n2209_), .B0(mai_mai_n108_), .Y(mai_mai_n2230_));
  NO3        m2181(.A(mai_mai_n1242_), .B(mai_mai_n147_), .C(mai_mai_n126_), .Y(mai_mai_n2231_));
  NO2        m2182(.A(mai_mai_n384_), .B(mai_mai_n55_), .Y(mai_mai_n2232_));
  NA2        m2183(.A(mai_mai_n2232_), .B(mai_mai_n116_), .Y(mai_mai_n2233_));
  OAI210     m2184(.A0(mai_mai_n638_), .A1(mai_mai_n595_), .B0(mai_mai_n821_), .Y(mai_mai_n2234_));
  NA2        m2185(.A(mai_mai_n2234_), .B(mai_mai_n2233_), .Y(mai_mai_n2235_));
  OAI210     m2186(.A0(mai_mai_n2235_), .A1(mai_mai_n2231_), .B0(x3), .Y(mai_mai_n2236_));
  OAI210     m2187(.A0(mai_mai_n904_), .A1(mai_mai_n275_), .B0(mai_mai_n50_), .Y(mai_mai_n2237_));
  AOI210     m2188(.A0(mai_mai_n62_), .A1(mai_mai_n110_), .B0(mai_mai_n2237_), .Y(mai_mai_n2238_));
  OAI210     m2189(.A0(mai_mai_n2238_), .A1(mai_mai_n1879_), .B0(mai_mai_n707_), .Y(mai_mai_n2239_));
  NO3        m2190(.A(mai_mai_n308_), .B(mai_mai_n175_), .C(mai_mai_n124_), .Y(mai_mai_n2240_));
  NO3        m2191(.A(mai_mai_n810_), .B(mai_mai_n367_), .C(mai_mai_n144_), .Y(mai_mai_n2241_));
  OAI210     m2192(.A0(mai_mai_n2241_), .A1(mai_mai_n2240_), .B0(mai_mai_n59_), .Y(mai_mai_n2242_));
  NA2        m2193(.A(mai_mai_n1164_), .B(mai_mai_n71_), .Y(mai_mai_n2243_));
  NO2        m2194(.A(mai_mai_n1950_), .B(mai_mai_n595_), .Y(mai_mai_n2244_));
  AOI210     m2195(.A0(mai_mai_n2244_), .A1(mai_mai_n1880_), .B0(mai_mai_n2243_), .Y(mai_mai_n2245_));
  NO2        m2196(.A(mai_mai_n278_), .B(mai_mai_n57_), .Y(mai_mai_n2246_));
  NO2        m2197(.A(mai_mai_n2246_), .B(mai_mai_n1017_), .Y(mai_mai_n2247_));
  NOi31      m2198(.An(mai_mai_n731_), .B(mai_mai_n2247_), .C(mai_mai_n284_), .Y(mai_mai_n2248_));
  NO3        m2199(.A(mai_mai_n1326_), .B(mai_mai_n219_), .C(mai_mai_n261_), .Y(mai_mai_n2249_));
  NO4        m2200(.A(mai_mai_n2249_), .B(mai_mai_n2248_), .C(mai_mai_n2245_), .D(x1), .Y(mai_mai_n2250_));
  NA4        m2201(.A(mai_mai_n2250_), .B(mai_mai_n2242_), .C(mai_mai_n2239_), .D(mai_mai_n2236_), .Y(mai_mai_n2251_));
  AO210      m2202(.A0(mai_mai_n1107_), .A1(mai_mai_n400_), .B0(mai_mai_n1020_), .Y(mai_mai_n2252_));
  NA3        m2203(.A(mai_mai_n1922_), .B(mai_mai_n559_), .C(mai_mai_n278_), .Y(mai_mai_n2253_));
  AOI210     m2204(.A0(mai_mai_n2253_), .A1(mai_mai_n2252_), .B0(mai_mai_n308_), .Y(mai_mai_n2254_));
  NA4        m2205(.A(mai_mai_n1279_), .B(mai_mai_n531_), .C(mai_mai_n389_), .D(mai_mai_n234_), .Y(mai_mai_n2255_));
  NO3        m2206(.A(mai_mai_n1447_), .B(mai_mai_n1020_), .C(x2), .Y(mai_mai_n2256_));
  NO2        m2207(.A(mai_mai_n1265_), .B(mai_mai_n387_), .Y(mai_mai_n2257_));
  NO2        m2208(.A(mai_mai_n1853_), .B(mai_mai_n64_), .Y(mai_mai_n2258_));
  NO4        m2209(.A(mai_mai_n2258_), .B(mai_mai_n2257_), .C(mai_mai_n2256_), .D(mai_mai_n53_), .Y(mai_mai_n2259_));
  NO3        m2210(.A(mai_mai_n470_), .B(mai_mai_n1101_), .C(mai_mai_n123_), .Y(mai_mai_n2260_));
  OAI220     m2211(.A0(mai_mai_n692_), .A1(mai_mai_n175_), .B0(mai_mai_n359_), .B1(mai_mai_n144_), .Y(mai_mai_n2261_));
  OAI210     m2212(.A0(mai_mai_n2261_), .A1(mai_mai_n2260_), .B0(mai_mai_n68_), .Y(mai_mai_n2262_));
  NO2        m2213(.A(mai_mai_n1997_), .B(mai_mai_n371_), .Y(mai_mai_n2263_));
  OAI210     m2214(.A0(mai_mai_n1885_), .A1(mai_mai_n613_), .B0(mai_mai_n2263_), .Y(mai_mai_n2264_));
  NA4        m2215(.A(mai_mai_n2264_), .B(mai_mai_n2262_), .C(mai_mai_n2259_), .D(mai_mai_n2255_), .Y(mai_mai_n2265_));
  OAI210     m2216(.A0(mai_mai_n2265_), .A1(mai_mai_n2254_), .B0(mai_mai_n2251_), .Y(mai_mai_n2266_));
  NO3        m2217(.A(mai_mai_n1229_), .B(mai_mai_n107_), .C(mai_mai_n71_), .Y(mai_mai_n2267_));
  NO2        m2218(.A(mai_mai_n568_), .B(mai_mai_n375_), .Y(mai_mai_n2268_));
  OAI210     m2219(.A0(mai_mai_n2267_), .A1(mai_mai_n1428_), .B0(mai_mai_n2268_), .Y(mai_mai_n2269_));
  NO3        m2220(.A(x8), .B(mai_mai_n71_), .C(x2), .Y(mai_mai_n2270_));
  OAI220     m2221(.A0(mai_mai_n2270_), .A1(mai_mai_n629_), .B0(mai_mai_n1438_), .B1(mai_mai_n91_), .Y(mai_mai_n2271_));
  AOI220     m2222(.A0(mai_mai_n560_), .A1(mai_mai_n821_), .B0(mai_mai_n682_), .B1(mai_mai_n259_), .Y(mai_mai_n2272_));
  AOI210     m2223(.A0(mai_mai_n2272_), .A1(mai_mai_n2271_), .B0(mai_mai_n269_), .Y(mai_mai_n2273_));
  NA2        m2224(.A(mai_mai_n1025_), .B(mai_mai_n1158_), .Y(mai_mai_n2274_));
  AOI210     m2225(.A0(mai_mai_n678_), .A1(mai_mai_n692_), .B0(mai_mai_n2274_), .Y(mai_mai_n2275_));
  AOI210     m2226(.A0(mai_mai_n593_), .A1(mai_mai_n629_), .B0(mai_mai_n698_), .Y(mai_mai_n2276_));
  NO2        m2227(.A(mai_mai_n2276_), .B(mai_mai_n1836_), .Y(mai_mai_n2277_));
  NO2        m2228(.A(mai_mai_n454_), .B(mai_mai_n435_), .Y(mai_mai_n2278_));
  NOi31      m2229(.An(mai_mai_n1516_), .B(mai_mai_n2278_), .C(mai_mai_n593_), .Y(mai_mai_n2279_));
  NO4        m2230(.A(mai_mai_n2279_), .B(mai_mai_n2277_), .C(mai_mai_n2275_), .D(mai_mai_n2273_), .Y(mai_mai_n2280_));
  NA4        m2231(.A(mai_mai_n2280_), .B(mai_mai_n2269_), .C(mai_mai_n2266_), .D(mai_mai_n2230_), .Y(mai33));
  OAI210     m2232(.A0(mai_mai_n817_), .A1(x1), .B0(mai_mai_n204_), .Y(mai_mai_n2282_));
  OAI210     m2233(.A0(mai_mai_n2102_), .A1(mai_mai_n180_), .B0(mai_mai_n333_), .Y(mai_mai_n2283_));
  OAI220     m2234(.A0(mai_mai_n1087_), .A1(mai_mai_n816_), .B0(mai_mai_n1689_), .B1(mai_mai_n358_), .Y(mai_mai_n2284_));
  NA3        m2235(.A(mai_mai_n2284_), .B(mai_mai_n2283_), .C(mai_mai_n641_), .Y(mai_mai_n2285_));
  AOI210     m2236(.A0(mai_mai_n2282_), .A1(x5), .B0(mai_mai_n2285_), .Y(mai_mai_n2286_));
  NA2        m2237(.A(mai_mai_n233_), .B(mai_mai_n76_), .Y(mai_mai_n2287_));
  NA4        m2238(.A(mai_mai_n1764_), .B(mai_mai_n569_), .C(mai_mai_n250_), .D(x4), .Y(mai_mai_n2288_));
  AOI210     m2239(.A0(mai_mai_n2288_), .A1(mai_mai_n2287_), .B0(mai_mai_n358_), .Y(mai_mai_n2289_));
  OAI210     m2240(.A0(mai_mai_n438_), .A1(mai_mai_n272_), .B0(mai_mai_n53_), .Y(mai_mai_n2290_));
  AOI210     m2241(.A0(mai_mai_n2290_), .A1(mai_mai_n440_), .B0(mai_mai_n64_), .Y(mai_mai_n2291_));
  NA2        m2242(.A(mai_mai_n1677_), .B(mai_mai_n71_), .Y(mai_mai_n2292_));
  NO3        m2243(.A(mai_mai_n2292_), .B(mai_mai_n2291_), .C(mai_mai_n2289_), .Y(mai_mai_n2293_));
  OAI210     m2244(.A0(mai_mai_n2286_), .A1(x4), .B0(mai_mai_n2293_), .Y(mai_mai_n2294_));
  OAI210     m2245(.A0(mai_mai_n145_), .A1(x5), .B0(mai_mai_n243_), .Y(mai_mai_n2295_));
  NA2        m2246(.A(mai_mai_n188_), .B(x4), .Y(mai_mai_n2296_));
  NA2        m2247(.A(mai_mai_n313_), .B(mai_mai_n290_), .Y(mai_mai_n2297_));
  NO2        m2248(.A(mai_mai_n971_), .B(mai_mai_n231_), .Y(mai_mai_n2298_));
  NA2        m2249(.A(mai_mai_n644_), .B(x7), .Y(mai_mai_n2299_));
  OAI220     m2250(.A0(mai_mai_n2299_), .A1(mai_mai_n2298_), .B0(mai_mai_n2297_), .B1(mai_mai_n2296_), .Y(mai_mai_n2300_));
  AOI210     m2251(.A0(mai_mai_n2295_), .A1(mai_mai_n1033_), .B0(mai_mai_n2300_), .Y(mai_mai_n2301_));
  NA2        m2252(.A(mai_mai_n215_), .B(mai_mai_n962_), .Y(mai_mai_n2302_));
  AOI210     m2253(.A0(mai_mai_n2302_), .A1(mai_mai_n2225_), .B0(mai_mai_n217_), .Y(mai_mai_n2303_));
  NO2        m2254(.A(mai_mai_n1663_), .B(mai_mai_n963_), .Y(mai_mai_n2304_));
  OAI210     m2255(.A0(mai_mai_n870_), .A1(mai_mai_n51_), .B0(x6), .Y(mai_mai_n2305_));
  NA3        m2256(.A(mai_mai_n927_), .B(mai_mai_n737_), .C(mai_mai_n55_), .Y(mai_mai_n2306_));
  OAI210     m2257(.A0(mai_mai_n623_), .A1(mai_mai_n508_), .B0(mai_mai_n2306_), .Y(mai_mai_n2307_));
  NO4        m2258(.A(mai_mai_n2307_), .B(mai_mai_n2305_), .C(mai_mai_n2304_), .D(mai_mai_n2303_), .Y(mai_mai_n2308_));
  OAI210     m2259(.A0(mai_mai_n2301_), .A1(mai_mai_n50_), .B0(mai_mai_n2308_), .Y(mai_mai_n2309_));
  NA3        m2260(.A(mai_mai_n2309_), .B(mai_mai_n2294_), .C(mai_mai_n59_), .Y(mai_mai_n2310_));
  NA2        m2261(.A(mai_mai_n538_), .B(mai_mai_n109_), .Y(mai_mai_n2311_));
  NO3        m2262(.A(mai_mai_n1582_), .B(mai_mai_n379_), .C(x4), .Y(mai_mai_n2312_));
  AOI210     m2263(.A0(mai_mai_n2312_), .A1(mai_mai_n2311_), .B0(mai_mai_n441_), .Y(mai_mai_n2313_));
  NA2        m2264(.A(mai_mai_n819_), .B(mai_mai_n108_), .Y(mai_mai_n2314_));
  NA2        m2265(.A(mai_mai_n504_), .B(mai_mai_n53_), .Y(mai_mai_n2315_));
  INV        m2266(.A(mai_mai_n2315_), .Y(mai_mai_n2316_));
  OAI210     m2267(.A0(mai_mai_n2313_), .A1(mai_mai_n59_), .B0(mai_mai_n2316_), .Y(mai_mai_n2317_));
  AOI220     m2268(.A0(mai_mai_n692_), .A1(mai_mai_n240_), .B0(mai_mai_n389_), .B1(mai_mai_n234_), .Y(mai_mai_n2318_));
  NA2        m2269(.A(mai_mai_n738_), .B(mai_mai_n983_), .Y(mai_mai_n2319_));
  OAI210     m2270(.A0(mai_mai_n2319_), .A1(mai_mai_n2318_), .B0(mai_mai_n307_), .Y(mai_mai_n2320_));
  AOI210     m2271(.A0(mai_mai_n2132_), .A1(mai_mai_n218_), .B0(mai_mai_n53_), .Y(mai_mai_n2321_));
  NO2        m2272(.A(mai_mai_n144_), .B(mai_mai_n343_), .Y(mai_mai_n2322_));
  AOI220     m2273(.A0(mai_mai_n2322_), .A1(mai_mai_n1003_), .B0(mai_mai_n677_), .B1(mai_mai_n358_), .Y(mai_mai_n2323_));
  NA2        m2274(.A(mai_mai_n449_), .B(mai_mai_n502_), .Y(mai_mai_n2324_));
  NO3        m2275(.A(mai_mai_n2324_), .B(mai_mai_n1039_), .C(mai_mai_n185_), .Y(mai_mai_n2325_));
  AOI210     m2276(.A0(mai_mai_n1812_), .A1(mai_mai_n1202_), .B0(mai_mai_n2325_), .Y(mai_mai_n2326_));
  NA4        m2277(.A(mai_mai_n2326_), .B(mai_mai_n2323_), .C(mai_mai_n2321_), .D(mai_mai_n2320_), .Y(mai_mai_n2327_));
  NA3        m2278(.A(mai_mai_n2327_), .B(mai_mai_n2317_), .C(mai_mai_n57_), .Y(mai_mai_n2328_));
  NAi21      m2279(.An(mai_mai_n1204_), .B(mai_mai_n493_), .Y(mai_mai_n2329_));
  NA4        m2280(.A(mai_mai_n644_), .B(mai_mai_n1315_), .C(mai_mai_n474_), .D(mai_mai_n50_), .Y(mai_mai_n2330_));
  OAI210     m2281(.A0(mai_mai_n2322_), .A1(mai_mai_n2076_), .B0(x2), .Y(mai_mai_n2331_));
  NA4        m2282(.A(mai_mai_n290_), .B(mai_mai_n158_), .C(mai_mai_n279_), .D(mai_mai_n123_), .Y(mai_mai_n2332_));
  NA3        m2283(.A(mai_mai_n2332_), .B(mai_mai_n2331_), .C(mai_mai_n2330_), .Y(mai_mai_n2333_));
  AO220      m2284(.A0(mai_mai_n2333_), .A1(x0), .B0(mai_mai_n2329_), .B1(mai_mai_n141_), .Y(mai_mai_n2334_));
  NA3        m2285(.A(mai_mai_n780_), .B(mai_mai_n358_), .C(mai_mai_n60_), .Y(mai_mai_n2335_));
  NO2        m2286(.A(mai_mai_n2270_), .B(mai_mai_n416_), .Y(mai_mai_n2336_));
  NA2        m2287(.A(mai_mai_n642_), .B(mai_mai_n520_), .Y(mai_mai_n2337_));
  OAI220     m2288(.A0(mai_mai_n2337_), .A1(mai_mai_n2336_), .B0(mai_mai_n2335_), .B1(mai_mai_n71_), .Y(mai_mai_n2338_));
  OAI210     m2289(.A0(mai_mai_n1546_), .A1(mai_mai_n354_), .B0(mai_mai_n111_), .Y(mai_mai_n2339_));
  AOI210     m2290(.A0(mai_mai_n593_), .A1(mai_mai_n470_), .B0(mai_mai_n141_), .Y(mai_mai_n2340_));
  OAI210     m2291(.A0(mai_mai_n2340_), .A1(mai_mai_n389_), .B0(mai_mai_n2339_), .Y(mai_mai_n2341_));
  OAI210     m2292(.A0(mai_mai_n2341_), .A1(mai_mai_n2338_), .B0(mai_mai_n102_), .Y(mai_mai_n2342_));
  NA3        m2293(.A(mai_mai_n1222_), .B(mai_mai_n134_), .C(mai_mai_n384_), .Y(mai_mai_n2343_));
  NA2        m2294(.A(mai_mai_n2343_), .B(mai_mai_n1840_), .Y(mai_mai_n2344_));
  NA2        m2295(.A(mai_mai_n1201_), .B(mai_mai_n716_), .Y(mai_mai_n2345_));
  AOI220     m2296(.A0(mai_mai_n2232_), .A1(mai_mai_n298_), .B0(mai_mai_n1371_), .B1(mai_mai_n1182_), .Y(mai_mai_n2346_));
  NA4        m2297(.A(mai_mai_n2346_), .B(mai_mai_n2345_), .C(mai_mai_n2344_), .D(mai_mai_n2342_), .Y(mai_mai_n2347_));
  AOI210     m2298(.A0(mai_mai_n2334_), .A1(x7), .B0(mai_mai_n2347_), .Y(mai_mai_n2348_));
  NA3        m2299(.A(mai_mai_n2348_), .B(mai_mai_n2328_), .C(mai_mai_n2310_), .Y(mai34));
  NA2        m2300(.A(mai_mai_n435_), .B(x4), .Y(mai_mai_n2350_));
  NO2        m2301(.A(mai_mai_n1975_), .B(mai_mai_n863_), .Y(mai_mai_n2351_));
  AOI210     m2302(.A0(mai_mai_n2351_), .A1(mai_mai_n2350_), .B0(mai_mai_n324_), .Y(mai_mai_n2352_));
  NA2        m2303(.A(mai_mai_n290_), .B(mai_mai_n124_), .Y(mai_mai_n2353_));
  NO2        m2304(.A(mai_mai_n981_), .B(mai_mai_n2353_), .Y(mai_mai_n2354_));
  AOI210     m2305(.A0(mai_mai_n2056_), .A1(mai_mai_n546_), .B0(mai_mai_n143_), .Y(mai_mai_n2355_));
  NA2        m2306(.A(mai_mai_n1975_), .B(x0), .Y(mai_mai_n2356_));
  OAI210     m2307(.A0(mai_mai_n1848_), .A1(mai_mai_n985_), .B0(mai_mai_n2356_), .Y(mai_mai_n2357_));
  NO4        m2308(.A(mai_mai_n2357_), .B(mai_mai_n2355_), .C(mai_mai_n2354_), .D(mai_mai_n2352_), .Y(mai_mai_n2358_));
  NO2        m2309(.A(mai_mai_n2358_), .B(mai_mai_n480_), .Y(mai_mai_n2359_));
  NA2        m2310(.A(mai_mai_n740_), .B(x8), .Y(mai_mai_n2360_));
  AO210      m2311(.A0(mai_mai_n2360_), .A1(mai_mai_n490_), .B0(mai_mai_n667_), .Y(mai_mai_n2361_));
  NA2        m2312(.A(mai_mai_n677_), .B(mai_mai_n634_), .Y(mai_mai_n2362_));
  AOI210     m2313(.A0(mai_mai_n2362_), .A1(mai_mai_n2361_), .B0(mai_mai_n269_), .Y(mai_mai_n2363_));
  OAI210     m2314(.A0(mai_mai_n123_), .A1(mai_mai_n1061_), .B0(mai_mai_n1481_), .Y(mai_mai_n2364_));
  OAI210     m2315(.A0(mai_mai_n1622_), .A1(mai_mai_n58_), .B0(mai_mai_n2364_), .Y(mai_mai_n2365_));
  NA3        m2316(.A(mai_mai_n2365_), .B(mai_mai_n344_), .C(x8), .Y(mai_mai_n2366_));
  NO3        m2317(.A(mai_mai_n1002_), .B(mai_mai_n713_), .C(mai_mai_n459_), .Y(mai_mai_n2367_));
  AOI210     m2318(.A0(mai_mai_n1604_), .A1(mai_mai_n332_), .B0(mai_mai_n2367_), .Y(mai_mai_n2368_));
  NA2        m2319(.A(mai_mai_n671_), .B(mai_mai_n324_), .Y(mai_mai_n2369_));
  NA2        m2320(.A(mai_mai_n137_), .B(x0), .Y(mai_mai_n2370_));
  NAi31      m2321(.An(mai_mai_n2370_), .B(mai_mai_n2369_), .C(mai_mai_n804_), .Y(mai_mai_n2371_));
  NA3        m2322(.A(mai_mai_n1617_), .B(mai_mai_n1413_), .C(mai_mai_n50_), .Y(mai_mai_n2372_));
  NA4        m2323(.A(mai_mai_n2372_), .B(mai_mai_n2371_), .C(mai_mai_n2368_), .D(mai_mai_n2366_), .Y(mai_mai_n2373_));
  NA2        m2324(.A(mai_mai_n1120_), .B(mai_mai_n756_), .Y(mai_mai_n2374_));
  NA3        m2325(.A(mai_mai_n1160_), .B(mai_mai_n169_), .C(mai_mai_n1104_), .Y(mai_mai_n2375_));
  AOI210     m2326(.A0(mai_mai_n2375_), .A1(mai_mai_n2374_), .B0(mai_mai_n766_), .Y(mai_mai_n2376_));
  AOI210     m2327(.A0(mai_mai_n1795_), .A1(mai_mai_n133_), .B0(mai_mai_n2376_), .Y(mai_mai_n2377_));
  AOI210     m2328(.A0(mai_mai_n560_), .A1(mai_mai_n821_), .B0(mai_mai_n258_), .Y(mai_mai_n2378_));
  OAI220     m2329(.A0(mai_mai_n2378_), .A1(mai_mai_n59_), .B0(mai_mai_n1131_), .B1(mai_mai_n55_), .Y(mai_mai_n2379_));
  NA3        m2330(.A(mai_mai_n2379_), .B(mai_mai_n740_), .C(mai_mai_n56_), .Y(mai_mai_n2380_));
  OAI210     m2331(.A0(mai_mai_n2377_), .A1(mai_mai_n144_), .B0(mai_mai_n2380_), .Y(mai_mai_n2381_));
  NO4        m2332(.A(mai_mai_n2381_), .B(mai_mai_n2373_), .C(mai_mai_n2363_), .D(mai_mai_n2359_), .Y(mai_mai_n2382_));
  NO2        m2333(.A(mai_mai_n314_), .B(mai_mai_n962_), .Y(mai_mai_n2383_));
  NO3        m2334(.A(mai_mai_n2383_), .B(mai_mai_n447_), .C(mai_mai_n332_), .Y(mai_mai_n2384_));
  NA2        m2335(.A(mai_mai_n789_), .B(mai_mai_n162_), .Y(mai_mai_n2385_));
  NO3        m2336(.A(mai_mai_n2246_), .B(mai_mai_n307_), .C(mai_mai_n1104_), .Y(mai_mai_n2386_));
  OAI220     m2337(.A0(mai_mai_n2386_), .A1(mai_mai_n1574_), .B0(mai_mai_n2385_), .B1(mai_mai_n1186_), .Y(mai_mai_n2387_));
  OAI210     m2338(.A0(mai_mai_n2387_), .A1(mai_mai_n2384_), .B0(x2), .Y(mai_mai_n2388_));
  OAI210     m2339(.A0(mai_mai_n873_), .A1(mai_mai_n375_), .B0(mai_mai_n2388_), .Y(mai_mai_n2389_));
  NA2        m2340(.A(mai_mai_n317_), .B(x4), .Y(mai_mai_n2390_));
  OAI220     m2341(.A0(mai_mai_n752_), .A1(mai_mai_n55_), .B0(mai_mai_n283_), .B1(mai_mai_n107_), .Y(mai_mai_n2391_));
  NO4        m2342(.A(mai_mai_n451_), .B(mai_mai_n77_), .C(x7), .D(x3), .Y(mai_mai_n2392_));
  NO2        m2343(.A(mai_mai_n1120_), .B(mai_mai_n291_), .Y(mai_mai_n2393_));
  NO4        m2344(.A(mai_mai_n2393_), .B(mai_mai_n2392_), .C(mai_mai_n2391_), .D(mai_mai_n2390_), .Y(mai_mai_n2394_));
  NA2        m2345(.A(mai_mai_n1256_), .B(mai_mai_n1059_), .Y(mai_mai_n2395_));
  NA4        m2346(.A(mai_mai_n740_), .B(mai_mai_n181_), .C(mai_mai_n57_), .D(mai_mai_n108_), .Y(mai_mai_n2396_));
  NA3        m2347(.A(mai_mai_n1410_), .B(mai_mai_n261_), .C(x7), .Y(mai_mai_n2397_));
  NA3        m2348(.A(mai_mai_n2397_), .B(mai_mai_n2396_), .C(mai_mai_n2395_), .Y(mai_mai_n2398_));
  OAI210     m2349(.A0(mai_mai_n2398_), .A1(mai_mai_n2394_), .B0(mai_mai_n166_), .Y(mai_mai_n2399_));
  NA3        m2350(.A(mai_mai_n868_), .B(mai_mai_n87_), .C(x0), .Y(mai_mai_n2400_));
  NA4        m2351(.A(mai_mai_n2400_), .B(mai_mai_n1164_), .C(mai_mai_n300_), .D(mai_mai_n591_), .Y(mai_mai_n2401_));
  NA2        m2352(.A(mai_mai_n1168_), .B(mai_mai_n682_), .Y(mai_mai_n2402_));
  OAI210     m2353(.A0(mai_mai_n2402_), .A1(mai_mai_n270_), .B0(mai_mai_n2184_), .Y(mai_mai_n2403_));
  AOI220     m2354(.A0(mai_mai_n2403_), .A1(x7), .B0(mai_mai_n1024_), .B1(mai_mai_n668_), .Y(mai_mai_n2404_));
  OAI210     m2355(.A0(mai_mai_n2069_), .A1(mai_mai_n266_), .B0(mai_mai_n744_), .Y(mai_mai_n2405_));
  AOI220     m2356(.A0(mai_mai_n412_), .A1(x8), .B0(mai_mai_n92_), .B1(x2), .Y(mai_mai_n2406_));
  AOI210     m2357(.A0(mai_mai_n273_), .A1(mai_mai_n53_), .B0(mai_mai_n659_), .Y(mai_mai_n2407_));
  OAI220     m2358(.A0(mai_mai_n2407_), .A1(mai_mai_n97_), .B0(mai_mai_n2406_), .B1(mai_mai_n1357_), .Y(mai_mai_n2408_));
  AOI220     m2359(.A0(mai_mai_n2408_), .A1(mai_mai_n1335_), .B0(mai_mai_n2405_), .B1(mai_mai_n1531_), .Y(mai_mai_n2409_));
  NA4        m2360(.A(mai_mai_n2409_), .B(mai_mai_n2404_), .C(mai_mai_n2401_), .D(mai_mai_n2399_), .Y(mai_mai_n2410_));
  AOI210     m2361(.A0(mai_mai_n2389_), .A1(mai_mai_n821_), .B0(mai_mai_n2410_), .Y(mai_mai_n2411_));
  OAI210     m2362(.A0(mai_mai_n2382_), .A1(x2), .B0(mai_mai_n2411_), .Y(mai35));
  NA2        m2363(.A(mai_mai_n508_), .B(mai_mai_n181_), .Y(mai_mai_n2413_));
  AOI220     m2364(.A0(mai_mai_n642_), .A1(mai_mai_n55_), .B0(mai_mai_n780_), .B1(mai_mai_n1236_), .Y(mai_mai_n2414_));
  AOI210     m2365(.A0(mai_mai_n2414_), .A1(mai_mai_n2413_), .B0(mai_mai_n71_), .Y(mai_mai_n2415_));
  NO3        m2366(.A(mai_mai_n516_), .B(mai_mai_n470_), .C(mai_mai_n343_), .Y(mai_mai_n2416_));
  OAI210     m2367(.A0(mai_mai_n2416_), .A1(mai_mai_n2415_), .B0(x2), .Y(mai_mai_n2417_));
  AOI210     m2368(.A0(mai_mai_n219_), .A1(x0), .B0(mai_mai_n277_), .Y(mai_mai_n2418_));
  OAI220     m2369(.A0(mai_mai_n2418_), .A1(mai_mai_n673_), .B0(mai_mai_n201_), .B1(x4), .Y(mai_mai_n2419_));
  NA2        m2370(.A(mai_mai_n2419_), .B(mai_mai_n141_), .Y(mai_mai_n2420_));
  NA3        m2371(.A(mai_mai_n412_), .B(x8), .C(mai_mai_n71_), .Y(mai_mai_n2421_));
  AOI210     m2372(.A0(mai_mai_n2421_), .A1(mai_mai_n1740_), .B0(mai_mai_n692_), .Y(mai_mai_n2422_));
  OAI210     m2373(.A0(mai_mai_n2335_), .A1(x6), .B0(mai_mai_n755_), .Y(mai_mai_n2423_));
  NO2        m2374(.A(mai_mai_n2423_), .B(mai_mai_n2422_), .Y(mai_mai_n2424_));
  NA3        m2375(.A(mai_mai_n2424_), .B(mai_mai_n2420_), .C(mai_mai_n2417_), .Y(mai_mai_n2425_));
  NAi21      m2376(.An(mai_mai_n1704_), .B(mai_mai_n1311_), .Y(mai_mai_n2426_));
  NA2        m2377(.A(mai_mai_n217_), .B(mai_mai_n578_), .Y(mai_mai_n2427_));
  NO2        m2378(.A(mai_mai_n435_), .B(mai_mai_n428_), .Y(mai_mai_n2428_));
  AOI220     m2379(.A0(mai_mai_n2428_), .A1(mai_mai_n2427_), .B0(mai_mai_n2426_), .B1(mai_mai_n56_), .Y(mai_mai_n2429_));
  NA2        m2380(.A(mai_mai_n769_), .B(mai_mai_n705_), .Y(mai_mai_n2430_));
  NO3        m2381(.A(mai_mai_n687_), .B(mai_mai_n55_), .C(x6), .Y(mai_mai_n2431_));
  OAI210     m2382(.A0(mai_mai_n2431_), .A1(mai_mai_n716_), .B0(mai_mai_n222_), .Y(mai_mai_n2432_));
  NA2        m2383(.A(mai_mai_n1343_), .B(mai_mai_n63_), .Y(mai_mai_n2433_));
  OAI210     m2384(.A0(mai_mai_n1083_), .A1(x6), .B0(mai_mai_n475_), .Y(mai_mai_n2434_));
  NA3        m2385(.A(mai_mai_n2434_), .B(mai_mai_n2433_), .C(mai_mai_n2432_), .Y(mai_mai_n2435_));
  NA3        m2386(.A(mai_mai_n1287_), .B(mai_mai_n758_), .C(x3), .Y(mai_mai_n2436_));
  NO3        m2387(.A(mai_mai_n2436_), .B(mai_mai_n689_), .C(mai_mai_n210_), .Y(mai_mai_n2437_));
  AOI210     m2388(.A0(mai_mai_n2435_), .A1(mai_mai_n50_), .B0(mai_mai_n2437_), .Y(mai_mai_n2438_));
  OAI210     m2389(.A0(mai_mai_n2430_), .A1(mai_mai_n2429_), .B0(mai_mai_n2438_), .Y(mai_mai_n2439_));
  AOI210     m2390(.A0(mai_mai_n2425_), .A1(mai_mai_n57_), .B0(mai_mai_n2439_), .Y(mai_mai_n2440_));
  NA2        m2391(.A(mai_mai_n971_), .B(mai_mai_n63_), .Y(mai_mai_n2441_));
  NO3        m2392(.A(mai_mai_n1083_), .B(mai_mai_n568_), .C(mai_mai_n124_), .Y(mai_mai_n2442_));
  OAI210     m2393(.A0(mai_mai_n159_), .A1(mai_mai_n67_), .B0(mai_mai_n2442_), .Y(mai_mai_n2443_));
  AOI210     m2394(.A0(mai_mai_n2443_), .A1(mai_mai_n2441_), .B0(mai_mai_n50_), .Y(mai_mai_n2444_));
  NA4        m2395(.A(mai_mai_n470_), .B(mai_mai_n234_), .C(mai_mai_n879_), .D(mai_mai_n104_), .Y(mai_mai_n2445_));
  OAI210     m2396(.A0(mai_mai_n971_), .A1(mai_mai_n259_), .B0(mai_mai_n759_), .Y(mai_mai_n2446_));
  OAI210     m2397(.A0(mai_mai_n259_), .A1(mai_mai_n590_), .B0(mai_mai_n2181_), .Y(mai_mai_n2447_));
  NA3        m2398(.A(mai_mai_n2447_), .B(mai_mai_n2446_), .C(mai_mai_n2445_), .Y(mai_mai_n2448_));
  OAI210     m2399(.A0(mai_mai_n2448_), .A1(mai_mai_n2444_), .B0(mai_mai_n59_), .Y(mai_mai_n2449_));
  AOI210     m2400(.A0(mai_mai_n868_), .A1(mai_mai_n537_), .B0(mai_mai_n1922_), .Y(mai_mai_n2450_));
  AOI210     m2401(.A0(mai_mai_n568_), .A1(mai_mai_n612_), .B0(mai_mai_n2450_), .Y(mai_mai_n2451_));
  NO4        m2402(.A(mai_mai_n963_), .B(mai_mai_n568_), .C(mai_mai_n367_), .D(mai_mai_n410_), .Y(mai_mai_n2452_));
  XN2        m2403(.A(x4), .B(x3), .Y(mai_mai_n2453_));
  NO3        m2404(.A(mai_mai_n2453_), .B(mai_mai_n672_), .C(mai_mai_n313_), .Y(mai_mai_n2454_));
  NO3        m2405(.A(mai_mai_n2454_), .B(mai_mai_n2452_), .C(mai_mai_n1477_), .Y(mai_mai_n2455_));
  OAI210     m2406(.A0(mai_mai_n2451_), .A1(x3), .B0(mai_mai_n2455_), .Y(mai_mai_n2456_));
  NO3        m2407(.A(mai_mai_n752_), .B(mai_mai_n870_), .C(mai_mai_n278_), .Y(mai_mai_n2457_));
  OAI210     m2408(.A0(mai_mai_n2457_), .A1(mai_mai_n1477_), .B0(mai_mai_n50_), .Y(mai_mai_n2458_));
  NA3        m2409(.A(mai_mai_n1091_), .B(mai_mai_n819_), .C(mai_mai_n258_), .Y(mai_mai_n2459_));
  NA2        m2410(.A(mai_mai_n2459_), .B(mai_mai_n2458_), .Y(mai_mai_n2460_));
  AOI210     m2411(.A0(mai_mai_n2456_), .A1(mai_mai_n593_), .B0(mai_mai_n2460_), .Y(mai_mai_n2461_));
  AOI210     m2412(.A0(mai_mai_n1447_), .A1(mai_mai_n649_), .B0(mai_mai_n689_), .Y(mai_mai_n2462_));
  NO2        m2413(.A(mai_mai_n879_), .B(mai_mai_n56_), .Y(mai_mai_n2463_));
  OAI210     m2414(.A0(mai_mai_n1978_), .A1(mai_mai_n612_), .B0(mai_mai_n2270_), .Y(mai_mai_n2464_));
  OAI210     m2415(.A0(mai_mai_n2360_), .A1(mai_mai_n2463_), .B0(mai_mai_n2464_), .Y(mai_mai_n2465_));
  OAI210     m2416(.A0(mai_mai_n2465_), .A1(mai_mai_n2462_), .B0(mai_mai_n92_), .Y(mai_mai_n2466_));
  NO2        m2417(.A(mai_mai_n861_), .B(mai_mai_n669_), .Y(mai_mai_n2467_));
  NO2        m2418(.A(mai_mai_n291_), .B(x6), .Y(mai_mai_n2468_));
  OAI210     m2419(.A0(mai_mai_n2467_), .A1(mai_mai_n1803_), .B0(mai_mai_n2468_), .Y(mai_mai_n2469_));
  NA4        m2420(.A(mai_mai_n2469_), .B(mai_mai_n2466_), .C(mai_mai_n2461_), .D(mai_mai_n2449_), .Y(mai_mai_n2470_));
  NA4        m2421(.A(mai_mai_n620_), .B(mai_mai_n692_), .C(mai_mai_n434_), .D(x6), .Y(mai_mai_n2471_));
  AOI210     m2422(.A0(mai_mai_n2471_), .A1(mai_mai_n429_), .B0(x1), .Y(mai_mai_n2472_));
  NO2        m2423(.A(mai_mai_n738_), .B(mai_mai_n689_), .Y(mai_mai_n2473_));
  OAI210     m2424(.A0(mai_mai_n470_), .A1(mai_mai_n170_), .B0(mai_mai_n801_), .Y(mai_mai_n2474_));
  AOI210     m2425(.A0(mai_mai_n2474_), .A1(mai_mai_n1029_), .B0(mai_mai_n53_), .Y(mai_mai_n2475_));
  NO3        m2426(.A(mai_mai_n2475_), .B(mai_mai_n2473_), .C(mai_mai_n2472_), .Y(mai_mai_n2476_));
  NA3        m2427(.A(mai_mai_n1449_), .B(mai_mai_n1288_), .C(mai_mai_n825_), .Y(mai_mai_n2477_));
  AOI220     m2428(.A0(mai_mai_n1965_), .A1(mai_mai_n141_), .B0(mai_mai_n421_), .B1(mai_mai_n128_), .Y(mai_mai_n2478_));
  AOI210     m2429(.A0(mai_mai_n2478_), .A1(mai_mai_n2477_), .B0(mai_mai_n1524_), .Y(mai_mai_n2479_));
  NO2        m2430(.A(mai_mai_n642_), .B(x3), .Y(mai_mai_n2480_));
  NO3        m2431(.A(mai_mai_n700_), .B(mai_mai_n1622_), .C(x2), .Y(mai_mai_n2481_));
  AOI220     m2432(.A0(mai_mai_n2481_), .A1(mai_mai_n2480_), .B0(mai_mai_n1938_), .B1(mai_mai_n776_), .Y(mai_mai_n2482_));
  NA3        m2433(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n2483_));
  OAI220     m2434(.A0(mai_mai_n2483_), .A1(mai_mai_n200_), .B0(mai_mai_n687_), .B1(mai_mai_n533_), .Y(mai_mai_n2484_));
  OAI220     m2435(.A0(mai_mai_n1324_), .A1(x8), .B0(mai_mai_n379_), .B1(mai_mai_n357_), .Y(mai_mai_n2485_));
  AOI220     m2436(.A0(mai_mai_n2485_), .A1(mai_mai_n421_), .B0(mai_mai_n2484_), .B1(mai_mai_n926_), .Y(mai_mai_n2486_));
  OAI210     m2437(.A0(mai_mai_n2482_), .A1(mai_mai_n1177_), .B0(mai_mai_n2486_), .Y(mai_mai_n2487_));
  NO2        m2438(.A(mai_mai_n2487_), .B(mai_mai_n2479_), .Y(mai_mai_n2488_));
  OAI210     m2439(.A0(mai_mai_n2476_), .A1(mai_mai_n317_), .B0(mai_mai_n2488_), .Y(mai_mai_n2489_));
  AOI210     m2440(.A0(mai_mai_n2470_), .A1(x5), .B0(mai_mai_n2489_), .Y(mai_mai_n2490_));
  OAI210     m2441(.A0(mai_mai_n2440_), .A1(x5), .B0(mai_mai_n2490_), .Y(mai36));
  NO2        m2442(.A(mai_mai_n870_), .B(mai_mai_n306_), .Y(mai_mai_n2492_));
  NO3        m2443(.A(mai_mai_n123_), .B(mai_mai_n1061_), .C(mai_mai_n55_), .Y(mai_mai_n2493_));
  NO3        m2444(.A(mai_mai_n2493_), .B(mai_mai_n1997_), .C(mai_mai_n1083_), .Y(mai_mai_n2494_));
  OAI210     m2445(.A0(mai_mai_n2494_), .A1(mai_mai_n2492_), .B0(mai_mai_n110_), .Y(mai_mai_n2495_));
  OR4        m2446(.A(mai_mai_n964_), .B(mai_mai_n812_), .C(mai_mai_n381_), .D(mai_mai_n497_), .Y(mai_mai_n2496_));
  INV        m2447(.A(mai_mai_n1014_), .Y(mai_mai_n2497_));
  OAI210     m2448(.A0(mai_mai_n2232_), .A1(mai_mai_n2497_), .B0(mai_mai_n283_), .Y(mai_mai_n2498_));
  NA3        m2449(.A(mai_mai_n449_), .B(mai_mai_n231_), .C(mai_mai_n122_), .Y(mai_mai_n2499_));
  NA4        m2450(.A(mai_mai_n2499_), .B(mai_mai_n2498_), .C(mai_mai_n2496_), .D(mai_mai_n2495_), .Y(mai_mai_n2500_));
  NO2        m2451(.A(mai_mai_n1003_), .B(x8), .Y(mai_mai_n2501_));
  NO3        m2452(.A(mai_mai_n2501_), .B(mai_mai_n999_), .C(mai_mai_n542_), .Y(mai_mai_n2502_));
  AOI220     m2453(.A0(mai_mai_n307_), .A1(x1), .B0(mai_mai_n140_), .B1(x6), .Y(mai_mai_n2503_));
  AOI210     m2454(.A0(mai_mai_n1104_), .A1(x6), .B0(mai_mai_n425_), .Y(mai_mai_n2504_));
  OAI220     m2455(.A0(mai_mai_n2504_), .A1(mai_mai_n366_), .B0(mai_mai_n2503_), .B1(mai_mai_n471_), .Y(mai_mai_n2505_));
  OAI210     m2456(.A0(mai_mai_n2505_), .A1(mai_mai_n2502_), .B0(mai_mai_n470_), .Y(mai_mai_n2506_));
  NA2        m2457(.A(mai_mai_n677_), .B(mai_mai_n497_), .Y(mai_mai_n2507_));
  AOI210     m2458(.A0(mai_mai_n2507_), .A1(mai_mai_n656_), .B0(mai_mai_n270_), .Y(mai_mai_n2508_));
  NO3        m2459(.A(mai_mai_n1895_), .B(mai_mai_n1621_), .C(mai_mai_n279_), .Y(mai_mai_n2509_));
  NO2        m2460(.A(mai_mai_n2441_), .B(mai_mai_n233_), .Y(mai_mai_n2510_));
  NO4        m2461(.A(mai_mai_n2510_), .B(mai_mai_n2509_), .C(mai_mai_n2508_), .D(mai_mai_n423_), .Y(mai_mai_n2511_));
  OAI210     m2462(.A0(mai_mai_n644_), .A1(mai_mai_n811_), .B0(mai_mai_n989_), .Y(mai_mai_n2512_));
  OAI220     m2463(.A0(mai_mai_n1668_), .A1(mai_mai_n1663_), .B0(mai_mai_n989_), .B1(mai_mai_n1104_), .Y(mai_mai_n2513_));
  AOI220     m2464(.A0(mai_mai_n2513_), .A1(mai_mai_n121_), .B0(mai_mai_n2512_), .B1(mai_mai_n634_), .Y(mai_mai_n2514_));
  NA3        m2465(.A(mai_mai_n2514_), .B(mai_mai_n2511_), .C(mai_mai_n2506_), .Y(mai_mai_n2515_));
  AOI210     m2466(.A0(mai_mai_n2500_), .A1(mai_mai_n344_), .B0(mai_mai_n2515_), .Y(mai_mai_n2516_));
  OAI210     m2467(.A0(mai_mai_n598_), .A1(mai_mai_n521_), .B0(mai_mai_n170_), .Y(mai_mai_n2517_));
  OAI210     m2468(.A0(mai_mai_n2012_), .A1(mai_mai_n70_), .B0(mai_mai_n2517_), .Y(mai_mai_n2518_));
  OAI210     m2469(.A0(mai_mai_n500_), .A1(mai_mai_n242_), .B0(mai_mai_n259_), .Y(mai_mai_n2519_));
  NO2        m2470(.A(mai_mai_n2021_), .B(mai_mai_n177_), .Y(mai_mai_n2520_));
  NA2        m2471(.A(mai_mai_n1223_), .B(mai_mai_n55_), .Y(mai_mai_n2521_));
  OAI210     m2472(.A0(mai_mai_n2521_), .A1(mai_mai_n2520_), .B0(mai_mai_n2519_), .Y(mai_mai_n2522_));
  OAI210     m2473(.A0(mai_mai_n2522_), .A1(mai_mai_n2518_), .B0(mai_mai_n904_), .Y(mai_mai_n2523_));
  AOI210     m2474(.A0(mai_mai_n107_), .A1(mai_mai_n110_), .B0(mai_mai_n346_), .Y(mai_mai_n2524_));
  NA2        m2475(.A(mai_mai_n677_), .B(mai_mai_n1622_), .Y(mai_mai_n2525_));
  OAI220     m2476(.A0(mai_mai_n2525_), .A1(mai_mai_n2524_), .B0(mai_mai_n755_), .B1(mai_mai_n1270_), .Y(mai_mai_n2526_));
  NO2        m2477(.A(mai_mai_n1413_), .B(mai_mai_n584_), .Y(mai_mai_n2527_));
  NO3        m2478(.A(mai_mai_n2527_), .B(mai_mai_n1811_), .C(mai_mai_n700_), .Y(mai_mai_n2528_));
  NOi31      m2479(.An(mai_mai_n2033_), .B(mai_mai_n2324_), .C(mai_mai_n765_), .Y(mai_mai_n2529_));
  NO3        m2480(.A(mai_mai_n2529_), .B(mai_mai_n2528_), .C(mai_mai_n2526_), .Y(mai_mai_n2530_));
  AOI210     m2481(.A0(mai_mai_n2530_), .A1(mai_mai_n2523_), .B0(x7), .Y(mai_mai_n2531_));
  AOI210     m2482(.A0(mai_mai_n593_), .A1(mai_mai_n629_), .B0(mai_mai_n1202_), .Y(mai_mai_n2532_));
  NA3        m2483(.A(mai_mai_n2532_), .B(mai_mai_n1002_), .C(mai_mai_n897_), .Y(mai_mai_n2533_));
  NA2        m2484(.A(mai_mai_n2533_), .B(mai_mai_n508_), .Y(mai_mai_n2534_));
  AOI220     m2485(.A0(mai_mai_n1764_), .A1(mai_mai_n262_), .B0(mai_mai_n1059_), .B1(mai_mai_n128_), .Y(mai_mai_n2535_));
  NO2        m2486(.A(mai_mai_n2535_), .B(mai_mai_n449_), .Y(mai_mai_n2536_));
  NO2        m2487(.A(mai_mai_n410_), .B(mai_mai_n231_), .Y(mai_mai_n2537_));
  NO3        m2488(.A(mai_mai_n2537_), .B(mai_mai_n1292_), .C(mai_mai_n59_), .Y(mai_mai_n2538_));
  AOI210     m2489(.A0(mai_mai_n1240_), .A1(mai_mai_n411_), .B0(x6), .Y(mai_mai_n2539_));
  NA3        m2490(.A(mai_mai_n1695_), .B(mai_mai_n283_), .C(mai_mai_n273_), .Y(mai_mai_n2540_));
  NA2        m2491(.A(mai_mai_n2540_), .B(mai_mai_n1648_), .Y(mai_mai_n2541_));
  NO4        m2492(.A(mai_mai_n2541_), .B(mai_mai_n2539_), .C(mai_mai_n2538_), .D(mai_mai_n2536_), .Y(mai_mai_n2542_));
  AOI210     m2493(.A0(mai_mai_n2542_), .A1(mai_mai_n2534_), .B0(mai_mai_n459_), .Y(mai_mai_n2543_));
  NO3        m2494(.A(mai_mai_n2453_), .B(mai_mai_n910_), .C(mai_mai_n507_), .Y(mai_mai_n2544_));
  AOI210     m2495(.A0(mai_mai_n1290_), .A1(mai_mai_n272_), .B0(mai_mai_n2544_), .Y(mai_mai_n2545_));
  OAI210     m2496(.A0(mai_mai_n877_), .A1(mai_mai_n278_), .B0(mai_mai_n400_), .Y(mai_mai_n2546_));
  NA2        m2497(.A(mai_mai_n1223_), .B(mai_mai_n175_), .Y(mai_mai_n2547_));
  NO2        m2498(.A(mai_mai_n619_), .B(mai_mai_n110_), .Y(mai_mai_n2548_));
  AO210      m2499(.A0(mai_mai_n2548_), .A1(mai_mai_n2547_), .B0(mai_mai_n1781_), .Y(mai_mai_n2549_));
  NO2        m2500(.A(mai_mai_n466_), .B(mai_mai_n422_), .Y(mai_mai_n2550_));
  AOI220     m2501(.A0(mai_mai_n2550_), .A1(mai_mai_n2549_), .B0(mai_mai_n2546_), .B1(mai_mai_n298_), .Y(mai_mai_n2551_));
  OAI210     m2502(.A0(mai_mai_n2545_), .A1(x1), .B0(mai_mai_n2551_), .Y(mai_mai_n2552_));
  NO3        m2503(.A(mai_mai_n2552_), .B(mai_mai_n2543_), .C(mai_mai_n2531_), .Y(mai_mai_n2553_));
  OAI210     m2504(.A0(mai_mai_n2516_), .A1(mai_mai_n57_), .B0(mai_mai_n2553_), .Y(mai37));
  NA3        m2505(.A(mai_mai_n1080_), .B(mai_mai_n143_), .C(x3), .Y(mai_mai_n2555_));
  NA3        m2506(.A(mai_mai_n789_), .B(mai_mai_n162_), .C(mai_mai_n50_), .Y(mai_mai_n2556_));
  AOI210     m2507(.A0(mai_mai_n2556_), .A1(mai_mai_n2555_), .B0(mai_mai_n693_), .Y(mai_mai_n2557_));
  NO3        m2508(.A(mai_mai_n1080_), .B(mai_mai_n381_), .C(mai_mai_n515_), .Y(mai_mai_n2558_));
  OAI210     m2509(.A0(mai_mai_n2558_), .A1(mai_mai_n2557_), .B0(mai_mai_n56_), .Y(mai_mai_n2559_));
  NA2        m2510(.A(mai_mai_n607_), .B(mai_mai_n756_), .Y(mai_mai_n2560_));
  AOI210     m2511(.A0(mai_mai_n2560_), .A1(mai_mai_n1060_), .B0(x3), .Y(mai_mai_n2561_));
  AOI220     m2512(.A0(mai_mai_n607_), .A1(mai_mai_n756_), .B0(mai_mai_n470_), .B1(mai_mai_n1059_), .Y(mai_mai_n2562_));
  NO2        m2513(.A(mai_mai_n672_), .B(mai_mai_n184_), .Y(mai_mai_n2563_));
  OAI220     m2514(.A0(mai_mai_n2563_), .A1(mai_mai_n846_), .B0(mai_mai_n2562_), .B1(mai_mai_n110_), .Y(mai_mai_n2564_));
  OAI210     m2515(.A0(mai_mai_n2564_), .A1(mai_mai_n2561_), .B0(mai_mai_n71_), .Y(mai_mai_n2565_));
  NA2        m2516(.A(mai_mai_n1204_), .B(mai_mai_n1083_), .Y(mai_mai_n2566_));
  OAI210     m2517(.A0(mai_mai_n1225_), .A1(mai_mai_n194_), .B0(mai_mai_n460_), .Y(mai_mai_n2567_));
  NA4        m2518(.A(mai_mai_n2567_), .B(mai_mai_n2566_), .C(mai_mai_n2565_), .D(mai_mai_n2559_), .Y(mai_mai_n2568_));
  NA2        m2519(.A(mai_mai_n428_), .B(mai_mai_n140_), .Y(mai_mai_n2569_));
  NO2        m2520(.A(mai_mai_n1726_), .B(mai_mai_n109_), .Y(mai_mai_n2570_));
  AOI210     m2521(.A0(mai_mai_n1999_), .A1(mai_mai_n871_), .B0(mai_mai_n2570_), .Y(mai_mai_n2571_));
  OAI220     m2522(.A0(mai_mai_n2571_), .A1(mai_mai_n51_), .B0(mai_mai_n1623_), .B1(mai_mai_n2569_), .Y(mai_mai_n2572_));
  AOI210     m2523(.A0(mai_mai_n2568_), .A1(mai_mai_n68_), .B0(mai_mai_n2572_), .Y(mai_mai_n2573_));
  OAI210     m2524(.A0(mai_mai_n273_), .A1(mai_mai_n1108_), .B0(mai_mai_n491_), .Y(mai_mai_n2574_));
  NA3        m2525(.A(mai_mai_n2574_), .B(mai_mai_n270_), .C(mai_mai_n1061_), .Y(mai_mai_n2575_));
  OAI210     m2526(.A0(mai_mai_n234_), .A1(mai_mai_n222_), .B0(mai_mai_n1740_), .Y(mai_mai_n2576_));
  NA2        m2527(.A(mai_mai_n352_), .B(mai_mai_n277_), .Y(mai_mai_n2577_));
  NA3        m2528(.A(mai_mai_n406_), .B(mai_mai_n825_), .C(mai_mai_n110_), .Y(mai_mai_n2578_));
  NO2        m2529(.A(mai_mai_n534_), .B(mai_mai_n56_), .Y(mai_mai_n2579_));
  NA3        m2530(.A(mai_mai_n2579_), .B(mai_mai_n2578_), .C(mai_mai_n2577_), .Y(mai_mai_n2580_));
  AOI210     m2531(.A0(mai_mai_n2576_), .A1(mai_mai_n515_), .B0(mai_mai_n2580_), .Y(mai_mai_n2581_));
  NO2        m2532(.A(mai_mai_n1195_), .B(mai_mai_n278_), .Y(mai_mai_n2582_));
  OAI210     m2533(.A0(mai_mai_n298_), .A1(mai_mai_n268_), .B0(mai_mai_n2582_), .Y(mai_mai_n2583_));
  OAI210     m2534(.A0(mai_mai_n674_), .A1(mai_mai_n141_), .B0(x3), .Y(mai_mai_n2584_));
  AOI210     m2535(.A0(mai_mai_n674_), .A1(mai_mai_n371_), .B0(mai_mai_n2584_), .Y(mai_mai_n2585_));
  AOI210     m2536(.A0(mai_mai_n1622_), .A1(mai_mai_n50_), .B0(mai_mai_n352_), .Y(mai_mai_n2586_));
  OAI210     m2537(.A0(mai_mai_n2586_), .A1(mai_mai_n405_), .B0(mai_mai_n56_), .Y(mai_mai_n2587_));
  NO2        m2538(.A(mai_mai_n2587_), .B(mai_mai_n2585_), .Y(mai_mai_n2588_));
  AOI220     m2539(.A0(mai_mai_n2588_), .A1(mai_mai_n2583_), .B0(mai_mai_n2581_), .B1(mai_mai_n2575_), .Y(mai_mai_n2589_));
  OAI210     m2540(.A0(mai_mai_n2589_), .A1(mai_mai_n1779_), .B0(mai_mai_n102_), .Y(mai_mai_n2590_));
  NA2        m2541(.A(mai_mai_n700_), .B(mai_mai_n1209_), .Y(mai_mai_n2591_));
  NOi21      m2542(.An(mai_mai_n1377_), .B(mai_mai_n111_), .Y(mai_mai_n2592_));
  AOI210     m2543(.A0(mai_mai_n2592_), .A1(mai_mai_n2591_), .B0(mai_mai_n438_), .Y(mai_mai_n2593_));
  NO2        m2544(.A(mai_mai_n2243_), .B(mai_mai_n55_), .Y(mai_mai_n2594_));
  OAI210     m2545(.A0(mai_mai_n2594_), .A1(mai_mai_n2593_), .B0(mai_mai_n1840_), .Y(mai_mai_n2595_));
  NA2        m2546(.A(mai_mai_n181_), .B(mai_mai_n108_), .Y(mai_mai_n2596_));
  NA2        m2547(.A(mai_mai_n692_), .B(x6), .Y(mai_mai_n2597_));
  AOI210     m2548(.A0(mai_mai_n2597_), .A1(mai_mai_n490_), .B0(mai_mai_n2596_), .Y(mai_mai_n2598_));
  AOI210     m2549(.A0(mai_mai_n359_), .A1(mai_mai_n143_), .B0(mai_mai_n144_), .Y(mai_mai_n2599_));
  OAI210     m2550(.A0(mai_mai_n2599_), .A1(mai_mai_n2598_), .B0(mai_mai_n352_), .Y(mai_mai_n2600_));
  AOI210     m2551(.A0(mai_mai_n620_), .A1(mai_mai_n438_), .B0(mai_mai_n1300_), .Y(mai_mai_n2601_));
  NO3        m2552(.A(mai_mai_n2601_), .B(mai_mai_n270_), .C(mai_mai_n63_), .Y(mai_mai_n2602_));
  OAI220     m2553(.A0(mai_mai_n2360_), .A1(mai_mai_n488_), .B0(mai_mai_n2115_), .B1(mai_mai_n389_), .Y(mai_mai_n2603_));
  OAI210     m2554(.A0(mai_mai_n2603_), .A1(mai_mai_n2602_), .B0(mai_mai_n53_), .Y(mai_mai_n2604_));
  NO4        m2555(.A(mai_mai_n2370_), .B(mai_mai_n942_), .C(mai_mai_n439_), .D(mai_mai_n225_), .Y(mai_mai_n2605_));
  NO4        m2556(.A(mai_mai_n740_), .B(mai_mai_n608_), .C(mai_mai_n447_), .D(mai_mai_n1069_), .Y(mai_mai_n2606_));
  NO3        m2557(.A(mai_mai_n2606_), .B(mai_mai_n2605_), .C(mai_mai_n1075_), .Y(mai_mai_n2607_));
  NA4        m2558(.A(mai_mai_n2607_), .B(mai_mai_n2604_), .C(mai_mai_n2600_), .D(mai_mai_n2595_), .Y(mai_mai_n2608_));
  NO3        m2559(.A(mai_mai_n254_), .B(mai_mai_n358_), .C(mai_mai_n84_), .Y(mai_mai_n2609_));
  NO2        m2560(.A(mai_mai_n281_), .B(mai_mai_n780_), .Y(mai_mai_n2610_));
  NO3        m2561(.A(mai_mai_n2610_), .B(mai_mai_n1223_), .C(mai_mai_n1242_), .Y(mai_mai_n2611_));
  OAI220     m2562(.A0(mai_mai_n2611_), .A1(mai_mai_n2609_), .B0(mai_mai_n470_), .B1(mai_mai_n85_), .Y(mai_mai_n2612_));
  OR2        m2563(.A(mai_mai_n948_), .B(mai_mai_n758_), .Y(mai_mai_n2613_));
  NA2        m2564(.A(mai_mai_n1236_), .B(mai_mai_n55_), .Y(mai_mai_n2614_));
  NOi21      m2565(.An(mai_mai_n2614_), .B(mai_mai_n390_), .Y(mai_mai_n2615_));
  AOI210     m2566(.A0(mai_mai_n2615_), .A1(mai_mai_n2613_), .B0(x1), .Y(mai_mai_n2616_));
  NA2        m2567(.A(mai_mai_n269_), .B(mai_mai_n84_), .Y(mai_mai_n2617_));
  AOI210     m2568(.A0(mai_mai_n1574_), .A1(mai_mai_n405_), .B0(mai_mai_n2617_), .Y(mai_mai_n2618_));
  NA2        m2569(.A(mai_mai_n1120_), .B(mai_mai_n62_), .Y(mai_mai_n2619_));
  NA2        m2570(.A(mai_mai_n1168_), .B(mai_mai_n177_), .Y(mai_mai_n2620_));
  OAI210     m2571(.A0(mai_mai_n2619_), .A1(mai_mai_n316_), .B0(mai_mai_n2620_), .Y(mai_mai_n2621_));
  NO3        m2572(.A(mai_mai_n2621_), .B(mai_mai_n2618_), .C(mai_mai_n2616_), .Y(mai_mai_n2622_));
  OAI210     m2573(.A0(mai_mai_n2622_), .A1(x6), .B0(mai_mai_n2612_), .Y(mai_mai_n2623_));
  AOI220     m2574(.A0(mai_mai_n2623_), .A1(mai_mai_n1481_), .B0(mai_mai_n2608_), .B1(mai_mai_n57_), .Y(mai_mai_n2624_));
  NA3        m2575(.A(mai_mai_n2624_), .B(mai_mai_n2590_), .C(mai_mai_n2573_), .Y(mai38));
  AOI210     m2576(.A0(mai_mai_n1680_), .A1(mai_mai_n190_), .B0(mai_mai_n983_), .Y(mai_mai_n2626_));
  AOI210     m2577(.A0(mai_mai_n1240_), .A1(mai_mai_n583_), .B0(mai_mai_n1101_), .Y(mai_mai_n2627_));
  AOI210     m2578(.A0(mai_mai_n2614_), .A1(mai_mai_n1871_), .B0(mai_mai_n233_), .Y(mai_mai_n2628_));
  NO3        m2579(.A(mai_mai_n2628_), .B(mai_mai_n2627_), .C(mai_mai_n2626_), .Y(mai_mai_n2629_));
  NO2        m2580(.A(mai_mai_n2629_), .B(x6), .Y(mai_mai_n2630_));
  NA4        m2581(.A(mai_mai_n383_), .B(mai_mai_n261_), .C(mai_mai_n193_), .D(x8), .Y(mai_mai_n2631_));
  NA2        m2582(.A(mai_mai_n404_), .B(mai_mai_n108_), .Y(mai_mai_n2632_));
  AOI210     m2583(.A0(mai_mai_n2632_), .A1(mai_mai_n2631_), .B0(mai_mai_n144_), .Y(mai_mai_n2633_));
  AOI210     m2584(.A0(mai_mai_n439_), .A1(mai_mai_n409_), .B0(mai_mai_n1750_), .Y(mai_mai_n2634_));
  NO2        m2585(.A(mai_mai_n819_), .B(mai_mai_n92_), .Y(mai_mai_n2635_));
  OAI210     m2586(.A0(mai_mai_n1033_), .A1(mai_mai_n150_), .B0(mai_mai_n365_), .Y(mai_mai_n2636_));
  OAI220     m2587(.A0(mai_mai_n2636_), .A1(mai_mai_n2635_), .B0(mai_mai_n2634_), .B1(mai_mai_n193_), .Y(mai_mai_n2637_));
  OAI210     m2588(.A0(mai_mai_n2637_), .A1(mai_mai_n2633_), .B0(x6), .Y(mai_mai_n2638_));
  NO2        m2589(.A(mai_mai_n251_), .B(mai_mai_n780_), .Y(mai_mai_n2639_));
  NO3        m2590(.A(mai_mai_n2639_), .B(mai_mai_n1704_), .C(mai_mai_n261_), .Y(mai_mai_n2640_));
  NO3        m2591(.A(x3), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n2641_));
  OAI210     m2592(.A0(mai_mai_n527_), .A1(x2), .B0(mai_mai_n2641_), .Y(mai_mai_n2642_));
  NA3        m2593(.A(mai_mai_n438_), .B(mai_mai_n428_), .C(mai_mai_n297_), .Y(mai_mai_n2643_));
  NA3        m2594(.A(mai_mai_n2643_), .B(mai_mai_n2642_), .C(mai_mai_n1830_), .Y(mai_mai_n2644_));
  OAI210     m2595(.A0(mai_mai_n2644_), .A1(mai_mai_n2640_), .B0(mai_mai_n821_), .Y(mai_mai_n2645_));
  NO2        m2596(.A(mai_mai_n608_), .B(mai_mai_n279_), .Y(mai_mai_n2646_));
  AN3        m2597(.A(mai_mai_n826_), .B(mai_mai_n789_), .C(x0), .Y(mai_mai_n2647_));
  OAI210     m2598(.A0(mai_mai_n2647_), .A1(mai_mai_n2646_), .B0(mai_mai_n333_), .Y(mai_mai_n2648_));
  OAI220     m2599(.A0(mai_mai_n608_), .A1(mai_mai_n279_), .B0(mai_mai_n825_), .B1(mai_mai_n93_), .Y(mai_mai_n2649_));
  OAI210     m2600(.A0(mai_mai_n692_), .A1(x0), .B0(mai_mai_n51_), .Y(mai_mai_n2650_));
  AOI210     m2601(.A0(mai_mai_n589_), .A1(x4), .B0(mai_mai_n232_), .Y(mai_mai_n2651_));
  AOI220     m2602(.A0(mai_mai_n2651_), .A1(mai_mai_n2650_), .B0(mai_mai_n2649_), .B1(mai_mai_n406_), .Y(mai_mai_n2652_));
  NA4        m2603(.A(mai_mai_n2652_), .B(mai_mai_n2648_), .C(mai_mai_n2645_), .D(mai_mai_n2638_), .Y(mai_mai_n2653_));
  OAI210     m2604(.A0(mai_mai_n2653_), .A1(mai_mai_n2630_), .B0(x7), .Y(mai_mai_n2654_));
  AOI210     m2605(.A0(mai_mai_n380_), .A1(x1), .B0(mai_mai_n1248_), .Y(mai_mai_n2655_));
  NO2        m2606(.A(mai_mai_n2655_), .B(mai_mai_n51_), .Y(mai_mai_n2656_));
  AOI210     m2607(.A0(mai_mai_n92_), .A1(mai_mai_n71_), .B0(mai_mai_n2270_), .Y(mai_mai_n2657_));
  NA2        m2608(.A(mai_mai_n389_), .B(x3), .Y(mai_mai_n2658_));
  NO2        m2609(.A(mai_mai_n1771_), .B(mai_mai_n534_), .Y(mai_mai_n2659_));
  OAI210     m2610(.A0(mai_mai_n2658_), .A1(mai_mai_n2657_), .B0(mai_mai_n2659_), .Y(mai_mai_n2660_));
  OAI210     m2611(.A0(mai_mai_n2660_), .A1(mai_mai_n2656_), .B0(x4), .Y(mai_mai_n2661_));
  NO2        m2612(.A(mai_mai_n1782_), .B(mai_mai_n464_), .Y(mai_mai_n2662_));
  NO3        m2613(.A(mai_mai_n2662_), .B(mai_mai_n405_), .C(mai_mai_n121_), .Y(mai_mai_n2663_));
  AOI210     m2614(.A0(mai_mai_n1069_), .A1(mai_mai_n245_), .B0(mai_mai_n398_), .Y(mai_mai_n2664_));
  AO210      m2615(.A0(mai_mai_n1316_), .A1(x6), .B0(mai_mai_n2664_), .Y(mai_mai_n2665_));
  NO2        m2616(.A(mai_mai_n1434_), .B(mai_mai_n141_), .Y(mai_mai_n2666_));
  NA2        m2617(.A(mai_mai_n1975_), .B(mai_mai_n327_), .Y(mai_mai_n2667_));
  OAI220     m2618(.A0(mai_mai_n2667_), .A1(mai_mai_n1088_), .B0(mai_mai_n2666_), .B1(mai_mai_n1853_), .Y(mai_mai_n2668_));
  NO3        m2619(.A(mai_mai_n2668_), .B(mai_mai_n2665_), .C(mai_mai_n2663_), .Y(mai_mai_n2669_));
  AOI210     m2620(.A0(mai_mai_n2669_), .A1(mai_mai_n2661_), .B0(mai_mai_n108_), .Y(mai_mai_n2670_));
  NA3        m2621(.A(mai_mai_n1965_), .B(mai_mai_n608_), .C(mai_mai_n166_), .Y(mai_mai_n2671_));
  AOI210     m2622(.A0(mai_mai_n2671_), .A1(mai_mai_n1443_), .B0(mai_mai_n234_), .Y(mai_mai_n2672_));
  AOI210     m2623(.A0(mai_mai_n508_), .A1(mai_mai_n497_), .B0(mai_mai_n688_), .Y(mai_mai_n2673_));
  OAI220     m2624(.A0(mai_mai_n2673_), .A1(mai_mai_n471_), .B0(mai_mai_n201_), .B1(mai_mai_n119_), .Y(mai_mai_n2674_));
  OAI210     m2625(.A0(mai_mai_n2674_), .A1(mai_mai_n2672_), .B0(x0), .Y(mai_mai_n2675_));
  NA3        m2626(.A(mai_mai_n409_), .B(mai_mai_n825_), .C(mai_mai_n279_), .Y(mai_mai_n2676_));
  AOI210     m2627(.A0(mai_mai_n2676_), .A1(mai_mai_n724_), .B0(mai_mai_n2227_), .Y(mai_mai_n2677_));
  NA2        m2628(.A(mai_mai_n1140_), .B(mai_mai_n962_), .Y(mai_mai_n2678_));
  NA4        m2629(.A(mai_mai_n687_), .B(mai_mai_n608_), .C(mai_mai_n181_), .D(x3), .Y(mai_mai_n2679_));
  AOI210     m2630(.A0(mai_mai_n2679_), .A1(mai_mai_n2678_), .B0(mai_mai_n502_), .Y(mai_mai_n2680_));
  NO4        m2631(.A(mai_mai_n1427_), .B(mai_mai_n523_), .C(mai_mai_n1242_), .D(mai_mai_n780_), .Y(mai_mai_n2681_));
  OAI220     m2632(.A0(mai_mai_n1801_), .A1(mai_mai_n2314_), .B0(mai_mai_n232_), .B1(mai_mai_n152_), .Y(mai_mai_n2682_));
  NO4        m2633(.A(mai_mai_n2682_), .B(mai_mai_n2681_), .C(mai_mai_n2680_), .D(mai_mai_n2677_), .Y(mai_mai_n2683_));
  NA2        m2634(.A(mai_mai_n2683_), .B(mai_mai_n2675_), .Y(mai_mai_n2684_));
  OAI210     m2635(.A0(mai_mai_n2684_), .A1(mai_mai_n2670_), .B0(mai_mai_n57_), .Y(mai_mai_n2685_));
  NO2        m2636(.A(mai_mai_n1841_), .B(mai_mai_n689_), .Y(mai_mai_n2686_));
  OAI210     m2637(.A0(mai_mai_n1778_), .A1(mai_mai_n217_), .B0(mai_mai_n499_), .Y(mai_mai_n2687_));
  OAI210     m2638(.A0(mai_mai_n2687_), .A1(mai_mai_n2686_), .B0(mai_mai_n636_), .Y(mai_mai_n2688_));
  OAI220     m2639(.A0(mai_mai_n1785_), .A1(mai_mai_n279_), .B0(mai_mai_n260_), .B1(mai_mai_n104_), .Y(mai_mai_n2689_));
  NA2        m2640(.A(mai_mai_n1889_), .B(mai_mai_n360_), .Y(mai_mai_n2690_));
  OAI220     m2641(.A0(mai_mai_n2690_), .A1(mai_mai_n644_), .B0(mai_mai_n699_), .B1(mai_mai_n152_), .Y(mai_mai_n2691_));
  AOI210     m2642(.A0(mai_mai_n2689_), .A1(mai_mai_n1003_), .B0(mai_mai_n2691_), .Y(mai_mai_n2692_));
  NA4        m2643(.A(mai_mai_n2692_), .B(mai_mai_n2688_), .C(mai_mai_n2685_), .D(mai_mai_n2654_), .Y(mai39));
  INV        m2644(.A(mai_mai_n498_), .Y(mai_mai_n2696_));
  INV        u0000(.A(x3), .Y(men_men_n50_));
  NA2        u0001(.A(men_men_n50_), .B(x2), .Y(men_men_n51_));
  NA2        u0002(.A(x7), .B(x0), .Y(men_men_n52_));
  INV        u0003(.A(x1), .Y(men_men_n53_));
  NA2        u0004(.A(x5), .B(men_men_n53_), .Y(men_men_n54_));
  INV        u0005(.A(x8), .Y(men_men_n55_));
  INV        u0006(.A(x4), .Y(men_men_n56_));
  INV        u0007(.A(x7), .Y(men_men_n57_));
  NA2        u0008(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0009(.A(x0), .Y(men_men_n59_));
  NA2        u0010(.A(x4), .B(men_men_n59_), .Y(men_men_n60_));
  NA4        u0011(.A(men_men_n60_), .B(men_men_n58_), .C(men_men_n55_), .D(x6), .Y(men_men_n61_));
  NA2        u0012(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n62_));
  NO2        u0013(.A(men_men_n55_), .B(x6), .Y(men_men_n63_));
  NA2        u0014(.A(men_men_n57_), .B(x4), .Y(men_men_n64_));
  NA3        u0015(.A(men_men_n64_), .B(men_men_n63_), .C(men_men_n62_), .Y(men_men_n65_));
  AOI210     u0016(.A0(men_men_n65_), .A1(men_men_n61_), .B0(men_men_n54_), .Y(men_men_n66_));
  NO2        u0017(.A(x8), .B(men_men_n57_), .Y(men_men_n67_));
  NO2        u0018(.A(x7), .B(men_men_n59_), .Y(men_men_n68_));
  NO2        u0019(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi21      u0020(.An(x5), .B(x1), .Y(men_men_n70_));
  INV        u0021(.A(x6), .Y(men_men_n71_));
  NA2        u0022(.A(men_men_n71_), .B(x4), .Y(men_men_n72_));
  NO3        u0023(.A(men_men_n72_), .B(men_men_n70_), .C(men_men_n69_), .Y(men_men_n73_));
  OAI210     u0024(.A0(men_men_n73_), .A1(men_men_n66_), .B0(men_men_n52_), .Y(men_men_n74_));
  NA2        u0025(.A(x7), .B(x4), .Y(men_men_n75_));
  NO2        u0026(.A(men_men_n75_), .B(x1), .Y(men_men_n76_));
  NO2        u0027(.A(men_men_n71_), .B(x5), .Y(men_men_n77_));
  NO2        u0028(.A(x8), .B(men_men_n59_), .Y(men_men_n78_));
  NA3        u0029(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n76_), .Y(men_men_n79_));
  AOI210     u0030(.A0(men_men_n79_), .A1(men_men_n74_), .B0(men_men_n51_), .Y(men_men_n80_));
  NA2        u0031(.A(x5), .B(x3), .Y(men_men_n81_));
  NO2        u0032(.A(x6), .B(x0), .Y(men_men_n82_));
  NO2        u0033(.A(men_men_n82_), .B(x4), .Y(men_men_n83_));
  NO2        u0034(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u0035(.A(men_men_n71_), .B(men_men_n59_), .Y(men_men_n85_));
  NO2        u0036(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n86_));
  NA2        u0037(.A(x8), .B(x1), .Y(men_men_n87_));
  NO2        u0038(.A(men_men_n87_), .B(x7), .Y(men_men_n88_));
  INV        u0039(.A(men_men_n88_), .Y(men_men_n89_));
  OR3        u0040(.A(men_men_n89_), .B(men_men_n86_), .C(men_men_n83_), .Y(men_men_n90_));
  NO3        u0041(.A(x8), .B(men_men_n57_), .C(x6), .Y(men_men_n91_));
  NO2        u0042(.A(x1), .B(men_men_n59_), .Y(men_men_n92_));
  NO2        u0043(.A(men_men_n56_), .B(x2), .Y(men_men_n93_));
  NA3        u0044(.A(men_men_n93_), .B(men_men_n92_), .C(men_men_n91_), .Y(men_men_n94_));
  AOI210     u0045(.A0(men_men_n94_), .A1(men_men_n90_), .B0(men_men_n81_), .Y(men_men_n95_));
  XO2        u0046(.A(x7), .B(x1), .Y(men_men_n96_));
  INV        u0047(.A(men_men_n96_), .Y(men_men_n97_));
  NO2        u0048(.A(men_men_n97_), .B(x6), .Y(men_men_n98_));
  NO2        u0049(.A(men_men_n50_), .B(x0), .Y(men_men_n99_));
  NA2        u0050(.A(men_men_n99_), .B(men_men_n55_), .Y(men_men_n100_));
  NO2        u0051(.A(x6), .B(x5), .Y(men_men_n101_));
  NO2        u0052(.A(men_men_n57_), .B(x5), .Y(men_men_n102_));
  NO2        u0053(.A(men_men_n102_), .B(men_men_n101_), .Y(men_men_n103_));
  NA2        u0054(.A(x6), .B(x1), .Y(men_men_n104_));
  NA2        u0055(.A(men_men_n104_), .B(men_men_n84_), .Y(men_men_n105_));
  NO4        u0056(.A(men_men_n105_), .B(men_men_n103_), .C(men_men_n100_), .D(men_men_n98_), .Y(men_men_n106_));
  NA2        u0057(.A(x3), .B(x0), .Y(men_men_n107_));
  INV        u0058(.A(x5), .Y(men_men_n108_));
  NA2        u0059(.A(men_men_n71_), .B(men_men_n108_), .Y(men_men_n109_));
  INV        u0060(.A(x2), .Y(men_men_n110_));
  NO2        u0061(.A(men_men_n56_), .B(men_men_n110_), .Y(men_men_n111_));
  NA2        u0062(.A(men_men_n57_), .B(men_men_n108_), .Y(men_men_n112_));
  NA3        u0063(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n109_), .Y(men_men_n113_));
  NO3        u0064(.A(men_men_n113_), .B(men_men_n107_), .C(men_men_n53_), .Y(men_men_n114_));
  NO4        u0065(.A(men_men_n114_), .B(men_men_n106_), .C(men_men_n95_), .D(men_men_n80_), .Y(men00));
  NO2        u0066(.A(x7), .B(x6), .Y(men_men_n116_));
  INV        u0067(.A(men_men_n116_), .Y(men_men_n117_));
  NO2        u0068(.A(men_men_n55_), .B(men_men_n53_), .Y(men_men_n118_));
  NA2        u0069(.A(men_men_n118_), .B(men_men_n56_), .Y(men_men_n119_));
  NO2        u0070(.A(men_men_n119_), .B(men_men_n117_), .Y(men_men_n120_));
  XN2        u0071(.A(x6), .B(x1), .Y(men_men_n121_));
  INV        u0072(.A(men_men_n121_), .Y(men_men_n122_));
  NO2        u0073(.A(x6), .B(x4), .Y(men_men_n123_));
  NA2        u0074(.A(x6), .B(x4), .Y(men_men_n124_));
  NAi21      u0075(.An(men_men_n123_), .B(men_men_n124_), .Y(men_men_n125_));
  XN2        u0076(.A(x7), .B(x6), .Y(men_men_n126_));
  NO4        u0077(.A(men_men_n126_), .B(men_men_n125_), .C(men_men_n122_), .D(x8), .Y(men_men_n127_));
  NO2        u0078(.A(x3), .B(men_men_n110_), .Y(men_men_n128_));
  NA2        u0079(.A(men_men_n128_), .B(men_men_n108_), .Y(men_men_n129_));
  NO2        u0080(.A(men_men_n129_), .B(men_men_n59_), .Y(men_men_n130_));
  OAI210     u0081(.A0(men_men_n127_), .A1(men_men_n120_), .B0(men_men_n130_), .Y(men_men_n131_));
  NA2        u0082(.A(x3), .B(men_men_n110_), .Y(men_men_n132_));
  NO2        u0083(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n133_));
  NA2        u0084(.A(men_men_n133_), .B(men_men_n56_), .Y(men_men_n134_));
  NA2        u0085(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n135_));
  NA2        u0086(.A(men_men_n135_), .B(x2), .Y(men_men_n136_));
  NA2        u0087(.A(x8), .B(x3), .Y(men_men_n137_));
  NA2        u0088(.A(men_men_n137_), .B(men_men_n75_), .Y(men_men_n138_));
  OAI220     u0089(.A0(men_men_n138_), .A1(men_men_n136_), .B0(men_men_n134_), .B1(men_men_n132_), .Y(men_men_n139_));
  NO2        u0090(.A(x5), .B(x0), .Y(men_men_n140_));
  NO2        u0091(.A(x6), .B(x1), .Y(men_men_n141_));
  NA3        u0092(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n139_), .Y(men_men_n142_));
  NA2        u0093(.A(x8), .B(men_men_n108_), .Y(men_men_n143_));
  NA2        u0094(.A(x4), .B(men_men_n50_), .Y(men_men_n144_));
  NO3        u0095(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n104_), .Y(men_men_n145_));
  NAi21      u0096(.An(x7), .B(x2), .Y(men_men_n146_));
  NO2        u0097(.A(men_men_n146_), .B(x0), .Y(men_men_n147_));
  XO2        u0098(.A(x8), .B(x7), .Y(men_men_n148_));
  NA2        u0099(.A(men_men_n148_), .B(men_men_n110_), .Y(men_men_n149_));
  NA2        u0100(.A(x6), .B(x5), .Y(men_men_n150_));
  NO2        u0101(.A(men_men_n56_), .B(x0), .Y(men_men_n151_));
  NO2        u0102(.A(men_men_n50_), .B(x1), .Y(men_men_n152_));
  NA2        u0103(.A(men_men_n152_), .B(men_men_n151_), .Y(men_men_n153_));
  NO3        u0104(.A(men_men_n153_), .B(men_men_n150_), .C(men_men_n149_), .Y(men_men_n154_));
  AOI210     u0105(.A0(men_men_n147_), .A1(men_men_n145_), .B0(men_men_n154_), .Y(men_men_n155_));
  NA3        u0106(.A(men_men_n155_), .B(men_men_n142_), .C(men_men_n131_), .Y(men01));
  NA2        u0107(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n157_));
  NO2        u0108(.A(x2), .B(x1), .Y(men_men_n158_));
  NA2        u0109(.A(x2), .B(x1), .Y(men_men_n159_));
  NOi21      u0110(.An(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  NA2        u0111(.A(men_men_n108_), .B(men_men_n53_), .Y(men_men_n161_));
  NO2        u0112(.A(men_men_n161_), .B(x8), .Y(men_men_n162_));
  NAi21      u0113(.An(x8), .B(x1), .Y(men_men_n163_));
  NO2        u0114(.A(men_men_n163_), .B(x3), .Y(men_men_n164_));
  OAI210     u0115(.A0(men_men_n164_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n165_));
  NO2        u0116(.A(x5), .B(men_men_n50_), .Y(men_men_n166_));
  NO2        u0117(.A(men_men_n110_), .B(x1), .Y(men_men_n167_));
  NA2        u0118(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  AOI210     u0119(.A0(men_men_n168_), .A1(men_men_n165_), .B0(men_men_n157_), .Y(men_men_n169_));
  NAi21      u0120(.An(x7), .B(x0), .Y(men_men_n170_));
  NO2        u0121(.A(men_men_n55_), .B(x2), .Y(men_men_n171_));
  NO2        u0122(.A(men_men_n81_), .B(x1), .Y(men_men_n172_));
  NA2        u0123(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  NA2        u0124(.A(x5), .B(men_men_n50_), .Y(men_men_n174_));
  NO2        u0125(.A(men_men_n174_), .B(men_men_n163_), .Y(men_men_n175_));
  NA2        u0126(.A(x8), .B(x5), .Y(men_men_n176_));
  NO2        u0127(.A(men_men_n176_), .B(men_men_n51_), .Y(men_men_n177_));
  NO3        u0128(.A(x3), .B(men_men_n110_), .C(men_men_n53_), .Y(men_men_n178_));
  NO3        u0129(.A(men_men_n178_), .B(men_men_n177_), .C(men_men_n175_), .Y(men_men_n179_));
  AOI210     u0130(.A0(men_men_n179_), .A1(men_men_n173_), .B0(men_men_n170_), .Y(men_men_n180_));
  NO2        u0131(.A(men_men_n57_), .B(x3), .Y(men_men_n181_));
  NO2        u0132(.A(men_men_n55_), .B(x0), .Y(men_men_n182_));
  NA3        u0133(.A(men_men_n108_), .B(men_men_n110_), .C(x1), .Y(men_men_n183_));
  NO2        u0134(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  NO2        u0135(.A(men_men_n87_), .B(men_men_n50_), .Y(men_men_n185_));
  NA2        u0136(.A(men_men_n108_), .B(x0), .Y(men_men_n186_));
  NO2        u0137(.A(men_men_n186_), .B(x2), .Y(men_men_n187_));
  AOI220     u0138(.A0(men_men_n187_), .A1(men_men_n185_), .B0(men_men_n184_), .B1(men_men_n181_), .Y(men_men_n188_));
  NA2        u0139(.A(x7), .B(men_men_n110_), .Y(men_men_n189_));
  NA2        u0140(.A(men_men_n166_), .B(x8), .Y(men_men_n190_));
  NA4        u0141(.A(x5), .B(x3), .C(x1), .D(x0), .Y(men_men_n191_));
  AO210      u0142(.A0(men_men_n191_), .A1(men_men_n190_), .B0(men_men_n189_), .Y(men_men_n192_));
  NO2        u0143(.A(men_men_n159_), .B(men_men_n50_), .Y(men_men_n193_));
  NAi21      u0144(.An(x1), .B(x2), .Y(men_men_n194_));
  NO2        u0145(.A(men_men_n174_), .B(men_men_n194_), .Y(men_men_n195_));
  NA2        u0146(.A(x8), .B(x7), .Y(men_men_n196_));
  NO2        u0147(.A(men_men_n196_), .B(x0), .Y(men_men_n197_));
  OAI210     u0148(.A0(men_men_n195_), .A1(men_men_n193_), .B0(men_men_n197_), .Y(men_men_n198_));
  NA3        u0149(.A(men_men_n198_), .B(men_men_n192_), .C(men_men_n188_), .Y(men_men_n199_));
  NO3        u0150(.A(men_men_n199_), .B(men_men_n180_), .C(men_men_n169_), .Y(men_men_n200_));
  NA2        u0151(.A(x3), .B(x1), .Y(men_men_n201_));
  NA2        u0152(.A(men_men_n50_), .B(men_men_n110_), .Y(men_men_n202_));
  NO2        u0153(.A(men_men_n202_), .B(men_men_n70_), .Y(men_men_n203_));
  OAI210     u0154(.A0(men_men_n203_), .A1(men_men_n195_), .B0(men_men_n67_), .Y(men_men_n204_));
  NA2        u0155(.A(men_men_n133_), .B(men_men_n110_), .Y(men_men_n205_));
  OAI210     u0156(.A0(men_men_n205_), .A1(men_men_n201_), .B0(men_men_n204_), .Y(men_men_n206_));
  XO2        u0157(.A(x5), .B(x3), .Y(men_men_n207_));
  NA2        u0158(.A(men_men_n207_), .B(x8), .Y(men_men_n208_));
  NA2        u0159(.A(x8), .B(men_men_n59_), .Y(men_men_n209_));
  NA2        u0160(.A(men_men_n209_), .B(men_men_n137_), .Y(men_men_n210_));
  NA2        u0161(.A(x7), .B(men_men_n71_), .Y(men_men_n211_));
  NO2        u0162(.A(men_men_n194_), .B(men_men_n211_), .Y(men_men_n212_));
  OA210      u0163(.A0(men_men_n210_), .A1(men_men_n207_), .B0(men_men_n212_), .Y(men_men_n213_));
  AOI220     u0164(.A0(men_men_n213_), .A1(men_men_n208_), .B0(men_men_n206_), .B1(x0), .Y(men_men_n214_));
  OAI210     u0165(.A0(men_men_n200_), .A1(men_men_n71_), .B0(men_men_n214_), .Y(men_men_n215_));
  NO2        u0166(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n216_));
  NA4        u0167(.A(men_men_n55_), .B(x5), .C(x3), .D(x2), .Y(men_men_n217_));
  NA2        u0168(.A(x8), .B(men_men_n50_), .Y(men_men_n218_));
  NA2        u0169(.A(men_men_n218_), .B(x2), .Y(men_men_n219_));
  NA2        u0170(.A(men_men_n55_), .B(x3), .Y(men_men_n220_));
  NA4        u0171(.A(men_men_n220_), .B(men_men_n219_), .C(men_men_n207_), .D(men_men_n82_), .Y(men_men_n221_));
  AOI210     u0172(.A0(men_men_n221_), .A1(men_men_n217_), .B0(men_men_n53_), .Y(men_men_n222_));
  NO2        u0173(.A(men_men_n110_), .B(men_men_n59_), .Y(men_men_n223_));
  NA2        u0174(.A(x5), .B(x1), .Y(men_men_n224_));
  NO2        u0175(.A(men_men_n224_), .B(x6), .Y(men_men_n225_));
  NO2        u0176(.A(x3), .B(x1), .Y(men_men_n226_));
  AOI210     u0177(.A0(men_men_n226_), .A1(men_men_n77_), .B0(men_men_n225_), .Y(men_men_n227_));
  NO2        u0178(.A(men_men_n81_), .B(men_men_n55_), .Y(men_men_n228_));
  NO2        u0179(.A(men_men_n104_), .B(men_men_n50_), .Y(men_men_n229_));
  NO2        u0180(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  OAI210     u0181(.A0(men_men_n227_), .A1(x8), .B0(men_men_n230_), .Y(men_men_n231_));
  NO2        u0182(.A(men_men_n55_), .B(x5), .Y(men_men_n232_));
  NA2        u0183(.A(men_men_n232_), .B(men_men_n71_), .Y(men_men_n233_));
  NAi21      u0184(.An(x2), .B(x5), .Y(men_men_n234_));
  NA2        u0185(.A(x8), .B(x6), .Y(men_men_n235_));
  OAI210     u0186(.A0(men_men_n235_), .A1(men_men_n234_), .B0(men_men_n233_), .Y(men_men_n236_));
  NA2        u0187(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n237_));
  NO2        u0188(.A(men_men_n237_), .B(men_men_n59_), .Y(men_men_n238_));
  AO220      u0189(.A0(men_men_n238_), .A1(men_men_n236_), .B0(men_men_n231_), .B1(men_men_n223_), .Y(men_men_n239_));
  OAI210     u0190(.A0(men_men_n239_), .A1(men_men_n222_), .B0(men_men_n216_), .Y(men_men_n240_));
  NA2        u0191(.A(men_men_n71_), .B(men_men_n56_), .Y(men_men_n241_));
  NO2        u0192(.A(men_men_n241_), .B(x7), .Y(men_men_n242_));
  NO2        u0193(.A(men_men_n108_), .B(men_men_n53_), .Y(men_men_n243_));
  NA2        u0194(.A(men_men_n243_), .B(men_men_n110_), .Y(men_men_n244_));
  AOI210     u0195(.A0(men_men_n244_), .A1(men_men_n168_), .B0(men_men_n59_), .Y(men_men_n245_));
  NA2        u0196(.A(x3), .B(men_men_n59_), .Y(men_men_n246_));
  NO2        u0197(.A(men_men_n183_), .B(men_men_n246_), .Y(men_men_n247_));
  OA210      u0198(.A0(men_men_n247_), .A1(men_men_n245_), .B0(x8), .Y(men_men_n248_));
  NO2        u0199(.A(x1), .B(x0), .Y(men_men_n249_));
  NA2        u0200(.A(men_men_n249_), .B(men_men_n110_), .Y(men_men_n250_));
  NA2        u0201(.A(men_men_n108_), .B(men_men_n50_), .Y(men_men_n251_));
  XN2        u0202(.A(x3), .B(x2), .Y(men_men_n252_));
  NA2        u0203(.A(men_men_n252_), .B(men_men_n160_), .Y(men_men_n253_));
  NO2        u0204(.A(men_men_n108_), .B(x0), .Y(men_men_n254_));
  NA2        u0205(.A(x8), .B(men_men_n53_), .Y(men_men_n255_));
  NA2        u0206(.A(men_men_n255_), .B(men_men_n254_), .Y(men_men_n256_));
  OAI220     u0207(.A0(men_men_n256_), .A1(men_men_n253_), .B0(men_men_n251_), .B1(men_men_n250_), .Y(men_men_n257_));
  OAI210     u0208(.A0(men_men_n257_), .A1(men_men_n248_), .B0(men_men_n242_), .Y(men_men_n258_));
  NO2        u0209(.A(x7), .B(x1), .Y(men_men_n259_));
  NOi21      u0210(.An(x8), .B(x3), .Y(men_men_n260_));
  NA2        u0211(.A(men_men_n260_), .B(men_men_n59_), .Y(men_men_n261_));
  NA2        u0212(.A(x5), .B(x0), .Y(men_men_n262_));
  NAi21      u0213(.An(men_men_n140_), .B(men_men_n262_), .Y(men_men_n263_));
  NA2        u0214(.A(men_men_n71_), .B(men_men_n50_), .Y(men_men_n264_));
  OAI210     u0215(.A0(men_men_n264_), .A1(men_men_n263_), .B0(men_men_n261_), .Y(men_men_n265_));
  NA3        u0216(.A(men_men_n265_), .B(men_men_n143_), .C(men_men_n259_), .Y(men_men_n266_));
  NA2        u0217(.A(x8), .B(men_men_n57_), .Y(men_men_n267_));
  NO2        u0218(.A(men_men_n267_), .B(x5), .Y(men_men_n268_));
  NO2        u0219(.A(men_men_n152_), .B(men_men_n71_), .Y(men_men_n269_));
  NA2        u0220(.A(x1), .B(x0), .Y(men_men_n270_));
  NA2        u0221(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n271_));
  NA4        u0222(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n269_), .D(men_men_n268_), .Y(men_men_n272_));
  NA3        u0223(.A(men_men_n272_), .B(men_men_n266_), .C(men_men_n191_), .Y(men_men_n273_));
  NO2        u0224(.A(men_men_n108_), .B(x3), .Y(men_men_n274_));
  NO2        u0225(.A(men_men_n110_), .B(x0), .Y(men_men_n275_));
  NA2        u0226(.A(men_men_n275_), .B(men_men_n274_), .Y(men_men_n276_));
  NO2        u0227(.A(men_men_n55_), .B(x7), .Y(men_men_n277_));
  NA2        u0228(.A(men_men_n277_), .B(men_men_n141_), .Y(men_men_n278_));
  NO3        u0229(.A(x8), .B(men_men_n50_), .C(x0), .Y(men_men_n279_));
  NAi21      u0230(.An(x8), .B(x0), .Y(men_men_n280_));
  NAi21      u0231(.An(x1), .B(x3), .Y(men_men_n281_));
  NO2        u0232(.A(men_men_n281_), .B(men_men_n280_), .Y(men_men_n282_));
  NO2        u0233(.A(x2), .B(men_men_n53_), .Y(men_men_n283_));
  AOI210     u0234(.A0(men_men_n283_), .A1(men_men_n279_), .B0(men_men_n282_), .Y(men_men_n284_));
  NOi21      u0235(.An(x5), .B(x6), .Y(men_men_n285_));
  NO2        u0236(.A(men_men_n57_), .B(x4), .Y(men_men_n286_));
  NA2        u0237(.A(men_men_n286_), .B(men_men_n285_), .Y(men_men_n287_));
  OAI220     u0238(.A0(men_men_n287_), .A1(men_men_n284_), .B0(men_men_n278_), .B1(men_men_n276_), .Y(men_men_n288_));
  AOI210     u0239(.A0(men_men_n273_), .A1(men_men_n111_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA3        u0240(.A(men_men_n289_), .B(men_men_n258_), .C(men_men_n240_), .Y(men_men_n290_));
  AOI210     u0241(.A0(men_men_n215_), .A1(men_men_n56_), .B0(men_men_n290_), .Y(men02));
  NO2        u0242(.A(x8), .B(men_men_n108_), .Y(men_men_n292_));
  XN2        u0243(.A(x7), .B(x3), .Y(men_men_n293_));
  INV        u0244(.A(men_men_n293_), .Y(men_men_n294_));
  NO2        u0245(.A(x2), .B(x0), .Y(men_men_n295_));
  NA2        u0246(.A(men_men_n295_), .B(men_men_n71_), .Y(men_men_n296_));
  NO2        u0247(.A(men_men_n57_), .B(x1), .Y(men_men_n297_));
  NO3        u0248(.A(men_men_n297_), .B(men_men_n296_), .C(men_men_n294_), .Y(men_men_n298_));
  NA2        u0249(.A(men_men_n53_), .B(x0), .Y(men_men_n299_));
  NO2        u0250(.A(men_men_n281_), .B(x6), .Y(men_men_n300_));
  XO2        u0251(.A(x7), .B(x0), .Y(men_men_n301_));
  NO2        u0252(.A(men_men_n301_), .B(men_men_n295_), .Y(men_men_n302_));
  NA2        u0253(.A(men_men_n302_), .B(men_men_n300_), .Y(men_men_n303_));
  AN2        u0254(.A(x7), .B(x2), .Y(men_men_n304_));
  NA2        u0255(.A(men_men_n304_), .B(men_men_n50_), .Y(men_men_n305_));
  OAI210     u0256(.A0(men_men_n305_), .A1(men_men_n299_), .B0(men_men_n303_), .Y(men_men_n306_));
  OAI210     u0257(.A0(men_men_n306_), .A1(men_men_n298_), .B0(men_men_n292_), .Y(men_men_n307_));
  NAi21      u0258(.An(x8), .B(x6), .Y(men_men_n308_));
  NO2        u0259(.A(men_men_n108_), .B(men_men_n59_), .Y(men_men_n309_));
  NA2        u0260(.A(x7), .B(x3), .Y(men_men_n310_));
  NO2        u0261(.A(men_men_n310_), .B(x2), .Y(men_men_n311_));
  NA2        u0262(.A(x2), .B(x0), .Y(men_men_n312_));
  NA2        u0263(.A(men_men_n110_), .B(men_men_n59_), .Y(men_men_n313_));
  NA2        u0264(.A(men_men_n313_), .B(men_men_n312_), .Y(men_men_n314_));
  NAi21      u0265(.An(x7), .B(x1), .Y(men_men_n315_));
  NO2        u0266(.A(men_men_n315_), .B(x3), .Y(men_men_n316_));
  AOI220     u0267(.A0(men_men_n316_), .A1(men_men_n314_), .B0(men_men_n311_), .B1(men_men_n309_), .Y(men_men_n317_));
  NA2        u0268(.A(men_men_n283_), .B(men_men_n50_), .Y(men_men_n318_));
  NA3        u0269(.A(x7), .B(men_men_n108_), .C(x0), .Y(men_men_n319_));
  NA2        u0270(.A(men_men_n166_), .B(men_men_n57_), .Y(men_men_n320_));
  NO2        u0271(.A(men_men_n317_), .B(men_men_n308_), .Y(men_men_n321_));
  INV        u0272(.A(men_men_n301_), .Y(men_men_n322_));
  NO2        u0273(.A(x7), .B(men_men_n71_), .Y(men_men_n323_));
  NA2        u0274(.A(men_men_n108_), .B(x3), .Y(men_men_n324_));
  NO2        u0275(.A(men_men_n324_), .B(men_men_n323_), .Y(men_men_n325_));
  NA2        u0276(.A(men_men_n325_), .B(men_men_n322_), .Y(men_men_n326_));
  NA2        u0277(.A(men_men_n50_), .B(x0), .Y(men_men_n327_));
  NO2        u0278(.A(men_men_n327_), .B(x7), .Y(men_men_n328_));
  NA2        u0279(.A(men_men_n328_), .B(men_men_n285_), .Y(men_men_n329_));
  NA2        u0280(.A(men_men_n171_), .B(x1), .Y(men_men_n330_));
  AOI210     u0281(.A0(men_men_n329_), .A1(men_men_n326_), .B0(men_men_n330_), .Y(men_men_n331_));
  NO2        u0282(.A(men_men_n57_), .B(men_men_n50_), .Y(men_men_n332_));
  NO2        u0283(.A(men_men_n55_), .B(men_men_n110_), .Y(men_men_n333_));
  NA3        u0284(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n59_), .Y(men_men_n334_));
  NO2        u0285(.A(men_men_n161_), .B(x6), .Y(men_men_n335_));
  NO2        u0286(.A(men_men_n104_), .B(men_men_n108_), .Y(men_men_n336_));
  NA2        u0287(.A(men_men_n57_), .B(men_men_n110_), .Y(men_men_n337_));
  NO2        u0288(.A(men_men_n337_), .B(men_men_n271_), .Y(men_men_n338_));
  OAI210     u0289(.A0(men_men_n336_), .A1(men_men_n335_), .B0(men_men_n338_), .Y(men_men_n339_));
  OAI210     u0290(.A0(men_men_n334_), .A1(men_men_n104_), .B0(men_men_n339_), .Y(men_men_n340_));
  NO3        u0291(.A(men_men_n340_), .B(men_men_n331_), .C(men_men_n321_), .Y(men_men_n341_));
  AOI210     u0292(.A0(men_men_n341_), .A1(men_men_n307_), .B0(x4), .Y(men_men_n342_));
  NA2        u0293(.A(x8), .B(men_men_n71_), .Y(men_men_n343_));
  NO2        u0294(.A(x3), .B(men_men_n59_), .Y(men_men_n344_));
  NA3        u0295(.A(men_men_n344_), .B(men_men_n108_), .C(men_men_n53_), .Y(men_men_n345_));
  NO2        u0296(.A(x3), .B(x0), .Y(men_men_n346_));
  NAi21      u0297(.An(men_men_n346_), .B(men_men_n107_), .Y(men_men_n347_));
  NA2        u0298(.A(x5), .B(x2), .Y(men_men_n348_));
  NO2        u0299(.A(men_men_n348_), .B(men_men_n226_), .Y(men_men_n349_));
  AOI210     u0300(.A0(men_men_n349_), .A1(men_men_n347_), .B0(men_men_n247_), .Y(men_men_n350_));
  AO210      u0301(.A0(men_men_n350_), .A1(men_men_n345_), .B0(men_men_n343_), .Y(men_men_n351_));
  NO2        u0302(.A(men_men_n110_), .B(men_men_n53_), .Y(men_men_n352_));
  NA2        u0303(.A(men_men_n352_), .B(x3), .Y(men_men_n353_));
  NO2        u0304(.A(men_men_n55_), .B(x1), .Y(men_men_n354_));
  NA2        u0305(.A(men_men_n354_), .B(men_men_n110_), .Y(men_men_n355_));
  OAI210     u0306(.A0(men_men_n355_), .A1(men_men_n174_), .B0(men_men_n353_), .Y(men_men_n356_));
  NAi32      u0307(.An(x3), .Bn(x0), .C(x2), .Y(men_men_n357_));
  NO2        u0308(.A(men_men_n50_), .B(x2), .Y(men_men_n358_));
  NAi21      u0309(.An(x6), .B(x5), .Y(men_men_n359_));
  NO2        u0310(.A(x2), .B(men_men_n59_), .Y(men_men_n360_));
  NO4        u0311(.A(men_men_n360_), .B(men_men_n359_), .C(men_men_n163_), .D(men_men_n358_), .Y(men_men_n361_));
  AOI220     u0312(.A0(men_men_n361_), .A1(men_men_n357_), .B0(men_men_n356_), .B1(men_men_n85_), .Y(men_men_n362_));
  AOI210     u0313(.A0(men_men_n362_), .A1(men_men_n351_), .B0(men_men_n75_), .Y(men_men_n363_));
  NA2        u0314(.A(men_men_n354_), .B(men_men_n56_), .Y(men_men_n364_));
  NO2        u0315(.A(men_men_n108_), .B(men_men_n50_), .Y(men_men_n365_));
  NO2        u0316(.A(men_men_n295_), .B(men_men_n223_), .Y(men_men_n366_));
  XO2        u0317(.A(x7), .B(x2), .Y(men_men_n367_));
  INV        u0318(.A(men_men_n367_), .Y(men_men_n368_));
  XO2        u0319(.A(x6), .B(x2), .Y(men_men_n369_));
  NA4        u0320(.A(men_men_n369_), .B(men_men_n368_), .C(men_men_n366_), .D(men_men_n365_), .Y(men_men_n370_));
  NAi21      u0321(.An(x0), .B(x6), .Y(men_men_n371_));
  AOI210     u0322(.A0(men_men_n371_), .A1(men_men_n146_), .B0(men_men_n275_), .Y(men_men_n372_));
  XN2        u0323(.A(x7), .B(x5), .Y(men_men_n373_));
  NA2        u0324(.A(men_men_n373_), .B(men_men_n71_), .Y(men_men_n374_));
  NA2        u0325(.A(x7), .B(x5), .Y(men_men_n375_));
  AOI210     u0326(.A0(men_men_n375_), .A1(x6), .B0(men_men_n357_), .Y(men_men_n376_));
  AOI220     u0327(.A0(men_men_n376_), .A1(men_men_n374_), .B0(men_men_n372_), .B1(men_men_n325_), .Y(men_men_n377_));
  AOI210     u0328(.A0(men_men_n377_), .A1(men_men_n370_), .B0(men_men_n364_), .Y(men_men_n378_));
  NO2        u0329(.A(x8), .B(x6), .Y(men_men_n379_));
  NAi21      u0330(.An(men_men_n379_), .B(men_men_n235_), .Y(men_men_n380_));
  AOI210     u0331(.A0(men_men_n380_), .A1(men_men_n92_), .B0(x3), .Y(men_men_n381_));
  NA2        u0332(.A(men_men_n108_), .B(x2), .Y(men_men_n382_));
  NO2        u0333(.A(men_men_n382_), .B(men_men_n64_), .Y(men_men_n383_));
  NA2        u0334(.A(x1), .B(men_men_n59_), .Y(men_men_n384_));
  NO2        u0335(.A(men_men_n384_), .B(men_men_n235_), .Y(men_men_n385_));
  OAI210     u0336(.A0(men_men_n385_), .A1(men_men_n50_), .B0(men_men_n383_), .Y(men_men_n386_));
  NA2        u0337(.A(x4), .B(x2), .Y(men_men_n387_));
  NO2        u0338(.A(men_men_n387_), .B(men_men_n108_), .Y(men_men_n388_));
  NAi21      u0339(.An(x1), .B(x6), .Y(men_men_n389_));
  NA2        u0340(.A(men_men_n346_), .B(men_men_n277_), .Y(men_men_n390_));
  OAI220     u0341(.A0(men_men_n390_), .A1(men_men_n389_), .B0(men_men_n107_), .B1(men_men_n53_), .Y(men_men_n391_));
  NA2        u0342(.A(x8), .B(x2), .Y(men_men_n392_));
  NO2        u0343(.A(men_men_n392_), .B(men_men_n50_), .Y(men_men_n393_));
  INV        u0344(.A(men_men_n225_), .Y(men_men_n394_));
  NO2        u0345(.A(men_men_n394_), .B(men_men_n52_), .Y(men_men_n395_));
  AOI220     u0346(.A0(men_men_n395_), .A1(men_men_n393_), .B0(men_men_n391_), .B1(men_men_n388_), .Y(men_men_n396_));
  OAI210     u0347(.A0(men_men_n386_), .A1(men_men_n381_), .B0(men_men_n396_), .Y(men_men_n397_));
  NO4        u0348(.A(men_men_n397_), .B(men_men_n378_), .C(men_men_n363_), .D(men_men_n342_), .Y(men03));
  NAi21      u0349(.An(x2), .B(x0), .Y(men_men_n399_));
  NO3        u0350(.A(x8), .B(x6), .C(x4), .Y(men_men_n400_));
  INV        u0351(.A(men_men_n400_), .Y(men_men_n401_));
  NO2        u0352(.A(men_men_n401_), .B(men_men_n399_), .Y(men_men_n402_));
  NA2        u0353(.A(men_men_n111_), .B(men_men_n59_), .Y(men_men_n403_));
  NO2        u0354(.A(men_men_n403_), .B(men_men_n55_), .Y(men_men_n404_));
  OAI210     u0355(.A0(men_men_n404_), .A1(men_men_n402_), .B0(men_men_n166_), .Y(men_men_n405_));
  NA2        u0356(.A(x3), .B(x2), .Y(men_men_n406_));
  NO2        u0357(.A(men_men_n163_), .B(x0), .Y(men_men_n407_));
  NA2        u0358(.A(x8), .B(x0), .Y(men_men_n408_));
  NO2        u0359(.A(men_men_n408_), .B(x6), .Y(men_men_n409_));
  AOI210     u0360(.A0(men_men_n409_), .A1(x5), .B0(men_men_n407_), .Y(men_men_n410_));
  NO2        u0361(.A(men_men_n410_), .B(men_men_n406_), .Y(men_men_n411_));
  NO2        u0362(.A(x5), .B(men_men_n59_), .Y(men_men_n412_));
  NO2        u0363(.A(x3), .B(x2), .Y(men_men_n413_));
  NA2        u0364(.A(men_men_n413_), .B(men_men_n412_), .Y(men_men_n414_));
  NO2        u0365(.A(men_men_n53_), .B(x0), .Y(men_men_n415_));
  NA2        u0366(.A(men_men_n415_), .B(x5), .Y(men_men_n416_));
  AOI210     u0367(.A0(men_men_n416_), .A1(men_men_n414_), .B0(men_men_n308_), .Y(men_men_n417_));
  NA2        u0368(.A(men_men_n261_), .B(men_men_n176_), .Y(men_men_n418_));
  NO2        u0369(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n419_));
  NO2        u0370(.A(men_men_n71_), .B(x0), .Y(men_men_n420_));
  NO4        u0371(.A(men_men_n420_), .B(men_men_n419_), .C(x2), .D(men_men_n53_), .Y(men_men_n421_));
  AO210      u0372(.A0(men_men_n421_), .A1(men_men_n418_), .B0(men_men_n417_), .Y(men_men_n422_));
  OAI210     u0373(.A0(men_men_n422_), .A1(men_men_n411_), .B0(x4), .Y(men_men_n423_));
  NO2        u0374(.A(x4), .B(men_men_n53_), .Y(men_men_n424_));
  NA2        u0375(.A(men_men_n424_), .B(men_men_n59_), .Y(men_men_n425_));
  NO3        u0376(.A(men_men_n425_), .B(men_men_n235_), .C(x5), .Y(men_men_n426_));
  NA2        u0377(.A(x7), .B(men_men_n108_), .Y(men_men_n427_));
  NO3        u0378(.A(x5), .B(men_men_n53_), .C(x0), .Y(men_men_n428_));
  INV        u0379(.A(men_men_n428_), .Y(men_men_n429_));
  NO2        u0380(.A(x6), .B(men_men_n56_), .Y(men_men_n430_));
  NO2        u0381(.A(x8), .B(men_men_n50_), .Y(men_men_n431_));
  NA2        u0382(.A(men_men_n431_), .B(men_men_n430_), .Y(men_men_n432_));
  OAI210     u0383(.A0(men_men_n432_), .A1(men_men_n429_), .B0(men_men_n427_), .Y(men_men_n433_));
  AOI210     u0384(.A0(men_men_n426_), .A1(x2), .B0(men_men_n433_), .Y(men_men_n434_));
  AOI220     u0385(.A0(men_men_n434_), .A1(men_men_n423_), .B0(men_men_n405_), .B1(x7), .Y(men_men_n435_));
  NA2        u0386(.A(x7), .B(men_men_n53_), .Y(men_men_n436_));
  NO2        u0387(.A(men_men_n260_), .B(men_men_n110_), .Y(men_men_n437_));
  NO2        u0388(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n438_));
  NO3        u0389(.A(men_men_n438_), .B(men_men_n437_), .C(men_men_n150_), .Y(men_men_n439_));
  AOI210     u0390(.A0(men_men_n210_), .A1(men_men_n101_), .B0(men_men_n439_), .Y(men_men_n440_));
  NO2        u0391(.A(x5), .B(x2), .Y(men_men_n441_));
  NO2        u0392(.A(x8), .B(x3), .Y(men_men_n442_));
  NA2        u0393(.A(men_men_n442_), .B(men_men_n441_), .Y(men_men_n443_));
  NO2        u0394(.A(men_men_n443_), .B(x6), .Y(men_men_n444_));
  NA2        u0395(.A(men_men_n209_), .B(x2), .Y(men_men_n445_));
  NO3        u0396(.A(men_men_n442_), .B(men_men_n347_), .C(men_men_n359_), .Y(men_men_n446_));
  AOI210     u0397(.A0(men_men_n446_), .A1(men_men_n445_), .B0(men_men_n444_), .Y(men_men_n447_));
  OAI210     u0398(.A0(men_men_n440_), .A1(men_men_n295_), .B0(men_men_n447_), .Y(men_men_n448_));
  NA2        u0399(.A(men_men_n448_), .B(x4), .Y(men_men_n449_));
  NA2        u0400(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n450_));
  NO2        u0401(.A(men_men_n450_), .B(x5), .Y(men_men_n451_));
  NAi21      u0402(.An(x4), .B(x6), .Y(men_men_n452_));
  NO2        u0403(.A(men_men_n452_), .B(men_men_n51_), .Y(men_men_n453_));
  NO2        u0404(.A(men_men_n55_), .B(men_men_n71_), .Y(men_men_n454_));
  NO2        u0405(.A(men_men_n50_), .B(men_men_n110_), .Y(men_men_n455_));
  NO2        u0406(.A(men_men_n235_), .B(x0), .Y(men_men_n456_));
  NO2        u0407(.A(men_men_n359_), .B(x8), .Y(men_men_n457_));
  OAI210     u0408(.A0(men_men_n457_), .A1(men_men_n456_), .B0(men_men_n455_), .Y(men_men_n458_));
  OAI210     u0409(.A0(men_men_n414_), .A1(men_men_n454_), .B0(men_men_n458_), .Y(men_men_n459_));
  AOI220     u0410(.A0(men_men_n459_), .A1(men_men_n56_), .B0(men_men_n453_), .B1(men_men_n451_), .Y(men_men_n460_));
  AOI210     u0411(.A0(men_men_n460_), .A1(men_men_n449_), .B0(men_men_n436_), .Y(men_men_n461_));
  NA2        u0412(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n462_));
  NO2        u0413(.A(men_men_n71_), .B(men_men_n56_), .Y(men_men_n463_));
  NA2        u0414(.A(men_men_n358_), .B(men_men_n59_), .Y(men_men_n464_));
  OAI220     u0415(.A0(men_men_n464_), .A1(men_men_n55_), .B0(men_men_n202_), .B1(men_men_n280_), .Y(men_men_n465_));
  NA2        u0416(.A(men_men_n465_), .B(men_men_n463_), .Y(men_men_n466_));
  NO3        u0417(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n467_));
  NA2        u0418(.A(men_men_n438_), .B(x5), .Y(men_men_n468_));
  NO2        u0419(.A(x8), .B(x5), .Y(men_men_n469_));
  NAi21      u0420(.An(men_men_n469_), .B(men_men_n176_), .Y(men_men_n470_));
  OAI210     u0421(.A0(men_men_n470_), .A1(men_men_n313_), .B0(men_men_n468_), .Y(men_men_n471_));
  NA2        u0422(.A(men_men_n366_), .B(men_men_n77_), .Y(men_men_n472_));
  NOi21      u0423(.An(x3), .B(x4), .Y(men_men_n473_));
  NA2        u0424(.A(men_men_n55_), .B(men_men_n110_), .Y(men_men_n474_));
  NA2        u0425(.A(men_men_n474_), .B(men_men_n473_), .Y(men_men_n475_));
  NO2        u0426(.A(men_men_n51_), .B(x6), .Y(men_men_n476_));
  NO2        u0427(.A(men_men_n150_), .B(men_men_n55_), .Y(men_men_n477_));
  NO3        u0428(.A(men_men_n56_), .B(x2), .C(x0), .Y(men_men_n478_));
  AOI220     u0429(.A0(men_men_n478_), .A1(men_men_n477_), .B0(men_men_n476_), .B1(men_men_n451_), .Y(men_men_n479_));
  OAI210     u0430(.A0(men_men_n475_), .A1(men_men_n472_), .B0(men_men_n479_), .Y(men_men_n480_));
  AOI210     u0431(.A0(men_men_n471_), .A1(men_men_n467_), .B0(men_men_n480_), .Y(men_men_n481_));
  AOI210     u0432(.A0(men_men_n481_), .A1(men_men_n466_), .B0(men_men_n462_), .Y(men_men_n482_));
  NA2        u0433(.A(x7), .B(x1), .Y(men_men_n483_));
  NO3        u0434(.A(x5), .B(x4), .C(x2), .Y(men_men_n484_));
  AN2        u0435(.A(men_men_n484_), .B(men_men_n379_), .Y(men_men_n485_));
  NO3        u0436(.A(men_men_n485_), .B(men_men_n477_), .C(men_men_n388_), .Y(men_men_n486_));
  OAI210     u0437(.A0(men_men_n379_), .A1(men_men_n84_), .B0(men_men_n346_), .Y(men_men_n487_));
  NO2        u0438(.A(men_men_n487_), .B(men_men_n486_), .Y(men_men_n488_));
  NO2        u0439(.A(x4), .B(men_men_n110_), .Y(men_men_n489_));
  NA2        u0440(.A(men_men_n489_), .B(x6), .Y(men_men_n490_));
  NA3        u0441(.A(men_men_n108_), .B(x4), .C(men_men_n110_), .Y(men_men_n491_));
  AOI210     u0442(.A0(men_men_n491_), .A1(men_men_n490_), .B0(men_men_n100_), .Y(men_men_n492_));
  NA2        u0443(.A(men_men_n473_), .B(men_men_n71_), .Y(men_men_n493_));
  NA2        u0444(.A(men_men_n171_), .B(men_men_n59_), .Y(men_men_n494_));
  NO2        u0445(.A(men_men_n494_), .B(men_men_n493_), .Y(men_men_n495_));
  NA2        u0446(.A(men_men_n455_), .B(x4), .Y(men_men_n496_));
  NO3        u0447(.A(men_men_n496_), .B(men_men_n379_), .C(men_men_n420_), .Y(men_men_n497_));
  NO4        u0448(.A(men_men_n497_), .B(men_men_n495_), .C(men_men_n492_), .D(men_men_n488_), .Y(men_men_n498_));
  NA2        u0449(.A(x5), .B(x4), .Y(men_men_n499_));
  NO2        u0450(.A(men_men_n71_), .B(men_men_n53_), .Y(men_men_n500_));
  NO3        u0451(.A(x8), .B(x3), .C(x2), .Y(men_men_n501_));
  NA3        u0452(.A(men_men_n501_), .B(men_men_n500_), .C(men_men_n59_), .Y(men_men_n502_));
  NO3        u0453(.A(x6), .B(x5), .C(x2), .Y(men_men_n503_));
  NA3        u0454(.A(men_men_n503_), .B(men_men_n297_), .C(men_men_n78_), .Y(men_men_n504_));
  OAI210     u0455(.A0(men_men_n502_), .A1(men_men_n499_), .B0(men_men_n504_), .Y(men_men_n505_));
  NA2        u0456(.A(men_men_n71_), .B(x2), .Y(men_men_n506_));
  NO3        u0457(.A(x4), .B(x3), .C(men_men_n59_), .Y(men_men_n507_));
  NA2        u0458(.A(men_men_n507_), .B(men_men_n232_), .Y(men_men_n508_));
  NO3        u0459(.A(men_men_n508_), .B(men_men_n506_), .C(men_men_n96_), .Y(men_men_n509_));
  XO2        u0460(.A(x4), .B(x0), .Y(men_men_n510_));
  NA2        u0461(.A(men_men_n271_), .B(x5), .Y(men_men_n511_));
  NO2        u0462(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n512_));
  NO2        u0463(.A(men_men_n512_), .B(men_men_n63_), .Y(men_men_n513_));
  NO4        u0464(.A(men_men_n513_), .B(men_men_n511_), .C(men_men_n510_), .D(men_men_n159_), .Y(men_men_n514_));
  NO3        u0465(.A(men_men_n514_), .B(men_men_n509_), .C(men_men_n505_), .Y(men_men_n515_));
  OAI210     u0466(.A0(men_men_n498_), .A1(men_men_n483_), .B0(men_men_n515_), .Y(men_men_n516_));
  NO4        u0467(.A(men_men_n516_), .B(men_men_n482_), .C(men_men_n461_), .D(men_men_n435_), .Y(men04));
  NO2        u0468(.A(x7), .B(x2), .Y(men_men_n518_));
  NO2        u0469(.A(x3), .B(men_men_n53_), .Y(men_men_n519_));
  NO2        u0470(.A(men_men_n519_), .B(men_men_n152_), .Y(men_men_n520_));
  XN2        u0471(.A(x8), .B(x1), .Y(men_men_n521_));
  NO2        u0472(.A(men_men_n521_), .B(men_men_n150_), .Y(men_men_n522_));
  NA2        u0473(.A(men_men_n522_), .B(men_men_n520_), .Y(men_men_n523_));
  NA2        u0474(.A(x6), .B(x3), .Y(men_men_n524_));
  NO2        u0475(.A(men_men_n524_), .B(x5), .Y(men_men_n525_));
  NA2        u0476(.A(men_men_n71_), .B(x1), .Y(men_men_n526_));
  NO2        u0477(.A(men_men_n469_), .B(men_men_n260_), .Y(men_men_n527_));
  NO3        u0478(.A(men_men_n527_), .B(men_men_n442_), .C(men_men_n526_), .Y(men_men_n528_));
  AOI210     u0479(.A0(men_men_n525_), .A1(men_men_n354_), .B0(men_men_n528_), .Y(men_men_n529_));
  AOI210     u0480(.A0(men_men_n529_), .A1(men_men_n523_), .B0(x0), .Y(men_men_n530_));
  NOi21      u0481(.An(men_men_n176_), .B(men_men_n469_), .Y(men_men_n531_));
  NA2        u0482(.A(men_men_n109_), .B(x1), .Y(men_men_n532_));
  NO3        u0483(.A(men_men_n532_), .B(men_men_n531_), .C(men_men_n327_), .Y(men_men_n533_));
  OAI210     u0484(.A0(men_men_n533_), .A1(men_men_n530_), .B0(men_men_n518_), .Y(men_men_n534_));
  NA2        u0485(.A(men_men_n137_), .B(men_men_n246_), .Y(men_men_n535_));
  OR4        u0486(.A(men_men_n535_), .B(men_men_n380_), .C(men_men_n82_), .D(men_men_n54_), .Y(men_men_n536_));
  OR2        u0487(.A(x6), .B(x0), .Y(men_men_n537_));
  NO3        u0488(.A(men_men_n537_), .B(x3), .C(x1), .Y(men_men_n538_));
  AOI220     u0489(.A0(men_men_n538_), .A1(men_men_n108_), .B0(men_men_n285_), .B1(men_men_n279_), .Y(men_men_n539_));
  AOI210     u0490(.A0(men_men_n539_), .A1(men_men_n536_), .B0(men_men_n189_), .Y(men_men_n540_));
  NA2        u0491(.A(x7), .B(x2), .Y(men_men_n541_));
  INV        u0492(.A(men_men_n137_), .Y(men_men_n542_));
  OAI210     u0493(.A0(men_men_n175_), .A1(men_men_n542_), .B0(men_men_n82_), .Y(men_men_n543_));
  NO2        u0494(.A(men_men_n324_), .B(men_men_n55_), .Y(men_men_n544_));
  NO3        u0495(.A(x3), .B(x1), .C(x0), .Y(men_men_n545_));
  OR2        u0496(.A(x6), .B(x1), .Y(men_men_n546_));
  NA2        u0497(.A(men_men_n546_), .B(x0), .Y(men_men_n547_));
  AOI220     u0498(.A0(men_men_n547_), .A1(men_men_n544_), .B0(men_men_n545_), .B1(men_men_n477_), .Y(men_men_n548_));
  AOI210     u0499(.A0(men_men_n548_), .A1(men_men_n543_), .B0(men_men_n541_), .Y(men_men_n549_));
  NA2        u0500(.A(men_men_n71_), .B(x0), .Y(men_men_n550_));
  NOi31      u0501(.An(men_men_n349_), .B(men_men_n550_), .C(men_men_n267_), .Y(men_men_n551_));
  NO4        u0502(.A(men_men_n551_), .B(men_men_n549_), .C(men_men_n540_), .D(men_men_n56_), .Y(men_men_n552_));
  NA2        u0503(.A(men_men_n552_), .B(men_men_n534_), .Y(men_men_n553_));
  NA3        u0504(.A(x8), .B(x7), .C(x0), .Y(men_men_n554_));
  INV        u0505(.A(men_men_n554_), .Y(men_men_n555_));
  AOI210     u0506(.A0(men_men_n277_), .A1(men_men_n99_), .B0(men_men_n555_), .Y(men_men_n556_));
  NO2        u0507(.A(men_men_n556_), .B(men_men_n159_), .Y(men_men_n557_));
  NA2        u0508(.A(men_men_n438_), .B(men_men_n57_), .Y(men_men_n558_));
  NO2        u0509(.A(x8), .B(x0), .Y(men_men_n559_));
  NA2        u0510(.A(men_men_n559_), .B(men_men_n368_), .Y(men_men_n560_));
  AOI210     u0511(.A0(men_men_n560_), .A1(men_men_n558_), .B0(men_men_n281_), .Y(men_men_n561_));
  OAI210     u0512(.A0(men_men_n561_), .A1(men_men_n557_), .B0(men_men_n285_), .Y(men_men_n562_));
  NO2        u0513(.A(men_men_n71_), .B(men_men_n110_), .Y(men_men_n563_));
  NO2        u0514(.A(men_men_n375_), .B(x8), .Y(men_men_n564_));
  NO2        u0515(.A(men_men_n564_), .B(men_men_n268_), .Y(men_men_n565_));
  NO3        u0516(.A(men_men_n565_), .B(men_men_n384_), .C(men_men_n274_), .Y(men_men_n566_));
  NO2        u0517(.A(men_men_n294_), .B(x8), .Y(men_men_n567_));
  OAI210     u0518(.A0(men_men_n469_), .A1(men_men_n332_), .B0(men_men_n249_), .Y(men_men_n568_));
  NA2        u0519(.A(men_men_n354_), .B(men_men_n181_), .Y(men_men_n569_));
  OAI220     u0520(.A0(men_men_n569_), .A1(men_men_n59_), .B0(men_men_n568_), .B1(men_men_n567_), .Y(men_men_n570_));
  OAI210     u0521(.A0(men_men_n570_), .A1(men_men_n566_), .B0(men_men_n563_), .Y(men_men_n571_));
  NO2        u0522(.A(x8), .B(x2), .Y(men_men_n572_));
  NO2        u0523(.A(men_men_n226_), .B(men_men_n57_), .Y(men_men_n573_));
  NA3        u0524(.A(men_men_n573_), .B(men_men_n572_), .C(men_men_n347_), .Y(men_men_n574_));
  NO2        u0525(.A(men_men_n250_), .B(men_men_n137_), .Y(men_men_n575_));
  AOI210     u0526(.A0(men_men_n328_), .A1(men_men_n167_), .B0(men_men_n575_), .Y(men_men_n576_));
  AOI210     u0527(.A0(men_men_n576_), .A1(men_men_n574_), .B0(men_men_n109_), .Y(men_men_n577_));
  NA2        u0528(.A(men_men_n344_), .B(x2), .Y(men_men_n578_));
  NO2        u0529(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n579_));
  NA2        u0530(.A(men_men_n579_), .B(men_men_n63_), .Y(men_men_n580_));
  AOI210     u0531(.A0(men_men_n578_), .A1(men_men_n464_), .B0(men_men_n580_), .Y(men_men_n581_));
  NA2        u0532(.A(men_men_n110_), .B(men_men_n53_), .Y(men_men_n582_));
  NO2        u0533(.A(men_men_n582_), .B(x8), .Y(men_men_n583_));
  NA2        u0534(.A(x7), .B(men_men_n50_), .Y(men_men_n584_));
  NO2        u0535(.A(men_men_n186_), .B(men_men_n584_), .Y(men_men_n585_));
  AN2        u0536(.A(men_men_n585_), .B(men_men_n583_), .Y(men_men_n586_));
  NA2        u0537(.A(men_men_n412_), .B(men_men_n152_), .Y(men_men_n587_));
  NO2        u0538(.A(men_men_n71_), .B(x2), .Y(men_men_n588_));
  NA2        u0539(.A(men_men_n588_), .B(men_men_n277_), .Y(men_men_n589_));
  OAI210     u0540(.A0(men_men_n589_), .A1(men_men_n587_), .B0(men_men_n56_), .Y(men_men_n590_));
  NO4        u0541(.A(men_men_n590_), .B(men_men_n586_), .C(men_men_n581_), .D(men_men_n577_), .Y(men_men_n591_));
  NA3        u0542(.A(men_men_n591_), .B(men_men_n571_), .C(men_men_n562_), .Y(men_men_n592_));
  NA2        u0543(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n593_));
  NOi21      u0544(.An(x2), .B(x7), .Y(men_men_n594_));
  NO2        u0545(.A(x6), .B(x3), .Y(men_men_n595_));
  NA2        u0546(.A(men_men_n595_), .B(men_men_n594_), .Y(men_men_n596_));
  NO2        u0547(.A(x6), .B(men_men_n59_), .Y(men_men_n597_));
  NO3        u0548(.A(men_men_n57_), .B(x2), .C(x1), .Y(men_men_n598_));
  NO3        u0549(.A(men_men_n57_), .B(x2), .C(x0), .Y(men_men_n599_));
  AOI220     u0550(.A0(men_men_n599_), .A1(men_men_n229_), .B0(men_men_n598_), .B1(men_men_n597_), .Y(men_men_n600_));
  OAI210     u0551(.A0(men_men_n596_), .A1(men_men_n593_), .B0(men_men_n600_), .Y(men_men_n601_));
  NO2        u0552(.A(men_men_n101_), .B(men_men_n53_), .Y(men_men_n602_));
  NA2        u0553(.A(men_men_n224_), .B(men_men_n57_), .Y(men_men_n603_));
  OAI210     u0554(.A0(men_men_n602_), .A1(men_men_n457_), .B0(men_men_n603_), .Y(men_men_n604_));
  NO3        u0555(.A(men_men_n604_), .B(men_men_n496_), .C(men_men_n59_), .Y(men_men_n605_));
  AO210      u0556(.A0(men_men_n601_), .A1(men_men_n469_), .B0(men_men_n605_), .Y(men_men_n606_));
  AOI210     u0557(.A0(men_men_n592_), .A1(men_men_n553_), .B0(men_men_n606_), .Y(men05));
  AOI210     u0558(.A0(men_men_n166_), .A1(men_men_n55_), .B0(men_men_n512_), .Y(men_men_n608_));
  OR2        u0559(.A(men_men_n608_), .B(men_men_n57_), .Y(men_men_n609_));
  NO2        u0560(.A(x7), .B(men_men_n108_), .Y(men_men_n610_));
  NO2        u0561(.A(x8), .B(men_men_n56_), .Y(men_men_n611_));
  NA2        u0562(.A(x5), .B(men_men_n56_), .Y(men_men_n612_));
  NO2        u0563(.A(men_men_n612_), .B(men_men_n584_), .Y(men_men_n613_));
  AOI210     u0564(.A0(men_men_n611_), .A1(men_men_n610_), .B0(men_men_n613_), .Y(men_men_n614_));
  AOI210     u0565(.A0(men_men_n614_), .A1(men_men_n609_), .B0(men_men_n110_), .Y(men_men_n615_));
  NO2        u0566(.A(x7), .B(x4), .Y(men_men_n616_));
  NO2        u0567(.A(men_men_n64_), .B(men_men_n55_), .Y(men_men_n617_));
  NO2        u0568(.A(men_men_n202_), .B(x5), .Y(men_men_n618_));
  NA2        u0569(.A(men_men_n108_), .B(men_men_n110_), .Y(men_men_n619_));
  NO2        u0570(.A(men_men_n619_), .B(men_men_n220_), .Y(men_men_n620_));
  AN2        u0571(.A(men_men_n620_), .B(men_men_n616_), .Y(men_men_n621_));
  OAI210     u0572(.A0(men_men_n621_), .A1(men_men_n615_), .B0(men_men_n500_), .Y(men_men_n622_));
  NO2        u0573(.A(x6), .B(men_men_n50_), .Y(men_men_n623_));
  NA2        u0574(.A(men_men_n55_), .B(x4), .Y(men_men_n624_));
  NO2        u0575(.A(men_men_n108_), .B(men_men_n110_), .Y(men_men_n625_));
  NA2        u0576(.A(men_men_n625_), .B(x7), .Y(men_men_n626_));
  NA2        u0577(.A(men_men_n441_), .B(men_men_n259_), .Y(men_men_n627_));
  AOI210     u0578(.A0(men_men_n627_), .A1(men_men_n626_), .B0(men_men_n624_), .Y(men_men_n628_));
  NA2        u0579(.A(men_men_n108_), .B(x4), .Y(men_men_n629_));
  XO2        u0580(.A(x7), .B(x5), .Y(men_men_n630_));
  NO2        u0581(.A(men_men_n630_), .B(men_men_n53_), .Y(men_men_n631_));
  NA3        u0582(.A(men_men_n631_), .B(men_men_n629_), .C(men_men_n333_), .Y(men_men_n632_));
  NO2        u0583(.A(men_men_n108_), .B(x2), .Y(men_men_n633_));
  NO2        u0584(.A(men_men_n75_), .B(men_men_n55_), .Y(men_men_n634_));
  NA2        u0585(.A(men_men_n634_), .B(men_men_n633_), .Y(men_men_n635_));
  NA2        u0586(.A(men_men_n635_), .B(men_men_n632_), .Y(men_men_n636_));
  OAI210     u0587(.A0(men_men_n636_), .A1(men_men_n628_), .B0(men_men_n623_), .Y(men_men_n637_));
  NO2        u0588(.A(men_men_n71_), .B(men_men_n50_), .Y(men_men_n638_));
  NO2        u0589(.A(men_men_n196_), .B(x4), .Y(men_men_n639_));
  NO2        u0590(.A(x5), .B(men_men_n56_), .Y(men_men_n640_));
  XO2        u0591(.A(x5), .B(x2), .Y(men_men_n641_));
  NO3        u0592(.A(x8), .B(x7), .C(men_men_n110_), .Y(men_men_n642_));
  AO220      u0593(.A0(men_men_n642_), .A1(men_men_n640_), .B0(men_men_n641_), .B1(men_men_n639_), .Y(men_men_n643_));
  NA3        u0594(.A(men_men_n643_), .B(men_men_n638_), .C(men_men_n53_), .Y(men_men_n644_));
  NA2        u0595(.A(men_men_n274_), .B(men_men_n594_), .Y(men_men_n645_));
  NOi21      u0596(.An(x4), .B(x1), .Y(men_men_n646_));
  NA2        u0597(.A(men_men_n646_), .B(men_men_n63_), .Y(men_men_n647_));
  NA2        u0598(.A(x4), .B(x1), .Y(men_men_n648_));
  NO2        u0599(.A(men_men_n648_), .B(men_men_n50_), .Y(men_men_n649_));
  AOI210     u0600(.A0(men_men_n649_), .A1(men_men_n625_), .B0(men_men_n59_), .Y(men_men_n650_));
  OA210      u0601(.A0(men_men_n647_), .A1(men_men_n645_), .B0(men_men_n650_), .Y(men_men_n651_));
  NA4        u0602(.A(men_men_n651_), .B(men_men_n644_), .C(men_men_n637_), .D(men_men_n622_), .Y(men_men_n652_));
  NA2        u0603(.A(men_men_n638_), .B(men_men_n56_), .Y(men_men_n653_));
  NA2        u0604(.A(men_men_n572_), .B(men_men_n610_), .Y(men_men_n654_));
  NO2        u0605(.A(men_men_n654_), .B(men_men_n653_), .Y(men_men_n655_));
  NA2        u0606(.A(men_men_n277_), .B(men_men_n123_), .Y(men_men_n656_));
  OAI210     u0607(.A0(men_men_n656_), .A1(men_men_n168_), .B0(men_men_n59_), .Y(men_men_n657_));
  NA2        u0608(.A(men_men_n57_), .B(x6), .Y(men_men_n658_));
  AOI210     u0609(.A0(men_men_n658_), .A1(x3), .B0(men_men_n91_), .Y(men_men_n659_));
  NA2        u0610(.A(men_men_n640_), .B(men_men_n158_), .Y(men_men_n660_));
  NO3        u0611(.A(men_men_n660_), .B(men_men_n659_), .C(men_men_n431_), .Y(men_men_n661_));
  NA2        u0612(.A(men_men_n286_), .B(men_men_n71_), .Y(men_men_n662_));
  NO2        u0613(.A(men_men_n392_), .B(x3), .Y(men_men_n663_));
  NA2        u0614(.A(men_men_n663_), .B(men_men_n243_), .Y(men_men_n664_));
  NO2        u0615(.A(men_men_n431_), .B(men_men_n639_), .Y(men_men_n665_));
  NO2        u0616(.A(men_men_n473_), .B(men_men_n108_), .Y(men_men_n666_));
  NO2        u0617(.A(men_men_n582_), .B(x6), .Y(men_men_n667_));
  NA2        u0618(.A(men_men_n667_), .B(men_men_n666_), .Y(men_men_n668_));
  OAI220     u0619(.A0(men_men_n668_), .A1(men_men_n665_), .B0(men_men_n664_), .B1(men_men_n662_), .Y(men_men_n669_));
  NO4        u0620(.A(men_men_n669_), .B(men_men_n661_), .C(men_men_n657_), .D(men_men_n655_), .Y(men_men_n670_));
  NA2        u0621(.A(men_men_n57_), .B(x5), .Y(men_men_n671_));
  NO2        u0622(.A(men_men_n671_), .B(x1), .Y(men_men_n672_));
  NA2        u0623(.A(x8), .B(men_men_n56_), .Y(men_men_n673_));
  NO2        u0624(.A(men_men_n673_), .B(men_men_n132_), .Y(men_men_n674_));
  NA2        u0625(.A(x8), .B(x4), .Y(men_men_n675_));
  NO2        u0626(.A(x8), .B(x4), .Y(men_men_n676_));
  NAi21      u0627(.An(men_men_n676_), .B(men_men_n675_), .Y(men_men_n677_));
  NAi21      u0628(.An(men_men_n572_), .B(men_men_n392_), .Y(men_men_n678_));
  NO4        u0629(.A(men_men_n678_), .B(men_men_n677_), .C(men_men_n431_), .D(men_men_n71_), .Y(men_men_n679_));
  OAI210     u0630(.A0(men_men_n679_), .A1(men_men_n674_), .B0(men_men_n672_), .Y(men_men_n680_));
  NO3        u0631(.A(x8), .B(men_men_n108_), .C(x4), .Y(men_men_n681_));
  INV        u0632(.A(men_men_n681_), .Y(men_men_n682_));
  NO2        u0633(.A(men_men_n682_), .B(men_men_n110_), .Y(men_men_n683_));
  NO2        u0634(.A(x5), .B(x4), .Y(men_men_n684_));
  NA3        u0635(.A(men_men_n684_), .B(men_men_n63_), .C(men_men_n110_), .Y(men_men_n685_));
  NO2        u0636(.A(x6), .B(men_men_n110_), .Y(men_men_n686_));
  NA2        u0637(.A(men_men_n673_), .B(men_men_n686_), .Y(men_men_n687_));
  OAI210     u0638(.A0(men_men_n687_), .A1(men_men_n531_), .B0(men_men_n685_), .Y(men_men_n688_));
  OAI210     u0639(.A0(men_men_n688_), .A1(men_men_n683_), .B0(men_men_n316_), .Y(men_men_n689_));
  NA3        u0640(.A(men_men_n689_), .B(men_men_n680_), .C(men_men_n670_), .Y(men_men_n690_));
  OR2        u0641(.A(x4), .B(x1), .Y(men_men_n691_));
  NO2        u0642(.A(men_men_n691_), .B(x3), .Y(men_men_n692_));
  NA2        u0643(.A(men_men_n55_), .B(x2), .Y(men_men_n693_));
  NO3        u0644(.A(men_men_n373_), .B(men_men_n693_), .C(x6), .Y(men_men_n694_));
  AOI220     u0645(.A0(men_men_n694_), .A1(men_men_n692_), .B0(men_men_n690_), .B1(men_men_n652_), .Y(men06));
  NA2        u0646(.A(men_men_n56_), .B(x3), .Y(men_men_n696_));
  NA2        u0647(.A(x6), .B(men_men_n110_), .Y(men_men_n697_));
  NA2        u0648(.A(men_men_n697_), .B(men_men_n55_), .Y(men_men_n698_));
  NA2        u0649(.A(x5), .B(men_men_n59_), .Y(men_men_n699_));
  NO2        u0650(.A(men_men_n699_), .B(men_men_n118_), .Y(men_men_n700_));
  NA3        u0651(.A(men_men_n700_), .B(men_men_n698_), .C(men_men_n506_), .Y(men_men_n701_));
  NO2        u0652(.A(men_men_n392_), .B(x0), .Y(men_men_n702_));
  NA2        u0653(.A(men_men_n343_), .B(x2), .Y(men_men_n703_));
  NOi21      u0654(.An(x6), .B(x8), .Y(men_men_n704_));
  NO2        u0655(.A(men_men_n704_), .B(x2), .Y(men_men_n705_));
  NO3        u0656(.A(men_men_n705_), .B(men_men_n70_), .C(men_men_n59_), .Y(men_men_n706_));
  AOI220     u0657(.A0(men_men_n706_), .A1(men_men_n703_), .B0(men_men_n702_), .B1(men_men_n335_), .Y(men_men_n707_));
  AOI210     u0658(.A0(men_men_n707_), .A1(men_men_n701_), .B0(men_men_n696_), .Y(men_men_n708_));
  NA2        u0659(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n709_));
  NA2        u0660(.A(men_men_n371_), .B(men_men_n359_), .Y(men_men_n710_));
  NO2        u0661(.A(men_men_n71_), .B(men_men_n108_), .Y(men_men_n711_));
  NO2        u0662(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n712_));
  NO4        u0663(.A(men_men_n712_), .B(men_men_n693_), .C(men_men_n711_), .D(men_men_n500_), .Y(men_men_n713_));
  AOI220     u0664(.A0(men_men_n713_), .A1(men_men_n710_), .B0(men_men_n428_), .B1(men_men_n63_), .Y(men_men_n714_));
  NO2        u0665(.A(men_men_n714_), .B(men_men_n709_), .Y(men_men_n715_));
  NO2        u0666(.A(men_men_n54_), .B(x0), .Y(men_men_n716_));
  NA2        u0667(.A(x4), .B(x3), .Y(men_men_n717_));
  NO2        u0668(.A(men_men_n104_), .B(men_men_n56_), .Y(men_men_n718_));
  INV        u0669(.A(men_men_n388_), .Y(men_men_n719_));
  NO2        u0670(.A(men_men_n415_), .B(x8), .Y(men_men_n720_));
  NO2        u0671(.A(men_men_n261_), .B(men_men_n526_), .Y(men_men_n721_));
  AOI210     u0672(.A0(men_men_n720_), .A1(men_men_n269_), .B0(men_men_n721_), .Y(men_men_n722_));
  NO2        u0673(.A(x5), .B(x3), .Y(men_men_n723_));
  NA3        u0674(.A(men_men_n559_), .B(men_men_n723_), .C(x1), .Y(men_men_n724_));
  NA2        u0675(.A(men_men_n611_), .B(men_men_n563_), .Y(men_men_n725_));
  OA220      u0676(.A0(men_men_n725_), .A1(men_men_n587_), .B0(men_men_n724_), .B1(men_men_n506_), .Y(men_men_n726_));
  OAI210     u0677(.A0(men_men_n722_), .A1(men_men_n719_), .B0(men_men_n726_), .Y(men_men_n727_));
  OR3        u0678(.A(men_men_n727_), .B(men_men_n715_), .C(men_men_n708_), .Y(men_men_n728_));
  NA2        u0679(.A(x7), .B(men_men_n56_), .Y(men_men_n729_));
  NO2        u0680(.A(men_men_n625_), .B(men_men_n59_), .Y(men_men_n730_));
  NA2        u0681(.A(men_men_n730_), .B(men_men_n638_), .Y(men_men_n731_));
  NO2        u0682(.A(men_men_n174_), .B(x6), .Y(men_men_n732_));
  NA2        u0683(.A(men_men_n732_), .B(men_men_n295_), .Y(men_men_n733_));
  AOI210     u0684(.A0(men_men_n733_), .A1(men_men_n731_), .B0(men_men_n729_), .Y(men_men_n734_));
  AN2        u0685(.A(men_men_n478_), .B(men_men_n325_), .Y(men_men_n735_));
  OAI210     u0686(.A0(men_men_n735_), .A1(men_men_n734_), .B0(men_men_n354_), .Y(men_men_n736_));
  NO2        u0687(.A(men_men_n312_), .B(men_men_n108_), .Y(men_men_n737_));
  NO2        u0688(.A(men_men_n56_), .B(x3), .Y(men_men_n738_));
  NA2        u0689(.A(men_men_n738_), .B(men_men_n71_), .Y(men_men_n739_));
  NO2        u0690(.A(men_men_n739_), .B(men_men_n255_), .Y(men_men_n740_));
  NO2        u0691(.A(men_men_n71_), .B(x3), .Y(men_men_n741_));
  NA3        u0692(.A(men_men_n741_), .B(men_men_n579_), .C(men_men_n56_), .Y(men_men_n742_));
  NO2        u0693(.A(men_men_n57_), .B(x6), .Y(men_men_n743_));
  NA2        u0694(.A(men_men_n185_), .B(men_men_n743_), .Y(men_men_n744_));
  NA3        u0695(.A(men_men_n611_), .B(men_men_n332_), .C(men_men_n71_), .Y(men_men_n745_));
  NA3        u0696(.A(men_men_n745_), .B(men_men_n744_), .C(men_men_n742_), .Y(men_men_n746_));
  OR3        u0697(.A(men_men_n746_), .B(men_men_n740_), .C(men_men_n649_), .Y(men_men_n747_));
  NA2        u0698(.A(men_men_n747_), .B(men_men_n737_), .Y(men_men_n748_));
  NA2        u0699(.A(men_men_n716_), .B(men_men_n638_), .Y(men_men_n749_));
  NA4        u0700(.A(men_men_n270_), .B(men_men_n595_), .C(men_men_n224_), .D(men_men_n262_), .Y(men_men_n750_));
  NA2        u0701(.A(men_men_n489_), .B(men_men_n67_), .Y(men_men_n751_));
  AOI210     u0702(.A0(men_men_n750_), .A1(men_men_n749_), .B0(men_men_n751_), .Y(men_men_n752_));
  NA2        u0703(.A(x7), .B(x6), .Y(men_men_n753_));
  NA3        u0704(.A(x2), .B(x1), .C(x0), .Y(men_men_n754_));
  NO3        u0705(.A(men_men_n754_), .B(men_men_n753_), .C(men_men_n608_), .Y(men_men_n755_));
  NA2        u0706(.A(men_men_n501_), .B(men_men_n151_), .Y(men_men_n756_));
  NO2        u0707(.A(x5), .B(x1), .Y(men_men_n757_));
  NA2        u0708(.A(men_men_n757_), .B(men_men_n743_), .Y(men_men_n758_));
  NA2        u0709(.A(x4), .B(x0), .Y(men_men_n759_));
  NO3        u0710(.A(men_men_n57_), .B(x6), .C(x2), .Y(men_men_n760_));
  NA2        u0711(.A(men_men_n760_), .B(men_men_n228_), .Y(men_men_n761_));
  OAI220     u0712(.A0(men_men_n761_), .A1(men_men_n759_), .B0(men_men_n758_), .B1(men_men_n756_), .Y(men_men_n762_));
  NO3        u0713(.A(men_men_n762_), .B(men_men_n755_), .C(men_men_n752_), .Y(men_men_n763_));
  NA3        u0714(.A(men_men_n763_), .B(men_men_n748_), .C(men_men_n736_), .Y(men_men_n764_));
  AOI210     u0715(.A0(men_men_n728_), .A1(men_men_n57_), .B0(men_men_n764_), .Y(men07));
  NA2        u0716(.A(men_men_n108_), .B(men_men_n59_), .Y(men_men_n766_));
  NOi21      u0717(.An(men_men_n753_), .B(men_men_n116_), .Y(men_men_n767_));
  NO4        u0718(.A(men_men_n767_), .B(men_men_n638_), .C(men_men_n255_), .D(men_men_n766_), .Y(men_men_n768_));
  NO3        u0719(.A(men_men_n57_), .B(x5), .C(x1), .Y(men_men_n769_));
  NA2        u0720(.A(men_men_n769_), .B(men_men_n379_), .Y(men_men_n770_));
  NO2        u0721(.A(men_men_n57_), .B(men_men_n71_), .Y(men_men_n771_));
  NO2        u0722(.A(men_men_n157_), .B(men_men_n109_), .Y(men_men_n772_));
  AOI210     u0723(.A0(men_men_n771_), .A1(men_men_n92_), .B0(men_men_n772_), .Y(men_men_n773_));
  NO2        u0724(.A(men_men_n773_), .B(men_men_n137_), .Y(men_men_n774_));
  OAI210     u0725(.A0(men_men_n774_), .A1(men_men_n768_), .B0(x2), .Y(men_men_n775_));
  NAi21      u0726(.An(men_men_n158_), .B(men_men_n159_), .Y(men_men_n776_));
  NA3        u0727(.A(men_men_n776_), .B(men_men_n91_), .C(x3), .Y(men_men_n777_));
  NO3        u0728(.A(men_men_n55_), .B(x3), .C(x1), .Y(men_men_n778_));
  NO2        u0729(.A(men_men_n519_), .B(x2), .Y(men_men_n779_));
  AOI210     u0730(.A0(men_men_n779_), .A1(men_men_n521_), .B0(men_men_n778_), .Y(men_men_n780_));
  OAI210     u0731(.A0(men_men_n780_), .A1(men_men_n658_), .B0(men_men_n777_), .Y(men_men_n781_));
  NO2        u0732(.A(x8), .B(men_men_n53_), .Y(men_men_n782_));
  NA2        u0733(.A(men_men_n782_), .B(men_men_n59_), .Y(men_men_n783_));
  NO2        u0734(.A(x7), .B(x3), .Y(men_men_n784_));
  NA2        u0735(.A(men_men_n784_), .B(men_men_n101_), .Y(men_men_n785_));
  NO2        u0736(.A(men_men_n783_), .B(men_men_n785_), .Y(men_men_n786_));
  AOI210     u0737(.A0(men_men_n781_), .A1(men_men_n254_), .B0(men_men_n786_), .Y(men_men_n787_));
  AOI210     u0738(.A0(men_men_n787_), .A1(men_men_n775_), .B0(x4), .Y(men_men_n788_));
  NA3        u0739(.A(men_men_n757_), .B(men_men_n323_), .C(men_men_n55_), .Y(men_men_n789_));
  AOI210     u0740(.A0(men_men_n789_), .A1(men_men_n604_), .B0(men_men_n110_), .Y(men_men_n790_));
  XO2        u0741(.A(x5), .B(x1), .Y(men_men_n791_));
  NO4        u0742(.A(men_men_n791_), .B(men_men_n167_), .C(men_men_n211_), .D(men_men_n55_), .Y(men_men_n792_));
  OAI210     u0743(.A0(men_men_n792_), .A1(men_men_n790_), .B0(men_men_n419_), .Y(men_men_n793_));
  NO3        u0744(.A(men_men_n50_), .B(x2), .C(x0), .Y(men_men_n794_));
  NO2        u0745(.A(men_men_n315_), .B(men_men_n108_), .Y(men_men_n795_));
  NA2        u0746(.A(x6), .B(x0), .Y(men_men_n796_));
  NO2        u0747(.A(men_men_n693_), .B(men_men_n796_), .Y(men_men_n797_));
  NO2        u0748(.A(men_men_n791_), .B(men_men_n704_), .Y(men_men_n798_));
  OAI210     u0749(.A0(men_men_n757_), .A1(men_men_n63_), .B0(men_men_n57_), .Y(men_men_n799_));
  OAI210     u0750(.A0(men_men_n799_), .A1(men_men_n798_), .B0(men_men_n770_), .Y(men_men_n800_));
  AOI220     u0751(.A0(men_men_n800_), .A1(men_men_n794_), .B0(men_men_n797_), .B1(men_men_n795_), .Y(men_men_n801_));
  AOI210     u0752(.A0(men_men_n801_), .A1(men_men_n793_), .B0(men_men_n56_), .Y(men_men_n802_));
  NOi21      u0753(.An(men_men_n235_), .B(men_men_n379_), .Y(men_men_n803_));
  NO3        u0754(.A(men_men_n803_), .B(men_men_n244_), .C(men_men_n67_), .Y(men_men_n804_));
  NO2        u0755(.A(men_men_n194_), .B(men_men_n71_), .Y(men_men_n805_));
  NO2        u0756(.A(men_men_n315_), .B(x6), .Y(men_men_n806_));
  AO220      u0757(.A0(men_men_n806_), .A1(men_men_n333_), .B0(men_men_n805_), .B1(men_men_n564_), .Y(men_men_n807_));
  OAI210     u0758(.A0(men_men_n807_), .A1(men_men_n804_), .B0(men_men_n59_), .Y(men_men_n808_));
  NA2        u0759(.A(men_men_n92_), .B(men_men_n71_), .Y(men_men_n809_));
  NO2        u0760(.A(men_men_n809_), .B(men_men_n654_), .Y(men_men_n810_));
  NAi21      u0761(.An(x8), .B(x7), .Y(men_men_n811_));
  NA2        u0762(.A(men_men_n803_), .B(men_men_n811_), .Y(men_men_n812_));
  NA2        u0763(.A(men_men_n412_), .B(men_men_n110_), .Y(men_men_n813_));
  NO2        u0764(.A(men_men_n704_), .B(x1), .Y(men_men_n814_));
  NO3        u0765(.A(men_men_n814_), .B(men_men_n813_), .C(men_men_n579_), .Y(men_men_n815_));
  AOI210     u0766(.A0(men_men_n815_), .A1(men_men_n812_), .B0(men_men_n810_), .Y(men_men_n816_));
  AOI210     u0767(.A0(men_men_n816_), .A1(men_men_n808_), .B0(men_men_n144_), .Y(men_men_n817_));
  NO2        u0768(.A(x8), .B(x7), .Y(men_men_n818_));
  NO2        u0769(.A(men_men_n818_), .B(x3), .Y(men_men_n819_));
  NA3        u0770(.A(men_men_n819_), .B(men_men_n368_), .C(x1), .Y(men_men_n820_));
  NO2        u0771(.A(x8), .B(men_men_n110_), .Y(men_men_n821_));
  AOI220     u0772(.A0(men_men_n332_), .A1(men_men_n354_), .B0(men_men_n821_), .B1(men_men_n259_), .Y(men_men_n822_));
  NO2        u0773(.A(men_men_n71_), .B(x4), .Y(men_men_n823_));
  NA2        u0774(.A(men_men_n823_), .B(men_men_n309_), .Y(men_men_n824_));
  AOI210     u0775(.A0(men_men_n822_), .A1(men_men_n820_), .B0(men_men_n824_), .Y(men_men_n825_));
  NO4        u0776(.A(men_men_n825_), .B(men_men_n817_), .C(men_men_n802_), .D(men_men_n788_), .Y(men08));
  NA2        u0777(.A(men_men_n50_), .B(x1), .Y(men_men_n827_));
  XN2        u0778(.A(x5), .B(x4), .Y(men_men_n828_));
  INV        u0779(.A(men_men_n828_), .Y(men_men_n829_));
  AOI220     u0780(.A0(men_men_n829_), .A1(men_men_n360_), .B0(men_men_n140_), .B1(men_men_n56_), .Y(men_men_n830_));
  NO2        u0781(.A(men_men_n246_), .B(men_men_n108_), .Y(men_men_n831_));
  AOI210     u0782(.A0(men_men_n831_), .A1(men_men_n283_), .B0(men_men_n195_), .Y(men_men_n832_));
  OAI220     u0783(.A0(men_men_n832_), .A1(x4), .B0(men_men_n830_), .B1(men_men_n827_), .Y(men_men_n833_));
  NA2        u0784(.A(men_men_n833_), .B(men_men_n277_), .Y(men_men_n834_));
  AOI210     u0785(.A0(men_men_n276_), .A1(men_men_n813_), .B0(men_men_n624_), .Y(men_men_n835_));
  NA2        u0786(.A(men_men_n619_), .B(men_men_n174_), .Y(men_men_n836_));
  OAI220     u0787(.A0(men_men_n836_), .A1(men_men_n673_), .B0(men_men_n491_), .B1(men_men_n50_), .Y(men_men_n837_));
  AO210      u0788(.A0(men_men_n837_), .A1(men_men_n347_), .B0(men_men_n835_), .Y(men_men_n838_));
  NA2        u0789(.A(men_men_n283_), .B(men_men_n151_), .Y(men_men_n839_));
  NA2        u0790(.A(men_men_n144_), .B(x7), .Y(men_men_n840_));
  OR3        u0791(.A(men_men_n754_), .B(men_men_n473_), .C(men_men_n723_), .Y(men_men_n841_));
  OAI220     u0792(.A0(men_men_n841_), .A1(men_men_n840_), .B0(men_men_n839_), .B1(men_men_n208_), .Y(men_men_n842_));
  AOI210     u0793(.A0(men_men_n838_), .A1(men_men_n297_), .B0(men_men_n842_), .Y(men_men_n843_));
  AOI210     u0794(.A0(men_men_n843_), .A1(men_men_n834_), .B0(men_men_n71_), .Y(men_men_n844_));
  NO2        u0795(.A(men_men_n818_), .B(men_men_n110_), .Y(men_men_n845_));
  NA2        u0796(.A(men_men_n845_), .B(men_men_n196_), .Y(men_men_n846_));
  OAI210     u0797(.A0(men_men_n415_), .A1(men_men_n309_), .B0(men_men_n347_), .Y(men_men_n847_));
  NA2        u0798(.A(men_men_n441_), .B(men_men_n237_), .Y(men_men_n848_));
  NA2        u0799(.A(men_men_n720_), .B(men_men_n107_), .Y(men_men_n849_));
  OAI220     u0800(.A0(men_men_n849_), .A1(men_men_n848_), .B0(men_men_n847_), .B1(men_men_n846_), .Y(men_men_n850_));
  NA2        u0801(.A(men_men_n850_), .B(men_men_n293_), .Y(men_men_n851_));
  NA2        u0802(.A(men_men_n337_), .B(men_men_n53_), .Y(men_men_n852_));
  NO3        u0803(.A(men_men_n415_), .B(men_men_n137_), .C(men_men_n68_), .Y(men_men_n853_));
  NO2        u0804(.A(men_men_n712_), .B(men_men_n249_), .Y(men_men_n854_));
  NO3        u0805(.A(men_men_n573_), .B(men_men_n474_), .C(men_men_n99_), .Y(men_men_n855_));
  AO220      u0806(.A0(men_men_n855_), .A1(men_men_n854_), .B0(men_men_n853_), .B1(men_men_n852_), .Y(men_men_n856_));
  NA2        u0807(.A(x7), .B(men_men_n59_), .Y(men_men_n857_));
  NO3        u0808(.A(men_men_n318_), .B(men_men_n857_), .C(men_men_n292_), .Y(men_men_n858_));
  AOI210     u0809(.A0(men_men_n856_), .A1(x5), .B0(men_men_n858_), .Y(men_men_n859_));
  AOI210     u0810(.A0(men_men_n859_), .A1(men_men_n851_), .B0(men_men_n72_), .Y(men_men_n860_));
  NO2        u0811(.A(men_men_n70_), .B(x3), .Y(men_men_n861_));
  OAI210     u0812(.A0(men_men_n861_), .A1(men_men_n268_), .B0(men_men_n149_), .Y(men_men_n862_));
  MUX2       u0813(.S(x3), .A(men_men_n167_), .B(men_men_n776_), .Y(men_men_n863_));
  NA2        u0814(.A(men_men_n863_), .B(men_men_n564_), .Y(men_men_n864_));
  NO3        u0815(.A(x6), .B(x4), .C(x0), .Y(men_men_n865_));
  INV        u0816(.A(men_men_n865_), .Y(men_men_n866_));
  AOI210     u0817(.A0(men_men_n864_), .A1(men_men_n862_), .B0(men_men_n866_), .Y(men_men_n867_));
  NO3        u0818(.A(x5), .B(x3), .C(men_men_n110_), .Y(men_men_n868_));
  AOI220     u0819(.A0(men_men_n829_), .A1(men_men_n314_), .B0(men_men_n868_), .B1(men_men_n59_), .Y(men_men_n869_));
  OR2        u0820(.A(x8), .B(x1), .Y(men_men_n870_));
  NO3        u0821(.A(men_men_n870_), .B(men_men_n869_), .C(men_men_n738_), .Y(men_men_n871_));
  NAi21      u0822(.An(x4), .B(x1), .Y(men_men_n872_));
  NO2        u0823(.A(men_men_n872_), .B(x0), .Y(men_men_n873_));
  NA2        u0824(.A(men_men_n618_), .B(men_men_n873_), .Y(men_men_n874_));
  NA3        u0825(.A(men_men_n55_), .B(x1), .C(x0), .Y(men_men_n875_));
  OAI210     u0826(.A0(men_men_n875_), .A1(men_men_n719_), .B0(men_men_n874_), .Y(men_men_n876_));
  OAI210     u0827(.A0(men_men_n876_), .A1(men_men_n871_), .B0(men_men_n323_), .Y(men_men_n877_));
  AO210      u0828(.A0(men_men_n295_), .A1(men_men_n268_), .B0(men_men_n737_), .Y(men_men_n878_));
  NA2        u0829(.A(men_men_n108_), .B(men_men_n56_), .Y(men_men_n879_));
  NO2        u0830(.A(men_men_n57_), .B(x2), .Y(men_men_n880_));
  NA2        u0831(.A(men_men_n878_), .B(men_men_n649_), .Y(men_men_n881_));
  NA2        u0832(.A(men_men_n881_), .B(men_men_n877_), .Y(men_men_n882_));
  NO4        u0833(.A(men_men_n882_), .B(men_men_n867_), .C(men_men_n860_), .D(men_men_n844_), .Y(men09));
  NO3        u0834(.A(men_men_n791_), .B(men_men_n121_), .C(men_men_n96_), .Y(men_men_n884_));
  AOI220     u0835(.A0(men_men_n304_), .A1(men_men_n70_), .B0(men_men_n594_), .B1(men_men_n546_), .Y(men_men_n885_));
  OAI210     u0836(.A0(men_men_n884_), .A1(x2), .B0(men_men_n885_), .Y(men_men_n886_));
  AOI210     u0837(.A0(men_men_n886_), .A1(men_men_n758_), .B0(men_men_n450_), .Y(men_men_n887_));
  NO2        u0838(.A(men_men_n593_), .B(men_men_n267_), .Y(men_men_n888_));
  NO2        u0839(.A(men_men_n757_), .B(men_men_n343_), .Y(men_men_n889_));
  NO3        u0840(.A(men_men_n610_), .B(men_men_n102_), .C(men_men_n110_), .Y(men_men_n890_));
  AO220      u0841(.A0(men_men_n890_), .A1(men_men_n889_), .B0(men_men_n888_), .B1(men_men_n625_), .Y(men_men_n891_));
  OAI210     u0842(.A0(men_men_n891_), .A1(men_men_n887_), .B0(x4), .Y(men_men_n892_));
  OAI220     u0843(.A0(men_men_n371_), .A1(men_men_n146_), .B0(men_men_n399_), .B1(men_men_n285_), .Y(men_men_n893_));
  NO2        u0844(.A(men_men_n194_), .B(men_men_n108_), .Y(men_men_n894_));
  AOI220     u0845(.A0(men_men_n894_), .A1(men_men_n126_), .B0(men_men_n893_), .B1(men_men_n631_), .Y(men_men_n895_));
  NO2        u0846(.A(men_men_n791_), .B(men_men_n96_), .Y(men_men_n896_));
  NAi21      u0847(.An(x0), .B(x2), .Y(men_men_n897_));
  NO2        u0848(.A(men_men_n308_), .B(men_men_n897_), .Y(men_men_n898_));
  OAI210     u0849(.A0(men_men_n483_), .A1(men_men_n280_), .B0(men_men_n194_), .Y(men_men_n899_));
  AOI210     u0850(.A0(men_men_n170_), .A1(men_men_n811_), .B0(men_men_n359_), .Y(men_men_n900_));
  AOI220     u0851(.A0(men_men_n900_), .A1(men_men_n899_), .B0(men_men_n898_), .B1(men_men_n896_), .Y(men_men_n901_));
  OAI210     u0852(.A0(men_men_n895_), .A1(men_men_n55_), .B0(men_men_n901_), .Y(men_men_n902_));
  NA2        u0853(.A(men_men_n902_), .B(men_men_n56_), .Y(men_men_n903_));
  NO2        u0854(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n904_));
  INV        u0855(.A(men_men_n126_), .Y(men_men_n905_));
  NA2        u0856(.A(men_men_n757_), .B(men_men_n55_), .Y(men_men_n906_));
  AOI210     u0857(.A0(x6), .A1(x1), .B0(x5), .Y(men_men_n907_));
  OAI210     u0858(.A0(men_men_n907_), .A1(men_men_n336_), .B0(x2), .Y(men_men_n908_));
  AOI210     u0859(.A0(men_men_n908_), .A1(men_men_n906_), .B0(men_men_n905_), .Y(men_men_n909_));
  NA2        u0860(.A(men_men_n563_), .B(men_men_n55_), .Y(men_men_n910_));
  NO4        u0861(.A(men_men_n57_), .B(x6), .C(x5), .D(x1), .Y(men_men_n911_));
  NO2        u0862(.A(men_men_n234_), .B(men_men_n389_), .Y(men_men_n912_));
  NO2        u0863(.A(men_men_n315_), .B(men_men_n150_), .Y(men_men_n913_));
  NO3        u0864(.A(men_men_n913_), .B(men_men_n912_), .C(men_men_n911_), .Y(men_men_n914_));
  OAI220     u0865(.A0(men_men_n914_), .A1(men_men_n55_), .B0(men_men_n910_), .B1(men_men_n462_), .Y(men_men_n915_));
  OAI210     u0866(.A0(men_men_n915_), .A1(men_men_n909_), .B0(men_men_n904_), .Y(men_men_n916_));
  NO2        u0867(.A(men_men_n408_), .B(men_men_n108_), .Y(men_men_n917_));
  NO2        u0868(.A(men_men_n337_), .B(men_men_n500_), .Y(men_men_n918_));
  AOI220     u0869(.A0(men_men_n918_), .A1(men_men_n917_), .B0(men_men_n212_), .B1(men_men_n232_), .Y(men_men_n919_));
  NA4        u0870(.A(men_men_n919_), .B(men_men_n916_), .C(men_men_n903_), .D(men_men_n892_), .Y(men_men_n920_));
  NA2        u0871(.A(men_men_n920_), .B(men_men_n50_), .Y(men_men_n921_));
  NO2        u0872(.A(men_men_n382_), .B(men_men_n163_), .Y(men_men_n922_));
  NA2        u0873(.A(men_men_n243_), .B(men_men_n594_), .Y(men_men_n923_));
  OAI210     u0874(.A0(men_men_n436_), .A1(men_men_n821_), .B0(men_men_n923_), .Y(men_men_n924_));
  OAI210     u0875(.A0(men_men_n924_), .A1(men_men_n922_), .B0(x0), .Y(men_men_n925_));
  NO3        u0876(.A(x8), .B(x7), .C(x2), .Y(men_men_n926_));
  NO3        u0877(.A(men_men_n57_), .B(x5), .C(x2), .Y(men_men_n927_));
  OAI210     u0878(.A0(men_men_n927_), .A1(men_men_n926_), .B0(men_men_n521_), .Y(men_men_n928_));
  AOI210     u0879(.A0(men_men_n928_), .A1(men_men_n925_), .B0(x4), .Y(men_men_n929_));
  NO2        u0880(.A(men_men_n429_), .B(men_men_n149_), .Y(men_men_n930_));
  NO2        u0881(.A(men_men_n52_), .B(x2), .Y(men_men_n931_));
  NO2        u0882(.A(men_men_n108_), .B(men_men_n56_), .Y(men_men_n932_));
  NA2        u0883(.A(men_men_n932_), .B(x8), .Y(men_men_n933_));
  NA2        u0884(.A(men_men_n933_), .B(men_men_n906_), .Y(men_men_n934_));
  AO210      u0885(.A0(men_men_n934_), .A1(men_men_n931_), .B0(men_men_n930_), .Y(men_men_n935_));
  OAI210     u0886(.A0(men_men_n935_), .A1(men_men_n929_), .B0(men_men_n623_), .Y(men_men_n936_));
  NO2        u0887(.A(men_men_n263_), .B(men_men_n119_), .Y(men_men_n937_));
  OAI210     u0888(.A0(x4), .A1(x2), .B0(x0), .Y(men_men_n938_));
  NA3        u0889(.A(men_men_n612_), .B(men_men_n624_), .C(men_men_n348_), .Y(men_men_n939_));
  OAI210     u0890(.A0(men_men_n938_), .A1(men_men_n292_), .B0(men_men_n53_), .Y(men_men_n940_));
  AOI210     u0891(.A0(men_men_n939_), .A1(men_men_n938_), .B0(men_men_n940_), .Y(men_men_n941_));
  OAI210     u0892(.A0(men_men_n941_), .A1(men_men_n937_), .B0(men_men_n332_), .Y(men_men_n942_));
  AOI220     u0893(.A0(men_men_n675_), .A1(men_men_n352_), .B0(men_men_n354_), .B1(men_men_n93_), .Y(men_men_n943_));
  NA2        u0894(.A(men_men_n93_), .B(x5), .Y(men_men_n944_));
  OAI220     u0895(.A0(men_men_n944_), .A1(men_men_n870_), .B0(men_men_n943_), .B1(men_men_n324_), .Y(men_men_n945_));
  NA2        u0896(.A(men_men_n945_), .B(men_men_n68_), .Y(men_men_n946_));
  NA2        u0897(.A(men_men_n412_), .B(men_men_n776_), .Y(men_men_n947_));
  NA2        u0898(.A(men_men_n254_), .B(men_men_n167_), .Y(men_men_n948_));
  AO210      u0899(.A0(men_men_n948_), .A1(men_men_n947_), .B0(men_men_n134_), .Y(men_men_n949_));
  NO2        u0900(.A(men_men_n442_), .B(x2), .Y(men_men_n950_));
  NO2        u0901(.A(x7), .B(men_men_n53_), .Y(men_men_n951_));
  NA2        u0902(.A(men_men_n951_), .B(x5), .Y(men_men_n952_));
  NO2        u0903(.A(men_men_n952_), .B(men_men_n60_), .Y(men_men_n953_));
  AOI220     u0904(.A0(men_men_n953_), .A1(men_men_n950_), .B0(men_men_n676_), .B1(men_men_n247_), .Y(men_men_n954_));
  NA4        u0905(.A(men_men_n954_), .B(men_men_n949_), .C(men_men_n946_), .D(men_men_n942_), .Y(men_men_n955_));
  NO4        u0906(.A(men_men_n939_), .B(men_men_n640_), .C(men_men_n462_), .D(men_men_n50_), .Y(men_men_n956_));
  AOI220     u0907(.A0(men_men_n611_), .A1(men_men_n610_), .B0(men_men_n286_), .B1(x5), .Y(men_men_n957_));
  NO2        u0908(.A(men_men_n684_), .B(men_men_n194_), .Y(men_men_n958_));
  NA3        u0909(.A(men_men_n958_), .B(men_men_n677_), .C(x7), .Y(men_men_n959_));
  OAI210     u0910(.A0(men_men_n957_), .A1(men_men_n353_), .B0(men_men_n959_), .Y(men_men_n960_));
  OAI210     u0911(.A0(men_men_n960_), .A1(men_men_n956_), .B0(men_men_n82_), .Y(men_men_n961_));
  NA2        u0912(.A(men_men_n782_), .B(x2), .Y(men_men_n962_));
  NO2        u0913(.A(men_men_n962_), .B(men_men_n58_), .Y(men_men_n963_));
  NO2        u0914(.A(x5), .B(men_men_n53_), .Y(men_men_n964_));
  NAi21      u0915(.An(x1), .B(x4), .Y(men_men_n965_));
  NA2        u0916(.A(men_men_n965_), .B(men_men_n872_), .Y(men_men_n966_));
  NO3        u0917(.A(men_men_n966_), .B(men_men_n205_), .C(men_men_n964_), .Y(men_men_n967_));
  OAI210     u0918(.A0(men_men_n967_), .A1(men_men_n963_), .B0(men_men_n419_), .Y(men_men_n968_));
  NA2        u0919(.A(men_men_n968_), .B(men_men_n961_), .Y(men_men_n969_));
  AOI210     u0920(.A0(men_men_n955_), .A1(x6), .B0(men_men_n969_), .Y(men_men_n970_));
  NA3        u0921(.A(men_men_n970_), .B(men_men_n936_), .C(men_men_n921_), .Y(men10));
  NO2        u0922(.A(x4), .B(x1), .Y(men_men_n972_));
  NO2        u0923(.A(men_men_n972_), .B(men_men_n151_), .Y(men_men_n973_));
  NA3        u0924(.A(x5), .B(x4), .C(x0), .Y(men_men_n974_));
  OAI220     u0925(.A0(men_men_n974_), .A1(men_men_n281_), .B0(men_men_n712_), .B1(men_men_n251_), .Y(men_men_n975_));
  NA2        u0926(.A(men_men_n975_), .B(men_men_n973_), .Y(men_men_n976_));
  NO3        u0927(.A(men_men_n360_), .B(men_men_n324_), .C(men_men_n92_), .Y(men_men_n977_));
  NA3        u0928(.A(men_men_n977_), .B(men_men_n387_), .C(men_men_n62_), .Y(men_men_n978_));
  AOI210     u0929(.A0(men_men_n978_), .A1(men_men_n976_), .B0(men_men_n308_), .Y(men_men_n979_));
  NOi21      u0930(.An(men_men_n262_), .B(men_men_n140_), .Y(men_men_n980_));
  AOI210     u0931(.A0(men_men_n507_), .A1(men_men_n625_), .B0(men_men_n333_), .Y(men_men_n981_));
  NO2        u0932(.A(men_men_n904_), .B(men_men_n346_), .Y(men_men_n982_));
  NOi31      u0933(.An(men_men_n982_), .B(men_men_n981_), .C(men_men_n980_), .Y(men_men_n983_));
  NA2        u0934(.A(x4), .B(men_men_n110_), .Y(men_men_n984_));
  NO2        u0935(.A(men_men_n327_), .B(men_men_n984_), .Y(men_men_n985_));
  NA2        u0936(.A(men_men_n99_), .B(x5), .Y(men_men_n986_));
  NO3        u0937(.A(men_men_n986_), .B(men_men_n111_), .C(men_men_n55_), .Y(men_men_n987_));
  NO3        u0938(.A(men_men_n987_), .B(men_men_n985_), .C(men_men_n983_), .Y(men_men_n988_));
  NA2        u0939(.A(men_men_n964_), .B(men_men_n50_), .Y(men_men_n989_));
  NA2        u0940(.A(men_men_n611_), .B(men_men_n275_), .Y(men_men_n990_));
  NO2        u0941(.A(men_men_n990_), .B(men_men_n989_), .Y(men_men_n991_));
  OAI220     u0942(.A0(men_men_n933_), .A1(men_men_n107_), .B0(men_men_n879_), .B1(men_men_n450_), .Y(men_men_n992_));
  AOI210     u0943(.A0(men_men_n992_), .A1(men_men_n283_), .B0(men_men_n991_), .Y(men_men_n993_));
  OAI210     u0944(.A0(men_men_n988_), .A1(men_men_n389_), .B0(men_men_n993_), .Y(men_men_n994_));
  OAI210     u0945(.A0(men_men_n994_), .A1(men_men_n979_), .B0(x7), .Y(men_men_n995_));
  NA2        u0946(.A(men_men_n55_), .B(men_men_n71_), .Y(men_men_n996_));
  AOI210     u0947(.A0(men_men_n450_), .A1(men_men_n359_), .B0(men_men_n984_), .Y(men_men_n997_));
  NO3        u0948(.A(men_men_n452_), .B(men_men_n897_), .C(x5), .Y(men_men_n998_));
  OAI210     u0949(.A0(men_men_n998_), .A1(men_men_n997_), .B0(men_men_n996_), .Y(men_men_n999_));
  NO2        u0950(.A(men_men_n360_), .B(men_men_n143_), .Y(men_men_n1000_));
  NA2        u0951(.A(men_men_n1000_), .B(men_men_n430_), .Y(men_men_n1001_));
  AOI210     u0952(.A0(men_men_n1001_), .A1(men_men_n999_), .B0(x3), .Y(men_men_n1002_));
  NA2        u0953(.A(men_men_n704_), .B(men_men_n254_), .Y(men_men_n1003_));
  NO2        u0954(.A(x5), .B(men_men_n110_), .Y(men_men_n1004_));
  OAI210     u0955(.A0(men_men_n1004_), .A1(men_men_n241_), .B0(men_men_n944_), .Y(men_men_n1005_));
  NA3        u0956(.A(men_men_n469_), .B(men_men_n132_), .C(men_men_n430_), .Y(men_men_n1006_));
  OAI210     u0957(.A0(men_men_n452_), .A1(men_men_n217_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  AOI210     u0958(.A0(men_men_n1005_), .A1(men_men_n260_), .B0(men_men_n1007_), .Y(men_men_n1008_));
  OAI220     u0959(.A0(men_men_n1008_), .A1(men_men_n59_), .B0(men_men_n1003_), .B1(men_men_n717_), .Y(men_men_n1009_));
  OAI210     u0960(.A0(men_men_n1009_), .A1(men_men_n1002_), .B0(men_men_n951_), .Y(men_men_n1010_));
  NO2        u0961(.A(x4), .B(x3), .Y(men_men_n1011_));
  NO3        u0962(.A(men_men_n1011_), .B(men_men_n347_), .C(men_men_n87_), .Y(men_men_n1012_));
  OAI210     u0963(.A0(men_men_n1012_), .A1(men_men_n282_), .B0(men_men_n441_), .Y(men_men_n1013_));
  AOI210     u0964(.A0(men_men_n403_), .A1(men_men_n129_), .B0(men_men_n255_), .Y(men_men_n1014_));
  NA2        u0965(.A(men_men_n972_), .B(men_men_n55_), .Y(men_men_n1015_));
  NO2        u0966(.A(men_men_n1015_), .B(men_men_n986_), .Y(men_men_n1016_));
  NO2        u0967(.A(men_men_n531_), .B(men_men_n365_), .Y(men_men_n1017_));
  NO3        u0968(.A(x4), .B(men_men_n110_), .C(men_men_n59_), .Y(men_men_n1018_));
  NO2        u0969(.A(men_men_n442_), .B(x1), .Y(men_men_n1019_));
  NOi31      u0970(.An(men_men_n1018_), .B(men_men_n1019_), .C(men_men_n1017_), .Y(men_men_n1020_));
  NA2        u0971(.A(men_men_n55_), .B(x5), .Y(men_men_n1021_));
  NO4        u0972(.A(men_men_n973_), .B(men_men_n520_), .C(men_men_n1021_), .D(x2), .Y(men_men_n1022_));
  NO4        u0973(.A(men_men_n1022_), .B(men_men_n1020_), .C(men_men_n1016_), .D(men_men_n1014_), .Y(men_men_n1023_));
  AOI210     u0974(.A0(men_men_n1023_), .A1(men_men_n1013_), .B0(men_men_n211_), .Y(men_men_n1024_));
  NO2        u0975(.A(men_men_n673_), .B(men_men_n506_), .Y(men_men_n1025_));
  NO2        u0976(.A(x6), .B(x2), .Y(men_men_n1026_));
  NO3        u0977(.A(men_men_n1026_), .B(men_men_n704_), .C(men_men_n60_), .Y(men_men_n1027_));
  OAI210     u0978(.A0(men_men_n1027_), .A1(men_men_n1025_), .B0(men_men_n274_), .Y(men_men_n1028_));
  NO2        u0979(.A(men_men_n879_), .B(men_men_n450_), .Y(men_men_n1029_));
  NA3        u0980(.A(x4), .B(x3), .C(men_men_n110_), .Y(men_men_n1030_));
  NO3        u0981(.A(men_men_n1030_), .B(men_men_n710_), .C(men_men_n469_), .Y(men_men_n1031_));
  AOI210     u0982(.A0(men_men_n1029_), .A1(men_men_n476_), .B0(men_men_n1031_), .Y(men_men_n1032_));
  AOI210     u0983(.A0(men_men_n1032_), .A1(men_men_n1028_), .B0(men_men_n462_), .Y(men_men_n1033_));
  NO2        u0984(.A(men_men_n55_), .B(men_men_n56_), .Y(men_men_n1034_));
  OAI220     u0985(.A0(men_men_n829_), .A1(men_men_n464_), .B0(men_men_n759_), .B1(men_men_n129_), .Y(men_men_n1035_));
  NOi21      u0986(.An(men_men_n124_), .B(men_men_n123_), .Y(men_men_n1036_));
  NO3        u0987(.A(men_men_n348_), .B(men_men_n327_), .C(men_men_n1036_), .Y(men_men_n1037_));
  AOI220     u0988(.A0(men_men_n1037_), .A1(men_men_n259_), .B0(men_men_n1035_), .B1(men_men_n116_), .Y(men_men_n1038_));
  NO2        u0989(.A(men_men_n1038_), .B(men_men_n1034_), .Y(men_men_n1039_));
  NA2        u0990(.A(men_men_n524_), .B(men_men_n264_), .Y(men_men_n1040_));
  NO2        u0991(.A(men_men_n491_), .B(men_men_n593_), .Y(men_men_n1041_));
  NA3        u0992(.A(men_men_n1041_), .B(men_men_n1040_), .C(men_men_n55_), .Y(men_men_n1042_));
  NO2        u0993(.A(men_men_n186_), .B(men_men_n110_), .Y(men_men_n1043_));
  NA3        u0994(.A(men_men_n1043_), .B(men_men_n185_), .C(men_men_n123_), .Y(men_men_n1044_));
  NA2        u0995(.A(men_men_n1044_), .B(men_men_n1042_), .Y(men_men_n1045_));
  NO4        u0996(.A(men_men_n1045_), .B(men_men_n1039_), .C(men_men_n1033_), .D(men_men_n1024_), .Y(men_men_n1046_));
  NA3        u0997(.A(men_men_n1046_), .B(men_men_n1010_), .C(men_men_n995_), .Y(men11));
  NA2        u0998(.A(men_men_n380_), .B(men_men_n92_), .Y(men_men_n1048_));
  INV        u0999(.A(men_men_n898_), .Y(men_men_n1049_));
  OAI220     u1000(.A0(men_men_n1049_), .A1(men_men_n53_), .B0(men_men_n1048_), .B1(men_men_n369_), .Y(men_men_n1050_));
  NO2        u1001(.A(men_men_n776_), .B(x5), .Y(men_men_n1051_));
  NO2        u1002(.A(men_men_n171_), .B(men_men_n537_), .Y(men_men_n1052_));
  AOI220     u1003(.A0(men_men_n1052_), .A1(men_men_n1051_), .B0(men_men_n1050_), .B1(x5), .Y(men_men_n1053_));
  OAI220     u1004(.A0(men_men_n980_), .A1(men_men_n220_), .B0(men_men_n218_), .B1(men_men_n186_), .Y(men_men_n1054_));
  NO2        u1005(.A(men_men_n344_), .B(men_men_n431_), .Y(men_men_n1055_));
  AOI220     u1006(.A0(men_men_n1055_), .A1(men_men_n184_), .B0(men_men_n1054_), .B1(men_men_n167_), .Y(men_men_n1056_));
  NO2        u1007(.A(men_men_n1056_), .B(men_men_n452_), .Y(men_men_n1057_));
  NO2        u1008(.A(men_men_n255_), .B(x2), .Y(men_men_n1058_));
  OAI210     u1009(.A0(men_men_n922_), .A1(men_men_n1058_), .B0(men_men_n420_), .Y(men_men_n1059_));
  NO2        u1010(.A(men_men_n55_), .B(men_men_n108_), .Y(men_men_n1060_));
  NA2        u1011(.A(men_men_n283_), .B(men_men_n1060_), .Y(men_men_n1061_));
  NO2        u1012(.A(men_men_n71_), .B(x1), .Y(men_men_n1062_));
  NA2        u1013(.A(men_men_n1062_), .B(men_men_n78_), .Y(men_men_n1063_));
  OA220      u1014(.A0(men_men_n1063_), .A1(men_men_n619_), .B0(men_men_n1061_), .B1(men_men_n537_), .Y(men_men_n1064_));
  AOI210     u1015(.A0(men_men_n1064_), .A1(men_men_n1059_), .B0(men_men_n717_), .Y(men_men_n1065_));
  NO2        u1016(.A(men_men_n309_), .B(men_men_n53_), .Y(men_men_n1066_));
  NO2        u1017(.A(men_men_n441_), .B(x3), .Y(men_men_n1067_));
  NA3        u1018(.A(men_men_n1067_), .B(men_men_n1066_), .C(men_men_n897_), .Y(men_men_n1068_));
  AOI210     u1019(.A0(men_men_n1068_), .A1(men_men_n948_), .B0(men_men_n401_), .Y(men_men_n1069_));
  NA2        u1020(.A(men_men_n110_), .B(x1), .Y(men_men_n1070_));
  NO2        u1021(.A(men_men_n625_), .B(men_men_n223_), .Y(men_men_n1071_));
  NA4        u1022(.A(men_men_n1071_), .B(men_men_n889_), .C(men_men_n473_), .D(men_men_n1070_), .Y(men_men_n1072_));
  NA3        u1023(.A(x6), .B(x5), .C(men_men_n110_), .Y(men_men_n1073_));
  NO2        u1024(.A(men_men_n1073_), .B(men_men_n281_), .Y(men_men_n1074_));
  NO2        u1025(.A(men_men_n452_), .B(x0), .Y(men_men_n1075_));
  NOi31      u1026(.An(men_men_n1075_), .B(men_men_n176_), .C(men_men_n51_), .Y(men_men_n1076_));
  AOI210     u1027(.A0(men_men_n1074_), .A1(men_men_n182_), .B0(men_men_n1076_), .Y(men_men_n1077_));
  NA2        u1028(.A(men_men_n1077_), .B(men_men_n1072_), .Y(men_men_n1078_));
  NO4        u1029(.A(men_men_n1078_), .B(men_men_n1069_), .C(men_men_n1065_), .D(men_men_n1057_), .Y(men_men_n1079_));
  OAI210     u1030(.A0(men_men_n1053_), .A1(men_men_n144_), .B0(men_men_n1079_), .Y(men_men_n1080_));
  NA2        u1031(.A(men_men_n870_), .B(men_men_n87_), .Y(men_men_n1081_));
  NO3        u1032(.A(men_men_n470_), .B(men_men_n782_), .C(men_men_n124_), .Y(men_men_n1082_));
  AOI210     u1033(.A0(men_men_n1081_), .A1(men_men_n101_), .B0(men_men_n1082_), .Y(men_men_n1083_));
  NO2        u1034(.A(x8), .B(x1), .Y(men_men_n1084_));
  NO3        u1035(.A(men_men_n1084_), .B(men_men_n696_), .C(men_men_n454_), .Y(men_men_n1085_));
  OAI210     u1036(.A0(men_men_n77_), .A1(men_men_n53_), .B0(men_men_n1085_), .Y(men_men_n1086_));
  OAI210     u1037(.A0(men_men_n1083_), .A1(x3), .B0(men_men_n1086_), .Y(men_men_n1087_));
  NO2        u1038(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n1088_));
  OAI210     u1039(.A0(men_men_n1088_), .A1(x2), .B0(men_men_n237_), .Y(men_men_n1089_));
  NO2        u1040(.A(men_men_n612_), .B(men_men_n235_), .Y(men_men_n1090_));
  NA2        u1041(.A(men_men_n1090_), .B(men_men_n1089_), .Y(men_men_n1091_));
  NO2        u1042(.A(men_men_n524_), .B(x4), .Y(men_men_n1092_));
  NO3        u1043(.A(men_men_n55_), .B(x6), .C(x1), .Y(men_men_n1093_));
  NOi21      u1044(.An(men_men_n1093_), .B(men_men_n491_), .Y(men_men_n1094_));
  AOI210     u1045(.A0(men_men_n1092_), .A1(men_men_n583_), .B0(men_men_n1094_), .Y(men_men_n1095_));
  NA2        u1046(.A(men_men_n1095_), .B(men_men_n1091_), .Y(men_men_n1096_));
  AOI210     u1047(.A0(men_men_n1087_), .A1(x2), .B0(men_men_n1096_), .Y(men_men_n1097_));
  NO2        u1048(.A(men_men_n235_), .B(x2), .Y(men_men_n1098_));
  NA2        u1049(.A(men_men_n1098_), .B(men_men_n1011_), .Y(men_men_n1099_));
  NOi21      u1050(.An(men_men_n392_), .B(men_men_n572_), .Y(men_men_n1100_));
  NO3        u1051(.A(men_men_n1100_), .B(men_men_n611_), .C(men_men_n327_), .Y(men_men_n1101_));
  NA2        u1052(.A(x8), .B(men_men_n110_), .Y(men_men_n1102_));
  OAI220     u1053(.A0(men_men_n717_), .A1(men_men_n1102_), .B0(men_men_n327_), .B1(men_men_n387_), .Y(men_men_n1103_));
  OAI210     u1054(.A0(men_men_n1103_), .A1(men_men_n1101_), .B0(men_men_n71_), .Y(men_men_n1104_));
  NO2        u1055(.A(men_men_n108_), .B(x1), .Y(men_men_n1105_));
  NA2        u1056(.A(men_men_n1105_), .B(x7), .Y(men_men_n1106_));
  AOI210     u1057(.A0(men_men_n1104_), .A1(men_men_n1099_), .B0(men_men_n1106_), .Y(men_men_n1107_));
  NA2        u1058(.A(men_men_n84_), .B(men_men_n71_), .Y(men_men_n1108_));
  INV        u1059(.A(men_men_n252_), .Y(men_men_n1109_));
  NA2        u1060(.A(men_men_n1109_), .B(men_men_n151_), .Y(men_men_n1110_));
  OAI220     u1061(.A0(men_men_n1110_), .A1(men_men_n369_), .B0(men_men_n1108_), .B1(men_men_n327_), .Y(men_men_n1111_));
  NO2        u1062(.A(men_men_n161_), .B(men_men_n55_), .Y(men_men_n1112_));
  AOI210     u1063(.A0(men_men_n1112_), .A1(men_men_n1111_), .B0(men_men_n1107_), .Y(men_men_n1113_));
  OAI210     u1064(.A0(men_men_n1097_), .A1(men_men_n857_), .B0(men_men_n1113_), .Y(men_men_n1114_));
  AO210      u1065(.A0(men_men_n1080_), .A1(men_men_n57_), .B0(men_men_n1114_), .Y(men12));
  NA2        u1066(.A(men_men_n888_), .B(men_men_n251_), .Y(men_men_n1116_));
  NO2        u1067(.A(men_men_n629_), .B(x7), .Y(men_men_n1117_));
  NA2        u1068(.A(men_men_n1117_), .B(men_men_n282_), .Y(men_men_n1118_));
  NA2        u1069(.A(men_men_n709_), .B(men_men_n879_), .Y(men_men_n1119_));
  AOI210     u1070(.A0(men_men_n1118_), .A1(men_men_n1116_), .B0(men_men_n1119_), .Y(men_men_n1120_));
  NOi21      u1071(.An(men_men_n408_), .B(men_men_n559_), .Y(men_men_n1121_));
  NO2        u1072(.A(x7), .B(men_men_n50_), .Y(men_men_n1122_));
  NO2        u1073(.A(men_men_n612_), .B(men_men_n1122_), .Y(men_men_n1123_));
  NO3        u1074(.A(men_men_n872_), .B(men_men_n112_), .C(men_men_n99_), .Y(men_men_n1124_));
  AOI210     u1075(.A0(men_men_n1123_), .A1(men_men_n1019_), .B0(men_men_n1124_), .Y(men_men_n1125_));
  NA2        u1076(.A(men_men_n1060_), .B(men_men_n56_), .Y(men_men_n1126_));
  OAI220     u1077(.A0(men_men_n1126_), .A1(men_men_n584_), .B0(men_men_n1125_), .B1(men_men_n1121_), .Y(men_men_n1127_));
  OAI210     u1078(.A0(men_men_n1127_), .A1(men_men_n1120_), .B0(men_men_n588_), .Y(men_men_n1128_));
  NA2        u1079(.A(men_men_n87_), .B(x5), .Y(men_men_n1129_));
  OAI210     u1080(.A0(men_men_n1129_), .A1(men_men_n327_), .B0(men_men_n724_), .Y(men_men_n1130_));
  AOI210     u1081(.A0(men_men_n831_), .A1(men_men_n118_), .B0(men_men_n1130_), .Y(men_men_n1131_));
  NA2        u1082(.A(men_men_n610_), .B(men_men_n53_), .Y(men_men_n1132_));
  NA2        u1083(.A(men_men_n292_), .B(men_men_n50_), .Y(men_men_n1133_));
  OAI220     u1084(.A0(men_men_n1133_), .A1(men_men_n315_), .B0(men_men_n1132_), .B1(men_men_n137_), .Y(men_men_n1134_));
  NO2        u1085(.A(men_men_n1081_), .B(men_men_n519_), .Y(men_men_n1135_));
  NO4        u1086(.A(men_men_n243_), .B(men_men_n274_), .C(men_men_n60_), .D(men_men_n57_), .Y(men_men_n1136_));
  AOI220     u1087(.A0(men_men_n1136_), .A1(men_men_n1135_), .B0(men_men_n1134_), .B1(men_men_n56_), .Y(men_men_n1137_));
  OAI210     u1088(.A0(men_men_n1131_), .A1(men_men_n64_), .B0(men_men_n1137_), .Y(men_men_n1138_));
  NO2        u1089(.A(men_men_n57_), .B(x0), .Y(men_men_n1139_));
  NO2        u1090(.A(men_men_n673_), .B(men_men_n324_), .Y(men_men_n1140_));
  NO2        u1091(.A(men_men_n759_), .B(x3), .Y(men_men_n1141_));
  NO2        u1092(.A(men_men_n671_), .B(x8), .Y(men_men_n1142_));
  AOI220     u1093(.A0(men_men_n1142_), .A1(men_men_n1141_), .B0(men_men_n1140_), .B1(men_men_n1139_), .Y(men_men_n1143_));
  AOI210     u1094(.A0(men_men_n696_), .A1(men_men_n251_), .B0(x7), .Y(men_men_n1144_));
  NO3        u1095(.A(men_men_n1144_), .B(men_men_n613_), .C(x8), .Y(men_men_n1145_));
  NA4        u1096(.A(men_men_n675_), .B(men_men_n667_), .C(men_men_n208_), .D(x0), .Y(men_men_n1146_));
  OAI220     u1097(.A0(men_men_n1146_), .A1(men_men_n1145_), .B0(men_men_n1143_), .B1(men_men_n582_), .Y(men_men_n1147_));
  AOI210     u1098(.A0(men_men_n1138_), .A1(men_men_n1026_), .B0(men_men_n1147_), .Y(men_men_n1148_));
  NO2        u1099(.A(men_men_n251_), .B(men_men_n55_), .Y(men_men_n1149_));
  NO2        u1100(.A(men_men_n259_), .B(x8), .Y(men_men_n1150_));
  NOi32      u1101(.An(men_men_n1150_), .Bn(men_men_n207_), .C(men_men_n573_), .Y(men_men_n1151_));
  NO2        u1102(.A(men_men_n88_), .B(men_men_n60_), .Y(men_men_n1152_));
  OAI210     u1103(.A0(men_men_n1151_), .A1(men_men_n1149_), .B0(men_men_n1152_), .Y(men_men_n1153_));
  NO2        u1104(.A(men_men_n951_), .B(men_men_n100_), .Y(men_men_n1154_));
  NO2        u1105(.A(men_men_n170_), .B(men_men_n53_), .Y(men_men_n1155_));
  AOI210     u1106(.A0(men_men_n344_), .A1(x8), .B0(men_men_n1155_), .Y(men_men_n1156_));
  AOI210     u1107(.A0(men_men_n220_), .A1(men_men_n96_), .B0(men_men_n1156_), .Y(men_men_n1157_));
  OAI210     u1108(.A0(men_men_n1157_), .A1(men_men_n1154_), .B0(men_men_n684_), .Y(men_men_n1158_));
  NO2        u1109(.A(x7), .B(x0), .Y(men_men_n1159_));
  NO3        u1110(.A(men_men_n161_), .B(men_men_n1159_), .C(men_men_n148_), .Y(men_men_n1160_));
  XN2        u1111(.A(x8), .B(x7), .Y(men_men_n1161_));
  NO3        u1112(.A(men_men_n1084_), .B(men_men_n262_), .C(men_men_n1161_), .Y(men_men_n1162_));
  OAI210     u1113(.A0(men_men_n1162_), .A1(men_men_n1160_), .B0(men_men_n738_), .Y(men_men_n1163_));
  NO2        u1114(.A(men_men_n271_), .B(men_men_n267_), .Y(men_men_n1164_));
  NO2        u1115(.A(men_men_n108_), .B(x4), .Y(men_men_n1165_));
  OAI210     u1116(.A0(men_men_n1164_), .A1(men_men_n282_), .B0(men_men_n1165_), .Y(men_men_n1166_));
  NA4        u1117(.A(men_men_n1166_), .B(men_men_n1163_), .C(men_men_n1158_), .D(men_men_n1153_), .Y(men_men_n1167_));
  NA2        u1118(.A(men_men_n1167_), .B(men_men_n563_), .Y(men_men_n1168_));
  NO2        u1119(.A(men_men_n55_), .B(x4), .Y(men_men_n1169_));
  NA2        u1120(.A(men_men_n1169_), .B(men_men_n166_), .Y(men_men_n1170_));
  NO2        u1121(.A(men_men_n677_), .B(men_men_n262_), .Y(men_men_n1171_));
  OAI210     u1122(.A0(men_men_n1171_), .A1(men_men_n1029_), .B0(men_men_n50_), .Y(men_men_n1172_));
  AOI210     u1123(.A0(men_men_n1172_), .A1(men_men_n1170_), .B0(men_men_n436_), .Y(men_men_n1173_));
  OAI220     u1124(.A0(men_men_n294_), .A1(men_men_n280_), .B0(men_men_n267_), .B1(men_men_n246_), .Y(men_men_n1174_));
  NA3        u1125(.A(men_men_n1174_), .B(men_men_n684_), .C(x1), .Y(men_men_n1175_));
  OAI210     u1126(.A0(x8), .A1(x0), .B0(x4), .Y(men_men_n1176_));
  NO2        u1127(.A(x7), .B(men_men_n56_), .Y(men_men_n1177_));
  NO2        u1128(.A(men_men_n68_), .B(men_men_n1177_), .Y(men_men_n1178_));
  NOi21      u1129(.An(men_men_n1176_), .B(men_men_n1178_), .Y(men_men_n1179_));
  NO2        u1130(.A(men_men_n675_), .B(men_men_n327_), .Y(men_men_n1180_));
  NO2        u1131(.A(men_men_n784_), .B(men_men_n224_), .Y(men_men_n1181_));
  OAI210     u1132(.A0(men_men_n1180_), .A1(men_men_n1179_), .B0(men_men_n1181_), .Y(men_men_n1182_));
  NO2        u1133(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n1183_));
  NO2        u1134(.A(men_men_n612_), .B(men_men_n450_), .Y(men_men_n1184_));
  OAI210     u1135(.A0(men_men_n1184_), .A1(men_men_n1183_), .B0(men_men_n259_), .Y(men_men_n1185_));
  NO2        u1136(.A(men_men_n827_), .B(men_men_n427_), .Y(men_men_n1186_));
  NA2        u1137(.A(men_men_n332_), .B(men_men_n59_), .Y(men_men_n1187_));
  NO2        u1138(.A(men_men_n1126_), .B(men_men_n1187_), .Y(men_men_n1188_));
  AOI210     u1139(.A0(men_men_n1186_), .A1(men_men_n182_), .B0(men_men_n1188_), .Y(men_men_n1189_));
  NA4        u1140(.A(men_men_n1189_), .B(men_men_n1185_), .C(men_men_n1182_), .D(men_men_n1175_), .Y(men_men_n1190_));
  OAI210     u1141(.A0(men_men_n1190_), .A1(men_men_n1173_), .B0(men_men_n686_), .Y(men_men_n1191_));
  NA4        u1142(.A(men_men_n1191_), .B(men_men_n1168_), .C(men_men_n1148_), .D(men_men_n1128_), .Y(men13));
  NO2        u1143(.A(men_men_n469_), .B(men_men_n354_), .Y(men_men_n1193_));
  NOi41      u1144(.An(men_men_n1193_), .B(men_men_n684_), .C(men_men_n296_), .D(men_men_n243_), .Y(men_men_n1194_));
  NO2        u1145(.A(men_men_n872_), .B(men_men_n186_), .Y(men_men_n1195_));
  NO2        u1146(.A(men_men_n160_), .B(men_men_n71_), .Y(men_men_n1196_));
  XN2        u1147(.A(x4), .B(x0), .Y(men_men_n1197_));
  NO3        u1148(.A(men_men_n1197_), .B(men_men_n111_), .C(men_men_n427_), .Y(men_men_n1198_));
  AO220      u1149(.A0(men_men_n1198_), .A1(men_men_n1196_), .B0(men_men_n1195_), .B1(men_men_n333_), .Y(men_men_n1199_));
  OAI210     u1150(.A0(men_men_n1199_), .A1(men_men_n1194_), .B0(x3), .Y(men_men_n1200_));
  NO2        u1151(.A(men_men_n872_), .B(x6), .Y(men_men_n1201_));
  NO2        u1152(.A(men_men_n1133_), .B(men_men_n399_), .Y(men_men_n1202_));
  NO3        u1153(.A(x8), .B(x5), .C(men_men_n110_), .Y(men_men_n1203_));
  NA2        u1154(.A(men_men_n1203_), .B(men_men_n649_), .Y(men_men_n1204_));
  NO2        u1155(.A(men_men_n612_), .B(men_men_n202_), .Y(men_men_n1205_));
  NA2        u1156(.A(men_men_n1205_), .B(men_men_n1093_), .Y(men_men_n1206_));
  NA2        u1157(.A(men_men_n454_), .B(men_men_n53_), .Y(men_men_n1207_));
  NO2        u1158(.A(men_men_n1207_), .B(men_men_n944_), .Y(men_men_n1208_));
  NA2        u1159(.A(men_men_n1126_), .B(men_men_n474_), .Y(men_men_n1209_));
  NA2        u1160(.A(men_men_n56_), .B(men_men_n110_), .Y(men_men_n1210_));
  NA2        u1161(.A(men_men_n1210_), .B(x1), .Y(men_men_n1211_));
  NO2        u1162(.A(men_men_n1211_), .B(men_men_n264_), .Y(men_men_n1212_));
  NO2        u1163(.A(men_men_n324_), .B(x6), .Y(men_men_n1213_));
  OAI210     u1164(.A0(men_men_n255_), .A1(men_men_n984_), .B0(men_men_n962_), .Y(men_men_n1214_));
  AOI220     u1165(.A0(men_men_n1214_), .A1(men_men_n1213_), .B0(men_men_n1212_), .B1(men_men_n1209_), .Y(men_men_n1215_));
  NAi41      u1166(.An(men_men_n1208_), .B(men_men_n1215_), .C(men_men_n1206_), .D(men_men_n1204_), .Y(men_men_n1216_));
  AOI220     u1167(.A0(men_men_n1216_), .A1(men_men_n68_), .B0(men_men_n1202_), .B1(men_men_n1201_), .Y(men_men_n1217_));
  NA2        u1168(.A(men_men_n71_), .B(x3), .Y(men_men_n1218_));
  NA2        u1169(.A(men_men_n1218_), .B(men_men_n906_), .Y(men_men_n1219_));
  OAI220     u1170(.A0(men_men_n308_), .A1(men_men_n827_), .B0(men_men_n87_), .B1(men_men_n77_), .Y(men_men_n1220_));
  AOI210     u1171(.A0(men_men_n1129_), .A1(men_men_n623_), .B0(men_men_n984_), .Y(men_men_n1221_));
  OA210      u1172(.A0(men_men_n1220_), .A1(men_men_n1219_), .B0(men_men_n1221_), .Y(men_men_n1222_));
  NA2        u1173(.A(men_men_n625_), .B(men_men_n55_), .Y(men_men_n1223_));
  NA2        u1174(.A(men_men_n512_), .B(men_men_n500_), .Y(men_men_n1224_));
  NA2        u1175(.A(x6), .B(men_men_n50_), .Y(men_men_n1225_));
  NA2        u1176(.A(men_men_n1225_), .B(men_men_n546_), .Y(men_men_n1226_));
  NO2        u1177(.A(men_men_n163_), .B(men_men_n132_), .Y(men_men_n1227_));
  AOI210     u1178(.A0(men_men_n1226_), .A1(men_men_n437_), .B0(men_men_n1227_), .Y(men_men_n1228_));
  OAI220     u1179(.A0(men_men_n1228_), .A1(men_men_n879_), .B0(men_men_n1224_), .B1(men_men_n1223_), .Y(men_men_n1229_));
  OAI210     u1180(.A0(men_men_n1229_), .A1(men_men_n1222_), .B0(men_men_n1159_), .Y(men_men_n1230_));
  NAi21      u1181(.An(men_men_n84_), .B(men_men_n387_), .Y(men_men_n1231_));
  NO2        u1182(.A(men_men_n1231_), .B(men_men_n71_), .Y(men_men_n1232_));
  AOI210     u1183(.A0(men_men_n166_), .A1(x4), .B0(men_men_n178_), .Y(men_men_n1233_));
  NO2        u1184(.A(men_men_n1233_), .B(x0), .Y(men_men_n1234_));
  NO2        u1185(.A(men_men_n174_), .B(men_men_n299_), .Y(men_men_n1235_));
  OAI210     u1186(.A0(men_men_n1235_), .A1(men_men_n1234_), .B0(men_men_n1232_), .Y(men_men_n1236_));
  NA3        u1187(.A(men_men_n1165_), .B(men_men_n193_), .C(men_men_n71_), .Y(men_men_n1237_));
  NO2        u1188(.A(x4), .B(x0), .Y(men_men_n1238_));
  NO3        u1189(.A(men_men_n1004_), .B(men_men_n252_), .C(men_men_n546_), .Y(men_men_n1239_));
  OAI210     u1190(.A0(men_men_n1239_), .A1(men_men_n203_), .B0(men_men_n1238_), .Y(men_men_n1240_));
  NA3        u1191(.A(men_men_n1240_), .B(men_men_n1237_), .C(men_men_n1236_), .Y(men_men_n1241_));
  NA2        u1192(.A(men_men_n254_), .B(men_men_n738_), .Y(men_men_n1242_));
  NO2        u1193(.A(men_men_n1242_), .B(men_men_n526_), .Y(men_men_n1243_));
  NA2        u1194(.A(men_men_n56_), .B(x0), .Y(men_men_n1244_));
  NO3        u1195(.A(men_men_n1244_), .B(men_men_n500_), .C(men_men_n81_), .Y(men_men_n1245_));
  OAI210     u1196(.A0(men_men_n1245_), .A1(men_men_n1243_), .B0(x2), .Y(men_men_n1246_));
  NO2        u1197(.A(men_men_n327_), .B(men_men_n387_), .Y(men_men_n1247_));
  NO2        u1198(.A(men_men_n696_), .B(x0), .Y(men_men_n1248_));
  OAI210     u1199(.A0(men_men_n1248_), .A1(men_men_n1247_), .B0(men_men_n336_), .Y(men_men_n1249_));
  NO2        u1200(.A(men_men_n796_), .B(x1), .Y(men_men_n1250_));
  AOI220     u1201(.A0(men_men_n1250_), .A1(men_men_n618_), .B0(men_men_n484_), .B1(men_men_n300_), .Y(men_men_n1251_));
  NA2        u1202(.A(men_men_n506_), .B(men_men_n50_), .Y(men_men_n1252_));
  AOI220     u1203(.A0(men_men_n1252_), .A1(men_men_n1195_), .B0(men_men_n985_), .B1(men_men_n101_), .Y(men_men_n1253_));
  NA4        u1204(.A(men_men_n1253_), .B(men_men_n1251_), .C(men_men_n1249_), .D(men_men_n1246_), .Y(men_men_n1254_));
  AOI220     u1205(.A0(men_men_n1254_), .A1(men_men_n133_), .B0(men_men_n1241_), .B1(men_men_n67_), .Y(men_men_n1255_));
  NA4        u1206(.A(men_men_n1255_), .B(men_men_n1230_), .C(men_men_n1217_), .D(men_men_n1200_), .Y(men14));
  NO2        u1207(.A(men_men_n375_), .B(men_men_n71_), .Y(men_men_n1257_));
  NO3        u1208(.A(x7), .B(x6), .C(x0), .Y(men_men_n1258_));
  OAI210     u1209(.A0(men_men_n1258_), .A1(men_men_n1257_), .B0(x8), .Y(men_men_n1259_));
  NA2        u1210(.A(men_men_n1142_), .B(men_men_n85_), .Y(men_men_n1260_));
  AOI210     u1211(.A0(men_men_n1260_), .A1(men_men_n1259_), .B0(men_men_n159_), .Y(men_men_n1261_));
  AOI220     u1212(.A0(men_men_n379_), .A1(men_men_n857_), .B0(men_men_n454_), .B1(men_men_n427_), .Y(men_men_n1262_));
  NA2        u1213(.A(men_men_n283_), .B(men_men_n980_), .Y(men_men_n1263_));
  OAI220     u1214(.A0(men_men_n1263_), .A1(men_men_n1262_), .B0(men_men_n472_), .B1(men_men_n811_), .Y(men_men_n1264_));
  OA210      u1215(.A0(men_men_n1264_), .A1(men_men_n1261_), .B0(x4), .Y(men_men_n1265_));
  NO2        u1216(.A(men_men_n143_), .B(men_men_n616_), .Y(men_men_n1266_));
  NA2        u1217(.A(x6), .B(x2), .Y(men_men_n1267_));
  NO2        u1218(.A(men_men_n634_), .B(men_men_n1267_), .Y(men_men_n1268_));
  OA210      u1219(.A0(men_men_n1266_), .A1(men_men_n216_), .B0(men_men_n1268_), .Y(men_men_n1269_));
  NO4        u1220(.A(men_men_n612_), .B(men_men_n380_), .C(men_men_n304_), .D(men_men_n116_), .Y(men_men_n1270_));
  OAI210     u1221(.A0(men_men_n1270_), .A1(men_men_n1269_), .B0(men_men_n59_), .Y(men_men_n1271_));
  NA2        u1222(.A(x6), .B(men_men_n108_), .Y(men_men_n1272_));
  NO2        u1223(.A(men_men_n673_), .B(men_men_n1272_), .Y(men_men_n1273_));
  NA2        u1224(.A(men_men_n1273_), .B(men_men_n931_), .Y(men_men_n1274_));
  AOI210     u1225(.A0(men_men_n1142_), .A1(men_men_n1018_), .B0(x1), .Y(men_men_n1275_));
  NO2        u1226(.A(men_men_n541_), .B(x5), .Y(men_men_n1276_));
  NA3        u1227(.A(men_men_n1276_), .B(men_men_n123_), .C(x0), .Y(men_men_n1277_));
  NA4        u1228(.A(men_men_n703_), .B(men_men_n932_), .C(men_men_n308_), .D(men_men_n68_), .Y(men_men_n1278_));
  AN4        u1229(.A(men_men_n1278_), .B(men_men_n1277_), .C(men_men_n1275_), .D(men_men_n1274_), .Y(men_men_n1279_));
  NO2        u1230(.A(men_men_n710_), .B(men_men_n1102_), .Y(men_men_n1280_));
  NO2        u1231(.A(men_men_n77_), .B(men_men_n58_), .Y(men_men_n1281_));
  OAI210     u1232(.A0(men_men_n1280_), .A1(men_men_n451_), .B0(men_men_n1281_), .Y(men_men_n1282_));
  AO210      u1233(.A0(men_men_n1257_), .A1(men_men_n1018_), .B0(men_men_n53_), .Y(men_men_n1283_));
  AOI210     u1234(.A0(men_men_n772_), .A1(men_men_n821_), .B0(men_men_n1283_), .Y(men_men_n1284_));
  AOI220     u1235(.A0(men_men_n1284_), .A1(men_men_n1282_), .B0(men_men_n1279_), .B1(men_men_n1271_), .Y(men_men_n1285_));
  NO2        u1236(.A(men_men_n1285_), .B(men_men_n1265_), .Y(men_men_n1286_));
  NO2        u1237(.A(men_men_n324_), .B(x2), .Y(men_men_n1287_));
  XN2        u1238(.A(x4), .B(x1), .Y(men_men_n1288_));
  NO2        u1239(.A(men_men_n1288_), .B(men_men_n308_), .Y(men_men_n1289_));
  NOi21      u1240(.An(men_men_n1289_), .B(men_men_n415_), .Y(men_men_n1290_));
  NO2        u1241(.A(men_men_n343_), .B(men_men_n60_), .Y(men_men_n1291_));
  OAI210     u1242(.A0(men_men_n1291_), .A1(men_men_n1290_), .B0(men_men_n1287_), .Y(men_men_n1292_));
  NA2        u1243(.A(men_men_n697_), .B(men_men_n56_), .Y(men_men_n1293_));
  OAI220     u1244(.A0(men_men_n1293_), .A1(men_men_n160_), .B0(men_men_n194_), .B1(men_men_n71_), .Y(men_men_n1294_));
  NO2        u1245(.A(men_men_n220_), .B(men_men_n262_), .Y(men_men_n1295_));
  AOI220     u1246(.A0(men_men_n140_), .A1(men_men_n56_), .B0(men_men_n93_), .B1(x5), .Y(men_men_n1296_));
  NA2        u1247(.A(men_men_n1093_), .B(men_men_n313_), .Y(men_men_n1297_));
  NA2        u1248(.A(men_men_n254_), .B(men_men_n358_), .Y(men_men_n1298_));
  NA2        u1249(.A(men_men_n648_), .B(men_men_n1036_), .Y(men_men_n1299_));
  OAI220     u1250(.A0(men_men_n1299_), .A1(men_men_n1298_), .B0(men_men_n1297_), .B1(men_men_n1296_), .Y(men_men_n1300_));
  AOI210     u1251(.A0(men_men_n1295_), .A1(men_men_n1294_), .B0(men_men_n1300_), .Y(men_men_n1301_));
  AOI210     u1252(.A0(men_men_n1301_), .A1(men_men_n1292_), .B0(x7), .Y(men_men_n1302_));
  NO2        u1253(.A(men_men_n499_), .B(x6), .Y(men_men_n1303_));
  AOI210     u1254(.A0(men_men_n823_), .A1(men_men_n964_), .B0(men_men_n1303_), .Y(men_men_n1304_));
  OAI220     u1255(.A0(men_men_n1304_), .A1(men_men_n55_), .B0(men_men_n499_), .B1(men_men_n104_), .Y(men_men_n1305_));
  NA2        u1256(.A(men_men_n1305_), .B(men_men_n360_), .Y(men_men_n1306_));
  NA3        u1257(.A(men_men_n619_), .B(men_men_n1070_), .C(men_men_n70_), .Y(men_men_n1307_));
  NO4        u1258(.A(men_men_n1307_), .B(men_men_n1244_), .C(men_men_n121_), .D(men_men_n55_), .Y(men_men_n1308_));
  NO3        u1259(.A(men_men_n1063_), .B(men_men_n829_), .C(men_men_n489_), .Y(men_men_n1309_));
  NO3        u1260(.A(men_men_n759_), .B(men_men_n506_), .C(men_men_n54_), .Y(men_men_n1310_));
  NO4        u1261(.A(men_men_n1310_), .B(men_men_n1309_), .C(men_men_n1308_), .D(men_men_n1041_), .Y(men_men_n1311_));
  AOI210     u1262(.A0(men_men_n1311_), .A1(men_men_n1306_), .B0(men_men_n310_), .Y(men_men_n1312_));
  NA2        u1263(.A(men_men_n904_), .B(men_men_n53_), .Y(men_men_n1313_));
  OAI210     u1264(.A0(men_men_n249_), .A1(men_men_n118_), .B0(x2), .Y(men_men_n1314_));
  NA2        u1265(.A(men_men_n371_), .B(men_men_n56_), .Y(men_men_n1315_));
  OA220      u1266(.A0(men_men_n1315_), .A1(men_men_n1314_), .B0(men_men_n1313_), .B1(men_men_n379_), .Y(men_men_n1316_));
  NA3        u1267(.A(men_men_n1041_), .B(men_men_n743_), .C(men_men_n55_), .Y(men_men_n1317_));
  NA2        u1268(.A(men_men_n56_), .B(x2), .Y(men_men_n1318_));
  NO2        u1269(.A(men_men_n1318_), .B(men_men_n201_), .Y(men_men_n1319_));
  NA4        u1270(.A(men_men_n1319_), .B(men_men_n371_), .C(men_men_n262_), .D(men_men_n67_), .Y(men_men_n1320_));
  NA3        u1271(.A(men_men_n1250_), .B(men_men_n625_), .C(men_men_n639_), .Y(men_men_n1321_));
  AN3        u1272(.A(men_men_n1321_), .B(men_men_n1320_), .C(men_men_n1317_), .Y(men_men_n1322_));
  OAI210     u1273(.A0(men_men_n1316_), .A1(men_men_n320_), .B0(men_men_n1322_), .Y(men_men_n1323_));
  NO3        u1274(.A(men_men_n1323_), .B(men_men_n1312_), .C(men_men_n1302_), .Y(men_men_n1324_));
  OAI210     u1275(.A0(men_men_n1286_), .A1(x3), .B0(men_men_n1324_), .Y(men15));
  NA2        u1276(.A(men_men_n594_), .B(men_men_n59_), .Y(men_men_n1326_));
  NAi41      u1277(.An(x2), .B(x7), .C(x6), .D(x0), .Y(men_men_n1327_));
  AOI210     u1278(.A0(men_men_n1327_), .A1(men_men_n1326_), .B0(men_men_n53_), .Y(men_men_n1328_));
  NA3        u1279(.A(men_men_n57_), .B(x6), .C(men_men_n110_), .Y(men_men_n1329_));
  NO2        u1280(.A(men_men_n1329_), .B(men_men_n299_), .Y(men_men_n1330_));
  OAI210     u1281(.A0(men_men_n1330_), .A1(men_men_n1328_), .B0(men_men_n1165_), .Y(men_men_n1331_));
  NA2        u1282(.A(men_men_n112_), .B(men_men_n110_), .Y(men_men_n1332_));
  NA4        u1283(.A(men_men_n1332_), .B(men_men_n646_), .C(men_men_n314_), .D(x6), .Y(men_men_n1333_));
  AOI210     u1284(.A0(men_men_n737_), .A1(men_men_n76_), .B0(x3), .Y(men_men_n1334_));
  NA3        u1285(.A(men_men_n1334_), .B(men_men_n1333_), .C(men_men_n1331_), .Y(men_men_n1335_));
  AOI210     u1286(.A0(men_men_n1075_), .A1(men_men_n598_), .B0(men_men_n50_), .Y(men_men_n1336_));
  NO2        u1287(.A(men_men_n299_), .B(men_men_n110_), .Y(men_men_n1337_));
  NO2        u1288(.A(men_men_n241_), .B(x5), .Y(men_men_n1338_));
  NA2        u1289(.A(men_men_n1338_), .B(men_men_n1337_), .Y(men_men_n1339_));
  NA3        u1290(.A(men_men_n1250_), .B(men_men_n633_), .C(men_men_n1177_), .Y(men_men_n1340_));
  NA4        u1291(.A(men_men_n1340_), .B(men_men_n1339_), .C(men_men_n1336_), .D(men_men_n1277_), .Y(men_men_n1341_));
  NA2        u1292(.A(men_men_n337_), .B(men_men_n346_), .Y(men_men_n1342_));
  AOI210     u1293(.A0(men_men_n1211_), .A1(men_men_n58_), .B0(men_men_n1342_), .Y(men_men_n1343_));
  NA4        u1294(.A(men_men_n1211_), .B(men_men_n709_), .C(men_men_n1139_), .D(men_men_n387_), .Y(men_men_n1344_));
  NA2        u1295(.A(men_men_n598_), .B(men_men_n473_), .Y(men_men_n1345_));
  NO2        u1296(.A(men_men_n759_), .B(men_men_n53_), .Y(men_men_n1346_));
  NO2        u1297(.A(men_men_n784_), .B(men_men_n304_), .Y(men_men_n1347_));
  NA2        u1298(.A(men_men_n1347_), .B(men_men_n1346_), .Y(men_men_n1348_));
  NA3        u1299(.A(men_men_n1348_), .B(men_men_n1345_), .C(men_men_n1344_), .Y(men_men_n1349_));
  OAI210     u1300(.A0(men_men_n1349_), .A1(men_men_n1343_), .B0(men_men_n77_), .Y(men_men_n1350_));
  NA2        u1301(.A(men_men_n373_), .B(men_men_n712_), .Y(men_men_n1351_));
  NA2        u1302(.A(men_men_n579_), .B(men_men_n56_), .Y(men_men_n1352_));
  NA3        u1303(.A(men_men_n1352_), .B(men_men_n346_), .C(men_men_n112_), .Y(men_men_n1353_));
  AOI210     u1304(.A0(men_men_n1353_), .A1(men_men_n1351_), .B0(men_men_n506_), .Y(men_men_n1354_));
  NO3        u1305(.A(men_men_n809_), .B(men_men_n630_), .C(men_men_n202_), .Y(men_men_n1355_));
  OAI210     u1306(.A0(men_men_n1355_), .A1(men_men_n1354_), .B0(men_men_n499_), .Y(men_men_n1356_));
  NO2        u1307(.A(men_men_n879_), .B(men_men_n50_), .Y(men_men_n1357_));
  NO2        u1308(.A(men_men_n251_), .B(men_men_n64_), .Y(men_men_n1358_));
  OA210      u1309(.A0(men_men_n1358_), .A1(men_men_n1357_), .B0(men_men_n415_), .Y(men_men_n1359_));
  NA2        u1310(.A(men_men_n57_), .B(x3), .Y(men_men_n1360_));
  AOI210     u1311(.A0(men_men_n986_), .A1(men_men_n1360_), .B0(men_men_n691_), .Y(men_men_n1361_));
  OAI210     u1312(.A0(men_men_n1361_), .A1(men_men_n1359_), .B0(men_men_n1026_), .Y(men_men_n1362_));
  NA2        u1313(.A(men_men_n1319_), .B(men_men_n68_), .Y(men_men_n1363_));
  NO2        u1314(.A(men_men_n1267_), .B(x0), .Y(men_men_n1364_));
  AOI210     u1315(.A0(men_men_n1364_), .A1(men_men_n613_), .B0(x8), .Y(men_men_n1365_));
  NO2        u1316(.A(men_men_n436_), .B(men_men_n81_), .Y(men_men_n1366_));
  NO2        u1317(.A(men_men_n938_), .B(men_men_n71_), .Y(men_men_n1367_));
  NA2        u1318(.A(men_men_n1367_), .B(men_men_n1366_), .Y(men_men_n1368_));
  NO2        u1319(.A(men_men_n984_), .B(x6), .Y(men_men_n1369_));
  NA4        u1320(.A(men_men_n1369_), .B(men_men_n603_), .C(men_men_n161_), .D(men_men_n419_), .Y(men_men_n1370_));
  AN4        u1321(.A(men_men_n1370_), .B(men_men_n1368_), .C(men_men_n1365_), .D(men_men_n1363_), .Y(men_men_n1371_));
  NA4        u1322(.A(men_men_n1371_), .B(men_men_n1362_), .C(men_men_n1356_), .D(men_men_n1350_), .Y(men_men_n1372_));
  NA2        u1323(.A(men_men_n167_), .B(men_men_n743_), .Y(men_men_n1373_));
  NO2        u1324(.A(men_men_n658_), .B(x2), .Y(men_men_n1374_));
  OAI210     u1325(.A0(men_men_n68_), .A1(men_men_n53_), .B0(men_men_n146_), .Y(men_men_n1375_));
  OAI210     u1326(.A0(men_men_n1374_), .A1(men_men_n85_), .B0(men_men_n1375_), .Y(men_men_n1376_));
  AOI210     u1327(.A0(men_men_n1376_), .A1(men_men_n1373_), .B0(men_men_n324_), .Y(men_men_n1377_));
  NO3        u1328(.A(men_men_n1329_), .B(men_men_n270_), .C(men_men_n251_), .Y(men_men_n1378_));
  NA3        u1329(.A(men_men_n57_), .B(x1), .C(x0), .Y(men_men_n1379_));
  NA3        u1330(.A(men_men_n71_), .B(x5), .C(x2), .Y(men_men_n1380_));
  NA4        u1331(.A(x7), .B(x3), .C(men_men_n53_), .D(x0), .Y(men_men_n1381_));
  OAI220     u1332(.A0(men_men_n1381_), .A1(x6), .B0(men_men_n1380_), .B1(men_men_n1379_), .Y(men_men_n1382_));
  NO2        u1333(.A(men_men_n1382_), .B(men_men_n1378_), .Y(men_men_n1383_));
  NAi21      u1334(.An(men_men_n116_), .B(men_men_n753_), .Y(men_men_n1384_));
  NA4        u1335(.A(men_men_n1384_), .B(men_men_n322_), .C(men_men_n294_), .D(men_men_n633_), .Y(men_men_n1385_));
  OAI220     u1336(.A0(men_men_n327_), .A1(x7), .B0(men_men_n132_), .B1(men_men_n71_), .Y(men_men_n1386_));
  NA3        u1337(.A(men_men_n1386_), .B(men_men_n796_), .C(men_men_n1105_), .Y(men_men_n1387_));
  NA2        u1338(.A(men_men_n82_), .B(men_men_n50_), .Y(men_men_n1388_));
  AO210      u1339(.A0(men_men_n1388_), .A1(men_men_n319_), .B0(men_men_n159_), .Y(men_men_n1389_));
  NA4        u1340(.A(men_men_n1389_), .B(men_men_n1387_), .C(men_men_n1385_), .D(men_men_n1383_), .Y(men_men_n1390_));
  OAI210     u1341(.A0(men_men_n1390_), .A1(men_men_n1377_), .B0(men_men_n56_), .Y(men_men_n1391_));
  AOI210     u1342(.A0(men_men_n699_), .A1(x4), .B0(men_men_n964_), .Y(men_men_n1392_));
  OAI220     u1343(.A0(men_men_n1392_), .A1(men_men_n305_), .B0(men_men_n1030_), .B1(men_men_n952_), .Y(men_men_n1393_));
  NA2        u1344(.A(men_men_n840_), .B(men_men_n412_), .Y(men_men_n1394_));
  OAI210     u1345(.A0(men_men_n1366_), .A1(men_men_n1358_), .B0(men_men_n295_), .Y(men_men_n1395_));
  OAI210     u1346(.A0(men_men_n1394_), .A1(men_men_n852_), .B0(men_men_n1395_), .Y(men_men_n1396_));
  OAI210     u1347(.A0(men_men_n1396_), .A1(men_men_n1393_), .B0(x6), .Y(men_men_n1397_));
  NO2        u1348(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n1398_));
  NO2        u1349(.A(x7), .B(x5), .Y(men_men_n1399_));
  AOI220     u1350(.A0(men_men_n861_), .A1(men_men_n1398_), .B0(men_men_n545_), .B1(men_men_n1399_), .Y(men_men_n1400_));
  NA2        u1351(.A(men_men_n769_), .B(men_men_n295_), .Y(men_men_n1401_));
  NA3        u1352(.A(men_men_n625_), .B(men_men_n297_), .C(men_men_n246_), .Y(men_men_n1402_));
  NA3        u1353(.A(men_men_n1402_), .B(men_men_n1401_), .C(men_men_n1400_), .Y(men_men_n1403_));
  NA2        u1354(.A(men_men_n1403_), .B(men_men_n430_), .Y(men_men_n1404_));
  AOI210     u1355(.A0(men_men_n383_), .A1(men_men_n344_), .B0(men_men_n55_), .Y(men_men_n1405_));
  NA4        u1356(.A(men_men_n1405_), .B(men_men_n1404_), .C(men_men_n1397_), .D(men_men_n1391_), .Y(men_men_n1406_));
  AO220      u1357(.A0(men_men_n1406_), .A1(men_men_n1372_), .B0(men_men_n1341_), .B1(men_men_n1335_), .Y(men16));
  NO2        u1358(.A(x4), .B(men_men_n59_), .Y(men_men_n1408_));
  NA2        u1359(.A(men_men_n672_), .B(men_men_n542_), .Y(men_men_n1409_));
  NA3        u1360(.A(men_men_n235_), .B(men_men_n437_), .C(men_men_n964_), .Y(men_men_n1410_));
  NA2        u1361(.A(men_men_n135_), .B(men_men_n211_), .Y(men_men_n1411_));
  AOI210     u1362(.A0(men_men_n1410_), .A1(men_men_n1409_), .B0(men_men_n1411_), .Y(men_men_n1412_));
  NO3        u1363(.A(x8), .B(x6), .C(men_men_n50_), .Y(men_men_n1413_));
  NO2        u1364(.A(men_men_n741_), .B(men_men_n189_), .Y(men_men_n1414_));
  OAI210     u1365(.A0(men_men_n1413_), .A1(men_men_n243_), .B0(men_men_n1414_), .Y(men_men_n1415_));
  NO2        u1366(.A(men_men_n163_), .B(x5), .Y(men_men_n1416_));
  NA2        u1367(.A(men_men_n1416_), .B(men_men_n1374_), .Y(men_men_n1417_));
  NA3        u1368(.A(men_men_n588_), .B(men_men_n544_), .C(men_men_n483_), .Y(men_men_n1418_));
  NA3        u1369(.A(men_men_n1418_), .B(men_men_n1417_), .C(men_men_n1415_), .Y(men_men_n1419_));
  OAI210     u1370(.A0(men_men_n1419_), .A1(men_men_n1412_), .B0(men_men_n1408_), .Y(men_men_n1420_));
  OAI210     u1371(.A0(men_men_n1287_), .A1(men_men_n931_), .B0(men_men_n427_), .Y(men_men_n1421_));
  NO2        u1372(.A(men_men_n324_), .B(x7), .Y(men_men_n1422_));
  NA2        u1373(.A(men_men_n1422_), .B(x0), .Y(men_men_n1423_));
  AOI210     u1374(.A0(men_men_n1423_), .A1(men_men_n1421_), .B0(men_men_n647_), .Y(men_men_n1424_));
  NA2        u1375(.A(men_men_n1084_), .B(men_men_n202_), .Y(men_men_n1425_));
  NA2        u1376(.A(men_men_n55_), .B(men_men_n108_), .Y(men_men_n1426_));
  NA2        u1377(.A(men_men_n1426_), .B(men_men_n693_), .Y(men_men_n1427_));
  NA2        u1378(.A(men_men_n382_), .B(men_men_n1088_), .Y(men_men_n1428_));
  OA220      u1379(.A0(men_men_n1428_), .A1(men_men_n1427_), .B0(men_men_n1425_), .B1(men_men_n641_), .Y(men_men_n1429_));
  OAI210     u1380(.A0(men_men_n1429_), .A1(men_men_n662_), .B0(men_men_n504_), .Y(men_men_n1430_));
  INV        u1381(.A(men_men_n1026_), .Y(men_men_n1431_));
  NO2        u1382(.A(men_men_n1431_), .B(men_men_n62_), .Y(men_men_n1432_));
  AOI220     u1383(.A0(men_men_n1432_), .A1(men_men_n274_), .B0(men_men_n1273_), .B1(men_men_n128_), .Y(men_men_n1433_));
  AOI220     u1384(.A0(men_men_n646_), .A1(men_men_n367_), .B0(men_men_n633_), .B1(men_men_n88_), .Y(men_men_n1434_));
  NA3        u1385(.A(men_men_n470_), .B(men_men_n595_), .C(men_men_n196_), .Y(men_men_n1435_));
  OAI220     u1386(.A0(men_men_n1435_), .A1(men_men_n1434_), .B0(men_men_n1433_), .B1(men_men_n315_), .Y(men_men_n1436_));
  NO3        u1387(.A(men_men_n1436_), .B(men_men_n1430_), .C(men_men_n1424_), .Y(men_men_n1437_));
  NO3        u1388(.A(x6), .B(x4), .C(x3), .Y(men_men_n1438_));
  NA2        u1389(.A(men_men_n1438_), .B(men_men_n541_), .Y(men_men_n1439_));
  NA4        u1390(.A(men_men_n717_), .B(men_men_n189_), .C(men_men_n58_), .D(x6), .Y(men_men_n1440_));
  AOI210     u1391(.A0(men_men_n1440_), .A1(men_men_n1439_), .B0(men_men_n54_), .Y(men_men_n1441_));
  NO2        u1392(.A(men_men_n729_), .B(x3), .Y(men_men_n1442_));
  AOI210     u1393(.A0(men_men_n671_), .A1(men_men_n150_), .B0(men_men_n1070_), .Y(men_men_n1443_));
  OA210      u1394(.A0(men_men_n1442_), .A1(men_men_n430_), .B0(men_men_n1443_), .Y(men_men_n1444_));
  NO3        u1395(.A(men_men_n506_), .B(men_men_n224_), .C(men_men_n75_), .Y(men_men_n1445_));
  NO2        u1396(.A(men_men_n769_), .B(men_men_n518_), .Y(men_men_n1446_));
  NO3        u1397(.A(men_men_n1446_), .B(men_men_n264_), .C(men_men_n158_), .Y(men_men_n1447_));
  NO4        u1398(.A(men_men_n1447_), .B(men_men_n1445_), .C(men_men_n1444_), .D(men_men_n1441_), .Y(men_men_n1448_));
  NA2        u1399(.A(men_men_n413_), .B(men_men_n964_), .Y(men_men_n1449_));
  NA4        u1400(.A(men_men_n489_), .B(men_men_n375_), .C(men_men_n226_), .D(x6), .Y(men_men_n1450_));
  OAI210     u1401(.A0(men_men_n729_), .A1(men_men_n1449_), .B0(men_men_n1450_), .Y(men_men_n1451_));
  NA2        u1402(.A(men_men_n913_), .B(men_men_n1318_), .Y(men_men_n1452_));
  NA2        u1403(.A(men_men_n738_), .B(x7), .Y(men_men_n1453_));
  OAI210     u1404(.A0(men_men_n1453_), .A1(men_men_n394_), .B0(men_men_n1452_), .Y(men_men_n1454_));
  NA2        u1405(.A(men_men_n281_), .B(x2), .Y(men_men_n1455_));
  NO3        u1406(.A(men_men_n1455_), .B(men_men_n603_), .C(men_men_n72_), .Y(men_men_n1456_));
  AOI210     u1407(.A0(men_men_n588_), .A1(men_men_n50_), .B0(men_men_n598_), .Y(men_men_n1457_));
  OAI210     u1408(.A0(men_men_n932_), .A1(men_men_n951_), .B0(men_men_n389_), .Y(men_men_n1458_));
  OAI220     u1409(.A0(men_men_n1458_), .A1(men_men_n1457_), .B0(men_men_n785_), .B1(men_men_n194_), .Y(men_men_n1459_));
  NO4        u1410(.A(men_men_n1459_), .B(men_men_n1456_), .C(men_men_n1454_), .D(men_men_n1451_), .Y(men_men_n1460_));
  OA220      u1411(.A0(men_men_n1460_), .A1(men_men_n450_), .B0(men_men_n1448_), .B1(men_men_n209_), .Y(men_men_n1461_));
  NO2        u1412(.A(men_men_n927_), .B(men_men_n55_), .Y(men_men_n1462_));
  NA2        u1413(.A(men_men_n424_), .B(men_men_n811_), .Y(men_men_n1463_));
  NO2        u1414(.A(men_men_n1463_), .B(men_men_n1462_), .Y(men_men_n1464_));
  NO3        u1415(.A(men_men_n965_), .B(men_men_n337_), .C(x8), .Y(men_men_n1465_));
  OAI210     u1416(.A0(men_men_n1465_), .A1(men_men_n1464_), .B0(x6), .Y(men_men_n1466_));
  NO2        u1417(.A(men_men_n1100_), .B(men_men_n1062_), .Y(men_men_n1467_));
  NA2        u1418(.A(men_men_n194_), .B(x7), .Y(men_men_n1468_));
  OAI220     u1419(.A0(men_men_n1468_), .A1(men_men_n1467_), .B0(men_men_n771_), .B1(men_men_n87_), .Y(men_men_n1469_));
  NA2        u1420(.A(men_men_n1469_), .B(men_men_n932_), .Y(men_men_n1470_));
  NA2        u1421(.A(men_men_n880_), .B(men_men_n71_), .Y(men_men_n1471_));
  OAI210     u1422(.A0(men_men_n1471_), .A1(men_men_n161_), .B0(men_men_n1015_), .Y(men_men_n1472_));
  AOI210     u1423(.A0(men_men_n506_), .A1(men_men_n57_), .B0(men_men_n641_), .Y(men_men_n1473_));
  NA3        u1424(.A(men_men_n232_), .B(men_men_n76_), .C(men_men_n71_), .Y(men_men_n1474_));
  OAI210     u1425(.A0(men_men_n923_), .A1(men_men_n235_), .B0(men_men_n1474_), .Y(men_men_n1475_));
  AOI210     u1426(.A0(men_men_n1473_), .A1(men_men_n1472_), .B0(men_men_n1475_), .Y(men_men_n1476_));
  NA3        u1427(.A(men_men_n1476_), .B(men_men_n1470_), .C(men_men_n1466_), .Y(men_men_n1477_));
  NO2        u1428(.A(men_men_n648_), .B(x6), .Y(men_men_n1478_));
  OAI210     u1429(.A0(men_men_n389_), .A1(men_men_n84_), .B0(men_men_n387_), .Y(men_men_n1479_));
  OA210      u1430(.A0(men_men_n1479_), .A1(men_men_n1478_), .B0(men_men_n133_), .Y(men_men_n1480_));
  NO3        u1431(.A(men_men_n452_), .B(men_men_n392_), .C(x7), .Y(men_men_n1481_));
  NO3        u1432(.A(men_men_n163_), .B(men_men_n75_), .C(x2), .Y(men_men_n1482_));
  NO3        u1433(.A(men_men_n1482_), .B(men_men_n1481_), .C(men_men_n1480_), .Y(men_men_n1483_));
  NO2        u1434(.A(men_men_n57_), .B(men_men_n108_), .Y(men_men_n1484_));
  AOI220     u1435(.A0(men_men_n771_), .A1(men_men_n782_), .B0(men_men_n521_), .B1(men_men_n285_), .Y(men_men_n1485_));
  NO2        u1436(.A(men_men_n1485_), .B(men_men_n1318_), .Y(men_men_n1486_));
  NO3        u1437(.A(men_men_n541_), .B(men_men_n176_), .C(men_men_n1062_), .Y(men_men_n1487_));
  NA2        u1438(.A(men_men_n951_), .B(x4), .Y(men_men_n1488_));
  OAI220     u1439(.A0(men_men_n1488_), .A1(men_men_n698_), .B0(men_men_n656_), .B1(men_men_n619_), .Y(men_men_n1489_));
  NO3        u1440(.A(men_men_n1489_), .B(men_men_n1487_), .C(men_men_n1486_), .Y(men_men_n1490_));
  OAI210     u1441(.A0(men_men_n1483_), .A1(x5), .B0(men_men_n1490_), .Y(men_men_n1491_));
  AOI220     u1442(.A0(men_men_n1491_), .A1(men_men_n99_), .B0(men_men_n1477_), .B1(men_men_n344_), .Y(men_men_n1492_));
  NA4        u1443(.A(men_men_n1492_), .B(men_men_n1461_), .C(men_men_n1437_), .D(men_men_n1420_), .Y(men17));
  NO4        u1444(.A(men_men_n610_), .B(men_men_n711_), .C(men_men_n102_), .D(men_men_n101_), .Y(men_men_n1494_));
  NO2        u1445(.A(men_men_n126_), .B(men_men_n1177_), .Y(men_men_n1495_));
  AOI220     u1446(.A0(men_men_n1495_), .A1(men_men_n723_), .B0(men_men_n1494_), .B1(men_men_n512_), .Y(men_men_n1496_));
  NA2        u1447(.A(men_men_n167_), .B(men_men_n78_), .Y(men_men_n1497_));
  NOi21      u1448(.An(men_men_n387_), .B(men_men_n84_), .Y(men_men_n1498_));
  OAI210     u1449(.A0(men_men_n633_), .A1(men_men_n55_), .B0(men_men_n1498_), .Y(men_men_n1499_));
  NA2        u1450(.A(men_men_n1231_), .B(men_men_n1021_), .Y(men_men_n1500_));
  NA4        u1451(.A(men_men_n1500_), .B(men_men_n1499_), .C(men_men_n741_), .D(men_men_n57_), .Y(men_men_n1501_));
  OAI210     u1452(.A0(men_men_n717_), .A1(x8), .B0(men_men_n1318_), .Y(men_men_n1502_));
  NA3        u1453(.A(men_men_n1502_), .B(men_men_n1257_), .C(men_men_n406_), .Y(men_men_n1503_));
  NA3        u1454(.A(men_men_n400_), .B(men_men_n274_), .C(men_men_n594_), .Y(men_men_n1504_));
  OA210      u1455(.A0(men_men_n1329_), .A1(men_men_n1170_), .B0(men_men_n761_), .Y(men_men_n1505_));
  NA4        u1456(.A(men_men_n1505_), .B(men_men_n1504_), .C(men_men_n1503_), .D(men_men_n1501_), .Y(men_men_n1506_));
  NA3        u1457(.A(men_men_n166_), .B(men_men_n639_), .C(men_men_n1062_), .Y(men_men_n1507_));
  AOI210     u1458(.A0(men_men_n1090_), .A1(men_men_n311_), .B0(men_men_n59_), .Y(men_men_n1508_));
  NA2        u1459(.A(men_men_n1508_), .B(men_men_n1507_), .Y(men_men_n1509_));
  AOI210     u1460(.A0(men_men_n1506_), .A1(x1), .B0(men_men_n1509_), .Y(men_men_n1510_));
  NO2        u1461(.A(men_men_n989_), .B(men_men_n506_), .Y(men_men_n1511_));
  OAI210     u1462(.A0(men_men_n1511_), .A1(men_men_n1074_), .B0(men_men_n616_), .Y(men_men_n1512_));
  NO3        u1463(.A(men_men_n641_), .B(men_men_n563_), .C(men_men_n532_), .Y(men_men_n1513_));
  OAI210     u1464(.A0(men_men_n1513_), .A1(men_men_n912_), .B0(men_men_n1442_), .Y(men_men_n1514_));
  AOI210     u1465(.A0(men_men_n1514_), .A1(men_men_n1512_), .B0(x8), .Y(men_men_n1515_));
  NA3        u1466(.A(men_men_n641_), .B(men_men_n277_), .C(men_men_n123_), .Y(men_men_n1516_));
  NO2        u1467(.A(men_men_n146_), .B(men_men_n144_), .Y(men_men_n1517_));
  NO3        u1468(.A(men_men_n907_), .B(men_men_n782_), .C(men_men_n711_), .Y(men_men_n1518_));
  AOI210     u1469(.A0(men_men_n1518_), .A1(men_men_n1517_), .B0(x0), .Y(men_men_n1519_));
  OAI210     u1470(.A0(men_men_n1516_), .A1(men_men_n253_), .B0(men_men_n1519_), .Y(men_men_n1520_));
  NO2        u1471(.A(men_men_n1520_), .B(men_men_n1515_), .Y(men_men_n1521_));
  OAI220     u1472(.A0(men_men_n1521_), .A1(men_men_n1510_), .B0(men_men_n1497_), .B1(men_men_n1496_), .Y(men18));
  AOI210     u1473(.A0(x8), .A1(x0), .B0(x5), .Y(men_men_n1523_));
  NOi31      u1474(.An(men_men_n311_), .B(men_men_n1523_), .C(men_men_n1060_), .Y(men_men_n1524_));
  NA2        u1475(.A(men_men_n610_), .B(men_men_n59_), .Y(men_men_n1525_));
  AOI210     u1476(.A0(men_men_n1425_), .A1(men_men_n355_), .B0(men_men_n1525_), .Y(men_men_n1526_));
  NO2        u1477(.A(men_men_n626_), .B(men_men_n783_), .Y(men_men_n1527_));
  NO4        u1478(.A(men_men_n260_), .B(men_men_n821_), .C(men_men_n157_), .D(men_men_n70_), .Y(men_men_n1528_));
  NO4        u1479(.A(men_men_n1528_), .B(men_men_n1527_), .C(men_men_n1526_), .D(men_men_n1524_), .Y(men_men_n1529_));
  NA3        u1480(.A(men_men_n527_), .B(men_men_n220_), .C(x0), .Y(men_men_n1530_));
  NAi21      u1481(.An(men_men_n393_), .B(men_men_n1530_), .Y(men_men_n1531_));
  NO2        u1482(.A(men_men_n897_), .B(x5), .Y(men_men_n1532_));
  AOI210     u1483(.A0(men_men_n1155_), .A1(x5), .B0(men_men_n1532_), .Y(men_men_n1533_));
  OA220      u1484(.A0(men_men_n527_), .A1(men_men_n337_), .B0(men_men_n406_), .B1(x5), .Y(men_men_n1534_));
  OAI220     u1485(.A0(men_men_n1534_), .A1(men_men_n299_), .B0(men_men_n1533_), .B1(men_men_n218_), .Y(men_men_n1535_));
  AOI210     u1486(.A0(men_men_n1531_), .A1(men_men_n297_), .B0(men_men_n1535_), .Y(men_men_n1536_));
  AOI210     u1487(.A0(men_men_n1536_), .A1(men_men_n1529_), .B0(x6), .Y(men_men_n1537_));
  NA3        u1488(.A(men_men_n531_), .B(men_men_n427_), .C(x2), .Y(men_men_n1538_));
  NA3        u1489(.A(men_men_n1060_), .B(men_men_n51_), .C(men_men_n57_), .Y(men_men_n1539_));
  AOI210     u1490(.A0(men_men_n1539_), .A1(men_men_n1538_), .B0(men_men_n796_), .Y(men_men_n1540_));
  AOI210     u1491(.A0(men_men_n431_), .A1(men_men_n140_), .B0(men_men_n794_), .Y(men_men_n1541_));
  NA2        u1492(.A(men_men_n274_), .B(x6), .Y(men_men_n1542_));
  OAI210     u1493(.A0(men_men_n182_), .A1(men_men_n110_), .B0(men_men_n1161_), .Y(men_men_n1543_));
  OAI220     u1494(.A0(men_men_n1543_), .A1(men_men_n1542_), .B0(men_men_n1541_), .B1(men_men_n753_), .Y(men_men_n1544_));
  OAI210     u1495(.A0(men_men_n1544_), .A1(men_men_n1540_), .B0(men_men_n53_), .Y(men_men_n1545_));
  NO2        u1496(.A(men_men_n697_), .B(men_men_n267_), .Y(men_men_n1546_));
  NO2        u1497(.A(men_men_n270_), .B(x3), .Y(men_men_n1547_));
  NO3        u1498(.A(men_men_n441_), .B(men_men_n610_), .C(men_men_n845_), .Y(men_men_n1548_));
  OAI210     u1499(.A0(men_men_n1548_), .A1(men_men_n1546_), .B0(men_men_n1547_), .Y(men_men_n1549_));
  AOI210     u1500(.A0(men_men_n1164_), .A1(men_men_n625_), .B0(x4), .Y(men_men_n1550_));
  OAI210     u1501(.A0(men_men_n563_), .A1(men_men_n610_), .B0(men_men_n59_), .Y(men_men_n1551_));
  OAI210     u1502(.A0(men_men_n633_), .A1(men_men_n658_), .B0(men_men_n1551_), .Y(men_men_n1552_));
  AO220      u1503(.A0(men_men_n1276_), .A1(men_men_n741_), .B0(men_men_n564_), .B1(men_men_n360_), .Y(men_men_n1553_));
  AOI220     u1504(.A0(men_men_n1553_), .A1(x1), .B0(men_men_n1552_), .B1(men_men_n164_), .Y(men_men_n1554_));
  NA4        u1505(.A(men_men_n1554_), .B(men_men_n1550_), .C(men_men_n1549_), .D(men_men_n1545_), .Y(men_men_n1555_));
  NO3        u1506(.A(men_men_n1081_), .B(men_men_n133_), .C(men_men_n132_), .Y(men_men_n1556_));
  OAI210     u1507(.A0(men_men_n1556_), .A1(men_men_n663_), .B0(men_men_n108_), .Y(men_men_n1557_));
  AOI210     u1508(.A0(men_men_n1557_), .A1(men_men_n569_), .B0(men_men_n796_), .Y(men_men_n1558_));
  NA3        u1509(.A(men_men_n1223_), .B(men_men_n194_), .C(men_men_n143_), .Y(men_men_n1559_));
  NA3        u1510(.A(men_men_n1084_), .B(men_men_n784_), .C(men_men_n348_), .Y(men_men_n1560_));
  NA2        u1511(.A(men_men_n174_), .B(men_men_n782_), .Y(men_men_n1561_));
  OAI210     u1512(.A0(men_men_n1561_), .A1(men_men_n1332_), .B0(men_men_n1560_), .Y(men_men_n1562_));
  AOI210     u1513(.A0(men_men_n1559_), .A1(men_men_n181_), .B0(men_men_n1562_), .Y(men_men_n1563_));
  OAI210     u1514(.A0(men_men_n1563_), .A1(men_men_n550_), .B0(x4), .Y(men_men_n1564_));
  OAI220     u1515(.A0(men_men_n1564_), .A1(men_men_n1558_), .B0(men_men_n1555_), .B1(men_men_n1537_), .Y(men_men_n1565_));
  NO2        u1516(.A(men_men_n149_), .B(men_men_n124_), .Y(men_men_n1566_));
  NO2        u1517(.A(men_men_n194_), .B(men_men_n811_), .Y(men_men_n1567_));
  AOI210     u1518(.A0(men_men_n611_), .A1(men_men_n518_), .B0(men_men_n1567_), .Y(men_men_n1568_));
  NO2        u1519(.A(men_men_n1568_), .B(x6), .Y(men_men_n1569_));
  NO2        u1520(.A(men_men_n392_), .B(men_men_n259_), .Y(men_men_n1570_));
  NO2        u1521(.A(men_men_n133_), .B(men_men_n743_), .Y(men_men_n1571_));
  NO2        u1522(.A(men_men_n965_), .B(men_men_n594_), .Y(men_men_n1572_));
  AO220      u1523(.A0(men_men_n1572_), .A1(men_men_n1571_), .B0(men_men_n1570_), .B1(men_men_n126_), .Y(men_men_n1573_));
  NO3        u1524(.A(men_men_n1573_), .B(men_men_n1569_), .C(men_men_n1566_), .Y(men_men_n1574_));
  NA2        u1525(.A(men_men_n1081_), .B(x3), .Y(men_men_n1575_));
  NA2        u1526(.A(men_men_n1369_), .B(men_men_n135_), .Y(men_men_n1576_));
  OAI220     u1527(.A0(men_men_n1576_), .A1(men_men_n1575_), .B0(men_men_n1574_), .B1(x3), .Y(men_men_n1577_));
  NO3        u1528(.A(men_men_n1011_), .B(men_men_n697_), .C(men_men_n332_), .Y(men_men_n1578_));
  AO210      u1529(.A0(men_men_n1040_), .A1(men_men_n304_), .B0(men_men_n1578_), .Y(men_men_n1579_));
  AOI220     u1530(.A0(men_men_n1579_), .A1(x8), .B0(men_men_n1369_), .B1(men_men_n442_), .Y(men_men_n1580_));
  NA2        u1531(.A(men_men_n757_), .B(men_men_n323_), .Y(men_men_n1581_));
  NO4        u1532(.A(men_men_n373_), .B(men_men_n207_), .C(men_men_n343_), .D(x2), .Y(men_men_n1582_));
  NA2        u1533(.A(men_men_n1426_), .B(men_men_n110_), .Y(men_men_n1583_));
  NO3        u1534(.A(men_men_n1225_), .B(men_men_n1004_), .C(men_men_n1161_), .Y(men_men_n1584_));
  AOI210     u1535(.A0(men_men_n1584_), .A1(men_men_n1583_), .B0(men_men_n1582_), .Y(men_men_n1585_));
  OA220      u1536(.A0(men_men_n1585_), .A1(men_men_n965_), .B0(men_men_n1581_), .B1(men_men_n578_), .Y(men_men_n1586_));
  OAI210     u1537(.A0(men_men_n1580_), .A1(men_men_n416_), .B0(men_men_n1586_), .Y(men_men_n1587_));
  AOI210     u1538(.A0(men_men_n1577_), .A1(men_men_n140_), .B0(men_men_n1587_), .Y(men_men_n1588_));
  NA2        u1539(.A(men_men_n1588_), .B(men_men_n1565_), .Y(men19));
  NO2        u1540(.A(men_men_n1471_), .B(men_men_n263_), .Y(men_men_n1590_));
  NA2        u1541(.A(men_men_n658_), .B(x3), .Y(men_men_n1591_));
  OAI210     u1542(.A0(men_men_n157_), .A1(men_men_n109_), .B0(men_men_n81_), .Y(men_men_n1592_));
  NA3        u1543(.A(men_men_n1592_), .B(men_men_n1591_), .C(men_men_n246_), .Y(men_men_n1593_));
  NO2        u1544(.A(men_men_n1327_), .B(men_men_n174_), .Y(men_men_n1594_));
  AOI210     u1545(.A0(men_men_n1494_), .A1(men_men_n358_), .B0(men_men_n1594_), .Y(men_men_n1595_));
  AOI210     u1546(.A0(men_men_n1595_), .A1(men_men_n1593_), .B0(men_men_n56_), .Y(men_men_n1596_));
  NO2        u1547(.A(men_men_n870_), .B(men_men_n1238_), .Y(men_men_n1597_));
  OAI210     u1548(.A0(men_men_n1596_), .A1(men_men_n1590_), .B0(men_men_n1597_), .Y(men_men_n1598_));
  NOi21      u1549(.An(men_men_n620_), .B(men_men_n662_), .Y(men_men_n1599_));
  AOI210     u1550(.A0(men_men_n358_), .A1(x6), .B0(men_men_n123_), .Y(men_men_n1600_));
  NO3        u1551(.A(men_men_n1600_), .B(men_men_n766_), .C(men_men_n128_), .Y(men_men_n1601_));
  NA2        u1552(.A(men_men_n1218_), .B(men_men_n124_), .Y(men_men_n1602_));
  NO4        u1553(.A(men_men_n1602_), .B(men_men_n1011_), .C(men_men_n897_), .D(men_men_n77_), .Y(men_men_n1603_));
  NO3        u1554(.A(men_men_n1603_), .B(men_men_n1601_), .C(men_men_n1037_), .Y(men_men_n1604_));
  NO2        u1555(.A(men_men_n550_), .B(men_men_n629_), .Y(men_men_n1605_));
  NA2        u1556(.A(men_men_n1272_), .B(men_men_n50_), .Y(men_men_n1606_));
  NO3        u1557(.A(men_men_n525_), .B(men_men_n313_), .C(men_men_n64_), .Y(men_men_n1607_));
  AOI220     u1558(.A0(men_men_n1607_), .A1(men_men_n1606_), .B0(men_men_n1605_), .B1(men_men_n784_), .Y(men_men_n1608_));
  OAI210     u1559(.A0(men_men_n1604_), .A1(men_men_n57_), .B0(men_men_n1608_), .Y(men_men_n1609_));
  AOI210     u1560(.A0(men_men_n1609_), .A1(men_men_n782_), .B0(men_men_n1599_), .Y(men_men_n1610_));
  AOI210     u1561(.A0(men_men_n831_), .A1(men_men_n743_), .B0(men_men_n772_), .Y(men_men_n1611_));
  NO2        u1562(.A(men_men_n1611_), .B(x4), .Y(men_men_n1612_));
  NA3        u1563(.A(men_men_n741_), .B(men_men_n262_), .C(x7), .Y(men_men_n1613_));
  AOI220     u1564(.A0(men_men_n1422_), .A1(men_men_n796_), .B0(men_men_n711_), .B1(men_men_n1177_), .Y(men_men_n1614_));
  AOI210     u1565(.A0(men_men_n1614_), .A1(men_men_n1613_), .B0(men_men_n510_), .Y(men_men_n1615_));
  OAI210     u1566(.A0(men_men_n1615_), .A1(men_men_n1612_), .B0(men_men_n821_), .Y(men_men_n1616_));
  NO2        u1567(.A(men_men_n753_), .B(men_men_n327_), .Y(men_men_n1617_));
  NO2        u1568(.A(men_men_n157_), .B(men_men_n1036_), .Y(men_men_n1618_));
  AOI220     u1569(.A0(men_men_n1618_), .A1(men_men_n1287_), .B0(men_men_n1617_), .B1(men_men_n484_), .Y(men_men_n1619_));
  AO210      u1570(.A0(men_men_n1619_), .A1(men_men_n1616_), .B0(x1), .Y(men_men_n1620_));
  NA3        u1571(.A(men_men_n641_), .B(men_men_n1062_), .C(men_men_n1210_), .Y(men_men_n1621_));
  NA2        u1572(.A(men_men_n150_), .B(men_men_n111_), .Y(men_men_n1622_));
  NOi21      u1573(.An(x1), .B(x6), .Y(men_men_n1623_));
  NA2        u1574(.A(men_men_n1623_), .B(men_men_n84_), .Y(men_men_n1624_));
  NA3        u1575(.A(men_men_n1624_), .B(men_men_n1622_), .C(men_men_n1621_), .Y(men_men_n1625_));
  AOI220     u1576(.A0(men_men_n1625_), .A1(x3), .B0(men_men_n1226_), .B1(men_men_n388_), .Y(men_men_n1626_));
  NA3        u1577(.A(men_men_n1231_), .B(men_men_n806_), .C(men_men_n612_), .Y(men_men_n1627_));
  AOI220     u1578(.A0(men_men_n1276_), .A1(men_men_n123_), .B0(men_men_n927_), .B1(men_men_n823_), .Y(men_men_n1628_));
  AOI210     u1579(.A0(men_men_n1628_), .A1(men_men_n1627_), .B0(men_men_n327_), .Y(men_men_n1629_));
  NA2        u1580(.A(men_men_n951_), .B(men_men_n50_), .Y(men_men_n1630_));
  NA3        u1581(.A(men_men_n1218_), .B(men_men_n389_), .C(men_men_n110_), .Y(men_men_n1631_));
  AOI210     u1582(.A0(men_men_n1631_), .A1(men_men_n1630_), .B0(men_men_n974_), .Y(men_men_n1632_));
  NO3        u1583(.A(men_men_n627_), .B(men_men_n524_), .C(men_men_n1244_), .Y(men_men_n1633_));
  NO3        u1584(.A(men_men_n1633_), .B(men_men_n1632_), .C(men_men_n1629_), .Y(men_men_n1634_));
  OAI210     u1585(.A0(men_men_n1626_), .A1(men_men_n857_), .B0(men_men_n1634_), .Y(men_men_n1635_));
  NO2        u1586(.A(men_men_n563_), .B(men_men_n68_), .Y(men_men_n1636_));
  OAI220     u1587(.A0(men_men_n1636_), .A1(men_men_n1591_), .B0(men_men_n312_), .B1(men_men_n905_), .Y(men_men_n1637_));
  AOI220     u1588(.A0(men_men_n1637_), .A1(men_men_n56_), .B0(men_men_n1374_), .B1(men_men_n738_), .Y(men_men_n1638_));
  NO2        u1589(.A(men_men_n54_), .B(men_men_n71_), .Y(men_men_n1639_));
  AO220      u1590(.A0(men_men_n1639_), .A1(men_men_n1011_), .B0(men_men_n823_), .B1(men_men_n964_), .Y(men_men_n1640_));
  NA2        u1591(.A(men_men_n1201_), .B(men_men_n365_), .Y(men_men_n1641_));
  NO2        u1592(.A(men_men_n1004_), .B(men_men_n1623_), .Y(men_men_n1642_));
  NA2        u1593(.A(men_men_n506_), .B(men_men_n738_), .Y(men_men_n1643_));
  OAI210     u1594(.A0(men_men_n1643_), .A1(men_men_n1642_), .B0(men_men_n1641_), .Y(men_men_n1644_));
  AOI210     u1595(.A0(men_men_n1640_), .A1(x2), .B0(men_men_n1644_), .Y(men_men_n1645_));
  OAI220     u1596(.A0(men_men_n1645_), .A1(men_men_n157_), .B0(men_men_n1638_), .B1(men_men_n54_), .Y(men_men_n1646_));
  OAI210     u1597(.A0(men_men_n1646_), .A1(men_men_n1635_), .B0(x8), .Y(men_men_n1647_));
  NA4        u1598(.A(men_men_n1647_), .B(men_men_n1620_), .C(men_men_n1610_), .D(men_men_n1598_), .Y(men20));
  NA4        u1599(.A(men_men_n399_), .B(men_men_n285_), .C(men_men_n387_), .D(men_men_n62_), .Y(men_men_n1649_));
  NA2        u1600(.A(men_men_n484_), .B(men_men_n420_), .Y(men_men_n1650_));
  AOI210     u1601(.A0(men_men_n1650_), .A1(men_men_n1649_), .B0(men_men_n87_), .Y(men_men_n1651_));
  AOI210     u1602(.A0(men_men_n1066_), .A1(men_men_n62_), .B0(men_men_n1605_), .Y(men_men_n1652_));
  AOI210     u1603(.A0(men_men_n998_), .A1(men_men_n354_), .B0(men_men_n1208_), .Y(men_men_n1653_));
  OAI210     u1604(.A0(men_men_n1652_), .A1(men_men_n693_), .B0(men_men_n1653_), .Y(men_men_n1654_));
  OAI210     u1605(.A0(men_men_n1654_), .A1(men_men_n1651_), .B0(men_men_n1122_), .Y(men_men_n1655_));
  NAi21      u1606(.An(men_men_n559_), .B(men_men_n408_), .Y(men_men_n1656_));
  NA3        u1607(.A(men_men_n1656_), .B(men_men_n996_), .C(men_men_n964_), .Y(men_men_n1657_));
  NA3        u1608(.A(men_men_n1121_), .B(men_men_n285_), .C(men_men_n593_), .Y(men_men_n1658_));
  AOI210     u1609(.A0(men_men_n1658_), .A1(men_men_n1657_), .B0(men_men_n1318_), .Y(men_men_n1659_));
  NO2        u1610(.A(men_men_n757_), .B(men_men_n984_), .Y(men_men_n1660_));
  NOi31      u1611(.An(men_men_n1660_), .B(men_men_n1193_), .C(men_men_n537_), .Y(men_men_n1661_));
  OAI210     u1612(.A0(men_men_n1661_), .A1(men_men_n1659_), .B0(men_men_n332_), .Y(men_men_n1662_));
  NO4        u1613(.A(men_men_n554_), .B(men_men_n241_), .C(x5), .D(x2), .Y(men_men_n1663_));
  NA2        u1614(.A(men_men_n323_), .B(men_men_n93_), .Y(men_men_n1664_));
  NA2        u1615(.A(men_men_n333_), .B(men_men_n108_), .Y(men_men_n1665_));
  NA2        u1616(.A(men_men_n430_), .B(men_men_n52_), .Y(men_men_n1666_));
  OAI220     u1617(.A0(men_men_n1666_), .A1(men_men_n1665_), .B0(men_men_n1664_), .B1(men_men_n280_), .Y(men_men_n1667_));
  OAI210     u1618(.A0(men_men_n1667_), .A1(men_men_n1663_), .B0(men_men_n226_), .Y(men_men_n1668_));
  NO2        u1619(.A(men_men_n677_), .B(men_men_n616_), .Y(men_men_n1669_));
  NA2        u1620(.A(men_men_n965_), .B(men_men_n50_), .Y(men_men_n1670_));
  NO3        u1621(.A(men_men_n1670_), .B(men_men_n371_), .C(men_men_n234_), .Y(men_men_n1671_));
  NA4        u1622(.A(men_men_n344_), .B(men_men_n243_), .C(men_men_n811_), .D(men_men_n64_), .Y(men_men_n1672_));
  OAI220     u1623(.A0(men_men_n1672_), .A1(men_men_n687_), .B0(men_men_n1488_), .B1(men_men_n1049_), .Y(men_men_n1673_));
  AOI210     u1624(.A0(men_men_n1671_), .A1(men_men_n1669_), .B0(men_men_n1673_), .Y(men_men_n1674_));
  NA4        u1625(.A(men_men_n1674_), .B(men_men_n1668_), .C(men_men_n1662_), .D(men_men_n1655_), .Y(men21));
  OAI210     u1626(.A0(men_men_n413_), .A1(men_men_n54_), .B0(x7), .Y(men_men_n1676_));
  OAI220     u1627(.A0(men_men_n1676_), .A1(men_men_n1307_), .B0(men_men_n1067_), .B1(men_men_n96_), .Y(men_men_n1677_));
  NA2        u1628(.A(men_men_n1677_), .B(men_men_n78_), .Y(men_men_n1678_));
  NA2        u1629(.A(men_men_n297_), .B(men_men_n868_), .Y(men_men_n1679_));
  AOI220     u1630(.A0(men_men_n1679_), .A1(men_men_n315_), .B0(men_men_n578_), .B1(men_men_n468_), .Y(men_men_n1680_));
  NA2        u1631(.A(men_men_n951_), .B(men_men_n279_), .Y(men_men_n1681_));
  NA2        u1632(.A(men_men_n545_), .B(men_men_n469_), .Y(men_men_n1682_));
  NA4        u1633(.A(men_men_n1682_), .B(men_men_n1681_), .C(men_men_n1401_), .D(men_men_n56_), .Y(men_men_n1683_));
  NO2        u1634(.A(men_men_n784_), .B(men_men_n441_), .Y(men_men_n1684_));
  NO3        u1635(.A(men_men_n1684_), .B(men_men_n730_), .C(men_men_n255_), .Y(men_men_n1685_));
  NOi31      u1636(.An(men_men_n197_), .B(men_men_n641_), .C(men_men_n1105_), .Y(men_men_n1686_));
  NO4        u1637(.A(men_men_n1686_), .B(men_men_n1685_), .C(men_men_n1683_), .D(men_men_n1680_), .Y(men_men_n1687_));
  NO3        u1638(.A(men_men_n441_), .B(men_men_n283_), .C(men_men_n52_), .Y(men_men_n1688_));
  OA210      u1639(.A0(men_men_n1688_), .A1(men_men_n894_), .B0(x3), .Y(men_men_n1689_));
  OAI210     u1640(.A0(men_men_n795_), .A1(men_men_n598_), .B0(men_men_n346_), .Y(men_men_n1690_));
  NO2        u1641(.A(men_men_n70_), .B(x2), .Y(men_men_n1691_));
  OAI210     u1642(.A0(men_men_n181_), .A1(x0), .B0(men_men_n1691_), .Y(men_men_n1692_));
  NA2        u1643(.A(men_men_n147_), .B(men_men_n108_), .Y(men_men_n1693_));
  NA3        u1644(.A(men_men_n1693_), .B(men_men_n1692_), .C(men_men_n1690_), .Y(men_men_n1694_));
  OAI210     u1645(.A0(men_men_n1694_), .A1(men_men_n1689_), .B0(x8), .Y(men_men_n1695_));
  NO3        u1646(.A(men_men_n783_), .B(men_men_n630_), .C(men_men_n594_), .Y(men_men_n1696_));
  NA2        u1647(.A(men_men_n55_), .B(men_men_n50_), .Y(men_men_n1697_));
  MUX2       u1648(.S(men_men_n610_), .A(men_men_n1697_), .B(men_men_n107_), .Y(men_men_n1698_));
  AOI210     u1649(.A0(men_men_n1379_), .A1(men_men_n244_), .B0(men_men_n1698_), .Y(men_men_n1699_));
  OAI210     u1650(.A0(men_men_n654_), .A1(men_men_n593_), .B0(x4), .Y(men_men_n1700_));
  NO3        u1651(.A(men_men_n1700_), .B(men_men_n1699_), .C(men_men_n1696_), .Y(men_men_n1701_));
  AO220      u1652(.A0(men_men_n1701_), .A1(men_men_n1695_), .B0(men_men_n1687_), .B1(men_men_n1678_), .Y(men_men_n1702_));
  AO220      u1653(.A0(men_men_n642_), .A1(men_men_n327_), .B0(men_men_n599_), .B1(x8), .Y(men_men_n1703_));
  NO2        u1654(.A(men_men_n870_), .B(x0), .Y(men_men_n1704_));
  NO3        u1655(.A(men_men_n1704_), .B(men_men_n555_), .C(men_men_n88_), .Y(men_men_n1705_));
  NO2        u1656(.A(men_men_n163_), .B(x2), .Y(men_men_n1706_));
  NO3        u1657(.A(men_men_n384_), .B(men_men_n260_), .C(men_men_n189_), .Y(men_men_n1707_));
  AOI210     u1658(.A0(men_men_n1706_), .A1(men_men_n68_), .B0(men_men_n1707_), .Y(men_men_n1708_));
  OAI210     u1659(.A0(men_men_n1705_), .A1(men_men_n406_), .B0(men_men_n1708_), .Y(men_men_n1709_));
  AOI220     u1660(.A0(men_men_n1709_), .A1(x5), .B0(men_men_n1703_), .B1(men_men_n757_), .Y(men_men_n1710_));
  AOI210     u1661(.A0(men_men_n1710_), .A1(men_men_n1702_), .B0(men_men_n71_), .Y(men_men_n1711_));
  NO2        u1662(.A(men_men_n917_), .B(men_men_n172_), .Y(men_men_n1712_));
  NOi41      u1663(.An(men_men_n1455_), .B(men_men_n1523_), .C(men_men_n1176_), .D(men_men_n861_), .Y(men_men_n1713_));
  NA2        u1664(.A(men_men_n1713_), .B(men_men_n1712_), .Y(men_men_n1714_));
  NO2        u1665(.A(men_men_n78_), .B(x4), .Y(men_men_n1715_));
  OAI210     u1666(.A0(men_men_n295_), .A1(men_men_n161_), .B0(men_men_n1715_), .Y(men_men_n1716_));
  OAI210     u1667(.A0(men_men_n415_), .A1(men_men_n431_), .B0(men_men_n234_), .Y(men_men_n1717_));
  NO2        u1668(.A(men_men_n262_), .B(men_men_n50_), .Y(men_men_n1718_));
  NO2        u1669(.A(men_men_n1718_), .B(men_men_n57_), .Y(men_men_n1719_));
  NA2        u1670(.A(men_men_n1719_), .B(men_men_n1717_), .Y(men_men_n1720_));
  AOI210     u1671(.A0(men_men_n1716_), .A1(men_men_n1714_), .B0(men_men_n1720_), .Y(men_men_n1721_));
  NA2        u1672(.A(men_men_n769_), .B(men_men_n559_), .Y(men_men_n1722_));
  AO210      u1673(.A0(men_men_n1722_), .A1(men_men_n974_), .B0(men_men_n50_), .Y(men_men_n1723_));
  NO2        u1674(.A(men_men_n1656_), .B(men_men_n1238_), .Y(men_men_n1724_));
  AOI220     u1675(.A0(men_men_n1724_), .A1(men_men_n1186_), .B0(men_men_n1346_), .B1(men_men_n1060_), .Y(men_men_n1725_));
  AOI210     u1676(.A0(men_men_n1725_), .A1(men_men_n1723_), .B0(men_men_n110_), .Y(men_men_n1726_));
  NA2        u1677(.A(men_men_n304_), .B(men_men_n108_), .Y(men_men_n1727_));
  NA2        u1678(.A(men_men_n904_), .B(men_men_n55_), .Y(men_men_n1728_));
  NO2        u1679(.A(men_men_n1728_), .B(men_men_n1727_), .Y(men_men_n1729_));
  NO2        u1680(.A(men_men_n682_), .B(men_men_n1070_), .Y(men_men_n1730_));
  NO4        u1681(.A(men_men_n1730_), .B(men_men_n1729_), .C(men_men_n1726_), .D(men_men_n1721_), .Y(men_men_n1731_));
  NO2        u1682(.A(men_men_n1731_), .B(x6), .Y(men_men_n1732_));
  AOI210     u1683(.A0(men_men_n619_), .A1(men_men_n1070_), .B0(men_men_n1523_), .Y(men_men_n1733_));
  OAI210     u1684(.A0(men_men_n1733_), .A1(men_men_n700_), .B0(men_men_n56_), .Y(men_men_n1734_));
  NO2        u1685(.A(men_men_n759_), .B(men_men_n54_), .Y(men_men_n1735_));
  NO4        u1686(.A(men_men_n972_), .B(men_men_n283_), .C(men_men_n782_), .D(men_men_n766_), .Y(men_men_n1736_));
  NO2        u1687(.A(men_men_n875_), .B(x5), .Y(men_men_n1737_));
  NO4        u1688(.A(men_men_n1737_), .B(men_men_n1736_), .C(men_men_n1735_), .D(men_men_n958_), .Y(men_men_n1738_));
  AOI210     u1689(.A0(men_men_n1738_), .A1(men_men_n1734_), .B0(men_men_n50_), .Y(men_men_n1739_));
  NA2        u1690(.A(men_men_n163_), .B(men_men_n108_), .Y(men_men_n1740_));
  OA220      u1691(.A0(men_men_n1740_), .A1(men_men_n445_), .B0(men_men_n474_), .B1(men_men_n757_), .Y(men_men_n1741_));
  NA3        u1692(.A(men_men_n55_), .B(x2), .C(x0), .Y(men_men_n1742_));
  AOI220     u1693(.A0(men_men_n1742_), .A1(men_men_n174_), .B0(men_men_n875_), .B1(men_men_n159_), .Y(men_men_n1743_));
  NO2        u1694(.A(men_men_n693_), .B(men_men_n262_), .Y(men_men_n1744_));
  NO3        u1695(.A(men_men_n250_), .B(men_men_n232_), .C(men_men_n365_), .Y(men_men_n1745_));
  NO3        u1696(.A(men_men_n1745_), .B(men_men_n1744_), .C(men_men_n1743_), .Y(men_men_n1746_));
  OAI220     u1697(.A0(men_men_n1746_), .A1(men_men_n56_), .B0(men_men_n1741_), .B1(men_men_n709_), .Y(men_men_n1747_));
  OAI210     u1698(.A0(men_men_n1747_), .A1(men_men_n1739_), .B0(men_men_n116_), .Y(men_men_n1748_));
  NO2        u1699(.A(men_men_n624_), .B(men_men_n310_), .Y(men_men_n1749_));
  AOI210     u1700(.A0(men_men_n617_), .A1(x5), .B0(men_men_n1749_), .Y(men_men_n1750_));
  NO2        u1701(.A(men_men_n1750_), .B(men_men_n110_), .Y(men_men_n1751_));
  NA2        u1702(.A(men_men_n717_), .B(men_men_n81_), .Y(men_men_n1752_));
  NA3        u1703(.A(men_men_n1752_), .B(men_men_n438_), .C(men_men_n57_), .Y(men_men_n1753_));
  OAI210     u1704(.A0(men_men_n1728_), .A1(men_men_n1727_), .B0(men_men_n1753_), .Y(men_men_n1754_));
  OAI210     u1705(.A0(men_men_n1754_), .A1(men_men_n1751_), .B0(x1), .Y(men_men_n1755_));
  NO4        u1706(.A(men_men_n424_), .B(men_men_n78_), .C(men_men_n151_), .D(x3), .Y(men_men_n1756_));
  NO2        u1707(.A(men_men_n333_), .B(men_men_n112_), .Y(men_men_n1757_));
  OAI210     u1708(.A0(men_men_n1756_), .A1(men_men_n1319_), .B0(men_men_n1757_), .Y(men_men_n1758_));
  NO2        u1709(.A(men_men_n60_), .B(men_men_n108_), .Y(men_men_n1759_));
  NO4        u1710(.A(men_men_n1727_), .B(men_men_n972_), .C(men_men_n677_), .D(men_men_n50_), .Y(men_men_n1760_));
  AOI210     u1711(.A0(men_men_n1759_), .A1(men_men_n1567_), .B0(men_men_n1760_), .Y(men_men_n1761_));
  NA4        u1712(.A(men_men_n1761_), .B(men_men_n1758_), .C(men_men_n1755_), .D(men_men_n1748_), .Y(men_men_n1762_));
  NO3        u1713(.A(men_men_n1762_), .B(men_men_n1732_), .C(men_men_n1711_), .Y(men22));
  AOI210     u1714(.A0(men_men_n531_), .A1(men_men_n71_), .B0(men_men_n477_), .Y(men_men_n1764_));
  NO2        u1715(.A(men_men_n1213_), .B(men_men_n563_), .Y(men_men_n1765_));
  AOI210     u1716(.A0(x5), .A1(x2), .B0(x8), .Y(men_men_n1766_));
  NA2        u1717(.A(men_men_n1766_), .B(men_men_n59_), .Y(men_men_n1767_));
  OAI220     u1718(.A0(men_men_n1767_), .A1(men_men_n1765_), .B0(men_men_n1764_), .B1(men_men_n406_), .Y(men_men_n1768_));
  NA2        u1719(.A(men_men_n593_), .B(men_men_n87_), .Y(men_men_n1769_));
  NA2        u1720(.A(men_men_n280_), .B(men_men_n77_), .Y(men_men_n1770_));
  OA220      u1721(.A0(men_men_n1770_), .A1(men_men_n1769_), .B0(men_men_n854_), .B1(men_men_n1021_), .Y(men_men_n1771_));
  NO4        u1722(.A(men_men_n392_), .B(men_men_n224_), .C(men_men_n71_), .D(x3), .Y(men_men_n1772_));
  NO3        u1723(.A(men_men_n1267_), .B(men_men_n87_), .C(x0), .Y(men_men_n1773_));
  OAI210     u1724(.A0(men_men_n406_), .A1(men_men_n209_), .B0(x4), .Y(men_men_n1774_));
  NO3        u1725(.A(men_men_n1774_), .B(men_men_n1773_), .C(men_men_n1772_), .Y(men_men_n1775_));
  OAI210     u1726(.A0(men_men_n1771_), .A1(men_men_n202_), .B0(men_men_n1775_), .Y(men_men_n1776_));
  AOI210     u1727(.A0(men_men_n1768_), .A1(men_men_n53_), .B0(men_men_n1776_), .Y(men_men_n1777_));
  NA2        u1728(.A(men_men_n308_), .B(men_men_n313_), .Y(men_men_n1778_));
  NA3        u1729(.A(men_men_n1778_), .B(men_men_n226_), .C(men_men_n312_), .Y(men_men_n1779_));
  NA2        u1730(.A(men_men_n588_), .B(men_men_n249_), .Y(men_men_n1780_));
  NO3        u1731(.A(men_men_n506_), .B(men_men_n270_), .C(men_men_n218_), .Y(men_men_n1781_));
  NAi31      u1732(.An(men_men_n1781_), .B(men_men_n1780_), .C(men_men_n1779_), .Y(men_men_n1782_));
  NO2        u1733(.A(men_men_n474_), .B(men_men_n264_), .Y(men_men_n1783_));
  NO2        u1734(.A(men_men_n1267_), .B(x3), .Y(men_men_n1784_));
  AOI210     u1735(.A0(men_men_n1784_), .A1(men_men_n354_), .B0(men_men_n1783_), .Y(men_men_n1785_));
  OAI210     u1736(.A0(men_men_n1100_), .A1(men_men_n191_), .B0(men_men_n56_), .Y(men_men_n1786_));
  NA3        u1737(.A(men_men_n55_), .B(men_men_n71_), .C(x0), .Y(men_men_n1787_));
  OAI220     u1738(.A0(men_men_n1787_), .A1(men_men_n1070_), .B0(men_men_n371_), .B1(men_men_n217_), .Y(men_men_n1788_));
  NO2        u1739(.A(men_men_n1788_), .B(men_men_n1786_), .Y(men_men_n1789_));
  OAI210     u1740(.A0(men_men_n1785_), .A1(men_men_n262_), .B0(men_men_n1789_), .Y(men_men_n1790_));
  AOI210     u1741(.A0(men_men_n1782_), .A1(men_men_n108_), .B0(men_men_n1790_), .Y(men_men_n1791_));
  NO2        u1742(.A(men_men_n962_), .B(men_men_n879_), .Y(men_men_n1792_));
  NO2        u1743(.A(men_men_n813_), .B(men_men_n163_), .Y(men_men_n1793_));
  OAI210     u1744(.A0(men_men_n1793_), .A1(men_men_n1792_), .B0(men_men_n623_), .Y(men_men_n1794_));
  OA210      u1745(.A0(men_men_n1791_), .A1(men_men_n1777_), .B0(men_men_n1794_), .Y(men_men_n1795_));
  OAI210     u1746(.A0(men_men_n1195_), .A1(men_men_n716_), .B0(men_men_n704_), .Y(men_men_n1796_));
  NO2        u1747(.A(men_men_n359_), .B(x0), .Y(men_men_n1797_));
  NA3        u1748(.A(men_men_n1797_), .B(men_men_n354_), .C(men_men_n56_), .Y(men_men_n1798_));
  AOI210     u1749(.A0(men_men_n1798_), .A1(men_men_n1796_), .B0(men_men_n406_), .Y(men_men_n1799_));
  NO3        u1750(.A(men_men_n174_), .B(men_men_n163_), .C(men_men_n62_), .Y(men_men_n1800_));
  OAI210     u1751(.A0(men_men_n1800_), .A1(men_men_n426_), .B0(men_men_n110_), .Y(men_men_n1801_));
  NA2        u1752(.A(men_men_n143_), .B(men_men_n796_), .Y(men_men_n1802_));
  NA2        u1753(.A(men_men_n424_), .B(x3), .Y(men_men_n1803_));
  NAi31      u1754(.An(men_men_n1803_), .B(men_men_n1802_), .C(men_men_n1583_), .Y(men_men_n1804_));
  NO3        u1755(.A(men_men_n870_), .B(men_men_n473_), .C(men_men_n110_), .Y(men_men_n1805_));
  NO2        u1756(.A(men_men_n1102_), .B(men_men_n144_), .Y(men_men_n1806_));
  NO3        u1757(.A(men_men_n907_), .B(men_men_n420_), .C(men_men_n309_), .Y(men_men_n1807_));
  AOI220     u1758(.A0(men_men_n1807_), .A1(men_men_n1806_), .B0(men_men_n1805_), .B1(men_men_n1797_), .Y(men_men_n1808_));
  NA3        u1759(.A(men_men_n420_), .B(men_men_n93_), .C(men_men_n81_), .Y(men_men_n1809_));
  AOI210     u1760(.A0(men_men_n619_), .A1(men_men_n463_), .B0(men_men_n503_), .Y(men_men_n1810_));
  NA2        u1761(.A(men_men_n1197_), .B(x3), .Y(men_men_n1811_));
  OAI210     u1762(.A0(men_men_n1811_), .A1(men_men_n1810_), .B0(men_men_n1809_), .Y(men_men_n1812_));
  NA3        u1763(.A(men_men_n56_), .B(men_men_n50_), .C(x0), .Y(men_men_n1813_));
  NOi21      u1764(.An(men_men_n83_), .B(men_men_n741_), .Y(men_men_n1814_));
  NA3        u1765(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n1815_));
  NA3        u1766(.A(men_men_n1815_), .B(men_men_n1004_), .C(men_men_n271_), .Y(men_men_n1816_));
  OAI220     u1767(.A0(men_men_n1816_), .A1(men_men_n1814_), .B0(men_men_n1073_), .B1(men_men_n1813_), .Y(men_men_n1817_));
  AOI220     u1768(.A0(men_men_n1817_), .A1(men_men_n1084_), .B0(men_men_n1812_), .B1(men_men_n354_), .Y(men_men_n1818_));
  NA4        u1769(.A(men_men_n1818_), .B(men_men_n1808_), .C(men_men_n1804_), .D(men_men_n1801_), .Y(men_men_n1819_));
  AOI210     u1770(.A0(men_men_n1819_), .A1(x7), .B0(men_men_n1799_), .Y(men_men_n1820_));
  OAI210     u1771(.A0(men_men_n1795_), .A1(x7), .B0(men_men_n1820_), .Y(men23));
  OR2        u1772(.A(men_men_n525_), .B(men_men_n226_), .Y(men_men_n1822_));
  AOI220     u1773(.A0(men_men_n1822_), .A1(men_men_n1660_), .B0(men_men_n625_), .B1(men_men_n300_), .Y(men_men_n1823_));
  NO3        u1774(.A(men_men_n854_), .B(men_men_n602_), .C(men_men_n496_), .Y(men_men_n1824_));
  NO3        u1775(.A(men_men_n966_), .B(men_men_n152_), .C(men_men_n117_), .Y(men_men_n1825_));
  AOI210     u1776(.A0(men_men_n1825_), .A1(men_men_n1043_), .B0(men_men_n1824_), .Y(men_men_n1826_));
  OAI210     u1777(.A0(men_men_n1823_), .A1(men_men_n157_), .B0(men_men_n1826_), .Y(men_men_n1827_));
  NA2        u1778(.A(men_men_n1827_), .B(men_men_n55_), .Y(men_men_n1828_));
  NO2        u1779(.A(men_men_n972_), .B(men_men_n523_), .Y(men_men_n1829_));
  AO220      u1780(.A0(men_men_n1303_), .A1(men_men_n185_), .B0(men_men_n1011_), .B1(men_men_n757_), .Y(men_men_n1830_));
  OAI210     u1781(.A0(men_men_n1830_), .A1(men_men_n1829_), .B0(men_men_n599_), .Y(men_men_n1831_));
  NA2        u1782(.A(men_men_n182_), .B(men_men_n172_), .Y(men_men_n1832_));
  NA2        u1783(.A(men_men_n412_), .B(men_men_n164_), .Y(men_men_n1833_));
  AOI210     u1784(.A0(men_men_n1833_), .A1(men_men_n1832_), .B0(men_men_n241_), .Y(men_men_n1834_));
  NA3        u1785(.A(men_men_n879_), .B(men_men_n431_), .C(men_men_n262_), .Y(men_men_n1835_));
  AOI210     u1786(.A0(men_men_n1835_), .A1(men_men_n508_), .B0(men_men_n389_), .Y(men_men_n1836_));
  OAI210     u1787(.A0(men_men_n1836_), .A1(men_men_n1834_), .B0(men_men_n304_), .Y(men_men_n1837_));
  NA3        u1788(.A(men_men_n57_), .B(x4), .C(x3), .Y(men_men_n1838_));
  NO3        u1789(.A(men_men_n1838_), .B(men_men_n754_), .C(men_men_n143_), .Y(men_men_n1839_));
  AOI210     u1790(.A0(men_men_n931_), .A1(men_men_n145_), .B0(men_men_n1839_), .Y(men_men_n1840_));
  NA4        u1791(.A(men_men_n1840_), .B(men_men_n1837_), .C(men_men_n1831_), .D(men_men_n1828_), .Y(men24));
  NO2        u1792(.A(men_men_n246_), .B(x1), .Y(men_men_n1842_));
  NA2        u1793(.A(men_men_n344_), .B(men_men_n500_), .Y(men_men_n1843_));
  NAi21      u1794(.An(men_men_n1842_), .B(men_men_n1843_), .Y(men_men_n1844_));
  NO3        u1795(.A(men_men_n550_), .B(men_men_n696_), .C(men_men_n159_), .Y(men_men_n1845_));
  AOI210     u1796(.A0(men_men_n1844_), .A1(men_men_n93_), .B0(men_men_n1845_), .Y(men_men_n1846_));
  NA2        u1797(.A(men_men_n102_), .B(x8), .Y(men_men_n1847_));
  NO3        u1798(.A(men_men_n1081_), .B(men_men_n1360_), .C(men_men_n1062_), .Y(men_men_n1848_));
  AOI210     u1799(.A0(men_men_n996_), .A1(men_men_n56_), .B0(men_men_n1478_), .Y(men_men_n1849_));
  AO220      u1800(.A0(men_men_n1849_), .A1(men_men_n1848_), .B0(men_men_n1289_), .B1(men_men_n332_), .Y(men_men_n1850_));
  NA2        u1801(.A(men_men_n463_), .B(x8), .Y(men_men_n1851_));
  NA2        u1802(.A(men_men_n678_), .B(men_men_n126_), .Y(men_men_n1852_));
  OAI220     u1803(.A0(men_men_n1852_), .A1(men_men_n1463_), .B0(men_men_n1851_), .B1(men_men_n852_), .Y(men_men_n1853_));
  AOI220     u1804(.A0(men_men_n1853_), .A1(men_men_n1718_), .B0(men_men_n1850_), .B1(men_men_n1043_), .Y(men_men_n1854_));
  OAI210     u1805(.A0(men_men_n1847_), .A1(men_men_n1846_), .B0(men_men_n1854_), .Y(men25));
  NA2        u1806(.A(men_men_n333_), .B(men_men_n59_), .Y(men_men_n1856_));
  NO2        u1807(.A(men_men_n1856_), .B(men_men_n324_), .Y(men_men_n1857_));
  OAI210     u1808(.A0(men_men_n1857_), .A1(men_men_n1202_), .B0(men_men_n116_), .Y(men_men_n1858_));
  INV        u1809(.A(men_men_n1298_), .Y(men_men_n1859_));
  NO2        u1810(.A(men_men_n753_), .B(men_men_n55_), .Y(men_men_n1860_));
  AOI220     u1811(.A0(men_men_n1860_), .A1(men_men_n1859_), .B0(men_men_n1617_), .B1(men_men_n1203_), .Y(men_men_n1861_));
  AOI210     u1812(.A0(men_men_n1861_), .A1(men_men_n1858_), .B0(men_men_n691_), .Y(men_men_n1862_));
  NO3        u1813(.A(men_men_n1055_), .B(men_men_n146_), .C(men_men_n78_), .Y(men_men_n1863_));
  OAI210     u1814(.A0(men_men_n202_), .A1(men_men_n280_), .B0(men_men_n334_), .Y(men_men_n1864_));
  OAI210     u1815(.A0(men_men_n1864_), .A1(men_men_n1863_), .B0(men_men_n1201_), .Y(men_men_n1865_));
  NO2        u1816(.A(men_men_n1413_), .B(men_men_n456_), .Y(men_men_n1866_));
  NO3        u1817(.A(men_men_n1866_), .B(men_men_n541_), .C(men_men_n99_), .Y(men_men_n1867_));
  NA2        u1818(.A(men_men_n518_), .B(men_men_n55_), .Y(men_men_n1868_));
  OAI220     u1819(.A0(men_men_n1868_), .A1(men_men_n246_), .B0(men_men_n596_), .B1(men_men_n280_), .Y(men_men_n1869_));
  OAI210     u1820(.A0(men_men_n1869_), .A1(men_men_n1867_), .B0(men_men_n646_), .Y(men_men_n1870_));
  AOI220     u1821(.A0(men_men_n1783_), .A1(men_men_n1155_), .B0(men_men_n1517_), .B1(men_men_n385_), .Y(men_men_n1871_));
  NA3        u1822(.A(men_men_n1871_), .B(men_men_n1870_), .C(men_men_n1865_), .Y(men_men_n1872_));
  AO210      u1823(.A0(men_men_n1872_), .A1(men_men_n108_), .B0(men_men_n1862_), .Y(men26));
  NA2        u1824(.A(men_men_n782_), .B(men_men_n50_), .Y(men_men_n1874_));
  OAI220     u1825(.A0(men_men_n310_), .A1(men_men_n255_), .B0(men_men_n1874_), .B1(x7), .Y(men_men_n1875_));
  AOI220     u1826(.A0(men_men_n1875_), .A1(men_men_n93_), .B0(men_men_n1319_), .B1(men_men_n1161_), .Y(men_men_n1876_));
  NA2        u1827(.A(men_men_n634_), .B(men_men_n588_), .Y(men_men_n1877_));
  OAI210     u1828(.A0(men_men_n642_), .A1(men_men_n634_), .B0(men_men_n757_), .Y(men_men_n1878_));
  AOI210     u1829(.A0(men_men_n1877_), .A1(men_men_n1225_), .B0(men_men_n1878_), .Y(men_men_n1879_));
  NA2        u1830(.A(men_men_n1034_), .B(men_men_n594_), .Y(men_men_n1880_));
  NO2        u1831(.A(men_men_n1880_), .B(men_men_n1272_), .Y(men_men_n1881_));
  AOI210     u1832(.A0(men_men_n1806_), .A1(men_men_n1484_), .B0(men_men_n1881_), .Y(men_men_n1882_));
  NO2        u1833(.A(men_men_n1102_), .B(men_men_n75_), .Y(men_men_n1883_));
  NA2        u1834(.A(men_men_n821_), .B(men_men_n181_), .Y(men_men_n1884_));
  NO2        u1835(.A(men_men_n1884_), .B(men_men_n546_), .Y(men_men_n1885_));
  AOI210     u1836(.A0(men_men_n1883_), .A1(men_men_n595_), .B0(men_men_n1885_), .Y(men_men_n1886_));
  OAI220     u1837(.A0(men_men_n1886_), .A1(men_men_n108_), .B0(men_men_n1882_), .B1(men_men_n53_), .Y(men_men_n1887_));
  NA2        u1838(.A(men_men_n611_), .B(men_men_n518_), .Y(men_men_n1888_));
  NO2        u1839(.A(men_men_n136_), .B(men_men_n133_), .Y(men_men_n1889_));
  NA2        u1840(.A(men_men_n1889_), .B(men_men_n123_), .Y(men_men_n1890_));
  NA2        u1841(.A(men_men_n757_), .B(x3), .Y(men_men_n1891_));
  AOI210     u1842(.A0(men_men_n1890_), .A1(men_men_n1888_), .B0(men_men_n1891_), .Y(men_men_n1892_));
  NO2        u1843(.A(men_men_n1021_), .B(x3), .Y(men_men_n1893_));
  AOI210     u1844(.A0(men_men_n454_), .A1(men_men_n108_), .B0(men_men_n1893_), .Y(men_men_n1894_));
  NA3        u1845(.A(men_men_n579_), .B(men_men_n51_), .C(men_men_n56_), .Y(men_men_n1895_));
  AOI210     u1846(.A0(men_men_n1669_), .A1(men_men_n1074_), .B0(x0), .Y(men_men_n1896_));
  OAI210     u1847(.A0(men_men_n1895_), .A1(men_men_n1894_), .B0(men_men_n1896_), .Y(men_men_n1897_));
  NO4        u1848(.A(men_men_n1897_), .B(men_men_n1892_), .C(men_men_n1887_), .D(men_men_n1879_), .Y(men_men_n1898_));
  AOI210     u1849(.A0(x8), .A1(x6), .B0(x5), .Y(men_men_n1899_));
  AO220      u1850(.A0(men_men_n1899_), .A1(men_men_n148_), .B0(men_men_n602_), .B1(men_men_n143_), .Y(men_men_n1900_));
  NA2        u1851(.A(men_men_n1900_), .B(men_men_n455_), .Y(men_men_n1901_));
  NO2        u1852(.A(men_men_n767_), .B(men_men_n148_), .Y(men_men_n1902_));
  NA3        u1853(.A(men_men_n1902_), .B(men_men_n1691_), .C(men_men_n137_), .Y(men_men_n1903_));
  NO2        u1854(.A(men_men_n406_), .B(men_men_n1399_), .Y(men_men_n1904_));
  NA2        u1855(.A(men_men_n1904_), .B(men_men_n454_), .Y(men_men_n1905_));
  NA3        u1856(.A(men_men_n379_), .B(men_men_n868_), .C(men_men_n259_), .Y(men_men_n1906_));
  NA4        u1857(.A(men_men_n1906_), .B(men_men_n1905_), .C(men_men_n1903_), .D(men_men_n1901_), .Y(men_men_n1907_));
  AOI210     u1858(.A0(men_men_n228_), .A1(x2), .B0(men_men_n501_), .Y(men_men_n1908_));
  NO2        u1859(.A(men_men_n1908_), .B(men_men_n117_), .Y(men_men_n1909_));
  NA3        u1860(.A(men_men_n823_), .B(men_men_n1021_), .C(x7), .Y(men_men_n1910_));
  AOI210     u1861(.A0(men_men_n348_), .A1(men_men_n220_), .B0(men_men_n1910_), .Y(men_men_n1911_));
  OAI220     u1862(.A0(men_men_n910_), .A1(men_men_n310_), .B0(men_men_n654_), .B1(men_men_n696_), .Y(men_men_n1912_));
  NO3        u1863(.A(men_men_n1912_), .B(men_men_n1911_), .C(men_men_n1909_), .Y(men_men_n1913_));
  NA3        u1864(.A(men_men_n678_), .B(men_men_n196_), .C(men_men_n964_), .Y(men_men_n1914_));
  NA2        u1865(.A(men_men_n1914_), .B(men_men_n654_), .Y(men_men_n1915_));
  NA2        u1866(.A(men_men_n143_), .B(men_men_n135_), .Y(men_men_n1916_));
  OAI210     u1867(.A0(men_men_n1916_), .A1(men_men_n1450_), .B0(x0), .Y(men_men_n1917_));
  AOI210     u1868(.A0(men_men_n1915_), .A1(men_men_n1438_), .B0(men_men_n1917_), .Y(men_men_n1918_));
  OAI210     u1869(.A0(men_men_n1913_), .A1(men_men_n53_), .B0(men_men_n1918_), .Y(men_men_n1919_));
  AOI210     u1870(.A0(men_men_n1907_), .A1(x4), .B0(men_men_n1919_), .Y(men_men_n1920_));
  OA220      u1871(.A0(men_men_n1920_), .A1(men_men_n1898_), .B0(men_men_n1876_), .B1(men_men_n109_), .Y(men27));
  NA2        u1872(.A(men_men_n1165_), .B(men_men_n454_), .Y(men_men_n1922_));
  NO2        u1873(.A(men_men_n1922_), .B(men_men_n305_), .Y(men_men_n1923_));
  NA2        u1874(.A(men_men_n927_), .B(men_men_n823_), .Y(men_men_n1924_));
  NA3        u1875(.A(men_men_n829_), .B(men_men_n368_), .C(men_men_n1036_), .Y(men_men_n1925_));
  AOI210     u1876(.A0(men_men_n1925_), .A1(men_men_n1924_), .B0(men_men_n220_), .Y(men_men_n1926_));
  OAI210     u1877(.A0(men_men_n1926_), .A1(men_men_n1923_), .B0(men_men_n712_), .Y(men_men_n1927_));
  XO2        u1878(.A(x8), .B(x4), .Y(men_men_n1928_));
  NO3        u1879(.A(men_men_n1928_), .B(men_men_n454_), .C(men_men_n174_), .Y(men_men_n1929_));
  OA210      u1880(.A0(men_men_n1929_), .A1(men_men_n1273_), .B0(men_men_n283_), .Y(men_men_n1930_));
  NO2        u1881(.A(men_men_n401_), .B(men_men_n168_), .Y(men_men_n1931_));
  OAI210     u1882(.A0(men_men_n1931_), .A1(men_men_n1930_), .B0(men_men_n1139_), .Y(men_men_n1932_));
  AOI210     u1883(.A0(men_men_n642_), .A1(men_men_n56_), .B0(men_men_n1883_), .Y(men_men_n1933_));
  OAI220     u1884(.A0(men_men_n1933_), .A1(men_men_n1272_), .B0(men_men_n1223_), .B1(men_men_n211_), .Y(men_men_n1934_));
  NO2        u1885(.A(men_men_n709_), .B(men_men_n146_), .Y(men_men_n1935_));
  NO2        u1886(.A(men_men_n1207_), .B(men_men_n262_), .Y(men_men_n1936_));
  AOI220     u1887(.A0(men_men_n1936_), .A1(men_men_n1935_), .B0(men_men_n1934_), .B1(men_men_n545_), .Y(men_men_n1937_));
  NA3        u1888(.A(men_men_n1937_), .B(men_men_n1932_), .C(men_men_n1927_), .Y(men28));
  NO3        u1889(.A(men_men_n1928_), .B(men_men_n1408_), .C(men_men_n150_), .Y(men_men_n1939_));
  OAI210     u1890(.A0(men_men_n1939_), .A1(men_men_n1291_), .B0(men_men_n594_), .Y(men_men_n1940_));
  NA3        u1891(.A(men_men_n1203_), .B(men_men_n904_), .C(x7), .Y(men_men_n1941_));
  NA3        u1892(.A(men_men_n503_), .B(men_men_n78_), .C(men_men_n616_), .Y(men_men_n1942_));
  NA3        u1893(.A(men_men_n1942_), .B(men_men_n1941_), .C(men_men_n1940_), .Y(men_men_n1943_));
  NA2        u1894(.A(men_men_n1267_), .B(men_men_n452_), .Y(men_men_n1944_));
  NA3        u1895(.A(men_men_n1944_), .B(men_men_n1427_), .C(men_men_n419_), .Y(men_men_n1945_));
  NO2        u1896(.A(men_men_n313_), .B(x4), .Y(men_men_n1946_));
  AOI220     u1897(.A0(men_men_n1946_), .A1(men_men_n1893_), .B0(men_men_n1140_), .B1(men_men_n686_), .Y(men_men_n1947_));
  NA2        u1898(.A(men_men_n1947_), .B(men_men_n1945_), .Y(men_men_n1948_));
  NO2        u1899(.A(men_men_n1267_), .B(men_men_n1244_), .Y(men_men_n1949_));
  NO4        u1900(.A(x6), .B(men_men_n56_), .C(x2), .D(x0), .Y(men_men_n1950_));
  OAI210     u1901(.A0(men_men_n1950_), .A1(men_men_n1949_), .B0(men_men_n1060_), .Y(men_men_n1951_));
  NA2        u1902(.A(men_men_n1197_), .B(men_men_n108_), .Y(men_men_n1952_));
  NA2        u1903(.A(men_men_n1098_), .B(men_men_n107_), .Y(men_men_n1953_));
  OAI210     u1904(.A0(men_men_n1953_), .A1(men_men_n1952_), .B0(men_men_n1951_), .Y(men_men_n1954_));
  OAI210     u1905(.A0(men_men_n1954_), .A1(men_men_n1948_), .B0(x7), .Y(men_men_n1955_));
  NO2        u1906(.A(men_men_n392_), .B(x7), .Y(men_men_n1956_));
  NO3        u1907(.A(men_men_n406_), .B(men_men_n277_), .C(men_men_n124_), .Y(men_men_n1957_));
  OAI210     u1908(.A0(men_men_n879_), .A1(men_men_n264_), .B0(men_men_n81_), .Y(men_men_n1958_));
  OAI220     u1909(.A0(men_men_n1958_), .A1(men_men_n1957_), .B0(men_men_n1956_), .B1(men_men_n111_), .Y(men_men_n1959_));
  NA2        u1910(.A(men_men_n1815_), .B(men_men_n666_), .Y(men_men_n1960_));
  NO2        u1911(.A(men_men_n1868_), .B(men_men_n77_), .Y(men_men_n1961_));
  AOI220     u1912(.A0(men_men_n1961_), .A1(men_men_n1960_), .B0(men_men_n485_), .B1(men_men_n50_), .Y(men_men_n1962_));
  AOI210     u1913(.A0(men_men_n1962_), .A1(men_men_n1959_), .B0(men_men_n59_), .Y(men_men_n1963_));
  AOI220     u1914(.A0(men_men_n1413_), .A1(men_men_n684_), .B0(men_men_n418_), .B1(men_men_n463_), .Y(men_men_n1964_));
  OAI210     u1915(.A0(men_men_n1964_), .A1(men_men_n146_), .B0(x1), .Y(men_men_n1965_));
  NO2        u1916(.A(men_men_n1965_), .B(men_men_n1963_), .Y(men_men_n1966_));
  AOI210     u1917(.A0(men_men_n1602_), .A1(men_men_n406_), .B0(men_men_n676_), .Y(men_men_n1967_));
  NO2        u1918(.A(men_men_n406_), .B(x5), .Y(men_men_n1968_));
  NO2        u1919(.A(men_men_n1968_), .B(men_men_n232_), .Y(men_men_n1969_));
  NO2        u1920(.A(men_men_n1969_), .B(men_men_n1967_), .Y(men_men_n1970_));
  NOi21      u1921(.An(men_men_n717_), .B(men_men_n1011_), .Y(men_men_n1971_));
  NA3        u1922(.A(men_men_n1971_), .B(men_men_n1098_), .C(men_men_n879_), .Y(men_men_n1972_));
  OAI210     u1923(.A0(men_men_n1380_), .A1(men_men_n1697_), .B0(men_men_n1972_), .Y(men_men_n1973_));
  OAI210     u1924(.A0(men_men_n1973_), .A1(men_men_n1970_), .B0(men_men_n1139_), .Y(men_men_n1974_));
  OAI210     u1925(.A0(men_men_n452_), .A1(men_men_n51_), .B0(men_men_n1030_), .Y(men_men_n1975_));
  AOI220     u1926(.A0(men_men_n1975_), .A1(men_men_n469_), .B0(men_men_n452_), .B1(men_men_n393_), .Y(men_men_n1976_));
  NO2        u1927(.A(men_men_n1976_), .B(men_men_n157_), .Y(men_men_n1977_));
  NA2        u1928(.A(men_men_n166_), .B(men_men_n71_), .Y(men_men_n1978_));
  OAI210     u1929(.A0(men_men_n1880_), .A1(men_men_n1978_), .B0(men_men_n53_), .Y(men_men_n1979_));
  OAI220     u1930(.A0(men_men_n697_), .A1(men_men_n267_), .B0(men_men_n693_), .B1(x6), .Y(men_men_n1980_));
  NO2        u1931(.A(men_men_n308_), .B(x4), .Y(men_men_n1981_));
  AOI220     u1932(.A0(men_men_n1981_), .A1(men_men_n368_), .B0(men_men_n1980_), .B1(x4), .Y(men_men_n1982_));
  NO3        u1933(.A(men_men_n1982_), .B(men_men_n327_), .C(x5), .Y(men_men_n1983_));
  NO2        u1934(.A(men_men_n717_), .B(men_men_n57_), .Y(men_men_n1984_));
  OAI210     u1935(.A0(men_men_n1984_), .A1(men_men_n1935_), .B0(men_men_n454_), .Y(men_men_n1985_));
  AOI220     u1936(.A0(men_men_n674_), .A1(men_men_n743_), .B0(men_men_n501_), .B1(men_men_n242_), .Y(men_men_n1986_));
  AOI210     u1937(.A0(men_men_n1986_), .A1(men_men_n1985_), .B0(men_men_n262_), .Y(men_men_n1987_));
  NO4        u1938(.A(men_men_n1987_), .B(men_men_n1983_), .C(men_men_n1979_), .D(men_men_n1977_), .Y(men_men_n1988_));
  AOI220     u1939(.A0(men_men_n1988_), .A1(men_men_n1974_), .B0(men_men_n1966_), .B1(men_men_n1955_), .Y(men_men_n1989_));
  AOI210     u1940(.A0(men_men_n1943_), .A1(x3), .B0(men_men_n1989_), .Y(men29));
  OAI210     u1941(.A0(men_men_n564_), .A1(men_men_n268_), .B0(men_men_n738_), .Y(men_men_n1991_));
  NA2        u1942(.A(men_men_n759_), .B(men_men_n1060_), .Y(men_men_n1992_));
  AO210      u1943(.A0(men_men_n1178_), .A1(men_men_n1187_), .B0(men_men_n1992_), .Y(men_men_n1993_));
  AOI210     u1944(.A0(men_men_n186_), .A1(men_men_n170_), .B0(men_men_n717_), .Y(men_men_n1994_));
  INV        u1945(.A(men_men_n1994_), .Y(men_men_n1995_));
  NA3        u1946(.A(men_men_n1995_), .B(men_men_n1993_), .C(men_men_n1991_), .Y(men_men_n1996_));
  NO3        u1947(.A(men_men_n676_), .B(men_men_n1161_), .C(men_men_n50_), .Y(men_men_n1997_));
  NO3        u1948(.A(men_men_n1997_), .B(men_men_n1266_), .C(men_men_n564_), .Y(men_men_n1998_));
  NO2        u1949(.A(men_men_n450_), .B(men_men_n58_), .Y(men_men_n1999_));
  AOI220     u1950(.A0(men_men_n1999_), .A1(men_men_n1225_), .B0(men_men_n681_), .B1(men_men_n1398_), .Y(men_men_n2000_));
  OAI210     u1951(.A0(men_men_n1998_), .A1(men_men_n550_), .B0(men_men_n2000_), .Y(men_men_n2001_));
  AOI210     u1952(.A0(men_men_n1996_), .A1(x6), .B0(men_men_n2001_), .Y(men_men_n2002_));
  OAI210     u1953(.A0(x8), .A1(x4), .B0(x5), .Y(men_men_n2003_));
  NA2        u1954(.A(men_men_n2003_), .B(men_men_n112_), .Y(men_men_n2004_));
  NA2        u1955(.A(men_men_n308_), .B(men_men_n150_), .Y(men_men_n2005_));
  NA4        u1956(.A(men_men_n2005_), .B(men_men_n2004_), .C(men_men_n675_), .D(men_men_n64_), .Y(men_men_n2006_));
  AOI210     u1957(.A0(men_men_n1338_), .A1(men_men_n277_), .B0(men_men_n1749_), .Y(men_men_n2007_));
  AOI210     u1958(.A0(men_men_n2007_), .A1(men_men_n2006_), .B0(men_men_n897_), .Y(men_men_n2008_));
  NA4        u1959(.A(men_men_n676_), .B(men_men_n313_), .C(men_men_n186_), .D(men_men_n170_), .Y(men_men_n2009_));
  NA3        u1960(.A(men_men_n640_), .B(men_men_n301_), .C(men_men_n811_), .Y(men_men_n2010_));
  AOI210     u1961(.A0(men_men_n2010_), .A1(men_men_n2009_), .B0(men_men_n1225_), .Y(men_men_n2011_));
  OAI210     u1962(.A0(men_men_n904_), .A1(x8), .B0(x7), .Y(men_men_n2012_));
  NO2        u1963(.A(men_men_n2012_), .B(men_men_n129_), .Y(men_men_n2013_));
  OA210      u1964(.A0(men_men_n879_), .A1(men_men_n280_), .B0(men_men_n2003_), .Y(men_men_n2014_));
  OAI220     u1965(.A0(men_men_n2014_), .A1(men_men_n596_), .B0(men_men_n1525_), .B1(men_men_n401_), .Y(men_men_n2015_));
  NO4        u1966(.A(men_men_n2015_), .B(men_men_n2013_), .C(men_men_n2011_), .D(men_men_n2008_), .Y(men_men_n2016_));
  OAI210     u1967(.A0(men_men_n2002_), .A1(x2), .B0(men_men_n2016_), .Y(men_men_n2017_));
  NA3        u1968(.A(x6), .B(men_men_n50_), .C(x2), .Y(men_men_n2018_));
  OAI210     u1969(.A0(men_men_n1244_), .A1(men_men_n358_), .B0(men_men_n2018_), .Y(men_men_n2019_));
  NO3        u1970(.A(men_men_n452_), .B(x3), .C(x0), .Y(men_men_n2020_));
  AO220      u1971(.A0(men_men_n2020_), .A1(x5), .B0(men_men_n1950_), .B1(men_men_n81_), .Y(men_men_n2021_));
  AOI210     u1972(.A0(men_men_n2019_), .A1(men_men_n348_), .B0(men_men_n2021_), .Y(men_men_n2022_));
  NO3        u1973(.A(men_men_n710_), .B(men_men_n369_), .C(men_men_n144_), .Y(men_men_n2023_));
  AOI210     u1974(.A0(men_men_n737_), .A1(men_men_n623_), .B0(men_men_n2023_), .Y(men_men_n2024_));
  OAI210     u1975(.A0(men_men_n2022_), .A1(x7), .B0(men_men_n2024_), .Y(men_men_n2025_));
  AOI210     u1976(.A0(men_men_n1108_), .A1(men_men_n406_), .B0(men_men_n1426_), .Y(men_men_n2026_));
  NO2        u1977(.A(men_men_n150_), .B(x2), .Y(men_men_n2027_));
  OA210      u1978(.A0(men_men_n2027_), .A1(men_men_n638_), .B0(men_men_n676_), .Y(men_men_n2028_));
  OAI210     u1979(.A0(men_men_n2028_), .A1(men_men_n2026_), .B0(men_men_n68_), .Y(men_men_n2029_));
  NO2        u1980(.A(men_men_n202_), .B(men_men_n85_), .Y(men_men_n2030_));
  OAI210     u1981(.A0(men_men_n2030_), .A1(men_men_n797_), .B0(men_men_n1117_), .Y(men_men_n2031_));
  NA3        u1982(.A(men_men_n1968_), .B(men_men_n235_), .C(men_men_n83_), .Y(men_men_n2032_));
  NA3        u1983(.A(men_men_n2032_), .B(men_men_n2031_), .C(men_men_n2029_), .Y(men_men_n2033_));
  AOI210     u1984(.A0(men_men_n2025_), .A1(x8), .B0(men_men_n2033_), .Y(men_men_n2034_));
  OAI210     u1985(.A0(men_men_n450_), .A1(men_men_n251_), .B0(men_men_n974_), .Y(men_men_n2035_));
  OAI210     u1986(.A0(men_men_n2035_), .A1(men_men_n1140_), .B0(men_men_n686_), .Y(men_men_n2036_));
  NO3        u1987(.A(men_men_n1034_), .B(men_men_n359_), .C(men_men_n151_), .Y(men_men_n2037_));
  NA3        u1988(.A(men_men_n2037_), .B(men_men_n1318_), .C(men_men_n50_), .Y(men_men_n2038_));
  NO2        u1989(.A(men_men_n137_), .B(men_men_n93_), .Y(men_men_n2039_));
  AOI220     u1990(.A0(men_men_n2039_), .A1(men_men_n597_), .B0(men_men_n1949_), .B1(men_men_n365_), .Y(men_men_n2040_));
  NOi31      u1991(.An(men_men_n1141_), .B(men_men_n1899_), .C(men_men_n633_), .Y(men_men_n2041_));
  NA2        u1992(.A(men_men_n176_), .B(x4), .Y(men_men_n2042_));
  NO3        u1993(.A(men_men_n1498_), .B(men_men_n246_), .C(men_men_n71_), .Y(men_men_n2043_));
  AOI210     u1994(.A0(men_men_n2043_), .A1(men_men_n2042_), .B0(men_men_n2041_), .Y(men_men_n2044_));
  NA4        u1995(.A(men_men_n2044_), .B(men_men_n2040_), .C(men_men_n2038_), .D(men_men_n2036_), .Y(men_men_n2045_));
  NO4        u1996(.A(men_men_n1244_), .B(men_men_n174_), .C(men_men_n55_), .D(men_men_n71_), .Y(men_men_n2046_));
  NO4        u1997(.A(men_men_n1218_), .B(men_men_n510_), .C(men_men_n1398_), .D(men_men_n108_), .Y(men_men_n2047_));
  OAI210     u1998(.A0(men_men_n2047_), .A1(men_men_n2046_), .B0(men_men_n110_), .Y(men_men_n2048_));
  AOI210     u1999(.A0(men_men_n312_), .A1(x4), .B0(men_men_n196_), .Y(men_men_n2049_));
  OAI210     u2000(.A0(men_men_n2049_), .A1(men_men_n1999_), .B0(men_men_n732_), .Y(men_men_n2050_));
  OR3        u2001(.A(men_men_n1770_), .B(men_men_n1453_), .C(men_men_n1100_), .Y(men_men_n2051_));
  NA2        u2002(.A(men_men_n1950_), .B(men_men_n818_), .Y(men_men_n2052_));
  OA220      u2003(.A0(men_men_n2052_), .A1(men_men_n251_), .B0(men_men_n589_), .B1(men_men_n1813_), .Y(men_men_n2053_));
  NA4        u2004(.A(men_men_n2053_), .B(men_men_n2051_), .C(men_men_n2050_), .D(men_men_n2048_), .Y(men_men_n2054_));
  AOI210     u2005(.A0(men_men_n2045_), .A1(men_men_n297_), .B0(men_men_n2054_), .Y(men_men_n2055_));
  OAI210     u2006(.A0(men_men_n2034_), .A1(x1), .B0(men_men_n2055_), .Y(men_men_n2056_));
  AO210      u2007(.A0(men_men_n2017_), .A1(x1), .B0(men_men_n2056_), .Y(men30));
  NO3        u2008(.A(men_men_n1797_), .B(men_men_n585_), .C(men_men_n99_), .Y(men_men_n2058_));
  NO3        u2009(.A(men_men_n1159_), .B(men_men_n140_), .C(men_men_n389_), .Y(men_men_n2059_));
  AOI210     u2010(.A0(men_men_n732_), .A1(men_men_n259_), .B0(men_men_n2059_), .Y(men_men_n2060_));
  AOI210     u2011(.A0(men_men_n2060_), .A1(men_men_n2058_), .B0(men_men_n56_), .Y(men_men_n2061_));
  NA2        u2012(.A(men_men_n823_), .B(men_men_n346_), .Y(men_men_n2062_));
  NA2        u2013(.A(men_men_n2062_), .B(men_men_n1381_), .Y(men_men_n2063_));
  OAI210     u2014(.A0(men_men_n2063_), .A1(men_men_n2061_), .B0(men_men_n110_), .Y(men_men_n2064_));
  OAI210     u2015(.A0(men_men_n1011_), .A1(men_men_n579_), .B0(men_men_n686_), .Y(men_men_n2065_));
  AOI220     u2016(.A0(men_men_n455_), .A1(men_men_n951_), .B0(men_men_n332_), .B1(men_men_n463_), .Y(men_men_n2066_));
  AOI210     u2017(.A0(men_men_n2066_), .A1(men_men_n2065_), .B0(men_men_n262_), .Y(men_men_n2067_));
  NO3        u2018(.A(men_men_n286_), .B(men_men_n125_), .C(x0), .Y(men_men_n2068_));
  AOI210     u2019(.A0(men_men_n512_), .A1(x6), .B0(men_men_n2068_), .Y(men_men_n2069_));
  AOI220     u2020(.A0(men_men_n1155_), .A1(men_men_n430_), .B0(men_men_n771_), .B1(men_men_n92_), .Y(men_men_n2070_));
  OAI220     u2021(.A0(men_men_n2070_), .A1(men_men_n251_), .B0(men_men_n2069_), .B1(men_men_n54_), .Y(men_men_n2071_));
  NA3        u2022(.A(men_men_n328_), .B(men_men_n167_), .C(men_men_n71_), .Y(men_men_n2072_));
  AO210      u2023(.A0(men_men_n578_), .A1(men_men_n526_), .B0(x5), .Y(men_men_n2073_));
  AOI210     u2024(.A0(men_men_n2072_), .A1(men_men_n729_), .B0(men_men_n2073_), .Y(men_men_n2074_));
  AOI210     u2025(.A0(men_men_n1623_), .A1(men_men_n50_), .B0(men_men_n463_), .Y(men_men_n2075_));
  NA2        u2026(.A(men_men_n201_), .B(x2), .Y(men_men_n2076_));
  OA220      u2027(.A0(men_men_n2076_), .A1(men_men_n2075_), .B0(men_men_n281_), .B1(x6), .Y(men_men_n2077_));
  OAI210     u2028(.A0(x7), .A1(x6), .B0(x1), .Y(men_men_n2078_));
  NA3        u2029(.A(men_men_n57_), .B(x4), .C(men_men_n59_), .Y(men_men_n2079_));
  AOI220     u2030(.A0(men_men_n2079_), .A1(men_men_n1388_), .B0(men_men_n2078_), .B1(men_men_n1838_), .Y(men_men_n2080_));
  NO3        u2031(.A(men_men_n1384_), .B(men_men_n348_), .C(men_men_n1036_), .Y(men_men_n2081_));
  NO2        u2032(.A(men_men_n524_), .B(men_men_n872_), .Y(men_men_n2082_));
  NOi21      u2033(.An(men_men_n2082_), .B(men_men_n857_), .Y(men_men_n2083_));
  NO3        u2034(.A(men_men_n1318_), .B(men_men_n237_), .C(men_men_n658_), .Y(men_men_n2084_));
  NO4        u2035(.A(men_men_n2084_), .B(men_men_n2083_), .C(men_men_n2081_), .D(men_men_n2080_), .Y(men_men_n2085_));
  OAI210     u2036(.A0(men_men_n2077_), .A1(men_men_n766_), .B0(men_men_n2085_), .Y(men_men_n2086_));
  NO4        u2037(.A(men_men_n2086_), .B(men_men_n2074_), .C(men_men_n2071_), .D(men_men_n2067_), .Y(men_men_n2087_));
  AOI210     u2038(.A0(men_men_n2087_), .A1(men_men_n2064_), .B0(x8), .Y(men_men_n2088_));
  NO3        u2039(.A(men_men_n499_), .B(men_men_n794_), .C(men_men_n53_), .Y(men_men_n2089_));
  OAI220     u2040(.A0(men_men_n1813_), .A1(men_men_n348_), .B0(men_men_n491_), .B1(men_men_n593_), .Y(men_men_n2090_));
  OAI210     u2041(.A0(men_men_n2090_), .A1(men_men_n2089_), .B0(x6), .Y(men_men_n2091_));
  OAI210     u2042(.A0(men_men_n1051_), .A1(men_men_n545_), .B0(men_men_n823_), .Y(men_men_n2092_));
  OAI210     u2043(.A0(men_men_n1759_), .A1(men_men_n335_), .B0(men_men_n128_), .Y(men_men_n2093_));
  AOI210     u2044(.A0(men_men_n384_), .A1(men_men_n234_), .B0(men_men_n72_), .Y(men_men_n2094_));
  AOI210     u2045(.A0(men_men_n1011_), .A1(men_men_n757_), .B0(men_men_n2094_), .Y(men_men_n2095_));
  NA4        u2046(.A(men_men_n2095_), .B(men_men_n2093_), .C(men_men_n2092_), .D(men_men_n2091_), .Y(men_men_n2096_));
  NA2        u2047(.A(men_men_n1105_), .B(men_men_n59_), .Y(men_men_n2097_));
  AOI210     u2048(.A0(men_men_n932_), .A1(men_men_n500_), .B0(men_men_n692_), .Y(men_men_n2098_));
  OAI220     u2049(.A0(men_men_n2098_), .A1(men_men_n312_), .B0(men_men_n2097_), .B1(men_men_n490_), .Y(men_men_n2099_));
  AOI210     u2050(.A0(men_men_n2096_), .A1(x8), .B0(men_men_n2099_), .Y(men_men_n2100_));
  NO2        u2051(.A(men_men_n2100_), .B(men_men_n57_), .Y(men_men_n2101_));
  NA2        u2052(.A(men_men_n441_), .B(men_men_n857_), .Y(men_men_n2102_));
  NO2        u2053(.A(men_men_n931_), .B(men_men_n672_), .Y(men_men_n2103_));
  AOI210     u2054(.A0(men_men_n2103_), .A1(men_men_n2102_), .B0(men_men_n452_), .Y(men_men_n2104_));
  NO3        u2055(.A(men_men_n646_), .B(men_men_n415_), .C(men_men_n1159_), .Y(men_men_n2105_));
  NO3        u2056(.A(men_men_n2105_), .B(men_men_n1272_), .C(men_men_n1398_), .Y(men_men_n2106_));
  AOI210     u2057(.A0(men_men_n309_), .A1(x1), .B0(men_men_n151_), .Y(men_men_n2107_));
  NO2        u2058(.A(men_men_n315_), .B(x5), .Y(men_men_n2108_));
  NO2        u2059(.A(men_men_n2108_), .B(men_men_n865_), .Y(men_men_n2109_));
  OAI220     u2060(.A0(men_men_n2109_), .A1(men_men_n1071_), .B0(men_men_n2107_), .B1(men_men_n211_), .Y(men_men_n2110_));
  NO3        u2061(.A(men_men_n2110_), .B(men_men_n2106_), .C(men_men_n2104_), .Y(men_men_n2111_));
  NA2        u2062(.A(men_men_n972_), .B(men_men_n82_), .Y(men_men_n2112_));
  AO210      u2063(.A0(men_men_n2112_), .A1(men_men_n1624_), .B0(x3), .Y(men_men_n2113_));
  NO2        u2064(.A(men_men_n223_), .B(men_men_n56_), .Y(men_men_n2114_));
  OAI220     u2065(.A0(men_men_n384_), .A1(men_men_n1272_), .B0(men_men_n359_), .B1(men_men_n237_), .Y(men_men_n2115_));
  AOI220     u2066(.A0(men_men_n2115_), .A1(x2), .B0(men_men_n2114_), .B1(men_men_n1639_), .Y(men_men_n2116_));
  AOI210     u2067(.A0(men_men_n2116_), .A1(men_men_n2113_), .B0(men_men_n267_), .Y(men_men_n2117_));
  NO3        u2068(.A(men_men_n828_), .B(men_men_n711_), .C(men_men_n170_), .Y(men_men_n2118_));
  OAI210     u2069(.A0(men_men_n2118_), .A1(men_men_n2696_), .B0(men_men_n158_), .Y(men_men_n2119_));
  NA3        u2070(.A(x5), .B(x4), .C(men_men_n59_), .Y(men_men_n2120_));
  AOI210     u2071(.A0(men_men_n2120_), .A1(men_men_n1326_), .B0(men_men_n546_), .Y(men_men_n2121_));
  AOI210     u2072(.A0(men_men_n1346_), .A1(x2), .B0(men_men_n2121_), .Y(men_men_n2122_));
  AOI210     u2073(.A0(men_men_n2122_), .A1(men_men_n2119_), .B0(men_men_n50_), .Y(men_men_n2123_));
  NA3        u2074(.A(men_men_n1495_), .B(men_men_n1150_), .C(men_men_n483_), .Y(men_men_n2124_));
  AOI210     u2075(.A0(men_men_n2124_), .A1(men_men_n2112_), .B0(men_men_n619_), .Y(men_men_n2125_));
  AOI210     u2076(.A0(men_men_n1036_), .A1(x1), .B0(men_men_n1338_), .Y(men_men_n2126_));
  OAI220     u2077(.A0(men_men_n313_), .A1(x4), .B0(men_men_n51_), .B1(x6), .Y(men_men_n2127_));
  NO2        u2078(.A(men_men_n123_), .B(men_men_n112_), .Y(men_men_n2128_));
  AOI220     u2079(.A0(men_men_n2128_), .A1(men_men_n2127_), .B0(men_men_n1180_), .B1(men_men_n633_), .Y(men_men_n2129_));
  OAI210     u2080(.A0(men_men_n2126_), .A1(men_men_n494_), .B0(men_men_n2129_), .Y(men_men_n2130_));
  NO4        u2081(.A(men_men_n2130_), .B(men_men_n2125_), .C(men_men_n2123_), .D(men_men_n2117_), .Y(men_men_n2131_));
  OAI210     u2082(.A0(men_men_n2111_), .A1(men_men_n137_), .B0(men_men_n2131_), .Y(men_men_n2132_));
  NO3        u2083(.A(men_men_n2132_), .B(men_men_n2101_), .C(men_men_n2088_), .Y(men31));
  NA2        u2084(.A(men_men_n996_), .B(men_men_n360_), .Y(men_men_n2134_));
  NO2        u2085(.A(men_men_n456_), .B(men_men_n686_), .Y(men_men_n2135_));
  AOI210     u2086(.A0(men_men_n2135_), .A1(men_men_n2134_), .B0(men_men_n58_), .Y(men_men_n2136_));
  NO2        u2087(.A(men_men_n796_), .B(men_men_n56_), .Y(men_men_n2137_));
  AOI220     u2088(.A0(men_men_n2137_), .A1(x2), .B0(men_men_n91_), .B1(x0), .Y(men_men_n2138_));
  NA3        u2089(.A(men_men_n2138_), .B(men_men_n2052_), .C(men_men_n1877_), .Y(men_men_n2139_));
  OAI210     u2090(.A0(men_men_n2139_), .A1(men_men_n2136_), .B0(men_men_n53_), .Y(men_men_n2140_));
  NO2        u2091(.A(men_men_n438_), .B(men_men_n686_), .Y(men_men_n2141_));
  NO3        u2092(.A(men_men_n1981_), .B(men_men_n1950_), .C(men_men_n898_), .Y(men_men_n2142_));
  OA220      u2093(.A0(men_men_n2142_), .A1(men_men_n483_), .B0(men_men_n2141_), .B1(men_men_n1488_), .Y(men_men_n2143_));
  AOI210     u2094(.A0(men_men_n2143_), .A1(men_men_n2140_), .B0(men_men_n108_), .Y(men_men_n2144_));
  NO2        u2095(.A(men_men_n506_), .B(men_men_n75_), .Y(men_men_n2145_));
  NA2        u2096(.A(men_men_n452_), .B(men_men_n57_), .Y(men_men_n2146_));
  AOI210     u2097(.A0(men_men_n312_), .A1(men_men_n86_), .B0(men_men_n2146_), .Y(men_men_n2147_));
  OAI210     u2098(.A0(men_men_n2147_), .A1(men_men_n2145_), .B0(men_men_n782_), .Y(men_men_n2148_));
  NO4        u2099(.A(men_men_n1176_), .B(men_men_n369_), .C(men_men_n1623_), .D(men_men_n67_), .Y(men_men_n2149_));
  AOI210     u2100(.A0(men_men_n1664_), .A1(men_men_n1373_), .B0(men_men_n450_), .Y(men_men_n2150_));
  NO2        u2101(.A(men_men_n1327_), .B(men_men_n965_), .Y(men_men_n2151_));
  NO3        u2102(.A(men_men_n2151_), .B(men_men_n2150_), .C(men_men_n2149_), .Y(men_men_n2152_));
  AOI210     u2103(.A0(men_men_n2152_), .A1(men_men_n2148_), .B0(x5), .Y(men_men_n2153_));
  AOI220     u2104(.A0(men_men_n454_), .A1(men_men_n633_), .B0(men_men_n579_), .B1(men_men_n63_), .Y(men_men_n2154_));
  AOI210     u2105(.A0(men_men_n2154_), .A1(men_men_n589_), .B0(men_men_n1244_), .Y(men_men_n2155_));
  AOI220     u2106(.A0(men_men_n973_), .A1(men_men_n743_), .B0(men_men_n1159_), .B1(men_men_n122_), .Y(men_men_n2156_));
  OAI220     u2107(.A0(men_men_n2156_), .A1(men_men_n392_), .B0(men_men_n490_), .B1(men_men_n783_), .Y(men_men_n2157_));
  NO4        u2108(.A(men_men_n2157_), .B(men_men_n2155_), .C(men_men_n2153_), .D(men_men_n2144_), .Y(men_men_n2158_));
  NA2        u2109(.A(men_men_n500_), .B(men_men_n59_), .Y(men_men_n2159_));
  AOI210     u2110(.A0(men_men_n550_), .A1(men_men_n2159_), .B0(men_men_n143_), .Y(men_men_n2160_));
  OAI210     u2111(.A0(men_men_n104_), .A1(men_men_n280_), .B0(men_men_n2097_), .Y(men_men_n2161_));
  OAI210     u2112(.A0(men_men_n2161_), .A1(men_men_n2160_), .B0(x7), .Y(men_men_n2162_));
  NO3        u2113(.A(men_men_n384_), .B(men_men_n55_), .C(x7), .Y(men_men_n2163_));
  OA210      u2114(.A0(men_men_n2163_), .A1(men_men_n1337_), .B0(men_men_n101_), .Y(men_men_n2164_));
  NA2        u2115(.A(men_men_n1102_), .B(men_men_n92_), .Y(men_men_n2165_));
  AOI210     u2116(.A0(men_men_n910_), .A1(men_men_n112_), .B0(men_men_n2165_), .Y(men_men_n2166_));
  NA2        u2117(.A(men_men_n1570_), .B(x6), .Y(men_men_n2167_));
  AOI210     u2118(.A0(men_men_n2167_), .A1(men_men_n296_), .B0(men_men_n108_), .Y(men_men_n2168_));
  NA2        u2119(.A(men_men_n1203_), .B(men_men_n323_), .Y(men_men_n2169_));
  AOI210     u2120(.A0(men_men_n2169_), .A1(men_men_n654_), .B0(men_men_n53_), .Y(men_men_n2170_));
  NO4        u2121(.A(men_men_n2170_), .B(men_men_n2168_), .C(men_men_n2166_), .D(men_men_n2164_), .Y(men_men_n2171_));
  AOI210     u2122(.A0(men_men_n2171_), .A1(men_men_n2162_), .B0(men_men_n696_), .Y(men_men_n2172_));
  NOi21      u2123(.An(men_men_n1787_), .B(men_men_n1075_), .Y(men_men_n2173_));
  OAI220     u2124(.A0(men_men_n2173_), .A1(men_men_n1952_), .B0(men_men_n933_), .B1(men_men_n2159_), .Y(men_men_n2174_));
  NA2        u2125(.A(men_men_n2174_), .B(x3), .Y(men_men_n2175_));
  AOI220     u2126(.A0(men_men_n1408_), .A1(x8), .B0(men_men_n60_), .B1(x1), .Y(men_men_n2176_));
  NO3        u2127(.A(men_men_n2176_), .B(men_men_n1129_), .C(x6), .Y(men_men_n2177_));
  NA2        u2128(.A(men_men_n623_), .B(men_men_n415_), .Y(men_men_n2178_));
  NA2        u2129(.A(men_men_n118_), .B(men_men_n537_), .Y(men_men_n2179_));
  OAI220     u2130(.A0(men_men_n2179_), .A1(men_men_n1952_), .B0(men_men_n2178_), .B1(x4), .Y(men_men_n2180_));
  NO2        u2131(.A(men_men_n2180_), .B(men_men_n2177_), .Y(men_men_n2181_));
  AOI210     u2132(.A0(men_men_n2181_), .A1(men_men_n2175_), .B0(men_men_n189_), .Y(men_men_n2182_));
  NO4        u2133(.A(men_men_n624_), .B(men_men_n597_), .C(men_men_n712_), .D(men_men_n711_), .Y(men_men_n2183_));
  OAI210     u2134(.A0(men_men_n2183_), .A1(men_men_n1093_), .B0(x3), .Y(men_men_n2184_));
  NO4        u2135(.A(men_men_n814_), .B(men_men_n1244_), .C(men_men_n782_), .D(x5), .Y(men_men_n2185_));
  NO3        u2136(.A(x6), .B(men_men_n56_), .C(x1), .Y(men_men_n2186_));
  NA2        u2137(.A(men_men_n2186_), .B(men_men_n292_), .Y(men_men_n2187_));
  OAI210     u2138(.A0(men_men_n1922_), .A1(men_men_n384_), .B0(men_men_n2187_), .Y(men_men_n2188_));
  NA4        u2139(.A(men_men_n646_), .B(men_men_n182_), .C(x6), .D(men_men_n108_), .Y(men_men_n2189_));
  NO2        u2140(.A(men_men_n866_), .B(men_men_n255_), .Y(men_men_n2190_));
  NOi41      u2141(.An(men_men_n2189_), .B(men_men_n2190_), .C(men_men_n2188_), .D(men_men_n2185_), .Y(men_men_n2191_));
  AOI210     u2142(.A0(men_men_n2191_), .A1(men_men_n2184_), .B0(men_men_n541_), .Y(men_men_n2192_));
  OAI210     u2143(.A0(men_men_n623_), .A1(men_men_n477_), .B0(men_men_n951_), .Y(men_men_n2193_));
  NO3        u2144(.A(men_men_n379_), .B(men_men_n77_), .C(men_men_n53_), .Y(men_men_n2194_));
  NO3        u2145(.A(men_men_n469_), .B(men_men_n354_), .C(men_men_n50_), .Y(men_men_n2195_));
  OAI210     u2146(.A0(men_men_n2195_), .A1(men_men_n2194_), .B0(men_men_n1177_), .Y(men_men_n2196_));
  AOI210     u2147(.A0(men_men_n2196_), .A1(men_men_n2193_), .B0(men_men_n399_), .Y(men_men_n2197_));
  NO2        u2148(.A(men_men_n220_), .B(men_men_n546_), .Y(men_men_n2198_));
  OAI210     u2149(.A0(men_men_n140_), .A1(x2), .B0(men_men_n2198_), .Y(men_men_n2199_));
  NA3        u2150(.A(men_men_n415_), .B(men_men_n333_), .C(men_men_n77_), .Y(men_men_n2200_));
  OA210      u2151(.A0(men_men_n250_), .A1(men_men_n233_), .B0(men_men_n2200_), .Y(men_men_n2201_));
  AOI210     u2152(.A0(men_men_n2201_), .A1(men_men_n2199_), .B0(men_men_n64_), .Y(men_men_n2202_));
  NA2        u2153(.A(men_men_n123_), .B(men_men_n57_), .Y(men_men_n2203_));
  AOI220     u2154(.A0(men_men_n1602_), .A1(men_men_n917_), .B0(men_men_n279_), .B1(x4), .Y(men_men_n2204_));
  AOI220     u2155(.A0(men_men_n1656_), .A1(men_men_n625_), .B0(men_men_n730_), .B1(men_men_n782_), .Y(men_men_n2205_));
  OAI220     u2156(.A0(men_men_n2205_), .A1(men_men_n2203_), .B0(men_men_n2204_), .B1(men_men_n194_), .Y(men_men_n2206_));
  OR3        u2157(.A(men_men_n2206_), .B(men_men_n2202_), .C(men_men_n2197_), .Y(men_men_n2207_));
  NO4        u2158(.A(men_men_n2207_), .B(men_men_n2192_), .C(men_men_n2182_), .D(men_men_n2172_), .Y(men_men_n2208_));
  OAI210     u2159(.A0(men_men_n2158_), .A1(x3), .B0(men_men_n2208_), .Y(men32));
  OAI210     u2160(.A0(men_men_n572_), .A1(men_men_n53_), .B0(men_men_n420_), .Y(men_men_n2210_));
  NA2        u2161(.A(men_men_n521_), .B(x2), .Y(men_men_n2211_));
  AOI210     u2162(.A0(men_men_n2211_), .A1(men_men_n2210_), .B0(men_men_n57_), .Y(men_men_n2212_));
  OAI210     u2163(.A0(men_men_n2212_), .A1(men_men_n797_), .B0(men_men_n56_), .Y(men_men_n2213_));
  OAI210     u2164(.A0(men_men_n1728_), .A1(men_men_n1471_), .B0(men_men_n1497_), .Y(men_men_n2214_));
  AOI210     u2165(.A0(men_men_n2137_), .A1(men_men_n283_), .B0(men_men_n2214_), .Y(men_men_n2215_));
  AOI210     u2166(.A0(men_men_n2215_), .A1(men_men_n2213_), .B0(men_men_n50_), .Y(men_men_n2216_));
  NA3        u2167(.A(men_men_n1571_), .B(men_men_n812_), .C(men_men_n295_), .Y(men_men_n2217_));
  NA2        u2168(.A(men_men_n754_), .B(men_men_n554_), .Y(men_men_n2218_));
  OAI220     u2169(.A0(men_men_n1070_), .A1(men_men_n235_), .B0(men_men_n693_), .B1(men_men_n211_), .Y(men_men_n2219_));
  NO3        u2170(.A(men_men_n380_), .B(men_men_n582_), .C(men_men_n818_), .Y(men_men_n2220_));
  NO3        u2171(.A(men_men_n1384_), .B(men_men_n593_), .C(men_men_n277_), .Y(men_men_n2221_));
  NO4        u2172(.A(men_men_n2221_), .B(men_men_n2220_), .C(men_men_n2219_), .D(men_men_n2218_), .Y(men_men_n2222_));
  AOI210     u2173(.A0(men_men_n2222_), .A1(men_men_n2217_), .B0(men_men_n144_), .Y(men_men_n2223_));
  OAI220     u2174(.A0(men_men_n408_), .A1(x7), .B0(men_men_n308_), .B1(men_men_n301_), .Y(men_men_n2224_));
  NA2        u2175(.A(men_men_n2224_), .B(men_men_n972_), .Y(men_men_n2225_));
  NO2        u2176(.A(men_men_n559_), .B(men_men_n872_), .Y(men_men_n2226_));
  AOI220     u2177(.A0(men_men_n2226_), .A1(men_men_n1902_), .B0(men_men_n538_), .B1(men_men_n133_), .Y(men_men_n2227_));
  AOI210     u2178(.A0(men_men_n2227_), .A1(men_men_n2225_), .B0(men_men_n110_), .Y(men_men_n2228_));
  NA3        u2179(.A(men_men_n1337_), .B(men_men_n1161_), .C(men_men_n117_), .Y(men_men_n2229_));
  AOI220     u2180(.A0(men_men_n1374_), .A1(men_men_n712_), .B0(men_men_n1258_), .B1(men_men_n1058_), .Y(men_men_n2230_));
  AOI210     u2181(.A0(men_men_n2230_), .A1(men_men_n2229_), .B0(men_men_n56_), .Y(men_men_n2231_));
  NA2        u2182(.A(men_men_n972_), .B(men_men_n57_), .Y(men_men_n2232_));
  NOi21      u2183(.An(men_men_n2232_), .B(men_men_n133_), .Y(men_men_n2233_));
  NA2        u2184(.A(men_men_n1026_), .B(men_men_n255_), .Y(men_men_n2234_));
  NO3        u2185(.A(men_men_n2234_), .B(men_men_n2233_), .C(men_men_n59_), .Y(men_men_n2235_));
  OR4        u2186(.A(men_men_n2235_), .B(men_men_n2231_), .C(men_men_n2228_), .D(men_men_n2223_), .Y(men_men_n2236_));
  OAI210     u2187(.A0(men_men_n2236_), .A1(men_men_n2216_), .B0(men_men_n108_), .Y(men_men_n2237_));
  NO3        u2188(.A(men_men_n1244_), .B(men_men_n148_), .C(men_men_n126_), .Y(men_men_n2238_));
  NO2        u2189(.A(men_men_n387_), .B(men_men_n55_), .Y(men_men_n2239_));
  NA2        u2190(.A(men_men_n2239_), .B(men_men_n116_), .Y(men_men_n2240_));
  OAI210     u2191(.A0(men_men_n642_), .A1(men_men_n599_), .B0(men_men_n823_), .Y(men_men_n2241_));
  NA2        u2192(.A(men_men_n2241_), .B(men_men_n2240_), .Y(men_men_n2242_));
  OAI210     u2193(.A0(men_men_n2242_), .A1(men_men_n2238_), .B0(x3), .Y(men_men_n2243_));
  OAI210     u2194(.A0(men_men_n904_), .A1(men_men_n277_), .B0(men_men_n50_), .Y(men_men_n2244_));
  AOI210     u2195(.A0(men_men_n62_), .A1(men_men_n110_), .B0(men_men_n2244_), .Y(men_men_n2245_));
  OAI210     u2196(.A0(men_men_n2245_), .A1(men_men_n1883_), .B0(men_men_n711_), .Y(men_men_n2246_));
  NO3        u2197(.A(men_men_n310_), .B(men_men_n176_), .C(men_men_n124_), .Y(men_men_n2247_));
  NO3        u2198(.A(men_men_n812_), .B(men_men_n367_), .C(men_men_n144_), .Y(men_men_n2248_));
  OAI210     u2199(.A0(men_men_n2248_), .A1(men_men_n2247_), .B0(men_men_n59_), .Y(men_men_n2249_));
  NA2        u2200(.A(men_men_n1165_), .B(men_men_n71_), .Y(men_men_n2250_));
  NO2        u2201(.A(men_men_n1956_), .B(men_men_n599_), .Y(men_men_n2251_));
  AOI210     u2202(.A0(men_men_n2251_), .A1(men_men_n1884_), .B0(men_men_n2250_), .Y(men_men_n2252_));
  NO2        u2203(.A(men_men_n280_), .B(men_men_n57_), .Y(men_men_n2253_));
  NO2        u2204(.A(men_men_n2253_), .B(men_men_n1018_), .Y(men_men_n2254_));
  NOi31      u2205(.An(men_men_n732_), .B(men_men_n2254_), .C(men_men_n286_), .Y(men_men_n2255_));
  NO3        u2206(.A(men_men_n1329_), .B(men_men_n220_), .C(men_men_n262_), .Y(men_men_n2256_));
  NO4        u2207(.A(men_men_n2256_), .B(men_men_n2255_), .C(men_men_n2252_), .D(x1), .Y(men_men_n2257_));
  NA4        u2208(.A(men_men_n2257_), .B(men_men_n2249_), .C(men_men_n2246_), .D(men_men_n2243_), .Y(men_men_n2258_));
  AO210      u2209(.A0(men_men_n1108_), .A1(men_men_n403_), .B0(men_men_n1021_), .Y(men_men_n2259_));
  NA3        u2210(.A(men_men_n1928_), .B(men_men_n563_), .C(men_men_n280_), .Y(men_men_n2260_));
  AOI210     u2211(.A0(men_men_n2260_), .A1(men_men_n2259_), .B0(men_men_n310_), .Y(men_men_n2261_));
  NA4        u2212(.A(men_men_n1281_), .B(men_men_n535_), .C(men_men_n392_), .D(men_men_n235_), .Y(men_men_n2262_));
  NO3        u2213(.A(men_men_n1453_), .B(men_men_n1021_), .C(x2), .Y(men_men_n2263_));
  NO2        u2214(.A(men_men_n1267_), .B(men_men_n390_), .Y(men_men_n2264_));
  NO2        u2215(.A(men_men_n1856_), .B(men_men_n64_), .Y(men_men_n2265_));
  NO4        u2216(.A(men_men_n2265_), .B(men_men_n2264_), .C(men_men_n2263_), .D(men_men_n53_), .Y(men_men_n2266_));
  NO3        u2217(.A(men_men_n473_), .B(men_men_n1102_), .C(men_men_n123_), .Y(men_men_n2267_));
  OAI220     u2218(.A0(men_men_n696_), .A1(men_men_n176_), .B0(men_men_n359_), .B1(men_men_n144_), .Y(men_men_n2268_));
  OAI210     u2219(.A0(men_men_n2268_), .A1(men_men_n2267_), .B0(men_men_n68_), .Y(men_men_n2269_));
  NO2        u2220(.A(men_men_n2003_), .B(men_men_n371_), .Y(men_men_n2270_));
  OAI210     u2221(.A0(men_men_n1889_), .A1(men_men_n617_), .B0(men_men_n2270_), .Y(men_men_n2271_));
  NA4        u2222(.A(men_men_n2271_), .B(men_men_n2269_), .C(men_men_n2266_), .D(men_men_n2262_), .Y(men_men_n2272_));
  OAI210     u2223(.A0(men_men_n2272_), .A1(men_men_n2261_), .B0(men_men_n2258_), .Y(men_men_n2273_));
  NO3        u2224(.A(men_men_n1231_), .B(men_men_n107_), .C(men_men_n71_), .Y(men_men_n2274_));
  NO2        u2225(.A(men_men_n572_), .B(men_men_n375_), .Y(men_men_n2275_));
  OAI210     u2226(.A0(men_men_n2274_), .A1(men_men_n1432_), .B0(men_men_n2275_), .Y(men_men_n2276_));
  NO3        u2227(.A(x8), .B(men_men_n71_), .C(x2), .Y(men_men_n2277_));
  OAI220     u2228(.A0(men_men_n2277_), .A1(men_men_n633_), .B0(men_men_n1442_), .B1(men_men_n91_), .Y(men_men_n2278_));
  AOI220     u2229(.A0(men_men_n564_), .A1(men_men_n823_), .B0(men_men_n686_), .B1(men_men_n260_), .Y(men_men_n2279_));
  AOI210     u2230(.A0(men_men_n2279_), .A1(men_men_n2278_), .B0(men_men_n270_), .Y(men_men_n2280_));
  NA2        u2231(.A(men_men_n1026_), .B(men_men_n1159_), .Y(men_men_n2281_));
  AOI210     u2232(.A0(men_men_n682_), .A1(men_men_n696_), .B0(men_men_n2281_), .Y(men_men_n2282_));
  AOI210     u2233(.A0(men_men_n597_), .A1(men_men_n633_), .B0(men_men_n702_), .Y(men_men_n2283_));
  NO2        u2234(.A(men_men_n2283_), .B(men_men_n1838_), .Y(men_men_n2284_));
  NO2        u2235(.A(men_men_n457_), .B(men_men_n438_), .Y(men_men_n2285_));
  NOi31      u2236(.An(men_men_n1517_), .B(men_men_n2285_), .C(men_men_n597_), .Y(men_men_n2286_));
  NO4        u2237(.A(men_men_n2286_), .B(men_men_n2284_), .C(men_men_n2282_), .D(men_men_n2280_), .Y(men_men_n2287_));
  NA4        u2238(.A(men_men_n2287_), .B(men_men_n2276_), .C(men_men_n2273_), .D(men_men_n2237_), .Y(men33));
  OAI210     u2239(.A0(men_men_n819_), .A1(x1), .B0(men_men_n205_), .Y(men_men_n2289_));
  OAI210     u2240(.A0(men_men_n2108_), .A1(men_men_n181_), .B0(men_men_n333_), .Y(men_men_n2290_));
  OAI220     u2241(.A0(men_men_n1088_), .A1(men_men_n818_), .B0(men_men_n1691_), .B1(men_men_n358_), .Y(men_men_n2291_));
  NA3        u2242(.A(men_men_n2291_), .B(men_men_n2290_), .C(men_men_n645_), .Y(men_men_n2292_));
  AOI210     u2243(.A0(men_men_n2289_), .A1(x5), .B0(men_men_n2292_), .Y(men_men_n2293_));
  NA2        u2244(.A(men_men_n234_), .B(men_men_n76_), .Y(men_men_n2294_));
  NA4        u2245(.A(men_men_n1766_), .B(men_men_n573_), .C(men_men_n251_), .D(x4), .Y(men_men_n2295_));
  AOI210     u2246(.A0(men_men_n2295_), .A1(men_men_n2294_), .B0(men_men_n358_), .Y(men_men_n2296_));
  OAI210     u2247(.A0(men_men_n441_), .A1(men_men_n274_), .B0(men_men_n53_), .Y(men_men_n2297_));
  AOI210     u2248(.A0(men_men_n2297_), .A1(men_men_n443_), .B0(men_men_n64_), .Y(men_men_n2298_));
  NA2        u2249(.A(men_men_n1679_), .B(men_men_n71_), .Y(men_men_n2299_));
  NO3        u2250(.A(men_men_n2299_), .B(men_men_n2298_), .C(men_men_n2296_), .Y(men_men_n2300_));
  OAI210     u2251(.A0(men_men_n2293_), .A1(x4), .B0(men_men_n2300_), .Y(men_men_n2301_));
  OAI210     u2252(.A0(men_men_n146_), .A1(x5), .B0(men_men_n244_), .Y(men_men_n2302_));
  NO2        u2253(.A(men_men_n972_), .B(men_men_n232_), .Y(men_men_n2303_));
  NA2        u2254(.A(men_men_n648_), .B(x7), .Y(men_men_n2304_));
  NO2        u2255(.A(men_men_n2304_), .B(men_men_n2303_), .Y(men_men_n2305_));
  AOI210     u2256(.A0(men_men_n2302_), .A1(men_men_n1034_), .B0(men_men_n2305_), .Y(men_men_n2306_));
  NA2        u2257(.A(men_men_n216_), .B(men_men_n964_), .Y(men_men_n2307_));
  AOI210     u2258(.A0(men_men_n2307_), .A1(men_men_n2232_), .B0(men_men_n218_), .Y(men_men_n2308_));
  NO2        u2259(.A(men_men_n1665_), .B(men_men_n965_), .Y(men_men_n2309_));
  OAI210     u2260(.A0(men_men_n872_), .A1(men_men_n51_), .B0(x6), .Y(men_men_n2310_));
  NA3        u2261(.A(men_men_n927_), .B(men_men_n738_), .C(men_men_n55_), .Y(men_men_n2311_));
  OAI210     u2262(.A0(men_men_n627_), .A1(men_men_n512_), .B0(men_men_n2311_), .Y(men_men_n2312_));
  NO4        u2263(.A(men_men_n2312_), .B(men_men_n2310_), .C(men_men_n2309_), .D(men_men_n2308_), .Y(men_men_n2313_));
  OAI210     u2264(.A0(men_men_n2306_), .A1(men_men_n50_), .B0(men_men_n2313_), .Y(men_men_n2314_));
  NA3        u2265(.A(men_men_n2314_), .B(men_men_n2301_), .C(men_men_n59_), .Y(men_men_n2315_));
  NO3        u2266(.A(men_men_n1583_), .B(men_men_n379_), .C(x4), .Y(men_men_n2316_));
  AOI210     u2267(.A0(men_men_n2316_), .A1(men_men_n137_), .B0(men_men_n444_), .Y(men_men_n2317_));
  NA2        u2268(.A(men_men_n821_), .B(men_men_n108_), .Y(men_men_n2318_));
  NA2        u2269(.A(men_men_n2318_), .B(men_men_n468_), .Y(men_men_n2319_));
  NO2        u2270(.A(men_men_n717_), .B(men_men_n380_), .Y(men_men_n2320_));
  NA2        u2271(.A(men_men_n508_), .B(men_men_n53_), .Y(men_men_n2321_));
  AOI210     u2272(.A0(men_men_n2320_), .A1(men_men_n2319_), .B0(men_men_n2321_), .Y(men_men_n2322_));
  OAI210     u2273(.A0(men_men_n2317_), .A1(men_men_n59_), .B0(men_men_n2322_), .Y(men_men_n2323_));
  AOI220     u2274(.A0(men_men_n696_), .A1(men_men_n241_), .B0(men_men_n392_), .B1(men_men_n235_), .Y(men_men_n2324_));
  NA2        u2275(.A(men_men_n739_), .B(men_men_n984_), .Y(men_men_n2325_));
  OAI210     u2276(.A0(men_men_n2325_), .A1(men_men_n2324_), .B0(men_men_n309_), .Y(men_men_n2326_));
  AOI210     u2277(.A0(men_men_n2137_), .A1(men_men_n219_), .B0(men_men_n53_), .Y(men_men_n2327_));
  NO2        u2278(.A(men_men_n144_), .B(men_men_n343_), .Y(men_men_n2328_));
  AOI220     u2279(.A0(men_men_n2328_), .A1(men_men_n1004_), .B0(men_men_n681_), .B1(men_men_n358_), .Y(men_men_n2329_));
  NA2        u2280(.A(men_men_n452_), .B(men_men_n506_), .Y(men_men_n2330_));
  NO3        u2281(.A(men_men_n2330_), .B(men_men_n1040_), .C(men_men_n186_), .Y(men_men_n2331_));
  AOI210     u2282(.A0(men_men_n1814_), .A1(men_men_n1203_), .B0(men_men_n2331_), .Y(men_men_n2332_));
  NA4        u2283(.A(men_men_n2332_), .B(men_men_n2329_), .C(men_men_n2327_), .D(men_men_n2326_), .Y(men_men_n2333_));
  NA3        u2284(.A(men_men_n2333_), .B(men_men_n2323_), .C(men_men_n57_), .Y(men_men_n2334_));
  NAi21      u2285(.An(men_men_n1205_), .B(men_men_n496_), .Y(men_men_n2335_));
  NA4        u2286(.A(men_men_n648_), .B(men_men_n1318_), .C(men_men_n477_), .D(men_men_n50_), .Y(men_men_n2336_));
  OAI210     u2287(.A0(men_men_n2328_), .A1(men_men_n2082_), .B0(x2), .Y(men_men_n2337_));
  NA4        u2288(.A(men_men_n292_), .B(men_men_n159_), .C(men_men_n281_), .D(men_men_n123_), .Y(men_men_n2338_));
  NA3        u2289(.A(men_men_n2338_), .B(men_men_n2337_), .C(men_men_n2336_), .Y(men_men_n2339_));
  AO220      u2290(.A0(men_men_n2339_), .A1(x0), .B0(men_men_n2335_), .B1(men_men_n141_), .Y(men_men_n2340_));
  NA3        u2291(.A(men_men_n782_), .B(men_men_n358_), .C(men_men_n60_), .Y(men_men_n2341_));
  NO2        u2292(.A(men_men_n2277_), .B(men_men_n419_), .Y(men_men_n2342_));
  NA2        u2293(.A(men_men_n646_), .B(men_men_n524_), .Y(men_men_n2343_));
  OAI220     u2294(.A0(men_men_n2343_), .A1(men_men_n2342_), .B0(men_men_n2341_), .B1(men_men_n71_), .Y(men_men_n2344_));
  OAI210     u2295(.A0(men_men_n1547_), .A1(men_men_n354_), .B0(men_men_n111_), .Y(men_men_n2345_));
  AOI210     u2296(.A0(men_men_n597_), .A1(men_men_n473_), .B0(men_men_n141_), .Y(men_men_n2346_));
  OAI210     u2297(.A0(men_men_n2346_), .A1(men_men_n392_), .B0(men_men_n2345_), .Y(men_men_n2347_));
  OAI210     u2298(.A0(men_men_n2347_), .A1(men_men_n2344_), .B0(men_men_n102_), .Y(men_men_n2348_));
  NA3        u2299(.A(men_men_n1223_), .B(men_men_n134_), .C(men_men_n387_), .Y(men_men_n2349_));
  NA2        u2300(.A(men_men_n2349_), .B(men_men_n1842_), .Y(men_men_n2350_));
  NA2        u2301(.A(men_men_n1202_), .B(men_men_n718_), .Y(men_men_n2351_));
  AOI220     u2302(.A0(men_men_n2239_), .A1(men_men_n300_), .B0(men_men_n1374_), .B1(men_men_n1183_), .Y(men_men_n2352_));
  NA4        u2303(.A(men_men_n2352_), .B(men_men_n2351_), .C(men_men_n2350_), .D(men_men_n2348_), .Y(men_men_n2353_));
  AOI210     u2304(.A0(men_men_n2340_), .A1(x7), .B0(men_men_n2353_), .Y(men_men_n2354_));
  NA3        u2305(.A(men_men_n2354_), .B(men_men_n2334_), .C(men_men_n2315_), .Y(men34));
  NA2        u2306(.A(men_men_n438_), .B(x4), .Y(men_men_n2356_));
  NO2        u2307(.A(men_men_n1981_), .B(men_men_n865_), .Y(men_men_n2357_));
  AOI210     u2308(.A0(men_men_n2357_), .A1(men_men_n2356_), .B0(men_men_n324_), .Y(men_men_n2358_));
  NA2        u2309(.A(men_men_n292_), .B(men_men_n124_), .Y(men_men_n2359_));
  NO2        u2310(.A(men_men_n982_), .B(men_men_n2359_), .Y(men_men_n2360_));
  AOI210     u2311(.A0(men_men_n2062_), .A1(men_men_n550_), .B0(men_men_n143_), .Y(men_men_n2361_));
  NO2        u2312(.A(men_men_n1851_), .B(men_men_n986_), .Y(men_men_n2362_));
  NO4        u2313(.A(men_men_n2362_), .B(men_men_n2361_), .C(men_men_n2360_), .D(men_men_n2358_), .Y(men_men_n2363_));
  NO2        u2314(.A(men_men_n2363_), .B(men_men_n483_), .Y(men_men_n2364_));
  NA2        u2315(.A(men_men_n741_), .B(x8), .Y(men_men_n2365_));
  AO210      u2316(.A0(men_men_n2365_), .A1(men_men_n493_), .B0(men_men_n671_), .Y(men_men_n2366_));
  NA2        u2317(.A(men_men_n681_), .B(men_men_n638_), .Y(men_men_n2367_));
  AOI210     u2318(.A0(men_men_n2367_), .A1(men_men_n2366_), .B0(men_men_n270_), .Y(men_men_n2368_));
  OAI210     u2319(.A0(men_men_n123_), .A1(men_men_n1062_), .B0(men_men_n1484_), .Y(men_men_n2369_));
  OAI210     u2320(.A0(men_men_n1623_), .A1(men_men_n58_), .B0(men_men_n2369_), .Y(men_men_n2370_));
  NA3        u2321(.A(men_men_n2370_), .B(men_men_n344_), .C(x8), .Y(men_men_n2371_));
  NA2        u2322(.A(men_men_n1605_), .B(men_men_n332_), .Y(men_men_n2372_));
  NA2        u2323(.A(men_men_n675_), .B(men_men_n324_), .Y(men_men_n2373_));
  NA2        u2324(.A(men_men_n137_), .B(x0), .Y(men_men_n2374_));
  NAi31      u2325(.An(men_men_n2374_), .B(men_men_n2373_), .C(men_men_n806_), .Y(men_men_n2375_));
  NA3        u2326(.A(men_men_n1618_), .B(men_men_n1416_), .C(men_men_n50_), .Y(men_men_n2376_));
  NA4        u2327(.A(men_men_n2376_), .B(men_men_n2375_), .C(men_men_n2372_), .D(men_men_n2371_), .Y(men_men_n2377_));
  NA2        u2328(.A(men_men_n1121_), .B(men_men_n757_), .Y(men_men_n2378_));
  NA3        u2329(.A(men_men_n1161_), .B(men_men_n170_), .C(men_men_n1105_), .Y(men_men_n2379_));
  AOI210     u2330(.A0(men_men_n2379_), .A1(men_men_n2378_), .B0(men_men_n767_), .Y(men_men_n2380_));
  AOI210     u2331(.A0(men_men_n1797_), .A1(men_men_n133_), .B0(men_men_n2380_), .Y(men_men_n2381_));
  AOI210     u2332(.A0(men_men_n564_), .A1(men_men_n823_), .B0(men_men_n259_), .Y(men_men_n2382_));
  OAI220     u2333(.A0(men_men_n2382_), .A1(men_men_n59_), .B0(men_men_n1132_), .B1(men_men_n55_), .Y(men_men_n2383_));
  NA3        u2334(.A(men_men_n2383_), .B(men_men_n741_), .C(men_men_n56_), .Y(men_men_n2384_));
  OAI210     u2335(.A0(men_men_n2381_), .A1(men_men_n144_), .B0(men_men_n2384_), .Y(men_men_n2385_));
  NO4        u2336(.A(men_men_n2385_), .B(men_men_n2377_), .C(men_men_n2368_), .D(men_men_n2364_), .Y(men_men_n2386_));
  NO2        u2337(.A(men_men_n316_), .B(men_men_n964_), .Y(men_men_n2387_));
  NO3        u2338(.A(men_men_n2387_), .B(men_men_n450_), .C(men_men_n332_), .Y(men_men_n2388_));
  NA2        u2339(.A(men_men_n791_), .B(men_men_n163_), .Y(men_men_n2389_));
  NO2        u2340(.A(men_men_n2253_), .B(men_men_n309_), .Y(men_men_n2390_));
  OAI220     u2341(.A0(men_men_n2390_), .A1(men_men_n1575_), .B0(men_men_n2389_), .B1(men_men_n1187_), .Y(men_men_n2391_));
  OAI210     u2342(.A0(men_men_n2391_), .A1(men_men_n2388_), .B0(x2), .Y(men_men_n2392_));
  OAI210     u2343(.A0(men_men_n875_), .A1(men_men_n375_), .B0(men_men_n2392_), .Y(men_men_n2393_));
  NA2        u2344(.A(men_men_n319_), .B(x4), .Y(men_men_n2394_));
  OAI220     u2345(.A0(men_men_n753_), .A1(men_men_n55_), .B0(men_men_n285_), .B1(men_men_n107_), .Y(men_men_n2395_));
  NO4        u2346(.A(men_men_n454_), .B(men_men_n77_), .C(x7), .D(x3), .Y(men_men_n2396_));
  NO2        u2347(.A(men_men_n1121_), .B(men_men_n293_), .Y(men_men_n2397_));
  NO4        u2348(.A(men_men_n2397_), .B(men_men_n2396_), .C(men_men_n2395_), .D(men_men_n2394_), .Y(men_men_n2398_));
  NA2        u2349(.A(men_men_n1258_), .B(men_men_n1060_), .Y(men_men_n2399_));
  NA4        u2350(.A(men_men_n741_), .B(men_men_n182_), .C(men_men_n57_), .D(men_men_n108_), .Y(men_men_n2400_));
  NA3        u2351(.A(men_men_n1413_), .B(men_men_n262_), .C(x7), .Y(men_men_n2401_));
  NA3        u2352(.A(men_men_n2401_), .B(men_men_n2400_), .C(men_men_n2399_), .Y(men_men_n2402_));
  OAI210     u2353(.A0(men_men_n2402_), .A1(men_men_n2398_), .B0(men_men_n167_), .Y(men_men_n2403_));
  NA3        u2354(.A(men_men_n870_), .B(men_men_n87_), .C(x0), .Y(men_men_n2404_));
  NA4        u2355(.A(men_men_n2404_), .B(men_men_n1165_), .C(men_men_n302_), .D(men_men_n595_), .Y(men_men_n2405_));
  NA2        u2356(.A(men_men_n1169_), .B(men_men_n686_), .Y(men_men_n2406_));
  OAI210     u2357(.A0(men_men_n2406_), .A1(men_men_n271_), .B0(men_men_n2189_), .Y(men_men_n2407_));
  AOI220     u2358(.A0(men_men_n2407_), .A1(x7), .B0(men_men_n1025_), .B1(men_men_n672_), .Y(men_men_n2408_));
  OAI210     u2359(.A0(men_men_n2075_), .A1(men_men_n267_), .B0(men_men_n745_), .Y(men_men_n2409_));
  AOI220     u2360(.A0(men_men_n415_), .A1(x8), .B0(men_men_n92_), .B1(x2), .Y(men_men_n2410_));
  AOI210     u2361(.A0(men_men_n275_), .A1(men_men_n53_), .B0(men_men_n663_), .Y(men_men_n2411_));
  OAI220     u2362(.A0(men_men_n2411_), .A1(men_men_n97_), .B0(men_men_n2410_), .B1(men_men_n1360_), .Y(men_men_n2412_));
  AOI220     u2363(.A0(men_men_n2412_), .A1(men_men_n1338_), .B0(men_men_n2409_), .B1(men_men_n1532_), .Y(men_men_n2413_));
  NA4        u2364(.A(men_men_n2413_), .B(men_men_n2408_), .C(men_men_n2405_), .D(men_men_n2403_), .Y(men_men_n2414_));
  AOI210     u2365(.A0(men_men_n2393_), .A1(men_men_n823_), .B0(men_men_n2414_), .Y(men_men_n2415_));
  OAI210     u2366(.A0(men_men_n2386_), .A1(x2), .B0(men_men_n2415_), .Y(men35));
  NA2        u2367(.A(men_men_n512_), .B(men_men_n182_), .Y(men_men_n2417_));
  AOI220     u2368(.A0(men_men_n646_), .A1(men_men_n55_), .B0(men_men_n782_), .B1(men_men_n1238_), .Y(men_men_n2418_));
  AOI210     u2369(.A0(men_men_n2418_), .A1(men_men_n2417_), .B0(men_men_n71_), .Y(men_men_n2419_));
  NO3        u2370(.A(men_men_n520_), .B(men_men_n473_), .C(men_men_n343_), .Y(men_men_n2420_));
  OAI210     u2371(.A0(men_men_n2420_), .A1(men_men_n2419_), .B0(x2), .Y(men_men_n2421_));
  AOI210     u2372(.A0(men_men_n220_), .A1(x0), .B0(men_men_n279_), .Y(men_men_n2422_));
  OAI220     u2373(.A0(men_men_n2422_), .A1(men_men_n677_), .B0(men_men_n202_), .B1(x4), .Y(men_men_n2423_));
  NA2        u2374(.A(men_men_n2423_), .B(men_men_n141_), .Y(men_men_n2424_));
  NA3        u2375(.A(men_men_n415_), .B(x8), .C(men_men_n71_), .Y(men_men_n2425_));
  AOI210     u2376(.A0(men_men_n2425_), .A1(men_men_n1742_), .B0(men_men_n696_), .Y(men_men_n2426_));
  OAI210     u2377(.A0(men_men_n2341_), .A1(x6), .B0(men_men_n756_), .Y(men_men_n2427_));
  NO2        u2378(.A(men_men_n2427_), .B(men_men_n2426_), .Y(men_men_n2428_));
  NA3        u2379(.A(men_men_n2428_), .B(men_men_n2424_), .C(men_men_n2421_), .Y(men_men_n2429_));
  NAi21      u2380(.An(men_men_n1706_), .B(men_men_n1314_), .Y(men_men_n2430_));
  NA2        u2381(.A(men_men_n218_), .B(men_men_n582_), .Y(men_men_n2431_));
  NO2        u2382(.A(men_men_n438_), .B(men_men_n431_), .Y(men_men_n2432_));
  AOI220     u2383(.A0(men_men_n2432_), .A1(men_men_n2431_), .B0(men_men_n2430_), .B1(men_men_n56_), .Y(men_men_n2433_));
  NA2        u2384(.A(men_men_n771_), .B(men_men_n709_), .Y(men_men_n2434_));
  NO3        u2385(.A(men_men_n691_), .B(men_men_n55_), .C(x6), .Y(men_men_n2435_));
  OAI210     u2386(.A0(men_men_n2435_), .A1(men_men_n718_), .B0(men_men_n223_), .Y(men_men_n2436_));
  NA2        u2387(.A(men_men_n1346_), .B(men_men_n63_), .Y(men_men_n2437_));
  OAI210     u2388(.A0(men_men_n1084_), .A1(x6), .B0(men_men_n478_), .Y(men_men_n2438_));
  NA3        u2389(.A(men_men_n2438_), .B(men_men_n2437_), .C(men_men_n2436_), .Y(men_men_n2439_));
  NA3        u2390(.A(men_men_n1288_), .B(men_men_n759_), .C(x3), .Y(men_men_n2440_));
  NO3        u2391(.A(men_men_n2440_), .B(men_men_n693_), .C(men_men_n211_), .Y(men_men_n2441_));
  AOI210     u2392(.A0(men_men_n2439_), .A1(men_men_n50_), .B0(men_men_n2441_), .Y(men_men_n2442_));
  OAI210     u2393(.A0(men_men_n2434_), .A1(men_men_n2433_), .B0(men_men_n2442_), .Y(men_men_n2443_));
  AOI210     u2394(.A0(men_men_n2429_), .A1(men_men_n57_), .B0(men_men_n2443_), .Y(men_men_n2444_));
  NA2        u2395(.A(men_men_n972_), .B(men_men_n63_), .Y(men_men_n2445_));
  NO3        u2396(.A(men_men_n1084_), .B(men_men_n572_), .C(men_men_n124_), .Y(men_men_n2446_));
  OAI210     u2397(.A0(men_men_n160_), .A1(men_men_n67_), .B0(men_men_n2446_), .Y(men_men_n2447_));
  AOI210     u2398(.A0(men_men_n2447_), .A1(men_men_n2445_), .B0(men_men_n50_), .Y(men_men_n2448_));
  NA4        u2399(.A(men_men_n473_), .B(men_men_n235_), .C(men_men_n880_), .D(men_men_n104_), .Y(men_men_n2449_));
  OAI210     u2400(.A0(men_men_n972_), .A1(men_men_n260_), .B0(men_men_n760_), .Y(men_men_n2450_));
  OAI210     u2401(.A0(men_men_n260_), .A1(men_men_n594_), .B0(men_men_n2186_), .Y(men_men_n2451_));
  NA3        u2402(.A(men_men_n2451_), .B(men_men_n2450_), .C(men_men_n2449_), .Y(men_men_n2452_));
  OAI210     u2403(.A0(men_men_n2452_), .A1(men_men_n2448_), .B0(men_men_n59_), .Y(men_men_n2453_));
  AOI210     u2404(.A0(men_men_n870_), .A1(men_men_n541_), .B0(men_men_n1928_), .Y(men_men_n2454_));
  AOI210     u2405(.A0(men_men_n572_), .A1(men_men_n616_), .B0(men_men_n2454_), .Y(men_men_n2455_));
  NO4        u2406(.A(men_men_n965_), .B(men_men_n572_), .C(men_men_n367_), .D(men_men_n413_), .Y(men_men_n2456_));
  XN2        u2407(.A(x4), .B(x3), .Y(men_men_n2457_));
  NO3        u2408(.A(men_men_n2457_), .B(men_men_n676_), .C(men_men_n315_), .Y(men_men_n2458_));
  NO3        u2409(.A(men_men_n2458_), .B(men_men_n2456_), .C(men_men_n1482_), .Y(men_men_n2459_));
  OAI210     u2410(.A0(men_men_n2455_), .A1(x3), .B0(men_men_n2459_), .Y(men_men_n2460_));
  NO3        u2411(.A(men_men_n753_), .B(men_men_n872_), .C(men_men_n280_), .Y(men_men_n2461_));
  OAI210     u2412(.A0(men_men_n2461_), .A1(men_men_n1482_), .B0(men_men_n50_), .Y(men_men_n2462_));
  INV        u2413(.A(men_men_n2462_), .Y(men_men_n2463_));
  AOI210     u2414(.A0(men_men_n2460_), .A1(men_men_n597_), .B0(men_men_n2463_), .Y(men_men_n2464_));
  AOI210     u2415(.A0(men_men_n1453_), .A1(men_men_n653_), .B0(men_men_n693_), .Y(men_men_n2465_));
  NO2        u2416(.A(men_men_n880_), .B(men_men_n56_), .Y(men_men_n2466_));
  OAI210     u2417(.A0(men_men_n1984_), .A1(men_men_n616_), .B0(men_men_n2277_), .Y(men_men_n2467_));
  OAI210     u2418(.A0(men_men_n2365_), .A1(men_men_n2466_), .B0(men_men_n2467_), .Y(men_men_n2468_));
  OAI210     u2419(.A0(men_men_n2468_), .A1(men_men_n2465_), .B0(men_men_n92_), .Y(men_men_n2469_));
  NO2        u2420(.A(men_men_n863_), .B(men_men_n673_), .Y(men_men_n2470_));
  NO2        u2421(.A(men_men_n293_), .B(x6), .Y(men_men_n2471_));
  OAI210     u2422(.A0(men_men_n2470_), .A1(men_men_n1805_), .B0(men_men_n2471_), .Y(men_men_n2472_));
  NA4        u2423(.A(men_men_n2472_), .B(men_men_n2469_), .C(men_men_n2464_), .D(men_men_n2453_), .Y(men_men_n2473_));
  NA4        u2424(.A(men_men_n624_), .B(men_men_n696_), .C(men_men_n437_), .D(x6), .Y(men_men_n2474_));
  AOI210     u2425(.A0(men_men_n2474_), .A1(men_men_n432_), .B0(x1), .Y(men_men_n2475_));
  NO2        u2426(.A(men_men_n739_), .B(men_men_n693_), .Y(men_men_n2476_));
  OAI210     u2427(.A0(men_men_n473_), .A1(men_men_n171_), .B0(men_men_n803_), .Y(men_men_n2477_));
  AOI210     u2428(.A0(men_men_n2477_), .A1(men_men_n1030_), .B0(men_men_n53_), .Y(men_men_n2478_));
  NO3        u2429(.A(men_men_n2478_), .B(men_men_n2476_), .C(men_men_n2475_), .Y(men_men_n2479_));
  NA3        u2430(.A(men_men_n1455_), .B(men_men_n1289_), .C(men_men_n827_), .Y(men_men_n2480_));
  AOI220     u2431(.A0(men_men_n1971_), .A1(men_men_n141_), .B0(men_men_n424_), .B1(men_men_n128_), .Y(men_men_n2481_));
  AOI210     u2432(.A0(men_men_n2481_), .A1(men_men_n2480_), .B0(men_men_n1525_), .Y(men_men_n2482_));
  NO2        u2433(.A(men_men_n646_), .B(x3), .Y(men_men_n2483_));
  NO3        u2434(.A(men_men_n704_), .B(men_men_n1623_), .C(x2), .Y(men_men_n2484_));
  AOI220     u2435(.A0(men_men_n2484_), .A1(men_men_n2483_), .B0(men_men_n1944_), .B1(men_men_n778_), .Y(men_men_n2485_));
  NA3        u2436(.A(x6), .B(x4), .C(x0), .Y(men_men_n2486_));
  OAI220     u2437(.A0(men_men_n2486_), .A1(men_men_n201_), .B0(men_men_n691_), .B1(men_men_n537_), .Y(men_men_n2487_));
  OAI220     u2438(.A0(men_men_n1327_), .A1(x8), .B0(men_men_n379_), .B1(men_men_n357_), .Y(men_men_n2488_));
  AOI220     u2439(.A0(men_men_n2488_), .A1(men_men_n424_), .B0(men_men_n2487_), .B1(men_men_n926_), .Y(men_men_n2489_));
  OAI210     u2440(.A0(men_men_n2485_), .A1(men_men_n1178_), .B0(men_men_n2489_), .Y(men_men_n2490_));
  NO2        u2441(.A(men_men_n2490_), .B(men_men_n2482_), .Y(men_men_n2491_));
  OAI210     u2442(.A0(men_men_n2479_), .A1(men_men_n319_), .B0(men_men_n2491_), .Y(men_men_n2492_));
  AOI210     u2443(.A0(men_men_n2473_), .A1(x5), .B0(men_men_n2492_), .Y(men_men_n2493_));
  OAI210     u2444(.A0(men_men_n2444_), .A1(x5), .B0(men_men_n2493_), .Y(men36));
  NO2        u2445(.A(men_men_n872_), .B(men_men_n308_), .Y(men_men_n2495_));
  NO3        u2446(.A(men_men_n123_), .B(men_men_n1062_), .C(men_men_n55_), .Y(men_men_n2496_));
  NO3        u2447(.A(men_men_n2496_), .B(men_men_n2003_), .C(men_men_n1084_), .Y(men_men_n2497_));
  OAI210     u2448(.A0(men_men_n2497_), .A1(men_men_n2495_), .B0(men_men_n110_), .Y(men_men_n2498_));
  OR4        u2449(.A(men_men_n966_), .B(men_men_n814_), .C(men_men_n382_), .D(men_men_n500_), .Y(men_men_n2499_));
  INV        u2450(.A(men_men_n1015_), .Y(men_men_n2500_));
  OAI210     u2451(.A0(men_men_n2239_), .A1(men_men_n2500_), .B0(men_men_n285_), .Y(men_men_n2501_));
  NA3        u2452(.A(men_men_n452_), .B(men_men_n232_), .C(men_men_n122_), .Y(men_men_n2502_));
  NA4        u2453(.A(men_men_n2502_), .B(men_men_n2501_), .C(men_men_n2499_), .D(men_men_n2498_), .Y(men_men_n2503_));
  NO2        u2454(.A(men_men_n1004_), .B(x8), .Y(men_men_n2504_));
  NO3        u2455(.A(men_men_n2504_), .B(men_men_n1000_), .C(men_men_n546_), .Y(men_men_n2505_));
  AOI220     u2456(.A0(men_men_n309_), .A1(x1), .B0(men_men_n140_), .B1(x6), .Y(men_men_n2506_));
  AOI210     u2457(.A0(men_men_n1105_), .A1(x6), .B0(men_men_n428_), .Y(men_men_n2507_));
  OAI220     u2458(.A0(men_men_n2507_), .A1(men_men_n366_), .B0(men_men_n2506_), .B1(men_men_n474_), .Y(men_men_n2508_));
  OAI210     u2459(.A0(men_men_n2508_), .A1(men_men_n2505_), .B0(men_men_n473_), .Y(men_men_n2509_));
  NA2        u2460(.A(men_men_n681_), .B(men_men_n500_), .Y(men_men_n2510_));
  AOI210     u2461(.A0(men_men_n2510_), .A1(men_men_n660_), .B0(men_men_n271_), .Y(men_men_n2511_));
  NO3        u2462(.A(men_men_n1899_), .B(men_men_n1622_), .C(men_men_n281_), .Y(men_men_n2512_));
  NO2        u2463(.A(men_men_n2445_), .B(men_men_n234_), .Y(men_men_n2513_));
  NO4        u2464(.A(men_men_n2513_), .B(men_men_n2512_), .C(men_men_n2511_), .D(men_men_n426_), .Y(men_men_n2514_));
  OAI210     u2465(.A0(men_men_n648_), .A1(men_men_n813_), .B0(men_men_n990_), .Y(men_men_n2515_));
  OAI220     u2466(.A0(men_men_n1670_), .A1(men_men_n1665_), .B0(men_men_n990_), .B1(men_men_n1105_), .Y(men_men_n2516_));
  AOI220     u2467(.A0(men_men_n2516_), .A1(men_men_n121_), .B0(men_men_n2515_), .B1(men_men_n638_), .Y(men_men_n2517_));
  NA3        u2468(.A(men_men_n2517_), .B(men_men_n2514_), .C(men_men_n2509_), .Y(men_men_n2518_));
  AOI210     u2469(.A0(men_men_n2503_), .A1(men_men_n344_), .B0(men_men_n2518_), .Y(men_men_n2519_));
  OAI210     u2470(.A0(men_men_n602_), .A1(men_men_n525_), .B0(men_men_n171_), .Y(men_men_n2520_));
  OAI210     u2471(.A0(men_men_n2018_), .A1(men_men_n70_), .B0(men_men_n2520_), .Y(men_men_n2521_));
  OAI210     u2472(.A0(men_men_n503_), .A1(men_men_n243_), .B0(men_men_n260_), .Y(men_men_n2522_));
  NO2        u2473(.A(men_men_n2027_), .B(men_men_n178_), .Y(men_men_n2523_));
  NA2        u2474(.A(men_men_n1225_), .B(men_men_n55_), .Y(men_men_n2524_));
  OAI210     u2475(.A0(men_men_n2524_), .A1(men_men_n2523_), .B0(men_men_n2522_), .Y(men_men_n2525_));
  OAI210     u2476(.A0(men_men_n2525_), .A1(men_men_n2521_), .B0(men_men_n904_), .Y(men_men_n2526_));
  AOI210     u2477(.A0(men_men_n107_), .A1(men_men_n110_), .B0(men_men_n346_), .Y(men_men_n2527_));
  NA2        u2478(.A(men_men_n681_), .B(men_men_n1623_), .Y(men_men_n2528_));
  OAI220     u2479(.A0(men_men_n2528_), .A1(men_men_n2527_), .B0(men_men_n756_), .B1(men_men_n1272_), .Y(men_men_n2529_));
  NO2        u2480(.A(men_men_n1416_), .B(men_men_n588_), .Y(men_men_n2530_));
  NO3        u2481(.A(men_men_n2530_), .B(men_men_n1813_), .C(men_men_n704_), .Y(men_men_n2531_));
  NOi31      u2482(.An(men_men_n2039_), .B(men_men_n2330_), .C(men_men_n766_), .Y(men_men_n2532_));
  NO3        u2483(.A(men_men_n2532_), .B(men_men_n2531_), .C(men_men_n2529_), .Y(men_men_n2533_));
  AOI210     u2484(.A0(men_men_n2533_), .A1(men_men_n2526_), .B0(x7), .Y(men_men_n2534_));
  NA2        u2485(.A(men_men_n140_), .B(men_men_n63_), .Y(men_men_n2535_));
  AOI210     u2486(.A0(men_men_n597_), .A1(men_men_n633_), .B0(men_men_n1203_), .Y(men_men_n2536_));
  NA3        u2487(.A(men_men_n2536_), .B(men_men_n2535_), .C(men_men_n897_), .Y(men_men_n2537_));
  NA2        u2488(.A(men_men_n2537_), .B(men_men_n512_), .Y(men_men_n2538_));
  AOI220     u2489(.A0(men_men_n1766_), .A1(men_men_n263_), .B0(men_men_n1060_), .B1(men_men_n128_), .Y(men_men_n2539_));
  NO2        u2490(.A(men_men_n2539_), .B(men_men_n452_), .Y(men_men_n2540_));
  NO2        u2491(.A(men_men_n413_), .B(men_men_n232_), .Y(men_men_n2541_));
  NO3        u2492(.A(men_men_n2541_), .B(men_men_n1293_), .C(men_men_n59_), .Y(men_men_n2542_));
  AOI210     u2493(.A0(men_men_n1242_), .A1(men_men_n414_), .B0(x6), .Y(men_men_n2543_));
  NA3        u2494(.A(men_men_n1697_), .B(men_men_n285_), .C(men_men_n275_), .Y(men_men_n2544_));
  NA2        u2495(.A(men_men_n2544_), .B(men_men_n1650_), .Y(men_men_n2545_));
  NO4        u2496(.A(men_men_n2545_), .B(men_men_n2543_), .C(men_men_n2542_), .D(men_men_n2540_), .Y(men_men_n2546_));
  AOI210     u2497(.A0(men_men_n2546_), .A1(men_men_n2538_), .B0(men_men_n462_), .Y(men_men_n2547_));
  NO3        u2498(.A(men_men_n2457_), .B(men_men_n910_), .C(men_men_n511_), .Y(men_men_n2548_));
  AOI210     u2499(.A0(men_men_n1291_), .A1(men_men_n274_), .B0(men_men_n2548_), .Y(men_men_n2549_));
  OAI210     u2500(.A0(men_men_n879_), .A1(men_men_n280_), .B0(men_men_n403_), .Y(men_men_n2550_));
  NA2        u2501(.A(men_men_n1225_), .B(men_men_n176_), .Y(men_men_n2551_));
  NO2        u2502(.A(men_men_n623_), .B(men_men_n110_), .Y(men_men_n2552_));
  AO210      u2503(.A0(men_men_n2552_), .A1(men_men_n2551_), .B0(men_men_n1783_), .Y(men_men_n2553_));
  NO2        u2504(.A(men_men_n469_), .B(men_men_n425_), .Y(men_men_n2554_));
  AOI220     u2505(.A0(men_men_n2554_), .A1(men_men_n2553_), .B0(men_men_n2550_), .B1(men_men_n300_), .Y(men_men_n2555_));
  OAI210     u2506(.A0(men_men_n2549_), .A1(x1), .B0(men_men_n2555_), .Y(men_men_n2556_));
  NO3        u2507(.A(men_men_n2556_), .B(men_men_n2547_), .C(men_men_n2534_), .Y(men_men_n2557_));
  OAI210     u2508(.A0(men_men_n2519_), .A1(men_men_n57_), .B0(men_men_n2557_), .Y(men37));
  NA3        u2509(.A(men_men_n1081_), .B(men_men_n143_), .C(x3), .Y(men_men_n2559_));
  NA3        u2510(.A(men_men_n791_), .B(men_men_n163_), .C(men_men_n50_), .Y(men_men_n2560_));
  AOI210     u2511(.A0(men_men_n2560_), .A1(men_men_n2559_), .B0(men_men_n697_), .Y(men_men_n2561_));
  NO3        u2512(.A(men_men_n1081_), .B(men_men_n382_), .C(men_men_n519_), .Y(men_men_n2562_));
  OAI210     u2513(.A0(men_men_n2562_), .A1(men_men_n2561_), .B0(men_men_n56_), .Y(men_men_n2563_));
  NA2        u2514(.A(men_men_n611_), .B(men_men_n757_), .Y(men_men_n2564_));
  AOI210     u2515(.A0(men_men_n2564_), .A1(men_men_n1061_), .B0(x3), .Y(men_men_n2565_));
  AOI220     u2516(.A0(men_men_n611_), .A1(men_men_n757_), .B0(men_men_n473_), .B1(men_men_n1060_), .Y(men_men_n2566_));
  NO2        u2517(.A(men_men_n676_), .B(men_men_n185_), .Y(men_men_n2567_));
  OAI220     u2518(.A0(men_men_n2567_), .A1(men_men_n848_), .B0(men_men_n2566_), .B1(men_men_n110_), .Y(men_men_n2568_));
  OAI210     u2519(.A0(men_men_n2568_), .A1(men_men_n2565_), .B0(men_men_n71_), .Y(men_men_n2569_));
  NA2        u2520(.A(men_men_n1205_), .B(men_men_n1084_), .Y(men_men_n2570_));
  OAI210     u2521(.A0(men_men_n1227_), .A1(men_men_n195_), .B0(men_men_n463_), .Y(men_men_n2571_));
  NA4        u2522(.A(men_men_n2571_), .B(men_men_n2570_), .C(men_men_n2569_), .D(men_men_n2563_), .Y(men_men_n2572_));
  NA2        u2523(.A(men_men_n431_), .B(men_men_n140_), .Y(men_men_n2573_));
  NO2        u2524(.A(men_men_n1728_), .B(men_men_n109_), .Y(men_men_n2574_));
  AOI210     u2525(.A0(men_men_n2005_), .A1(men_men_n873_), .B0(men_men_n2574_), .Y(men_men_n2575_));
  OAI220     u2526(.A0(men_men_n2575_), .A1(men_men_n51_), .B0(men_men_n1624_), .B1(men_men_n2573_), .Y(men_men_n2576_));
  AOI210     u2527(.A0(men_men_n2572_), .A1(men_men_n68_), .B0(men_men_n2576_), .Y(men_men_n2577_));
  OAI210     u2528(.A0(men_men_n275_), .A1(men_men_n1109_), .B0(men_men_n494_), .Y(men_men_n2578_));
  NA3        u2529(.A(men_men_n2578_), .B(men_men_n271_), .C(men_men_n1062_), .Y(men_men_n2579_));
  OAI210     u2530(.A0(men_men_n235_), .A1(men_men_n223_), .B0(men_men_n1742_), .Y(men_men_n2580_));
  NA2        u2531(.A(men_men_n352_), .B(men_men_n279_), .Y(men_men_n2581_));
  NA3        u2532(.A(men_men_n409_), .B(men_men_n827_), .C(men_men_n110_), .Y(men_men_n2582_));
  NO2        u2533(.A(men_men_n538_), .B(men_men_n56_), .Y(men_men_n2583_));
  NA3        u2534(.A(men_men_n2583_), .B(men_men_n2582_), .C(men_men_n2581_), .Y(men_men_n2584_));
  AOI210     u2535(.A0(men_men_n2580_), .A1(men_men_n519_), .B0(men_men_n2584_), .Y(men_men_n2585_));
  NO2        u2536(.A(men_men_n1196_), .B(men_men_n280_), .Y(men_men_n2586_));
  OAI210     u2537(.A0(men_men_n300_), .A1(men_men_n269_), .B0(men_men_n2586_), .Y(men_men_n2587_));
  OAI210     u2538(.A0(men_men_n678_), .A1(men_men_n141_), .B0(x3), .Y(men_men_n2588_));
  AOI210     u2539(.A0(men_men_n678_), .A1(men_men_n371_), .B0(men_men_n2588_), .Y(men_men_n2589_));
  AOI210     u2540(.A0(men_men_n1623_), .A1(men_men_n50_), .B0(men_men_n352_), .Y(men_men_n2590_));
  OAI210     u2541(.A0(men_men_n2590_), .A1(men_men_n408_), .B0(men_men_n56_), .Y(men_men_n2591_));
  NO2        u2542(.A(men_men_n2591_), .B(men_men_n2589_), .Y(men_men_n2592_));
  AOI220     u2543(.A0(men_men_n2592_), .A1(men_men_n2587_), .B0(men_men_n2585_), .B1(men_men_n2579_), .Y(men_men_n2593_));
  OAI210     u2544(.A0(men_men_n2593_), .A1(men_men_n1781_), .B0(men_men_n102_), .Y(men_men_n2594_));
  NO2        u2545(.A(men_men_n2250_), .B(men_men_n55_), .Y(men_men_n2595_));
  OAI210     u2546(.A0(men_men_n2595_), .A1(men_men_n111_), .B0(men_men_n1842_), .Y(men_men_n2596_));
  NA2        u2547(.A(men_men_n182_), .B(men_men_n108_), .Y(men_men_n2597_));
  NA2        u2548(.A(men_men_n696_), .B(x6), .Y(men_men_n2598_));
  AOI210     u2549(.A0(men_men_n2598_), .A1(men_men_n493_), .B0(men_men_n2597_), .Y(men_men_n2599_));
  AOI210     u2550(.A0(men_men_n359_), .A1(men_men_n143_), .B0(men_men_n144_), .Y(men_men_n2600_));
  OAI210     u2551(.A0(men_men_n2600_), .A1(men_men_n2599_), .B0(men_men_n352_), .Y(men_men_n2601_));
  AOI210     u2552(.A0(men_men_n624_), .A1(men_men_n441_), .B0(men_men_n1303_), .Y(men_men_n2602_));
  NO3        u2553(.A(men_men_n2602_), .B(men_men_n271_), .C(men_men_n63_), .Y(men_men_n2603_));
  OAI220     u2554(.A0(men_men_n2365_), .A1(men_men_n491_), .B0(men_men_n2120_), .B1(men_men_n392_), .Y(men_men_n2604_));
  OAI210     u2555(.A0(men_men_n2604_), .A1(men_men_n2603_), .B0(men_men_n53_), .Y(men_men_n2605_));
  NO4        u2556(.A(men_men_n2374_), .B(men_men_n944_), .C(men_men_n442_), .D(men_men_n226_), .Y(men_men_n2606_));
  NO4        u2557(.A(men_men_n741_), .B(men_men_n612_), .C(men_men_n450_), .D(men_men_n1070_), .Y(men_men_n2607_));
  NO3        u2558(.A(men_men_n2607_), .B(men_men_n2606_), .C(men_men_n1076_), .Y(men_men_n2608_));
  NA4        u2559(.A(men_men_n2608_), .B(men_men_n2605_), .C(men_men_n2601_), .D(men_men_n2596_), .Y(men_men_n2609_));
  NO3        u2560(.A(men_men_n255_), .B(men_men_n358_), .C(men_men_n84_), .Y(men_men_n2610_));
  NO2        u2561(.A(men_men_n283_), .B(men_men_n782_), .Y(men_men_n2611_));
  NO3        u2562(.A(men_men_n2611_), .B(men_men_n1225_), .C(men_men_n1244_), .Y(men_men_n2612_));
  OAI220     u2563(.A0(men_men_n2612_), .A1(men_men_n2610_), .B0(men_men_n473_), .B1(men_men_n85_), .Y(men_men_n2613_));
  OR2        u2564(.A(men_men_n950_), .B(men_men_n759_), .Y(men_men_n2614_));
  NA2        u2565(.A(men_men_n1238_), .B(men_men_n55_), .Y(men_men_n2615_));
  NOi21      u2566(.An(men_men_n2615_), .B(men_men_n393_), .Y(men_men_n2616_));
  AOI210     u2567(.A0(men_men_n2616_), .A1(men_men_n2614_), .B0(x1), .Y(men_men_n2617_));
  NA2        u2568(.A(men_men_n270_), .B(men_men_n84_), .Y(men_men_n2618_));
  AOI210     u2569(.A0(men_men_n1575_), .A1(men_men_n408_), .B0(men_men_n2618_), .Y(men_men_n2619_));
  NA2        u2570(.A(men_men_n1121_), .B(men_men_n62_), .Y(men_men_n2620_));
  NA2        u2571(.A(men_men_n1169_), .B(men_men_n178_), .Y(men_men_n2621_));
  OAI210     u2572(.A0(men_men_n2620_), .A1(men_men_n318_), .B0(men_men_n2621_), .Y(men_men_n2622_));
  NO3        u2573(.A(men_men_n2622_), .B(men_men_n2619_), .C(men_men_n2617_), .Y(men_men_n2623_));
  OAI210     u2574(.A0(men_men_n2623_), .A1(x6), .B0(men_men_n2613_), .Y(men_men_n2624_));
  AOI220     u2575(.A0(men_men_n2624_), .A1(men_men_n1484_), .B0(men_men_n2609_), .B1(men_men_n57_), .Y(men_men_n2625_));
  NA3        u2576(.A(men_men_n2625_), .B(men_men_n2594_), .C(men_men_n2577_), .Y(men38));
  AOI210     u2577(.A0(men_men_n1682_), .A1(men_men_n191_), .B0(men_men_n984_), .Y(men_men_n2627_));
  AOI210     u2578(.A0(men_men_n1242_), .A1(men_men_n587_), .B0(men_men_n1102_), .Y(men_men_n2628_));
  AOI210     u2579(.A0(men_men_n2615_), .A1(men_men_n1874_), .B0(men_men_n234_), .Y(men_men_n2629_));
  NO3        u2580(.A(men_men_n1313_), .B(men_men_n324_), .C(x8), .Y(men_men_n2630_));
  NO4        u2581(.A(men_men_n2630_), .B(men_men_n2629_), .C(men_men_n2628_), .D(men_men_n2627_), .Y(men_men_n2631_));
  NO2        u2582(.A(men_men_n2631_), .B(x6), .Y(men_men_n2632_));
  NA4        u2583(.A(men_men_n384_), .B(men_men_n262_), .C(men_men_n194_), .D(x8), .Y(men_men_n2633_));
  NA2        u2584(.A(men_men_n407_), .B(men_men_n108_), .Y(men_men_n2634_));
  AOI210     u2585(.A0(men_men_n2634_), .A1(men_men_n2633_), .B0(men_men_n144_), .Y(men_men_n2635_));
  AOI210     u2586(.A0(men_men_n442_), .A1(men_men_n412_), .B0(men_men_n1752_), .Y(men_men_n2636_));
  NO2        u2587(.A(men_men_n2636_), .B(men_men_n194_), .Y(men_men_n2637_));
  OAI210     u2588(.A0(men_men_n2637_), .A1(men_men_n2635_), .B0(x6), .Y(men_men_n2638_));
  NO2        u2589(.A(men_men_n252_), .B(men_men_n782_), .Y(men_men_n2639_));
  NO3        u2590(.A(men_men_n2639_), .B(men_men_n1706_), .C(men_men_n262_), .Y(men_men_n2640_));
  NO3        u2591(.A(x3), .B(men_men_n53_), .C(x0), .Y(men_men_n2641_));
  OAI210     u2592(.A0(men_men_n531_), .A1(x2), .B0(men_men_n2641_), .Y(men_men_n2642_));
  NA3        u2593(.A(men_men_n441_), .B(men_men_n431_), .C(men_men_n299_), .Y(men_men_n2643_));
  NA3        u2594(.A(men_men_n2643_), .B(men_men_n2642_), .C(men_men_n1832_), .Y(men_men_n2644_));
  OAI210     u2595(.A0(men_men_n2644_), .A1(men_men_n2640_), .B0(men_men_n823_), .Y(men_men_n2645_));
  NO2        u2596(.A(men_men_n612_), .B(men_men_n281_), .Y(men_men_n2646_));
  AN3        u2597(.A(men_men_n828_), .B(men_men_n791_), .C(x0), .Y(men_men_n2647_));
  OAI210     u2598(.A0(men_men_n2647_), .A1(men_men_n2646_), .B0(men_men_n333_), .Y(men_men_n2648_));
  OAI220     u2599(.A0(men_men_n612_), .A1(men_men_n281_), .B0(men_men_n827_), .B1(men_men_n93_), .Y(men_men_n2649_));
  OAI210     u2600(.A0(men_men_n696_), .A1(x0), .B0(men_men_n51_), .Y(men_men_n2650_));
  AOI210     u2601(.A0(men_men_n593_), .A1(x4), .B0(men_men_n233_), .Y(men_men_n2651_));
  AOI220     u2602(.A0(men_men_n2651_), .A1(men_men_n2650_), .B0(men_men_n2649_), .B1(men_men_n409_), .Y(men_men_n2652_));
  NA4        u2603(.A(men_men_n2652_), .B(men_men_n2648_), .C(men_men_n2645_), .D(men_men_n2638_), .Y(men_men_n2653_));
  OAI210     u2604(.A0(men_men_n2653_), .A1(men_men_n2632_), .B0(x7), .Y(men_men_n2654_));
  AOI210     u2605(.A0(men_men_n380_), .A1(x1), .B0(men_men_n1250_), .Y(men_men_n2655_));
  NO2        u2606(.A(men_men_n2655_), .B(men_men_n51_), .Y(men_men_n2656_));
  AOI210     u2607(.A0(men_men_n92_), .A1(men_men_n71_), .B0(men_men_n2277_), .Y(men_men_n2657_));
  NA2        u2608(.A(men_men_n392_), .B(x3), .Y(men_men_n2658_));
  NO2        u2609(.A(men_men_n1773_), .B(men_men_n538_), .Y(men_men_n2659_));
  OAI210     u2610(.A0(men_men_n2658_), .A1(men_men_n2657_), .B0(men_men_n2659_), .Y(men_men_n2660_));
  OAI210     u2611(.A0(men_men_n2660_), .A1(men_men_n2656_), .B0(x4), .Y(men_men_n2661_));
  NO2        u2612(.A(men_men_n1784_), .B(men_men_n467_), .Y(men_men_n2662_));
  NO3        u2613(.A(men_men_n2662_), .B(men_men_n408_), .C(men_men_n121_), .Y(men_men_n2663_));
  AOI210     u2614(.A0(men_men_n1070_), .A1(men_men_n246_), .B0(men_men_n401_), .Y(men_men_n2664_));
  AO210      u2615(.A0(men_men_n1319_), .A1(x6), .B0(men_men_n2664_), .Y(men_men_n2665_));
  NO2        u2616(.A(men_men_n1438_), .B(men_men_n141_), .Y(men_men_n2666_));
  NA2        u2617(.A(men_men_n1981_), .B(men_men_n327_), .Y(men_men_n2667_));
  OAI220     u2618(.A0(men_men_n2667_), .A1(men_men_n1089_), .B0(men_men_n2666_), .B1(men_men_n1856_), .Y(men_men_n2668_));
  NO3        u2619(.A(men_men_n2668_), .B(men_men_n2665_), .C(men_men_n2663_), .Y(men_men_n2669_));
  AOI210     u2620(.A0(men_men_n2669_), .A1(men_men_n2661_), .B0(men_men_n108_), .Y(men_men_n2670_));
  NA3        u2621(.A(men_men_n1971_), .B(men_men_n612_), .C(men_men_n167_), .Y(men_men_n2671_));
  AOI210     u2622(.A0(men_men_n2671_), .A1(men_men_n1449_), .B0(men_men_n235_), .Y(men_men_n2672_));
  AOI210     u2623(.A0(men_men_n512_), .A1(men_men_n500_), .B0(men_men_n692_), .Y(men_men_n2673_));
  OAI220     u2624(.A0(men_men_n2673_), .A1(men_men_n474_), .B0(men_men_n202_), .B1(men_men_n119_), .Y(men_men_n2674_));
  OAI210     u2625(.A0(men_men_n2674_), .A1(men_men_n2672_), .B0(x0), .Y(men_men_n2675_));
  NA3        u2626(.A(men_men_n412_), .B(men_men_n827_), .C(men_men_n281_), .Y(men_men_n2676_));
  AOI210     u2627(.A0(men_men_n2676_), .A1(men_men_n724_), .B0(men_men_n2234_), .Y(men_men_n2677_));
  NA2        u2628(.A(men_men_n1141_), .B(men_men_n964_), .Y(men_men_n2678_));
  NA4        u2629(.A(men_men_n691_), .B(men_men_n612_), .C(men_men_n182_), .D(x3), .Y(men_men_n2679_));
  AOI210     u2630(.A0(men_men_n2679_), .A1(men_men_n2678_), .B0(men_men_n506_), .Y(men_men_n2680_));
  NO4        u2631(.A(men_men_n1431_), .B(men_men_n527_), .C(men_men_n1244_), .D(men_men_n782_), .Y(men_men_n2681_));
  OAI220     u2632(.A0(men_men_n1803_), .A1(men_men_n2318_), .B0(men_men_n233_), .B1(men_men_n153_), .Y(men_men_n2682_));
  NO4        u2633(.A(men_men_n2682_), .B(men_men_n2681_), .C(men_men_n2680_), .D(men_men_n2677_), .Y(men_men_n2683_));
  NA2        u2634(.A(men_men_n2683_), .B(men_men_n2675_), .Y(men_men_n2684_));
  OAI210     u2635(.A0(men_men_n2684_), .A1(men_men_n2670_), .B0(men_men_n57_), .Y(men_men_n2685_));
  AOI210     u2636(.A0(men_men_n1843_), .A1(men_men_n281_), .B0(men_men_n693_), .Y(men_men_n2686_));
  OAI210     u2637(.A0(men_men_n1780_), .A1(men_men_n218_), .B0(men_men_n502_), .Y(men_men_n2687_));
  OAI210     u2638(.A0(men_men_n2687_), .A1(men_men_n2686_), .B0(men_men_n640_), .Y(men_men_n2688_));
  OAI220     u2639(.A0(men_men_n1787_), .A1(men_men_n281_), .B0(men_men_n261_), .B1(men_men_n104_), .Y(men_men_n2689_));
  NA2        u2640(.A(men_men_n1893_), .B(men_men_n360_), .Y(men_men_n2690_));
  OAI220     u2641(.A0(men_men_n2690_), .A1(men_men_n648_), .B0(men_men_n703_), .B1(men_men_n153_), .Y(men_men_n2691_));
  AOI210     u2642(.A0(men_men_n2689_), .A1(men_men_n1004_), .B0(men_men_n2691_), .Y(men_men_n2692_));
  NA4        u2643(.A(men_men_n2692_), .B(men_men_n2688_), .C(men_men_n2685_), .D(men_men_n2654_), .Y(men39));
  INV        u2644(.A(men_men_n124_), .Y(men_men_n2696_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
  VOTADOR g14(.A(ori14), .B(mai14), .C(men14), .Y(z14));
  VOTADOR g15(.A(ori15), .B(mai15), .C(men15), .Y(z15));
  VOTADOR g16(.A(ori16), .B(mai16), .C(men16), .Y(z16));
  VOTADOR g17(.A(ori17), .B(mai17), .C(men17), .Y(z17));
  VOTADOR g18(.A(ori18), .B(mai18), .C(men18), .Y(z18));
  VOTADOR g19(.A(ori19), .B(mai19), .C(men19), .Y(z19));
  VOTADOR g20(.A(ori20), .B(mai20), .C(men20), .Y(z20));
  VOTADOR g21(.A(ori21), .B(mai21), .C(men21), .Y(z21));
  VOTADOR g22(.A(ori22), .B(mai22), .C(men22), .Y(z22));
  VOTADOR g23(.A(ori23), .B(mai23), .C(men23), .Y(z23));
  VOTADOR g24(.A(ori24), .B(mai24), .C(men24), .Y(z24));
  VOTADOR g25(.A(ori25), .B(mai25), .C(men25), .Y(z25));
  VOTADOR g26(.A(ori26), .B(mai26), .C(men26), .Y(z26));
  VOTADOR g27(.A(ori27), .B(mai27), .C(men27), .Y(z27));
  VOTADOR g28(.A(ori28), .B(mai28), .C(men28), .Y(z28));
  VOTADOR g29(.A(ori29), .B(mai29), .C(men29), .Y(z29));
  VOTADOR g30(.A(ori30), .B(mai30), .C(men30), .Y(z30));
  VOTADOR g31(.A(ori31), .B(mai31), .C(men31), .Y(z31));
  VOTADOR g32(.A(ori32), .B(mai32), .C(men32), .Y(z32));
  VOTADOR g33(.A(ori33), .B(mai33), .C(men33), .Y(z33));
  VOTADOR g34(.A(ori34), .B(mai34), .C(men34), .Y(z34));
  VOTADOR g35(.A(ori35), .B(mai35), .C(men35), .Y(z35));
  VOTADOR g36(.A(ori36), .B(mai36), .C(men36), .Y(z36));
  VOTADOR g37(.A(ori37), .B(mai37), .C(men37), .Y(z37));
  VOTADOR g38(.A(ori38), .B(mai38), .C(men38), .Y(z38));
  VOTADOR g39(.A(ori39), .B(mai39), .C(men39), .Y(z39));
endmodule