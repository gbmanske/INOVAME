// Benchmark "top" written by ABC on Fri Jun 21 17:49:20 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n537_, new_new_n538_,
    new_new_n539_, new_new_n540_, new_new_n541_, new_new_n542_,
    new_new_n543_, new_new_n544_, new_new_n545_, new_new_n546_,
    new_new_n547_, new_new_n548_, new_new_n549_, new_new_n550_,
    new_new_n551_, new_new_n552_, new_new_n553_, new_new_n554_,
    new_new_n555_, new_new_n556_, new_new_n557_, new_new_n558_,
    new_new_n559_, new_new_n560_, new_new_n561_, new_new_n562_,
    new_new_n563_, new_new_n564_, new_new_n565_, new_new_n566_,
    new_new_n567_, new_new_n568_, new_new_n569_, new_new_n570_,
    new_new_n571_, new_new_n572_, new_new_n573_, new_new_n574_,
    new_new_n575_, new_new_n576_, new_new_n577_, new_new_n578_,
    new_new_n579_, new_new_n580_, new_new_n581_, new_new_n582_,
    new_new_n583_, new_new_n584_, new_new_n586_, new_new_n587_,
    new_new_n588_, new_new_n589_, new_new_n590_, new_new_n591_,
    new_new_n592_, new_new_n593_, new_new_n594_, new_new_n595_,
    new_new_n596_, new_new_n597_, new_new_n598_, new_new_n599_,
    new_new_n600_, new_new_n601_, new_new_n602_, new_new_n603_,
    new_new_n604_, new_new_n605_, new_new_n606_, new_new_n607_,
    new_new_n608_, new_new_n609_, new_new_n610_, new_new_n611_,
    new_new_n612_, new_new_n613_, new_new_n614_, new_new_n615_,
    new_new_n616_, new_new_n617_, new_new_n618_, new_new_n619_,
    new_new_n620_, new_new_n621_, new_new_n622_, new_new_n623_,
    new_new_n624_, new_new_n625_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n771_,
    new_new_n772_, new_new_n773_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  OAI210     g033(.A0(new_new_n55_), .A1(new_new_n52_), .B0(new_new_n45_), .Y(new_new_n56_));
  NA3        g034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g040(.A(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO2        g062(.A(new_new_n83_), .B(new_new_n63_), .Y(new_new_n85_));
  INV        g063(.A(i_6_), .Y(new_new_n86_));
  NO2        g064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n87_), .Y(new_new_n88_));
  OAI210     g066(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n88_), .Y(new_new_n89_));
  NAi21      g067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n63_), .Y(new_new_n92_));
  NA2        g070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  NO3        g071(.A(new_new_n93_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n94_), .B(new_new_n92_), .Y(new_new_n95_));
  AOI210     g073(.A0(new_new_n95_), .A1(new_new_n89_), .B0(new_new_n80_), .Y(new_new_n96_));
  AN3        g074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n97_));
  NAi21      g075(.An(i_6_), .B(i_11_), .Y(new_new_n98_));
  NO2        g076(.A(i_5_), .B(i_8_), .Y(new_new_n99_));
  NOi21      g077(.An(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  AOI220     g078(.A0(new_new_n100_), .A1(new_new_n62_), .B0(new_new_n97_), .B1(new_new_n32_), .Y(new_new_n101_));
  INV        g079(.A(i_7_), .Y(new_new_n102_));
  NA2        g080(.A(new_new_n46_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(new_new_n86_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  INV        g084(.A(new_new_n106_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n103_), .Y(new_new_n108_));
  NAi21      g086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n90_), .C(new_new_n53_), .Y(new_new_n110_));
  AN2        g088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g090(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n113_));
  NO2        g091(.A(i_8_), .B(new_new_n102_), .Y(new_new_n114_));
  NO3        g092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NAi41      g099(.An(new_new_n110_), .B(new_new_n121_), .C(new_new_n108_), .D(new_new_n101_), .Y(new_new_n122_));
  NOi21      g100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g105(.A(new_new_n127_), .B(new_new_n46_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n129_));
  NAi21      g107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n62_), .Y(new_new_n131_));
  NOi31      g109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g110(.A(i_1_), .B(new_new_n86_), .Y(new_new_n133_));
  NO2        g111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g113(.A0(new_new_n135_), .A1(new_new_n47_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g114(.A0(new_new_n136_), .A1(new_new_n109_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n96_), .Y(new_new_n138_));
  NA3        g116(.A(new_new_n138_), .B(new_new_n79_), .C(new_new_n56_), .Y(ori2));
  NO2        g117(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n140_));
  NA2        g118(.A(new_new_n772_), .B(new_new_n140_), .Y(new_new_n141_));
  NA4        g119(.A(new_new_n141_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(ori0));
  AN2        g120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  AN2        g128(.A(new_new_n145_), .B(new_new_n83_), .Y(new_new_n151_));
  NA2        g129(.A(i_1_), .B(i_5_), .Y(new_new_n152_));
  OR2        g130(.A(i_0_), .B(i_1_), .Y(new_new_n153_));
  NO3        g131(.A(new_new_n153_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n154_));
  NAi32      g132(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n155_));
  NAi21      g133(.An(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  NOi21      g134(.An(i_4_), .B(i_10_), .Y(new_new_n157_));
  NA2        g135(.A(new_new_n157_), .B(new_new_n40_), .Y(new_new_n158_));
  NOi21      g136(.An(i_4_), .B(i_9_), .Y(new_new_n159_));
  NOi21      g137(.An(i_11_), .B(i_13_), .Y(new_new_n160_));
  NA2        g138(.A(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NAi21      g139(.An(i_12_), .B(i_11_), .Y(new_new_n162_));
  NO2        g140(.A(new_new_n162_), .B(i_13_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n164_));
  NO2        g142(.A(new_new_n73_), .B(i_5_), .Y(new_new_n165_));
  NO2        g143(.A(i_13_), .B(i_10_), .Y(new_new_n166_));
  NA3        g144(.A(new_new_n166_), .B(new_new_n165_), .C(new_new_n44_), .Y(new_new_n167_));
  NO2        g145(.A(i_2_), .B(i_1_), .Y(new_new_n168_));
  NAi21      g146(.An(i_4_), .B(i_12_), .Y(new_new_n169_));
  INV        g147(.A(i_8_), .Y(new_new_n170_));
  NO3        g148(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n171_));
  NO2        g149(.A(i_3_), .B(i_8_), .Y(new_new_n172_));
  NO3        g150(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n173_));
  NA3        g151(.A(new_new_n173_), .B(new_new_n172_), .C(new_new_n40_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n104_), .B(new_new_n58_), .Y(new_new_n175_));
  NA2        g153(.A(new_new_n175_), .B(new_new_n153_), .Y(new_new_n176_));
  NO2        g154(.A(i_13_), .B(i_9_), .Y(new_new_n177_));
  NAi21      g155(.An(i_12_), .B(i_3_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n44_), .B(i_5_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n176_), .B(new_new_n174_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(i_7_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n181_), .B(i_4_), .Y(new_new_n182_));
  NAi21      g160(.An(i_12_), .B(i_7_), .Y(new_new_n183_));
  NA3        g161(.A(i_13_), .B(new_new_n170_), .C(i_10_), .Y(new_new_n184_));
  NA2        g162(.A(i_0_), .B(i_5_), .Y(new_new_n185_));
  NAi31      g163(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n36_), .B(i_13_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n189_));
  INV        g167(.A(i_13_), .Y(new_new_n190_));
  NO2        g168(.A(i_12_), .B(new_new_n190_), .Y(new_new_n191_));
  NO2        g169(.A(i_12_), .B(new_new_n37_), .Y(new_new_n192_));
  OR2        g170(.A(i_8_), .B(i_7_), .Y(new_new_n193_));
  INV        g171(.A(i_12_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n44_), .B(new_new_n194_), .Y(new_new_n195_));
  NO3        g173(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n196_));
  NA2        g174(.A(i_2_), .B(i_1_), .Y(new_new_n197_));
  NO3        g175(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n198_));
  NAi21      g176(.An(i_4_), .B(i_3_), .Y(new_new_n199_));
  NO2        g177(.A(i_0_), .B(i_6_), .Y(new_new_n200_));
  NOi41      g178(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n201_), .B(new_new_n200_), .Y(new_new_n202_));
  NO2        g180(.A(i_11_), .B(new_new_n190_), .Y(new_new_n203_));
  NOi21      g181(.An(i_1_), .B(i_6_), .Y(new_new_n204_));
  NAi21      g182(.An(i_3_), .B(i_7_), .Y(new_new_n205_));
  NA2        g183(.A(new_new_n194_), .B(i_9_), .Y(new_new_n206_));
  OR4        g184(.A(new_new_n206_), .B(new_new_n205_), .C(new_new_n204_), .D(new_new_n165_), .Y(new_new_n207_));
  NA2        g185(.A(new_new_n73_), .B(i_5_), .Y(new_new_n208_));
  NA2        g186(.A(i_3_), .B(i_9_), .Y(new_new_n209_));
  NAi21      g187(.An(i_7_), .B(i_10_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n210_), .B(new_new_n209_), .Y(new_new_n211_));
  NA3        g189(.A(new_new_n211_), .B(new_new_n208_), .C(new_new_n64_), .Y(new_new_n212_));
  NA2        g190(.A(new_new_n212_), .B(new_new_n207_), .Y(new_new_n213_));
  INV        g191(.A(new_new_n144_), .Y(new_new_n214_));
  NA2        g192(.A(new_new_n194_), .B(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n215_), .B(new_new_n75_), .Y(new_new_n216_));
  AOI220     g194(.A0(new_new_n216_), .A1(new_new_n214_), .B0(new_new_n213_), .B1(new_new_n203_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n193_), .B(new_new_n37_), .Y(new_new_n218_));
  NA2        g196(.A(i_12_), .B(i_6_), .Y(new_new_n219_));
  OR2        g197(.A(i_13_), .B(i_9_), .Y(new_new_n220_));
  NO3        g198(.A(new_new_n220_), .B(new_new_n219_), .C(new_new_n48_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n199_), .B(i_2_), .Y(new_new_n222_));
  NA3        g200(.A(new_new_n222_), .B(new_new_n221_), .C(new_new_n44_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n203_), .B(i_9_), .Y(new_new_n224_));
  NA3        g202(.A(new_new_n208_), .B(new_new_n153_), .C(new_new_n64_), .Y(new_new_n225_));
  OAI210     g203(.A0(new_new_n225_), .A1(new_new_n224_), .B0(new_new_n223_), .Y(new_new_n226_));
  NO3        g204(.A(i_11_), .B(new_new_n190_), .C(new_new_n25_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n205_), .B(i_8_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n226_), .B(new_new_n218_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n217_), .Y(new_new_n230_));
  NO3        g208(.A(i_12_), .B(new_new_n190_), .C(new_new_n37_), .Y(new_new_n231_));
  NO2        g209(.A(i_2_), .B(new_new_n102_), .Y(new_new_n232_));
  AN2        g210(.A(i_3_), .B(i_10_), .Y(new_new_n233_));
  NO2        g211(.A(i_5_), .B(new_new_n37_), .Y(new_new_n234_));
  NO2        g212(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n230_), .B(new_new_n182_), .Y(new_new_n236_));
  NO3        g214(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n237_));
  NO2        g215(.A(i_2_), .B(i_3_), .Y(new_new_n238_));
  OR2        g216(.A(i_0_), .B(i_5_), .Y(new_new_n239_));
  NO2        g217(.A(i_12_), .B(i_10_), .Y(new_new_n240_));
  NOi21      g218(.An(i_5_), .B(i_0_), .Y(new_new_n241_));
  NA4        g219(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n242_));
  NO2        g220(.A(i_1_), .B(i_7_), .Y(new_new_n243_));
  NOi21      g221(.An(new_new_n152_), .B(new_new_n105_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n244_), .B(new_new_n126_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n245_), .B(i_3_), .Y(new_new_n246_));
  NO2        g224(.A(new_new_n170_), .B(i_9_), .Y(new_new_n247_));
  NA3        g225(.A(new_new_n247_), .B(new_new_n175_), .C(new_new_n153_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n248_), .B(new_new_n46_), .Y(new_new_n249_));
  INV        g227(.A(new_new_n249_), .Y(new_new_n250_));
  AOI210     g228(.A0(new_new_n250_), .A1(new_new_n246_), .B0(new_new_n158_), .Y(new_new_n251_));
  INV        g229(.A(new_new_n251_), .Y(new_new_n252_));
  NOi32      g230(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n253_));
  INV        g231(.A(new_new_n253_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n186_), .B(new_new_n155_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n155_), .B(new_new_n153_), .Y(new_new_n256_));
  NOi32      g234(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n257_));
  NAi21      g235(.An(i_6_), .B(i_1_), .Y(new_new_n258_));
  NA3        g236(.A(new_new_n258_), .B(new_new_n257_), .C(new_new_n46_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n259_), .B(i_0_), .Y(new_new_n260_));
  OR3        g238(.A(new_new_n260_), .B(new_new_n256_), .C(new_new_n255_), .Y(new_new_n261_));
  NO2        g239(.A(i_1_), .B(new_new_n102_), .Y(new_new_n262_));
  NAi21      g240(.An(i_3_), .B(i_4_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n263_), .B(i_9_), .Y(new_new_n264_));
  AN2        g242(.A(i_6_), .B(i_7_), .Y(new_new_n265_));
  OAI210     g243(.A0(new_new_n265_), .A1(new_new_n262_), .B0(new_new_n264_), .Y(new_new_n266_));
  NA2        g244(.A(i_2_), .B(i_7_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n263_), .B(i_10_), .Y(new_new_n268_));
  NA3        g246(.A(new_new_n268_), .B(new_new_n267_), .C(new_new_n200_), .Y(new_new_n269_));
  AOI210     g247(.A0(new_new_n269_), .A1(new_new_n266_), .B0(new_new_n165_), .Y(new_new_n270_));
  AOI210     g248(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n271_));
  OAI210     g249(.A0(new_new_n271_), .A1(new_new_n168_), .B0(new_new_n268_), .Y(new_new_n272_));
  AOI220     g250(.A0(new_new_n268_), .A1(new_new_n243_), .B0(new_new_n196_), .B1(new_new_n168_), .Y(new_new_n273_));
  AOI210     g251(.A0(new_new_n273_), .A1(new_new_n272_), .B0(i_5_), .Y(new_new_n274_));
  NO4        g252(.A(new_new_n274_), .B(new_new_n270_), .C(new_new_n261_), .D(new_new_n773_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n275_), .B(new_new_n254_), .Y(new_new_n276_));
  AN2        g254(.A(i_12_), .B(i_5_), .Y(new_new_n277_));
  NO2        g255(.A(i_11_), .B(i_6_), .Y(new_new_n278_));
  NO2        g256(.A(i_5_), .B(i_10_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n280_));
  NO3        g258(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n281_));
  NO2        g259(.A(i_11_), .B(i_12_), .Y(new_new_n282_));
  NAi21      g260(.An(i_13_), .B(i_0_), .Y(new_new_n283_));
  NO3        g261(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n284_));
  NO2        g262(.A(i_0_), .B(i_11_), .Y(new_new_n285_));
  AN2        g263(.A(i_1_), .B(i_6_), .Y(new_new_n286_));
  NOi21      g264(.An(i_2_), .B(i_12_), .Y(new_new_n287_));
  NAi21      g265(.An(i_9_), .B(i_4_), .Y(new_new_n288_));
  OR2        g266(.A(i_13_), .B(i_10_), .Y(new_new_n289_));
  NO3        g267(.A(new_new_n289_), .B(new_new_n119_), .C(new_new_n288_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n161_), .B(new_new_n125_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n231_), .B(new_new_n292_), .Y(new_new_n293_));
  NO2        g271(.A(new_new_n293_), .B(new_new_n244_), .Y(new_new_n294_));
  INV        g272(.A(new_new_n294_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n295_), .B(new_new_n26_), .Y(new_new_n296_));
  NA2        g274(.A(new_new_n170_), .B(i_10_), .Y(new_new_n297_));
  NA3        g275(.A(new_new_n208_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n298_), .B(new_new_n297_), .Y(new_new_n299_));
  INV        g277(.A(new_new_n299_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n300_), .B(new_new_n224_), .Y(new_new_n301_));
  NO3        g279(.A(new_new_n301_), .B(new_new_n296_), .C(new_new_n276_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n73_), .B(i_13_), .Y(new_new_n303_));
  NO2        g281(.A(i_10_), .B(i_9_), .Y(new_new_n304_));
  NAi21      g282(.An(i_12_), .B(i_8_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n305_), .B(i_3_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n235_), .B(i_0_), .Y(new_new_n307_));
  NO3        g285(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n219_), .B(new_new_n98_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n309_), .B(new_new_n308_), .Y(new_new_n310_));
  NA2        g288(.A(i_8_), .B(i_9_), .Y(new_new_n311_));
  AOI210     g289(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n312_));
  OR2        g290(.A(new_new_n312_), .B(new_new_n311_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n231_), .B(new_new_n175_), .Y(new_new_n314_));
  OAI220     g292(.A0(new_new_n314_), .A1(new_new_n313_), .B0(new_new_n310_), .B1(new_new_n307_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n203_), .B(new_new_n234_), .Y(new_new_n316_));
  NO3        g294(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n317_));
  INV        g295(.A(new_new_n317_), .Y(new_new_n318_));
  NA3        g296(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n319_));
  NA4        g297(.A(new_new_n146_), .B(new_new_n117_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n320_));
  OAI220     g298(.A0(new_new_n320_), .A1(new_new_n319_), .B0(new_new_n318_), .B1(new_new_n316_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n321_), .B(new_new_n315_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n97_), .B(i_13_), .Y(new_new_n323_));
  NO2        g301(.A(i_2_), .B(i_13_), .Y(new_new_n324_));
  NO3        g302(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n325_));
  NO2        g303(.A(i_6_), .B(i_7_), .Y(new_new_n326_));
  NO2        g304(.A(i_11_), .B(i_1_), .Y(new_new_n327_));
  NOi21      g305(.An(i_2_), .B(i_7_), .Y(new_new_n328_));
  NO2        g306(.A(i_3_), .B(new_new_n170_), .Y(new_new_n329_));
  NO2        g307(.A(i_6_), .B(i_10_), .Y(new_new_n330_));
  NA3        g308(.A(new_new_n201_), .B(new_new_n160_), .C(new_new_n134_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n153_), .B(i_3_), .Y(new_new_n333_));
  NAi31      g311(.An(new_new_n332_), .B(new_new_n333_), .C(new_new_n191_), .Y(new_new_n334_));
  NA3        g312(.A(new_new_n280_), .B(new_new_n164_), .C(new_new_n150_), .Y(new_new_n335_));
  NA3        g313(.A(new_new_n335_), .B(new_new_n334_), .C(new_new_n331_), .Y(new_new_n336_));
  INV        g314(.A(new_new_n336_), .Y(new_new_n337_));
  NA2        g315(.A(new_new_n308_), .B(new_new_n277_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n317_), .B(new_new_n279_), .Y(new_new_n339_));
  NAi21      g317(.An(new_new_n184_), .B(new_new_n282_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n243_), .B(new_new_n185_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n27_), .B(i_10_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n237_), .B(new_new_n196_), .Y(new_new_n344_));
  OAI220     g322(.A0(new_new_n344_), .A1(new_new_n298_), .B0(new_new_n343_), .B1(new_new_n323_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n345_), .B(new_new_n342_), .Y(new_new_n346_));
  NA3        g324(.A(new_new_n346_), .B(new_new_n337_), .C(new_new_n322_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n277_), .B(new_new_n190_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n265_), .B(new_new_n257_), .Y(new_new_n349_));
  OR2        g327(.A(new_new_n348_), .B(new_new_n349_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n36_), .B(i_8_), .Y(new_new_n351_));
  AOI210     g329(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n290_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n352_), .B(new_new_n350_), .Y(new_new_n353_));
  INV        g331(.A(new_new_n353_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n208_), .B(new_new_n64_), .Y(new_new_n355_));
  OAI210     g333(.A0(i_8_), .A1(new_new_n355_), .B0(new_new_n136_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n356_), .B(new_new_n291_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n357_), .B(new_new_n354_), .Y(new_new_n358_));
  NO2        g336(.A(i_12_), .B(new_new_n170_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n44_), .B(i_10_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n360_), .B(i_6_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n153_), .B(i_5_), .Y(new_new_n362_));
  NA3        g340(.A(new_new_n185_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n231_), .B(new_new_n84_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n363_), .B(new_new_n364_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n189_), .B(new_new_n188_), .Y(new_new_n366_));
  NA2        g344(.A(new_new_n304_), .B(new_new_n187_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n366_), .B(new_new_n367_), .Y(new_new_n368_));
  AOI210     g346(.A0(new_new_n258_), .A1(new_new_n46_), .B0(new_new_n262_), .Y(new_new_n369_));
  NA2        g347(.A(i_0_), .B(new_new_n48_), .Y(new_new_n370_));
  NA3        g348(.A(new_new_n359_), .B(new_new_n227_), .C(new_new_n370_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n369_), .B(new_new_n371_), .Y(new_new_n372_));
  NO3        g350(.A(new_new_n372_), .B(new_new_n368_), .C(new_new_n365_), .Y(new_new_n373_));
  NO4        g351(.A(new_new_n204_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n374_));
  NO3        g352(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n289_), .B(i_1_), .Y(new_new_n376_));
  NOi31      g354(.An(new_new_n376_), .B(new_new_n309_), .C(new_new_n73_), .Y(new_new_n377_));
  NOi21      g355(.An(i_10_), .B(i_6_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n379_));
  AOI220     g357(.A0(new_new_n231_), .A1(new_new_n379_), .B0(new_new_n227_), .B1(new_new_n378_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n380_), .B(new_new_n307_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n382_));
  NOi31      g360(.An(new_new_n147_), .B(i_10_), .C(new_new_n242_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n381_), .Y(new_new_n384_));
  INV        g362(.A(new_new_n238_), .Y(new_new_n385_));
  NO2        g363(.A(i_12_), .B(new_new_n86_), .Y(new_new_n386_));
  NA3        g364(.A(new_new_n386_), .B(new_new_n227_), .C(new_new_n370_), .Y(new_new_n387_));
  NA3        g365(.A(new_new_n278_), .B(new_new_n231_), .C(new_new_n185_), .Y(new_new_n388_));
  AOI210     g366(.A0(new_new_n388_), .A1(new_new_n387_), .B0(new_new_n385_), .Y(new_new_n389_));
  OR2        g367(.A(i_2_), .B(i_5_), .Y(new_new_n390_));
  OR2        g368(.A(new_new_n390_), .B(new_new_n286_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n267_), .B(new_new_n200_), .Y(new_new_n392_));
  AOI210     g370(.A0(new_new_n392_), .A1(new_new_n391_), .B0(new_new_n340_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n393_), .B(new_new_n389_), .Y(new_new_n394_));
  NA3        g372(.A(new_new_n394_), .B(new_new_n384_), .C(new_new_n373_), .Y(new_new_n395_));
  NO3        g373(.A(new_new_n395_), .B(new_new_n358_), .C(new_new_n347_), .Y(new_new_n396_));
  NA4        g374(.A(new_new_n396_), .B(new_new_n302_), .C(new_new_n252_), .D(new_new_n236_), .Y(ori7));
  NO2        g375(.A(new_new_n93_), .B(new_new_n54_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n330_), .B(new_new_n84_), .Y(new_new_n399_));
  NA2        g377(.A(i_11_), .B(new_new_n170_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n145_), .B(new_new_n400_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n401_), .B(new_new_n399_), .Y(new_new_n402_));
  NA3        g380(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n194_), .B(i_4_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n404_), .B(i_8_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n106_), .B(new_new_n403_), .Y(new_new_n406_));
  NA2        g384(.A(i_2_), .B(new_new_n86_), .Y(new_new_n407_));
  OAI210     g385(.A0(new_new_n87_), .A1(new_new_n172_), .B0(new_new_n173_), .Y(new_new_n408_));
  NO2        g386(.A(i_7_), .B(new_new_n37_), .Y(new_new_n409_));
  NA2        g387(.A(i_4_), .B(i_8_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n410_), .A1(new_new_n233_), .B0(new_new_n409_), .Y(new_new_n411_));
  OAI220     g389(.A0(new_new_n411_), .A1(new_new_n407_), .B0(new_new_n408_), .B1(i_13_), .Y(new_new_n412_));
  NO4        g390(.A(new_new_n412_), .B(new_new_n406_), .C(new_new_n402_), .D(new_new_n398_), .Y(new_new_n413_));
  AOI210     g391(.A0(new_new_n130_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n414_));
  AOI210     g392(.A0(new_new_n414_), .A1(new_new_n194_), .B0(new_new_n157_), .Y(new_new_n415_));
  OR2        g393(.A(i_6_), .B(i_10_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n416_), .B(new_new_n23_), .Y(new_new_n417_));
  OR3        g395(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n418_));
  INV        g396(.A(new_new_n171_), .Y(new_new_n419_));
  INV        g397(.A(new_new_n417_), .Y(new_new_n420_));
  OA220      g398(.A0(new_new_n420_), .A1(new_new_n385_), .B0(new_new_n415_), .B1(new_new_n220_), .Y(new_new_n421_));
  AOI210     g399(.A0(new_new_n421_), .A1(new_new_n413_), .B0(new_new_n63_), .Y(new_new_n422_));
  NOi21      g400(.An(i_11_), .B(i_7_), .Y(new_new_n423_));
  AO210      g401(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n424_), .B(new_new_n423_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n425_), .B(new_new_n177_), .Y(new_new_n426_));
  NA3        g404(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n427_));
  NO2        g405(.A(new_new_n426_), .B(new_new_n63_), .Y(new_new_n428_));
  OR2        g406(.A(new_new_n273_), .B(new_new_n41_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n210_), .B(new_new_n178_), .C(new_new_n400_), .Y(new_new_n430_));
  OAI210     g408(.A0(new_new_n430_), .A1(new_new_n191_), .B0(new_new_n63_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n287_), .B(new_new_n31_), .Y(new_new_n432_));
  OR2        g410(.A(new_new_n178_), .B(new_new_n109_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n433_), .B(new_new_n432_), .Y(new_new_n434_));
  NO2        g412(.A(i_1_), .B(i_4_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n435_), .B(new_new_n434_), .Y(new_new_n436_));
  NO2        g414(.A(i_1_), .B(i_12_), .Y(new_new_n437_));
  NA3        g415(.A(new_new_n437_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n438_));
  BUFFER     g416(.A(new_new_n438_), .Y(new_new_n439_));
  NA4        g417(.A(new_new_n439_), .B(new_new_n436_), .C(new_new_n431_), .D(new_new_n429_), .Y(new_new_n440_));
  OAI210     g418(.A0(new_new_n440_), .A1(new_new_n428_), .B0(i_6_), .Y(new_new_n441_));
  NO2        g419(.A(new_new_n427_), .B(new_new_n109_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n442_), .B(new_new_n386_), .Y(new_new_n443_));
  NO2        g421(.A(i_6_), .B(i_11_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n443_), .B(new_new_n310_), .Y(new_new_n445_));
  NO3        g423(.A(new_new_n416_), .B(new_new_n193_), .C(new_new_n23_), .Y(new_new_n446_));
  AOI210     g424(.A0(i_1_), .A1(new_new_n211_), .B0(new_new_n446_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n447_), .B(new_new_n44_), .Y(new_new_n448_));
  INV        g426(.A(i_2_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n140_), .B(i_9_), .Y(new_new_n450_));
  NA3        g428(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n46_), .B(i_1_), .Y(new_new_n452_));
  NA3        g430(.A(new_new_n452_), .B(new_new_n219_), .C(new_new_n44_), .Y(new_new_n453_));
  OAI220     g431(.A0(new_new_n453_), .A1(new_new_n451_), .B0(new_new_n450_), .B1(new_new_n449_), .Y(new_new_n454_));
  AOI210     g432(.A0(new_new_n327_), .A1(new_new_n292_), .B0(new_new_n198_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n455_), .B(new_new_n407_), .Y(new_new_n456_));
  NO2        g434(.A(i_11_), .B(new_new_n37_), .Y(new_new_n457_));
  OR2        g435(.A(new_new_n456_), .B(new_new_n454_), .Y(new_new_n458_));
  NO3        g436(.A(new_new_n458_), .B(new_new_n448_), .C(new_new_n445_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n194_), .B(new_new_n102_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n460_), .B(new_new_n423_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n461_), .B(i_1_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n418_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n288_), .B(new_new_n86_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n463_), .B(new_new_n46_), .Y(new_new_n465_));
  NA2        g443(.A(i_3_), .B(new_new_n170_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n466_), .B(new_new_n116_), .Y(new_new_n467_));
  AN2        g445(.A(new_new_n467_), .B(new_new_n361_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n193_), .B(new_new_n44_), .Y(new_new_n469_));
  NO3        g447(.A(new_new_n469_), .B(new_new_n235_), .C(new_new_n195_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n471_), .B(i_6_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n86_), .B(i_9_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n473_), .B(new_new_n63_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n437_), .Y(new_new_n475_));
  NO4        g453(.A(new_new_n475_), .B(new_new_n472_), .C(new_new_n470_), .D(i_4_), .Y(new_new_n476_));
  NA2        g454(.A(i_1_), .B(i_3_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n311_), .B(new_new_n93_), .Y(new_new_n478_));
  AOI210     g456(.A0(new_new_n469_), .A1(new_new_n378_), .B0(new_new_n478_), .Y(new_new_n479_));
  NO2        g457(.A(new_new_n479_), .B(new_new_n477_), .Y(new_new_n480_));
  NO3        g458(.A(new_new_n480_), .B(new_new_n476_), .C(new_new_n468_), .Y(new_new_n481_));
  NA4        g459(.A(new_new_n481_), .B(new_new_n465_), .C(new_new_n459_), .D(new_new_n441_), .Y(new_new_n482_));
  AN2        g460(.A(new_new_n201_), .B(new_new_n86_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n484_));
  NO3        g462(.A(new_new_n328_), .B(new_new_n410_), .C(new_new_n86_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n485_), .B(new_new_n25_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(new_new_n484_), .Y(new_new_n487_));
  OAI210     g465(.A0(new_new_n487_), .A1(new_new_n483_), .B0(i_1_), .Y(new_new_n488_));
  AOI210     g466(.A0(new_new_n219_), .A1(new_new_n98_), .B0(i_1_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n263_), .B(i_2_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(new_new_n489_), .Y(new_new_n491_));
  AOI210     g469(.A0(new_new_n491_), .A1(new_new_n488_), .B0(i_13_), .Y(new_new_n492_));
  OR2        g470(.A(i_11_), .B(i_7_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n54_), .B(i_12_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n328_), .B(new_new_n24_), .Y(new_new_n495_));
  AOI220     g473(.A0(new_new_n495_), .A1(new_new_n464_), .B0(new_new_n201_), .B1(new_new_n133_), .Y(new_new_n496_));
  OAI220     g474(.A0(new_new_n496_), .A1(new_new_n41_), .B0(new_new_n771_), .B1(new_new_n93_), .Y(new_new_n497_));
  INV        g475(.A(new_new_n497_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n116_), .Y(new_new_n499_));
  AOI220     g477(.A0(new_new_n499_), .A1(new_new_n72_), .B0(new_new_n278_), .B1(new_new_n452_), .Y(new_new_n500_));
  NO2        g478(.A(new_new_n500_), .B(new_new_n199_), .Y(new_new_n501_));
  AOI210     g479(.A0(new_new_n305_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n502_));
  NOi31      g480(.An(new_new_n502_), .B(new_new_n399_), .C(new_new_n44_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n129_), .B(i_13_), .Y(new_new_n504_));
  NO2        g482(.A(new_new_n451_), .B(new_new_n116_), .Y(new_new_n505_));
  INV        g483(.A(new_new_n505_), .Y(new_new_n506_));
  OAI220     g484(.A0(new_new_n506_), .A1(new_new_n71_), .B0(new_new_n504_), .B1(new_new_n489_), .Y(new_new_n507_));
  NO3        g485(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n102_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n26_), .B(new_new_n170_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n509_), .B(i_7_), .Y(new_new_n510_));
  NO3        g488(.A(new_new_n328_), .B(new_new_n194_), .C(new_new_n86_), .Y(new_new_n511_));
  AOI210     g489(.A0(new_new_n511_), .A1(new_new_n510_), .B0(new_new_n508_), .Y(new_new_n512_));
  AOI220     g490(.A0(new_new_n278_), .A1(new_new_n452_), .B0(new_new_n92_), .B1(new_new_n103_), .Y(new_new_n513_));
  OAI220     g491(.A0(new_new_n513_), .A1(new_new_n405_), .B0(new_new_n512_), .B1(new_new_n419_), .Y(new_new_n514_));
  NO4        g492(.A(new_new_n514_), .B(new_new_n507_), .C(new_new_n503_), .D(new_new_n501_), .Y(new_new_n515_));
  OR2        g493(.A(i_11_), .B(i_6_), .Y(new_new_n516_));
  NA3        g494(.A(new_new_n404_), .B(new_new_n509_), .C(i_7_), .Y(new_new_n517_));
  AOI210     g495(.A0(new_new_n517_), .A1(new_new_n506_), .B0(new_new_n516_), .Y(new_new_n518_));
  NA3        g496(.A(new_new_n287_), .B(new_new_n409_), .C(new_new_n98_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n444_), .B(i_13_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n103_), .B(new_new_n509_), .Y(new_new_n521_));
  NAi21      g499(.An(i_11_), .B(i_12_), .Y(new_new_n522_));
  NOi41      g500(.An(new_new_n112_), .B(new_new_n522_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n523_));
  NO3        g501(.A(new_new_n328_), .B(new_new_n386_), .C(new_new_n410_), .Y(new_new_n524_));
  AOI220     g502(.A0(new_new_n524_), .A1(new_new_n237_), .B0(new_new_n523_), .B1(new_new_n521_), .Y(new_new_n525_));
  NA3        g503(.A(new_new_n525_), .B(new_new_n520_), .C(new_new_n519_), .Y(new_new_n526_));
  OAI210     g504(.A0(new_new_n526_), .A1(new_new_n518_), .B0(new_new_n63_), .Y(new_new_n527_));
  NO2        g505(.A(i_2_), .B(i_12_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n262_), .B(new_new_n528_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n264_), .B(new_new_n262_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n130_), .B(i_2_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n531_), .B(new_new_n437_), .Y(new_new_n532_));
  NA3        g510(.A(new_new_n532_), .B(new_new_n530_), .C(new_new_n529_), .Y(new_new_n533_));
  NA3        g511(.A(new_new_n533_), .B(new_new_n45_), .C(new_new_n190_), .Y(new_new_n534_));
  NA4        g512(.A(new_new_n534_), .B(new_new_n527_), .C(new_new_n515_), .D(new_new_n498_), .Y(new_new_n535_));
  OR4        g513(.A(new_new_n535_), .B(new_new_n492_), .C(new_new_n482_), .D(new_new_n422_), .Y(ori5));
  NA2        g514(.A(new_new_n461_), .B(new_new_n222_), .Y(new_new_n537_));
  AN2        g515(.A(new_new_n24_), .B(i_10_), .Y(new_new_n538_));
  NA3        g516(.A(new_new_n538_), .B(new_new_n528_), .C(new_new_n109_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n405_), .B(i_11_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n87_), .B(new_new_n540_), .Y(new_new_n541_));
  NA3        g519(.A(new_new_n541_), .B(new_new_n539_), .C(new_new_n537_), .Y(new_new_n542_));
  NO3        g520(.A(i_11_), .B(new_new_n194_), .C(i_13_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n544_));
  NA2        g522(.A(i_12_), .B(i_8_), .Y(new_new_n545_));
  OAI210     g523(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n545_), .Y(new_new_n546_));
  INV        g524(.A(new_new_n304_), .Y(new_new_n547_));
  AOI220     g525(.A0(new_new_n238_), .A1(new_new_n382_), .B0(new_new_n546_), .B1(new_new_n544_), .Y(new_new_n548_));
  INV        g526(.A(new_new_n548_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n549_), .B(new_new_n542_), .Y(new_new_n550_));
  INV        g528(.A(new_new_n160_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n201_), .Y(new_new_n552_));
  OAI210     g530(.A0(new_new_n490_), .A1(new_new_n306_), .B0(new_new_n112_), .Y(new_new_n553_));
  AOI210     g531(.A0(new_new_n553_), .A1(new_new_n552_), .B0(new_new_n551_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n311_), .B(new_new_n26_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n555_), .B(new_new_n292_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n556_), .B(i_2_), .Y(new_new_n557_));
  INV        g535(.A(new_new_n557_), .Y(new_new_n558_));
  AOI210     g536(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n289_), .Y(new_new_n559_));
  AOI210     g537(.A0(new_new_n559_), .A1(new_new_n558_), .B0(new_new_n554_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n169_), .B(new_new_n127_), .Y(new_new_n561_));
  OAI210     g539(.A0(new_new_n561_), .A1(new_new_n544_), .B0(i_2_), .Y(new_new_n562_));
  INV        g540(.A(new_new_n161_), .Y(new_new_n563_));
  NO3        g541(.A(new_new_n424_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n563_), .A1(new_new_n87_), .B0(new_new_n564_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n565_), .A1(new_new_n562_), .B0(new_new_n170_), .Y(new_new_n566_));
  OA210      g544(.A0(new_new_n425_), .A1(new_new_n128_), .B0(i_13_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n171_), .B(new_new_n172_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n151_), .B(new_new_n400_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n569_), .A1(new_new_n568_), .B0(new_new_n267_), .Y(new_new_n570_));
  AOI210     g548(.A0(new_new_n178_), .A1(new_new_n149_), .B0(new_new_n351_), .Y(new_new_n571_));
  OAI210     g549(.A0(new_new_n571_), .A1(new_new_n191_), .B0(new_new_n292_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n103_), .B(new_new_n44_), .Y(new_new_n573_));
  INV        g551(.A(new_new_n232_), .Y(new_new_n574_));
  NA4        g552(.A(new_new_n574_), .B(new_new_n233_), .C(new_new_n126_), .D(new_new_n42_), .Y(new_new_n575_));
  OAI210     g553(.A0(new_new_n575_), .A1(new_new_n573_), .B0(new_new_n572_), .Y(new_new_n576_));
  NO4        g554(.A(new_new_n576_), .B(new_new_n570_), .C(new_new_n567_), .D(new_new_n566_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n382_), .B(new_new_n28_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n543_), .B(new_new_n228_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n579_), .B(new_new_n578_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n62_), .B(i_12_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n581_), .B(new_new_n128_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n582_), .B(new_new_n400_), .Y(new_new_n583_));
  AOI220     g561(.A0(new_new_n583_), .A1(new_new_n36_), .B0(new_new_n580_), .B1(new_new_n46_), .Y(new_new_n584_));
  NA4        g562(.A(new_new_n584_), .B(new_new_n577_), .C(new_new_n560_), .D(new_new_n550_), .Y(ori6));
  NA4        g563(.A(new_new_n279_), .B(new_new_n329_), .C(new_new_n71_), .D(new_new_n102_), .Y(new_new_n586_));
  INV        g564(.A(new_new_n586_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n186_), .B(new_new_n332_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n587_), .B(new_new_n241_), .Y(new_new_n589_));
  OR2        g567(.A(new_new_n589_), .B(i_12_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n386_), .B(new_new_n63_), .Y(new_new_n591_));
  INV        g569(.A(new_new_n591_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n592_), .B(new_new_n73_), .Y(new_new_n593_));
  INV        g571(.A(new_new_n240_), .Y(new_new_n594_));
  NA2        g572(.A(new_new_n75_), .B(new_new_n133_), .Y(new_new_n595_));
  INV        g573(.A(new_new_n126_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n596_), .B(new_new_n46_), .Y(new_new_n597_));
  AOI210     g575(.A0(new_new_n597_), .A1(new_new_n595_), .B0(new_new_n594_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n204_), .B(i_9_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n599_), .B(new_new_n581_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n600_), .A1(new_new_n349_), .B0(new_new_n165_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n32_), .B(i_11_), .Y(new_new_n602_));
  NAi32      g580(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n516_), .B(new_new_n603_), .Y(new_new_n604_));
  OR3        g582(.A(new_new_n604_), .B(new_new_n601_), .C(new_new_n598_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n493_), .B(i_2_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n607_), .B(new_new_n286_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n608_), .B(new_new_n606_), .Y(new_new_n609_));
  OR2        g587(.A(new_new_n425_), .B(new_new_n306_), .Y(new_new_n610_));
  NA3        g588(.A(new_new_n610_), .B(new_new_n148_), .C(new_new_n69_), .Y(new_new_n611_));
  AO210      g589(.A0(new_new_n339_), .A1(new_new_n547_), .B0(new_new_n36_), .Y(new_new_n612_));
  NA3        g590(.A(new_new_n612_), .B(new_new_n611_), .C(new_new_n609_), .Y(new_new_n613_));
  NO2        g591(.A(i_6_), .B(i_11_), .Y(new_new_n614_));
  AOI220     g592(.A0(new_new_n614_), .A1(new_new_n375_), .B0(new_new_n588_), .B1(new_new_n510_), .Y(new_new_n615_));
  NA3        g593(.A(new_new_n267_), .B(new_new_n196_), .C(new_new_n148_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n281_), .B(new_new_n70_), .Y(new_new_n617_));
  NA4        g595(.A(new_new_n617_), .B(new_new_n616_), .C(new_new_n615_), .D(new_new_n408_), .Y(new_new_n618_));
  AOI210     g596(.A0(new_new_n306_), .A1(new_new_n304_), .B0(new_new_n374_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n416_), .B(new_new_n103_), .Y(new_new_n620_));
  OAI210     g598(.A0(new_new_n620_), .A1(new_new_n113_), .B0(new_new_n285_), .Y(new_new_n621_));
  INV        g599(.A(new_new_n391_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n622_), .B(new_new_n240_), .C(i_7_), .Y(new_new_n623_));
  NA3        g601(.A(new_new_n623_), .B(new_new_n621_), .C(new_new_n619_), .Y(new_new_n624_));
  NO4        g602(.A(new_new_n624_), .B(new_new_n618_), .C(new_new_n613_), .D(new_new_n605_), .Y(new_new_n625_));
  NA4        g603(.A(new_new_n625_), .B(new_new_n593_), .C(new_new_n590_), .D(new_new_n275_), .Y(ori3));
  NA2        g604(.A(i_12_), .B(i_10_), .Y(new_new_n627_));
  NO2        g605(.A(i_11_), .B(new_new_n194_), .Y(new_new_n628_));
  NA3        g606(.A(new_new_n616_), .B(new_new_n408_), .C(new_new_n266_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n629_), .B(new_new_n40_), .Y(new_new_n630_));
  NOi21      g608(.An(new_new_n97_), .B(new_new_n556_), .Y(new_new_n631_));
  NO3        g609(.A(new_new_n433_), .B(new_new_n311_), .C(new_new_n133_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n287_), .B(new_new_n45_), .Y(new_new_n633_));
  AN2        g611(.A(new_new_n309_), .B(new_new_n55_), .Y(new_new_n634_));
  NO3        g612(.A(new_new_n634_), .B(new_new_n632_), .C(new_new_n631_), .Y(new_new_n635_));
  AOI210     g613(.A0(new_new_n635_), .A1(new_new_n630_), .B0(new_new_n48_), .Y(new_new_n636_));
  NO4        g614(.A(new_new_n271_), .B(new_new_n277_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n165_), .B(new_new_n378_), .Y(new_new_n638_));
  NOi31      g616(.An(new_new_n638_), .B(new_new_n637_), .C(new_new_n39_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n639_), .B(new_new_n63_), .Y(new_new_n640_));
  NOi21      g618(.An(i_5_), .B(i_9_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(new_new_n303_), .Y(new_new_n642_));
  BUFFER     g620(.A(new_new_n219_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n643_), .A1(new_new_n327_), .B0(new_new_n485_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n642_), .Y(new_new_n645_));
  NO3        g623(.A(new_new_n645_), .B(new_new_n640_), .C(new_new_n636_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n165_), .B(new_new_n24_), .Y(new_new_n647_));
  INV        g625(.A(new_new_n471_), .Y(new_new_n648_));
  NO2        g626(.A(new_new_n648_), .B(new_new_n647_), .Y(new_new_n649_));
  INV        g627(.A(new_new_n649_), .Y(new_new_n650_));
  NA2        g628(.A(new_new_n379_), .B(i_0_), .Y(new_new_n651_));
  NO4        g629(.A(new_new_n390_), .B(new_new_n183_), .C(new_new_n289_), .D(new_new_n286_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n652_), .B(i_11_), .Y(new_new_n653_));
  NA2        g631(.A(new_new_n543_), .B(new_new_n241_), .Y(new_new_n654_));
  AOI210     g632(.A0(new_new_n330_), .A1(new_new_n87_), .B0(new_new_n58_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n655_), .B(new_new_n654_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n206_), .B(new_new_n152_), .Y(new_new_n657_));
  NA2        g635(.A(i_0_), .B(i_10_), .Y(new_new_n658_));
  INV        g636(.A(new_new_n360_), .Y(new_new_n659_));
  NO4        g637(.A(new_new_n116_), .B(new_new_n58_), .C(new_new_n466_), .D(i_5_), .Y(new_new_n660_));
  AO220      g638(.A0(new_new_n660_), .A1(new_new_n659_), .B0(new_new_n657_), .B1(i_6_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n661_), .B(new_new_n656_), .Y(new_new_n662_));
  NA3        g640(.A(new_new_n662_), .B(new_new_n653_), .C(new_new_n650_), .Y(new_new_n663_));
  NO2        g641(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n664_));
  NA2        g642(.A(i_11_), .B(i_9_), .Y(new_new_n665_));
  NO3        g643(.A(i_12_), .B(new_new_n665_), .C(new_new_n407_), .Y(new_new_n666_));
  AN2        g644(.A(new_new_n666_), .B(new_new_n664_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n280_), .B(new_new_n164_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n668_), .B(new_new_n156_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n665_), .B(new_new_n73_), .Y(new_new_n670_));
  NO2        g648(.A(new_new_n162_), .B(i_0_), .Y(new_new_n671_));
  INV        g649(.A(new_new_n284_), .Y(new_new_n672_));
  NO2        g650(.A(new_new_n672_), .B(new_new_n642_), .Y(new_new_n673_));
  NO3        g651(.A(new_new_n673_), .B(new_new_n669_), .C(new_new_n667_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n457_), .B(new_new_n123_), .Y(new_new_n675_));
  NO2        g653(.A(i_6_), .B(new_new_n675_), .Y(new_new_n676_));
  AOI210     g654(.A0(new_new_n305_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n160_), .B(new_new_n104_), .Y(new_new_n678_));
  NOi32      g656(.An(new_new_n677_), .Bn(new_new_n168_), .C(new_new_n678_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n409_), .B(new_new_n241_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n680_), .B(new_new_n633_), .Y(new_new_n681_));
  NO3        g659(.A(new_new_n681_), .B(new_new_n679_), .C(new_new_n676_), .Y(new_new_n682_));
  NOi21      g660(.An(i_7_), .B(i_5_), .Y(new_new_n683_));
  INV        g661(.A(new_new_n239_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n682_), .B(new_new_n674_), .Y(new_new_n685_));
  NO2        g663(.A(new_new_n627_), .B(new_new_n238_), .Y(new_new_n686_));
  OA210      g664(.A0(new_new_n326_), .A1(new_new_n189_), .B0(new_new_n325_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n686_), .B(new_new_n670_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n670_), .B(new_new_n233_), .Y(new_new_n689_));
  OAI210     g667(.A0(i_2_), .A1(new_new_n167_), .B0(new_new_n689_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n690_), .B(new_new_n326_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n75_), .B(new_new_n545_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n692_), .B(i_11_), .Y(new_new_n693_));
  NO2        g671(.A(new_new_n693_), .B(new_new_n47_), .Y(new_new_n694_));
  NA2        g672(.A(new_new_n495_), .B(new_new_n362_), .Y(new_new_n695_));
  NAi21      g673(.An(i_9_), .B(i_5_), .Y(new_new_n696_));
  NO2        g674(.A(new_new_n696_), .B(new_new_n283_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n403_), .B(new_new_n106_), .Y(new_new_n698_));
  AOI220     g676(.A0(new_new_n698_), .A1(i_0_), .B0(new_new_n697_), .B1(new_new_n425_), .Y(new_new_n699_));
  OAI220     g677(.A0(new_new_n699_), .A1(new_new_n86_), .B0(new_new_n695_), .B1(new_new_n161_), .Y(new_new_n700_));
  NO3        g678(.A(new_new_n700_), .B(new_new_n694_), .C(new_new_n353_), .Y(new_new_n701_));
  NA3        g679(.A(new_new_n701_), .B(new_new_n691_), .C(new_new_n688_), .Y(new_new_n702_));
  NO3        g680(.A(new_new_n702_), .B(new_new_n685_), .C(new_new_n663_), .Y(new_new_n703_));
  NO2        g681(.A(i_0_), .B(new_new_n522_), .Y(new_new_n704_));
  AOI210     g682(.A0(new_new_n591_), .A1(new_new_n484_), .B0(new_new_n678_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n705_), .Y(new_new_n706_));
  OAI210     g684(.A0(new_new_n200_), .A1(i_9_), .B0(new_new_n192_), .Y(new_new_n707_));
  AOI210     g685(.A0(new_new_n707_), .A1(new_new_n651_), .B0(new_new_n152_), .Y(new_new_n708_));
  INV        g686(.A(new_new_n708_), .Y(new_new_n709_));
  NA2        g687(.A(new_new_n709_), .B(new_new_n706_), .Y(new_new_n710_));
  NO3        g688(.A(new_new_n658_), .B(new_new_n641_), .C(new_new_n169_), .Y(new_new_n711_));
  AOI220     g689(.A0(new_new_n711_), .A1(i_11_), .B0(new_new_n377_), .B1(new_new_n75_), .Y(new_new_n712_));
  NO3        g690(.A(new_new_n179_), .B(new_new_n277_), .C(i_0_), .Y(new_new_n713_));
  OAI210     g691(.A0(new_new_n713_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n714_), .B(new_new_n712_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n199_), .B(new_new_n93_), .Y(new_new_n716_));
  AOI210     g694(.A0(new_new_n716_), .A1(new_new_n704_), .B0(new_new_n110_), .Y(new_new_n717_));
  OR2        g695(.A(new_new_n717_), .B(i_5_), .Y(new_new_n718_));
  AOI210     g696(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n162_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n719_), .B(new_new_n687_), .Y(new_new_n720_));
  NO3        g698(.A(new_new_n633_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n338_), .B(new_new_n331_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n722_), .B(new_new_n721_), .Y(new_new_n723_));
  NA3        g701(.A(new_new_n279_), .B(new_new_n160_), .C(new_new_n159_), .Y(new_new_n724_));
  INV        g702(.A(new_new_n724_), .Y(new_new_n725_));
  NO3        g703(.A(new_new_n665_), .B(new_new_n185_), .C(new_new_n169_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n726_), .B(new_new_n725_), .Y(new_new_n727_));
  NA4        g705(.A(new_new_n727_), .B(new_new_n723_), .C(new_new_n720_), .D(new_new_n718_), .Y(new_new_n728_));
  NO2        g706(.A(new_new_n86_), .B(i_5_), .Y(new_new_n729_));
  NA3        g707(.A(new_new_n628_), .B(new_new_n111_), .C(new_new_n126_), .Y(new_new_n730_));
  INV        g708(.A(new_new_n730_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n731_), .B(new_new_n729_), .Y(new_new_n732_));
  NAi21      g710(.An(new_new_n198_), .B(new_new_n199_), .Y(new_new_n733_));
  NO4        g711(.A(new_new_n197_), .B(new_new_n179_), .C(i_0_), .D(i_12_), .Y(new_new_n734_));
  AOI220     g712(.A0(new_new_n734_), .A1(new_new_n733_), .B0(new_new_n587_), .B1(new_new_n163_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n683_), .B(new_new_n324_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n736_), .B(new_new_n474_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n737_), .B(new_new_n671_), .Y(new_new_n738_));
  NA3        g716(.A(new_new_n738_), .B(new_new_n735_), .C(new_new_n732_), .Y(new_new_n739_));
  NO4        g717(.A(new_new_n739_), .B(new_new_n728_), .C(new_new_n715_), .D(new_new_n710_), .Y(new_new_n740_));
  OAI210     g718(.A0(new_new_n606_), .A1(new_new_n602_), .B0(new_new_n37_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n741_), .B(new_new_n415_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n742_), .B(new_new_n177_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n166_), .B(new_new_n168_), .Y(new_new_n744_));
  AO210      g722(.A0(new_new_n493_), .A1(new_new_n33_), .B0(new_new_n744_), .Y(new_new_n745_));
  NAi31      g723(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n746_));
  AOI210     g724(.A0(new_new_n119_), .A1(new_new_n70_), .B0(new_new_n746_), .Y(new_new_n747_));
  NO2        g725(.A(new_new_n747_), .B(new_new_n446_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n748_), .B(new_new_n745_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n319_), .B(new_new_n219_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n750_), .B(new_new_n652_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n751_), .Y(new_new_n752_));
  AOI210     g730(.A0(new_new_n749_), .A1(new_new_n48_), .B0(new_new_n752_), .Y(new_new_n753_));
  AOI210     g731(.A0(new_new_n753_), .A1(new_new_n743_), .B0(new_new_n73_), .Y(new_new_n754_));
  INV        g732(.A(new_new_n274_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n755_), .B(new_new_n551_), .Y(new_new_n756_));
  OAI210     g734(.A0(new_new_n221_), .A1(new_new_n154_), .B0(new_new_n87_), .Y(new_new_n757_));
  NO2        g735(.A(new_new_n757_), .B(i_11_), .Y(new_new_n758_));
  NO3        g736(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n759_));
  OAI210     g737(.A0(new_new_n684_), .A1(new_new_n234_), .B0(new_new_n759_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n760_), .B(new_new_n522_), .Y(new_new_n761_));
  INV        g739(.A(new_new_n374_), .Y(new_new_n762_));
  NO2        g740(.A(new_new_n604_), .B(new_new_n255_), .Y(new_new_n763_));
  AOI210     g741(.A0(new_new_n763_), .A1(new_new_n762_), .B0(new_new_n41_), .Y(new_new_n764_));
  NO3        g742(.A(new_new_n764_), .B(new_new_n761_), .C(new_new_n758_), .Y(new_new_n765_));
  INV        g743(.A(new_new_n765_), .Y(new_new_n766_));
  NO3        g744(.A(new_new_n766_), .B(new_new_n756_), .C(new_new_n754_), .Y(new_new_n767_));
  NA4        g745(.A(new_new_n767_), .B(new_new_n740_), .C(new_new_n703_), .D(new_new_n646_), .Y(ori4));
  INV        g746(.A(new_new_n494_), .Y(new_new_n771_));
  INV        g747(.A(i_6_), .Y(new_new_n772_));
  INV        g748(.A(new_new_n202_), .Y(new_new_n773_));
endmodule


