//Benchmark atmr_alu4_1266_0.125

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n124_, ori_ori_n125_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NOi21      o016(.An(i_12_), .B(i_13_), .Y(ori_ori_n39_));
  INV        o017(.A(ori_ori_n39_), .Y(ori_ori_n40_));
  NAi31      o018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n41_));
  INV        o019(.A(ori_ori_n35_), .Y(ori1));
  INV        o020(.A(i_11_), .Y(ori_ori_n43_));
  NO2        o021(.A(ori_ori_n43_), .B(i_6_), .Y(ori_ori_n44_));
  INV        o022(.A(i_2_), .Y(ori_ori_n45_));
  NA2        o023(.A(i_0_), .B(i_3_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_5_), .A1(ori_ori_n46_), .B0(ori_ori_n45_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_0_), .B(i_2_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NA2        o031(.A(ori_ori_n50_), .B(ori_ori_n44_), .Y(ori_ori_n54_));
  NO2        o032(.A(i_1_), .B(i_6_), .Y(ori_ori_n55_));
  NA2        o033(.A(i_8_), .B(i_7_), .Y(ori_ori_n56_));
  NAi21      o034(.An(i_2_), .B(i_7_), .Y(ori_ori_n57_));
  INV        o035(.A(i_1_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(i_6_), .Y(ori_ori_n59_));
  NA3        o037(.A(ori_ori_n59_), .B(ori_ori_n57_), .C(ori_ori_n31_), .Y(ori_ori_n60_));
  INV        o038(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n62_));
  AOI210     o040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_1_), .B(i_6_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(ori_ori_n25_), .Y(ori_ori_n65_));
  INV        o043(.A(i_0_), .Y(ori_ori_n66_));
  NAi21      o044(.An(i_5_), .B(i_10_), .Y(ori_ori_n67_));
  NA2        o045(.A(i_5_), .B(i_9_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n67_), .B0(ori_ori_n66_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n65_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n63_), .A1(ori_ori_n62_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n61_), .B0(i_0_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_12_), .B(i_5_), .Y(ori_ori_n73_));
  NO2        o051(.A(i_3_), .B(i_7_), .Y(ori_ori_n74_));
  INV        o052(.A(i_6_), .Y(ori_ori_n75_));
  OR4        o053(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n76_));
  INV        o054(.A(ori_ori_n76_), .Y(ori_ori_n77_));
  NO2        o055(.A(i_2_), .B(i_7_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n77_), .B(ori_ori_n78_), .Y(ori_ori_n79_));
  OAI210     o057(.A0(i_1_), .A1(i_6_), .B0(ori_ori_n79_), .Y(ori_ori_n80_));
  NAi21      o058(.An(i_6_), .B(i_10_), .Y(ori_ori_n81_));
  NA2        o059(.A(i_6_), .B(i_9_), .Y(ori_ori_n82_));
  AOI210     o060(.A0(ori_ori_n82_), .A1(ori_ori_n81_), .B0(ori_ori_n58_), .Y(ori_ori_n83_));
  NA2        o061(.A(i_2_), .B(i_6_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n83_), .Y(ori_ori_n85_));
  AOI210     o063(.A0(ori_ori_n85_), .A1(ori_ori_n80_), .B0(ori_ori_n73_), .Y(ori_ori_n86_));
  AN3        o064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n87_));
  NAi21      o065(.An(i_6_), .B(i_11_), .Y(ori_ori_n88_));
  NA2        o066(.A(ori_ori_n87_), .B(ori_ori_n32_), .Y(ori_ori_n89_));
  INV        o067(.A(i_7_), .Y(ori_ori_n90_));
  NA2        o068(.A(ori_ori_n45_), .B(ori_ori_n90_), .Y(ori_ori_n91_));
  NO2        o069(.A(i_0_), .B(i_5_), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(ori_ori_n75_), .Y(ori_ori_n93_));
  NA2        o071(.A(i_12_), .B(i_3_), .Y(ori_ori_n94_));
  INV        o072(.A(ori_ori_n94_), .Y(ori_ori_n95_));
  NAi21      o073(.An(i_7_), .B(i_11_), .Y(ori_ori_n96_));
  NO3        o074(.A(ori_ori_n96_), .B(ori_ori_n81_), .C(ori_ori_n51_), .Y(ori_ori_n97_));
  NO2        o075(.A(i_2_), .B(i_7_), .Y(ori_ori_n98_));
  OR2        o076(.A(ori_ori_n73_), .B(ori_ori_n55_), .Y(ori_ori_n99_));
  NA2        o077(.A(i_12_), .B(i_7_), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n58_), .B(ori_ori_n26_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n101_), .B(i_0_), .Y(ori_ori_n102_));
  NA2        o080(.A(i_11_), .B(i_12_), .Y(ori_ori_n103_));
  OAI210     o081(.A0(ori_ori_n102_), .A1(ori_ori_n100_), .B0(ori_ori_n103_), .Y(ori_ori_n104_));
  INV        o082(.A(ori_ori_n104_), .Y(ori_ori_n105_));
  NAi31      o083(.An(ori_ori_n97_), .B(ori_ori_n105_), .C(ori_ori_n89_), .Y(ori_ori_n106_));
  NOi21      o084(.An(i_1_), .B(i_5_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n107_), .B(i_11_), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n90_), .B(ori_ori_n37_), .Y(ori_ori_n109_));
  NA2        o087(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n110_), .B(ori_ori_n109_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(ori_ori_n45_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n113_));
  NAi21      o091(.An(i_3_), .B(i_8_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(ori_ori_n57_), .Y(ori_ori_n115_));
  NOi31      o093(.An(ori_ori_n115_), .B(ori_ori_n113_), .C(ori_ori_n112_), .Y(ori_ori_n116_));
  NO2        o094(.A(i_1_), .B(ori_ori_n75_), .Y(ori_ori_n117_));
  NO2        o095(.A(i_6_), .B(i_5_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(i_3_), .Y(ori_ori_n119_));
  AO210      o097(.A0(ori_ori_n119_), .A1(ori_ori_n46_), .B0(ori_ori_n117_), .Y(ori_ori_n120_));
  OAI220     o098(.A0(ori_ori_n120_), .A1(ori_ori_n96_), .B0(ori_ori_n116_), .B1(ori_ori_n108_), .Y(ori_ori_n121_));
  NO3        o099(.A(ori_ori_n121_), .B(ori_ori_n106_), .C(ori_ori_n86_), .Y(ori_ori_n122_));
  NA3        o100(.A(ori_ori_n122_), .B(ori_ori_n72_), .C(ori_ori_n54_), .Y(ori2));
  NO2        o101(.A(ori_ori_n58_), .B(ori_ori_n37_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n707_), .B(ori_ori_n124_), .Y(ori_ori_n125_));
  NA4        o103(.A(ori_ori_n125_), .B(ori_ori_n70_), .C(ori_ori_n62_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o104(.A(i_12_), .B(i_13_), .Y(ori_ori_n127_));
  NAi21      o105(.An(i_5_), .B(i_11_), .Y(ori_ori_n128_));
  NO2        o106(.A(i_0_), .B(i_1_), .Y(ori_ori_n129_));
  NA2        o107(.A(i_2_), .B(i_3_), .Y(ori_ori_n130_));
  NA2        o108(.A(i_1_), .B(i_5_), .Y(ori_ori_n131_));
  OR2        o109(.A(i_0_), .B(i_1_), .Y(ori_ori_n132_));
  NO3        o110(.A(ori_ori_n132_), .B(ori_ori_n73_), .C(i_13_), .Y(ori_ori_n133_));
  NAi32      o111(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n134_));
  NOi21      o112(.An(i_4_), .B(i_10_), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n135_), .B(ori_ori_n39_), .Y(ori_ori_n136_));
  NOi21      o114(.An(i_4_), .B(i_9_), .Y(ori_ori_n137_));
  NOi21      o115(.An(i_11_), .B(i_13_), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n139_));
  NO2        o117(.A(i_4_), .B(i_5_), .Y(ori_ori_n140_));
  NAi21      o118(.An(i_12_), .B(i_11_), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n141_), .B(i_13_), .Y(ori_ori_n142_));
  NO2        o120(.A(ori_ori_n66_), .B(ori_ori_n58_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n66_), .B(i_5_), .Y(ori_ori_n144_));
  NO2        o122(.A(i_13_), .B(i_10_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_2_), .B(i_1_), .Y(ori_ori_n146_));
  NAi21      o124(.An(i_4_), .B(i_12_), .Y(ori_ori_n147_));
  INV        o125(.A(i_8_), .Y(ori_ori_n148_));
  NO3        o126(.A(i_3_), .B(ori_ori_n75_), .C(ori_ori_n47_), .Y(ori_ori_n149_));
  NA2        o127(.A(ori_ori_n149_), .B(i_7_), .Y(ori_ori_n150_));
  NO3        o128(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n151_));
  NO2        o129(.A(i_3_), .B(i_8_), .Y(ori_ori_n152_));
  NO3        o130(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n153_));
  NA3        o131(.A(ori_ori_n153_), .B(ori_ori_n152_), .C(ori_ori_n39_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n92_), .B(ori_ori_n55_), .Y(ori_ori_n155_));
  INV        o133(.A(ori_ori_n155_), .Y(ori_ori_n156_));
  NO2        o134(.A(i_13_), .B(i_9_), .Y(ori_ori_n157_));
  NAi21      o135(.An(i_12_), .B(i_3_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n43_), .B(i_5_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n156_), .B(ori_ori_n154_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(i_7_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n161_), .B(i_4_), .Y(ori_ori_n162_));
  NA3        o140(.A(i_13_), .B(ori_ori_n148_), .C(i_10_), .Y(ori_ori_n163_));
  NA2        o141(.A(i_0_), .B(i_5_), .Y(ori_ori_n164_));
  NAi31      o142(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n66_), .B(ori_ori_n26_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n45_), .B(ori_ori_n58_), .Y(ori_ori_n168_));
  INV        o146(.A(i_13_), .Y(ori_ori_n169_));
  NO2        o147(.A(i_12_), .B(ori_ori_n169_), .Y(ori_ori_n170_));
  NO2        o148(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n171_));
  OR2        o149(.A(i_8_), .B(i_7_), .Y(ori_ori_n172_));
  INV        o150(.A(i_12_), .Y(ori_ori_n173_));
  NO3        o151(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n174_));
  NA2        o152(.A(i_2_), .B(i_1_), .Y(ori_ori_n175_));
  NO3        o153(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n176_));
  NAi21      o154(.An(i_4_), .B(i_3_), .Y(ori_ori_n177_));
  NO2        o155(.A(i_0_), .B(i_6_), .Y(ori_ori_n178_));
  NOi41      o156(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n179_));
  NO2        o157(.A(i_11_), .B(ori_ori_n169_), .Y(ori_ori_n180_));
  NOi21      o158(.An(i_1_), .B(i_6_), .Y(ori_ori_n181_));
  NAi21      o159(.An(i_3_), .B(i_7_), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n173_), .B(i_9_), .Y(ori_ori_n183_));
  OR4        o161(.A(ori_ori_n183_), .B(ori_ori_n182_), .C(ori_ori_n181_), .D(ori_ori_n144_), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n66_), .B(i_5_), .Y(ori_ori_n185_));
  NA2        o163(.A(i_3_), .B(i_9_), .Y(ori_ori_n186_));
  NAi21      o164(.An(i_7_), .B(i_10_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NA3        o166(.A(ori_ori_n188_), .B(ori_ori_n185_), .C(ori_ori_n59_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n189_), .B(ori_ori_n184_), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n190_), .B(ori_ori_n180_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n172_), .B(ori_ori_n37_), .Y(ori_ori_n192_));
  NA2        o170(.A(i_12_), .B(i_6_), .Y(ori_ori_n193_));
  OR2        o171(.A(i_13_), .B(i_9_), .Y(ori_ori_n194_));
  NO3        o172(.A(ori_ori_n194_), .B(ori_ori_n193_), .C(ori_ori_n47_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n177_), .B(i_2_), .Y(ori_ori_n196_));
  NA3        o174(.A(ori_ori_n196_), .B(ori_ori_n195_), .C(ori_ori_n43_), .Y(ori_ori_n197_));
  NA2        o175(.A(ori_ori_n180_), .B(i_9_), .Y(ori_ori_n198_));
  OAI210     o176(.A0(ori_ori_n66_), .A1(ori_ori_n198_), .B0(ori_ori_n197_), .Y(ori_ori_n199_));
  NO3        o177(.A(i_11_), .B(ori_ori_n169_), .C(ori_ori_n25_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n182_), .B(i_8_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n199_), .B(ori_ori_n192_), .Y(ori_ori_n202_));
  NA2        o180(.A(ori_ori_n202_), .B(ori_ori_n191_), .Y(ori_ori_n203_));
  NO3        o181(.A(i_12_), .B(ori_ori_n169_), .C(ori_ori_n37_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n175_), .B(i_0_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_3_), .B(i_10_), .Y(ori_ori_n206_));
  NO2        o184(.A(i_2_), .B(ori_ori_n90_), .Y(ori_ori_n207_));
  AN2        o185(.A(i_3_), .B(i_10_), .Y(ori_ori_n208_));
  NO2        o186(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n45_), .B(ori_ori_n26_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n203_), .B(ori_ori_n162_), .Y(ori_ori_n211_));
  NO3        o189(.A(ori_ori_n43_), .B(i_13_), .C(i_9_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_2_), .B(i_3_), .Y(ori_ori_n213_));
  OR2        o191(.A(i_0_), .B(i_5_), .Y(ori_ori_n214_));
  NO2        o192(.A(i_12_), .B(i_10_), .Y(ori_ori_n215_));
  NOi21      o193(.An(i_5_), .B(i_0_), .Y(ori_ori_n216_));
  NO2        o194(.A(i_2_), .B(ori_ori_n90_), .Y(ori_ori_n217_));
  NO4        o195(.A(ori_ori_n217_), .B(i_4_), .C(ori_ori_n216_), .D(ori_ori_n114_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n215_), .Y(ori_ori_n219_));
  INV        o197(.A(i_6_), .Y(ori_ori_n220_));
  NO2        o198(.A(i_1_), .B(i_7_), .Y(ori_ori_n221_));
  INV        o199(.A(ori_ori_n219_), .Y(ori_ori_n222_));
  NOi21      o200(.An(ori_ori_n131_), .B(ori_ori_n93_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(ori_ori_n110_), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n224_), .B(i_3_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n148_), .B(i_9_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n226_), .B(ori_ori_n155_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n45_), .Y(ori_ori_n228_));
  INV        o206(.A(ori_ori_n228_), .Y(ori_ori_n229_));
  AOI210     o207(.A0(ori_ori_n229_), .A1(ori_ori_n225_), .B0(ori_ori_n136_), .Y(ori_ori_n230_));
  AOI210     o208(.A0(ori_ori_n222_), .A1(ori_ori_n212_), .B0(ori_ori_n230_), .Y(ori_ori_n231_));
  NOi32      o209(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n232_));
  INV        o210(.A(ori_ori_n232_), .Y(ori_ori_n233_));
  NAi21      o211(.An(i_0_), .B(i_6_), .Y(ori_ori_n234_));
  NAi21      o212(.An(i_1_), .B(i_5_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n235_), .B(ori_ori_n234_), .Y(ori_ori_n236_));
  NA2        o214(.A(ori_ori_n236_), .B(ori_ori_n25_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n237_), .B(ori_ori_n134_), .Y(ori_ori_n238_));
  NAi41      o216(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n239_));
  OAI220     o217(.A0(ori_ori_n239_), .A1(ori_ori_n235_), .B0(ori_ori_n165_), .B1(ori_ori_n134_), .Y(ori_ori_n240_));
  AOI210     o218(.A0(ori_ori_n239_), .A1(ori_ori_n134_), .B0(ori_ori_n132_), .Y(ori_ori_n241_));
  NOi32      o219(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n242_));
  NAi21      o220(.An(i_6_), .B(i_1_), .Y(ori_ori_n243_));
  NA3        o221(.A(ori_ori_n243_), .B(ori_ori_n242_), .C(ori_ori_n45_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(i_0_), .Y(ori_ori_n245_));
  OR3        o223(.A(ori_ori_n245_), .B(ori_ori_n241_), .C(ori_ori_n240_), .Y(ori_ori_n246_));
  NAi21      o224(.An(i_3_), .B(i_4_), .Y(ori_ori_n247_));
  NO2        o225(.A(ori_ori_n247_), .B(i_9_), .Y(ori_ori_n248_));
  AN2        o226(.A(i_6_), .B(i_7_), .Y(ori_ori_n249_));
  NA2        o227(.A(i_2_), .B(i_7_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n247_), .B(i_10_), .Y(ori_ori_n251_));
  AOI210     o229(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n252_), .A1(ori_ori_n146_), .B0(ori_ori_n251_), .Y(ori_ori_n253_));
  AOI220     o231(.A0(ori_ori_n251_), .A1(ori_ori_n221_), .B0(ori_ori_n174_), .B1(ori_ori_n146_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n254_), .A1(ori_ori_n253_), .B0(i_5_), .Y(ori_ori_n255_));
  NO3        o233(.A(ori_ori_n255_), .B(ori_ori_n246_), .C(ori_ori_n238_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n256_), .B(ori_ori_n233_), .Y(ori_ori_n257_));
  AN2        o235(.A(i_12_), .B(i_5_), .Y(ori_ori_n258_));
  NA2        o236(.A(i_3_), .B(ori_ori_n258_), .Y(ori_ori_n259_));
  NO2        o237(.A(i_11_), .B(i_6_), .Y(ori_ori_n260_));
  NO2        o238(.A(i_5_), .B(i_10_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n262_));
  NA4        o240(.A(ori_ori_n206_), .B(ori_ori_n82_), .C(ori_ori_n68_), .D(ori_ori_n52_), .Y(ori_ori_n263_));
  NO2        o241(.A(i_11_), .B(i_12_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n36_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n263_), .B(ori_ori_n265_), .Y(ori_ori_n266_));
  NAi21      o244(.An(i_13_), .B(i_0_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n267_), .B(ori_ori_n175_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n266_), .B(ori_ori_n268_), .Y(ori_ori_n269_));
  NO2        o247(.A(i_0_), .B(i_11_), .Y(ori_ori_n270_));
  NOi21      o248(.An(i_2_), .B(i_12_), .Y(ori_ori_n271_));
  NAi21      o249(.An(i_9_), .B(i_4_), .Y(ori_ori_n272_));
  OR2        o250(.A(i_13_), .B(i_10_), .Y(ori_ori_n273_));
  NO3        o251(.A(ori_ori_n273_), .B(ori_ori_n103_), .C(ori_ori_n272_), .Y(ori_ori_n274_));
  NO2        o252(.A(ori_ori_n139_), .B(ori_ori_n109_), .Y(ori_ori_n275_));
  NO2        o253(.A(ori_ori_n90_), .B(ori_ori_n25_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n204_), .B(ori_ori_n276_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n277_), .B(ori_ori_n223_), .Y(ori_ori_n278_));
  NA2        o256(.A(ori_ori_n148_), .B(i_10_), .Y(ori_ori_n279_));
  NA3        o257(.A(ori_ori_n185_), .B(ori_ori_n59_), .C(i_2_), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n280_), .B(ori_ori_n279_), .Y(ori_ori_n281_));
  INV        o259(.A(ori_ori_n281_), .Y(ori_ori_n282_));
  NO2        o260(.A(ori_ori_n282_), .B(ori_ori_n198_), .Y(ori_ori_n283_));
  NO4        o261(.A(ori_ori_n283_), .B(ori_ori_n278_), .C(ori_ori_n708_), .D(ori_ori_n257_), .Y(ori_ori_n284_));
  NO2        o262(.A(ori_ori_n66_), .B(i_13_), .Y(ori_ori_n285_));
  NO2        o263(.A(i_10_), .B(i_9_), .Y(ori_ori_n286_));
  NAi21      o264(.An(i_12_), .B(i_8_), .Y(ori_ori_n287_));
  NO2        o265(.A(ori_ori_n287_), .B(i_3_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n45_), .B(i_4_), .Y(ori_ori_n289_));
  NA2        o267(.A(ori_ori_n289_), .B(ori_ori_n93_), .Y(ori_ori_n290_));
  NO2        o268(.A(ori_ori_n290_), .B(ori_ori_n154_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n210_), .B(i_0_), .Y(ori_ori_n292_));
  NO3        o270(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n293_));
  NA2        o271(.A(ori_ori_n193_), .B(ori_ori_n88_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n294_), .B(ori_ori_n293_), .Y(ori_ori_n295_));
  NA2        o273(.A(i_8_), .B(i_9_), .Y(ori_ori_n296_));
  NO2        o274(.A(i_7_), .B(i_2_), .Y(ori_ori_n297_));
  OR2        o275(.A(ori_ori_n297_), .B(ori_ori_n296_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n204_), .B(ori_ori_n155_), .Y(ori_ori_n299_));
  OAI220     o277(.A0(ori_ori_n299_), .A1(ori_ori_n298_), .B0(ori_ori_n295_), .B1(ori_ori_n292_), .Y(ori_ori_n300_));
  NA2        o278(.A(ori_ori_n180_), .B(ori_ori_n209_), .Y(ori_ori_n301_));
  NO3        o279(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n302_));
  INV        o280(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  NA3        o281(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n304_));
  NA4        o282(.A(ori_ori_n128_), .B(ori_ori_n101_), .C(ori_ori_n73_), .D(ori_ori_n23_), .Y(ori_ori_n305_));
  OAI220     o283(.A0(ori_ori_n305_), .A1(ori_ori_n304_), .B0(ori_ori_n303_), .B1(ori_ori_n301_), .Y(ori_ori_n306_));
  NO3        o284(.A(ori_ori_n306_), .B(ori_ori_n300_), .C(ori_ori_n291_), .Y(ori_ori_n307_));
  OR2        o285(.A(ori_ori_n227_), .B(ori_ori_n90_), .Y(ori_ori_n308_));
  OR2        o286(.A(ori_ori_n308_), .B(ori_ori_n136_), .Y(ori_ori_n309_));
  NA2        o287(.A(ori_ori_n87_), .B(i_13_), .Y(ori_ori_n310_));
  NO2        o288(.A(i_2_), .B(i_13_), .Y(ori_ori_n311_));
  NO3        o289(.A(i_4_), .B(ori_ori_n47_), .C(i_8_), .Y(ori_ori_n312_));
  NO2        o290(.A(i_6_), .B(i_7_), .Y(ori_ori_n313_));
  NO2        o291(.A(i_11_), .B(i_1_), .Y(ori_ori_n314_));
  NOi21      o292(.An(i_2_), .B(i_7_), .Y(ori_ori_n315_));
  NO2        o293(.A(i_3_), .B(ori_ori_n148_), .Y(ori_ori_n316_));
  NO2        o294(.A(i_6_), .B(i_10_), .Y(ori_ori_n317_));
  NA3        o295(.A(ori_ori_n179_), .B(ori_ori_n138_), .C(ori_ori_n118_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n45_), .B(ori_ori_n43_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n132_), .B(i_3_), .Y(ori_ori_n320_));
  NAi31      o298(.An(ori_ori_n319_), .B(ori_ori_n320_), .C(ori_ori_n170_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n293_), .B(ori_ori_n258_), .Y(ori_ori_n322_));
  NAi21      o300(.An(ori_ori_n163_), .B(ori_ori_n264_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n221_), .B(ori_ori_n164_), .Y(ori_ori_n324_));
  NO2        o302(.A(ori_ori_n324_), .B(ori_ori_n323_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n212_), .B(ori_ori_n174_), .Y(ori_ori_n327_));
  OAI220     o305(.A0(ori_ori_n327_), .A1(ori_ori_n280_), .B0(ori_ori_n326_), .B1(ori_ori_n310_), .Y(ori_ori_n328_));
  NO2        o306(.A(ori_ori_n328_), .B(ori_ori_n325_), .Y(ori_ori_n329_));
  NA4        o307(.A(ori_ori_n329_), .B(ori_ori_n321_), .C(ori_ori_n309_), .D(ori_ori_n307_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n108_), .B(ori_ori_n99_), .Y(ori_ori_n331_));
  AN2        o309(.A(ori_ori_n331_), .B(ori_ori_n293_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n332_), .B(ori_ori_n210_), .Y(ori_ori_n333_));
  NA2        o311(.A(ori_ori_n258_), .B(ori_ori_n169_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n232_), .B(ori_ori_n66_), .Y(ori_ori_n335_));
  NA2        o313(.A(ori_ori_n249_), .B(ori_ori_n242_), .Y(ori_ori_n336_));
  OR2        o314(.A(ori_ori_n334_), .B(ori_ori_n336_), .Y(ori_ori_n337_));
  NO2        o315(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n338_));
  INV        o316(.A(ori_ori_n274_), .Y(ori_ori_n339_));
  NA2        o317(.A(ori_ori_n339_), .B(ori_ori_n337_), .Y(ori_ori_n340_));
  INV        o318(.A(ori_ori_n340_), .Y(ori_ori_n341_));
  INV        o319(.A(ori_ori_n185_), .Y(ori_ori_n342_));
  OAI210     o320(.A0(i_8_), .A1(ori_ori_n342_), .B0(ori_ori_n120_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n343_), .B(ori_ori_n275_), .Y(ori_ori_n344_));
  NA3        o322(.A(ori_ori_n344_), .B(ori_ori_n341_), .C(ori_ori_n333_), .Y(ori_ori_n345_));
  NO2        o323(.A(i_12_), .B(ori_ori_n148_), .Y(ori_ori_n346_));
  NO2        o324(.A(i_8_), .B(i_7_), .Y(ori_ori_n347_));
  NA2        o325(.A(ori_ori_n43_), .B(i_10_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(i_6_), .Y(ori_ori_n349_));
  NA3        o327(.A(ori_ori_n208_), .B(ori_ori_n140_), .C(ori_ori_n87_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n132_), .B(i_5_), .Y(ori_ori_n351_));
  INV        o329(.A(ori_ori_n350_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n352_), .B(ori_ori_n302_), .Y(ori_ori_n353_));
  INV        o331(.A(ori_ori_n353_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n168_), .B(ori_ori_n167_), .Y(ori_ori_n355_));
  NA2        o333(.A(ori_ori_n286_), .B(ori_ori_n166_), .Y(ori_ori_n356_));
  NO2        o334(.A(ori_ori_n355_), .B(ori_ori_n356_), .Y(ori_ori_n357_));
  NO2        o335(.A(ori_ori_n45_), .B(i_7_), .Y(ori_ori_n358_));
  NA2        o336(.A(i_0_), .B(ori_ori_n47_), .Y(ori_ori_n359_));
  NA3        o337(.A(ori_ori_n346_), .B(ori_ori_n200_), .C(ori_ori_n359_), .Y(ori_ori_n360_));
  NO2        o338(.A(ori_ori_n358_), .B(ori_ori_n360_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n361_), .B(ori_ori_n357_), .Y(ori_ori_n362_));
  NO4        o340(.A(ori_ori_n181_), .B(ori_ori_n41_), .C(i_2_), .D(ori_ori_n47_), .Y(ori_ori_n363_));
  NO3        o341(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n364_));
  NOi21      o342(.An(i_10_), .B(i_6_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n75_), .B(ori_ori_n25_), .Y(ori_ori_n366_));
  AOI220     o344(.A0(ori_ori_n204_), .A1(ori_ori_n366_), .B0(ori_ori_n200_), .B1(ori_ori_n365_), .Y(ori_ori_n367_));
  NO2        o345(.A(ori_ori_n367_), .B(ori_ori_n292_), .Y(ori_ori_n368_));
  NO2        o346(.A(ori_ori_n100_), .B(ori_ori_n23_), .Y(ori_ori_n369_));
  INV        o347(.A(ori_ori_n368_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n335_), .B(ori_ori_n254_), .Y(ori_ori_n371_));
  INV        o349(.A(ori_ori_n213_), .Y(ori_ori_n372_));
  NO2        o350(.A(i_12_), .B(ori_ori_n75_), .Y(ori_ori_n373_));
  NA2        o351(.A(ori_ori_n373_), .B(ori_ori_n200_), .Y(ori_ori_n374_));
  NA3        o352(.A(ori_ori_n260_), .B(ori_ori_n204_), .C(ori_ori_n164_), .Y(ori_ori_n375_));
  AOI210     o353(.A0(ori_ori_n375_), .A1(ori_ori_n374_), .B0(ori_ori_n372_), .Y(ori_ori_n376_));
  OR2        o354(.A(i_2_), .B(i_5_), .Y(ori_ori_n377_));
  NA2        o355(.A(ori_ori_n250_), .B(ori_ori_n178_), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n378_), .B(ori_ori_n323_), .Y(ori_ori_n379_));
  NO3        o357(.A(ori_ori_n379_), .B(ori_ori_n376_), .C(ori_ori_n371_), .Y(ori_ori_n380_));
  NA3        o358(.A(ori_ori_n380_), .B(ori_ori_n370_), .C(ori_ori_n362_), .Y(ori_ori_n381_));
  NO4        o359(.A(ori_ori_n381_), .B(ori_ori_n354_), .C(ori_ori_n345_), .D(ori_ori_n330_), .Y(ori_ori_n382_));
  NA4        o360(.A(ori_ori_n382_), .B(ori_ori_n284_), .C(ori_ori_n231_), .D(ori_ori_n211_), .Y(ori7));
  NO2        o361(.A(ori_ori_n84_), .B(ori_ori_n52_), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n96_), .B(ori_ori_n81_), .Y(ori_ori_n385_));
  NA2        o363(.A(i_3_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  NA2        o364(.A(ori_ori_n317_), .B(ori_ori_n74_), .Y(ori_ori_n387_));
  NA2        o365(.A(i_11_), .B(ori_ori_n148_), .Y(ori_ori_n388_));
  NA2        o366(.A(ori_ori_n127_), .B(ori_ori_n388_), .Y(ori_ori_n389_));
  OAI210     o367(.A0(ori_ori_n389_), .A1(ori_ori_n387_), .B0(ori_ori_n386_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n173_), .B(i_4_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n391_), .B(i_8_), .Y(ori_ori_n392_));
  NA2        o370(.A(i_2_), .B(ori_ori_n75_), .Y(ori_ori_n393_));
  OAI210     o371(.A0(ori_ori_n78_), .A1(ori_ori_n152_), .B0(ori_ori_n153_), .Y(ori_ori_n394_));
  NO2        o372(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n395_));
  NA2        o373(.A(i_4_), .B(i_8_), .Y(ori_ori_n396_));
  NO2        o374(.A(ori_ori_n394_), .B(i_13_), .Y(ori_ori_n397_));
  NO3        o375(.A(ori_ori_n397_), .B(ori_ori_n390_), .C(ori_ori_n384_), .Y(ori_ori_n398_));
  AOI210     o376(.A0(ori_ori_n114_), .A1(ori_ori_n57_), .B0(i_10_), .Y(ori_ori_n399_));
  AOI210     o377(.A0(ori_ori_n399_), .A1(ori_ori_n173_), .B0(ori_ori_n135_), .Y(ori_ori_n400_));
  OR2        o378(.A(i_6_), .B(i_10_), .Y(ori_ori_n401_));
  INV        o379(.A(ori_ori_n151_), .Y(ori_ori_n402_));
  OR2        o380(.A(ori_ori_n400_), .B(ori_ori_n194_), .Y(ori_ori_n403_));
  AOI210     o381(.A0(ori_ori_n403_), .A1(ori_ori_n398_), .B0(ori_ori_n58_), .Y(ori_ori_n404_));
  NOi21      o382(.An(i_11_), .B(i_7_), .Y(ori_ori_n405_));
  AO210      o383(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n406_));
  NO2        o384(.A(ori_ori_n406_), .B(ori_ori_n405_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n407_), .B(ori_ori_n157_), .Y(ori_ori_n408_));
  NA3        o386(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n409_));
  NAi31      o387(.An(ori_ori_n409_), .B(i_12_), .C(i_11_), .Y(ori_ori_n410_));
  AOI210     o388(.A0(ori_ori_n410_), .A1(ori_ori_n408_), .B0(ori_ori_n58_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n77_), .B(ori_ori_n58_), .Y(ori_ori_n412_));
  AO210      o390(.A0(ori_ori_n412_), .A1(ori_ori_n254_), .B0(ori_ori_n40_), .Y(ori_ori_n413_));
  NO3        o391(.A(ori_ori_n187_), .B(ori_ori_n158_), .C(ori_ori_n388_), .Y(ori_ori_n414_));
  OAI210     o392(.A0(ori_ori_n414_), .A1(ori_ori_n170_), .B0(ori_ori_n58_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n271_), .B(ori_ori_n31_), .Y(ori_ori_n416_));
  OR2        o394(.A(ori_ori_n158_), .B(ori_ori_n96_), .Y(ori_ori_n417_));
  NA2        o395(.A(ori_ori_n417_), .B(ori_ori_n416_), .Y(ori_ori_n418_));
  NO2        o396(.A(i_1_), .B(i_4_), .Y(ori_ori_n419_));
  NA2        o397(.A(ori_ori_n419_), .B(ori_ori_n418_), .Y(ori_ori_n420_));
  NO2        o398(.A(i_1_), .B(i_12_), .Y(ori_ori_n421_));
  NA3        o399(.A(ori_ori_n421_), .B(i_2_), .C(ori_ori_n24_), .Y(ori_ori_n422_));
  BUFFER     o400(.A(ori_ori_n422_), .Y(ori_ori_n423_));
  NA4        o401(.A(ori_ori_n423_), .B(ori_ori_n420_), .C(ori_ori_n415_), .D(ori_ori_n413_), .Y(ori_ori_n424_));
  OAI210     o402(.A0(ori_ori_n424_), .A1(ori_ori_n411_), .B0(i_6_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n409_), .B(ori_ori_n96_), .Y(ori_ori_n426_));
  NA2        o404(.A(ori_ori_n426_), .B(ori_ori_n373_), .Y(ori_ori_n427_));
  NO2        o405(.A(i_6_), .B(i_11_), .Y(ori_ori_n428_));
  NA2        o406(.A(ori_ori_n427_), .B(ori_ori_n295_), .Y(ori_ori_n429_));
  NO3        o407(.A(ori_ori_n401_), .B(ori_ori_n172_), .C(ori_ori_n23_), .Y(ori_ori_n430_));
  AOI210     o408(.A0(i_1_), .A1(ori_ori_n188_), .B0(ori_ori_n430_), .Y(ori_ori_n431_));
  NO2        o409(.A(ori_ori_n431_), .B(ori_ori_n43_), .Y(ori_ori_n432_));
  NA3        o410(.A(ori_ori_n347_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n433_));
  INV        o411(.A(i_2_), .Y(ori_ori_n434_));
  NA2        o412(.A(ori_ori_n124_), .B(i_9_), .Y(ori_ori_n435_));
  NA3        o413(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n45_), .B(i_1_), .Y(ori_ori_n437_));
  NA3        o415(.A(ori_ori_n437_), .B(ori_ori_n193_), .C(ori_ori_n43_), .Y(ori_ori_n438_));
  OAI220     o416(.A0(ori_ori_n438_), .A1(ori_ori_n436_), .B0(ori_ori_n435_), .B1(ori_ori_n434_), .Y(ori_ori_n439_));
  AOI210     o417(.A0(ori_ori_n314_), .A1(ori_ori_n276_), .B0(ori_ori_n176_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n440_), .B(ori_ori_n393_), .Y(ori_ori_n441_));
  NAi21      o419(.An(ori_ori_n433_), .B(ori_ori_n83_), .Y(ori_ori_n442_));
  INV        o420(.A(ori_ori_n442_), .Y(ori_ori_n443_));
  OR3        o421(.A(ori_ori_n443_), .B(ori_ori_n441_), .C(ori_ori_n439_), .Y(ori_ori_n444_));
  NO3        o422(.A(ori_ori_n444_), .B(ori_ori_n432_), .C(ori_ori_n429_), .Y(ori_ori_n445_));
  NO2        o423(.A(ori_ori_n173_), .B(ori_ori_n90_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n446_), .B(ori_ori_n405_), .Y(ori_ori_n447_));
  NO2        o425(.A(ori_ori_n709_), .B(ori_ori_n100_), .Y(ori_ori_n448_));
  AN2        o426(.A(ori_ori_n448_), .B(ori_ori_n349_), .Y(ori_ori_n449_));
  NO2        o427(.A(ori_ori_n103_), .B(ori_ori_n37_), .Y(ori_ori_n450_));
  NA2        o428(.A(i_1_), .B(i_3_), .Y(ori_ori_n451_));
  NO2        o429(.A(ori_ori_n296_), .B(ori_ori_n84_), .Y(ori_ori_n452_));
  INV        o430(.A(ori_ori_n452_), .Y(ori_ori_n453_));
  NO2        o431(.A(ori_ori_n453_), .B(ori_ori_n451_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n454_), .B(ori_ori_n449_), .Y(ori_ori_n455_));
  NA3        o433(.A(ori_ori_n455_), .B(ori_ori_n445_), .C(ori_ori_n425_), .Y(ori_ori_n456_));
  NA2        o434(.A(ori_ori_n249_), .B(ori_ori_n248_), .Y(ori_ori_n457_));
  NO3        o435(.A(ori_ori_n315_), .B(ori_ori_n396_), .C(ori_ori_n75_), .Y(ori_ori_n458_));
  NA2        o436(.A(ori_ori_n458_), .B(ori_ori_n25_), .Y(ori_ori_n459_));
  NA2        o437(.A(ori_ori_n459_), .B(ori_ori_n457_), .Y(ori_ori_n460_));
  NA2        o438(.A(ori_ori_n460_), .B(i_1_), .Y(ori_ori_n461_));
  AOI210     o439(.A0(ori_ori_n193_), .A1(ori_ori_n88_), .B0(i_1_), .Y(ori_ori_n462_));
  NO2        o440(.A(ori_ori_n247_), .B(i_2_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n463_), .B(ori_ori_n462_), .Y(ori_ori_n464_));
  AOI210     o442(.A0(ori_ori_n464_), .A1(ori_ori_n461_), .B0(i_13_), .Y(ori_ori_n465_));
  OR2        o443(.A(i_11_), .B(i_7_), .Y(ori_ori_n466_));
  NA3        o444(.A(ori_ori_n466_), .B(ori_ori_n95_), .C(ori_ori_n124_), .Y(ori_ori_n467_));
  AOI220     o445(.A0(ori_ori_n311_), .A1(ori_ori_n135_), .B0(ori_ori_n289_), .B1(ori_ori_n124_), .Y(ori_ori_n468_));
  OAI210     o446(.A0(ori_ori_n468_), .A1(ori_ori_n43_), .B0(ori_ori_n467_), .Y(ori_ori_n469_));
  NA2        o447(.A(ori_ori_n469_), .B(ori_ori_n220_), .Y(ori_ori_n470_));
  INV        o448(.A(ori_ori_n100_), .Y(ori_ori_n471_));
  AOI220     o449(.A0(ori_ori_n471_), .A1(ori_ori_n65_), .B0(ori_ori_n260_), .B1(ori_ori_n437_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n472_), .B(ori_ori_n177_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n113_), .B(i_13_), .Y(ori_ori_n474_));
  NO2        o452(.A(ori_ori_n436_), .B(ori_ori_n100_), .Y(ori_ori_n475_));
  INV        o453(.A(ori_ori_n475_), .Y(ori_ori_n476_));
  OAI220     o454(.A0(ori_ori_n476_), .A1(ori_ori_n64_), .B0(ori_ori_n474_), .B1(ori_ori_n462_), .Y(ori_ori_n477_));
  NO3        o455(.A(ori_ori_n64_), .B(ori_ori_n32_), .C(ori_ori_n90_), .Y(ori_ori_n478_));
  NA2        o456(.A(i_3_), .B(i_7_), .Y(ori_ori_n479_));
  NO3        o457(.A(ori_ori_n315_), .B(ori_ori_n173_), .C(ori_ori_n75_), .Y(ori_ori_n480_));
  AOI210     o458(.A0(ori_ori_n480_), .A1(ori_ori_n479_), .B0(ori_ori_n478_), .Y(ori_ori_n481_));
  AOI220     o459(.A0(ori_ori_n260_), .A1(ori_ori_n437_), .B0(ori_ori_n83_), .B1(ori_ori_n91_), .Y(ori_ori_n482_));
  OAI220     o460(.A0(ori_ori_n482_), .A1(ori_ori_n392_), .B0(ori_ori_n481_), .B1(ori_ori_n402_), .Y(ori_ori_n483_));
  NO3        o461(.A(ori_ori_n483_), .B(ori_ori_n477_), .C(ori_ori_n473_), .Y(ori_ori_n484_));
  OR2        o462(.A(i_11_), .B(i_6_), .Y(ori_ori_n485_));
  NO2        o463(.A(ori_ori_n476_), .B(ori_ori_n485_), .Y(ori_ori_n486_));
  NA3        o464(.A(ori_ori_n271_), .B(ori_ori_n395_), .C(ori_ori_n88_), .Y(ori_ori_n487_));
  NA2        o465(.A(ori_ori_n428_), .B(i_13_), .Y(ori_ori_n488_));
  NAi21      o466(.An(i_11_), .B(i_12_), .Y(ori_ori_n489_));
  NO3        o467(.A(ori_ori_n315_), .B(ori_ori_n373_), .C(ori_ori_n396_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n490_), .B(ori_ori_n212_), .Y(ori_ori_n491_));
  NA3        o469(.A(ori_ori_n491_), .B(ori_ori_n488_), .C(ori_ori_n487_), .Y(ori_ori_n492_));
  OAI210     o470(.A0(ori_ori_n492_), .A1(ori_ori_n486_), .B0(ori_ori_n58_), .Y(ori_ori_n493_));
  NA2        o471(.A(ori_ori_n710_), .B(ori_ori_n421_), .Y(ori_ori_n494_));
  INV        o472(.A(ori_ori_n494_), .Y(ori_ori_n495_));
  NA3        o473(.A(ori_ori_n495_), .B(ori_ori_n44_), .C(ori_ori_n169_), .Y(ori_ori_n496_));
  NA4        o474(.A(ori_ori_n496_), .B(ori_ori_n493_), .C(ori_ori_n484_), .D(ori_ori_n470_), .Y(ori_ori_n497_));
  OR4        o475(.A(ori_ori_n497_), .B(ori_ori_n465_), .C(ori_ori_n456_), .D(ori_ori_n404_), .Y(ori5));
  NA2        o476(.A(ori_ori_n447_), .B(ori_ori_n196_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n392_), .B(i_11_), .Y(ori_ori_n500_));
  NA2        o478(.A(ori_ori_n78_), .B(ori_ori_n500_), .Y(ori_ori_n501_));
  NA2        o479(.A(ori_ori_n501_), .B(ori_ori_n499_), .Y(ori_ori_n502_));
  NO3        o480(.A(i_11_), .B(ori_ori_n173_), .C(i_13_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n110_), .B(ori_ori_n23_), .Y(ori_ori_n504_));
  INV        o482(.A(ori_ori_n286_), .Y(ori_ori_n505_));
  NA2        o483(.A(ori_ori_n213_), .B(ori_ori_n369_), .Y(ori_ori_n506_));
  INV        o484(.A(ori_ori_n506_), .Y(ori_ori_n507_));
  NO2        o485(.A(ori_ori_n507_), .B(ori_ori_n502_), .Y(ori_ori_n508_));
  INV        o486(.A(ori_ori_n138_), .Y(ori_ori_n509_));
  INV        o487(.A(ori_ori_n179_), .Y(ori_ori_n510_));
  OAI210     o488(.A0(ori_ori_n463_), .A1(ori_ori_n288_), .B0(ori_ori_n98_), .Y(ori_ori_n511_));
  AOI210     o489(.A0(ori_ori_n511_), .A1(ori_ori_n510_), .B0(ori_ori_n509_), .Y(ori_ori_n512_));
  NO2        o490(.A(ori_ori_n296_), .B(ori_ori_n26_), .Y(ori_ori_n513_));
  NO2        o491(.A(ori_ori_n513_), .B(ori_ori_n276_), .Y(ori_ori_n514_));
  NA2        o492(.A(ori_ori_n514_), .B(i_2_), .Y(ori_ori_n515_));
  INV        o493(.A(ori_ori_n515_), .Y(ori_ori_n516_));
  AOI210     o494(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n273_), .Y(ori_ori_n517_));
  AOI210     o495(.A0(ori_ori_n517_), .A1(ori_ori_n516_), .B0(ori_ori_n512_), .Y(ori_ori_n518_));
  NO2        o496(.A(ori_ori_n147_), .B(ori_ori_n111_), .Y(ori_ori_n519_));
  OAI210     o497(.A0(ori_ori_n519_), .A1(ori_ori_n504_), .B0(i_2_), .Y(ori_ori_n520_));
  INV        o498(.A(ori_ori_n139_), .Y(ori_ori_n521_));
  NO3        o499(.A(ori_ori_n406_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n522_));
  AOI210     o500(.A0(ori_ori_n521_), .A1(ori_ori_n78_), .B0(ori_ori_n522_), .Y(ori_ori_n523_));
  AOI210     o501(.A0(ori_ori_n523_), .A1(ori_ori_n520_), .B0(ori_ori_n148_), .Y(ori_ori_n524_));
  OA210      o502(.A0(ori_ori_n407_), .A1(ori_ori_n112_), .B0(i_13_), .Y(ori_ori_n525_));
  NA2        o503(.A(ori_ori_n151_), .B(ori_ori_n152_), .Y(ori_ori_n526_));
  NO2        o504(.A(ori_ori_n526_), .B(ori_ori_n250_), .Y(ori_ori_n527_));
  AOI210     o505(.A0(ori_ori_n158_), .A1(ori_ori_n130_), .B0(ori_ori_n338_), .Y(ori_ori_n528_));
  NA2        o506(.A(ori_ori_n528_), .B(ori_ori_n276_), .Y(ori_ori_n529_));
  NO2        o507(.A(ori_ori_n91_), .B(ori_ori_n43_), .Y(ori_ori_n530_));
  INV        o508(.A(ori_ori_n207_), .Y(ori_ori_n531_));
  NA4        o509(.A(ori_ori_n531_), .B(ori_ori_n208_), .C(ori_ori_n110_), .D(ori_ori_n41_), .Y(ori_ori_n532_));
  OAI210     o510(.A0(ori_ori_n532_), .A1(ori_ori_n530_), .B0(ori_ori_n529_), .Y(ori_ori_n533_));
  NO4        o511(.A(ori_ori_n533_), .B(ori_ori_n527_), .C(ori_ori_n525_), .D(ori_ori_n524_), .Y(ori_ori_n534_));
  NA2        o512(.A(ori_ori_n369_), .B(ori_ori_n28_), .Y(ori_ori_n535_));
  NA2        o513(.A(ori_ori_n503_), .B(ori_ori_n201_), .Y(ori_ori_n536_));
  NA2        o514(.A(ori_ori_n536_), .B(ori_ori_n535_), .Y(ori_ori_n537_));
  NO2        o515(.A(ori_ori_n57_), .B(i_12_), .Y(ori_ori_n538_));
  NO2        o516(.A(ori_ori_n538_), .B(ori_ori_n112_), .Y(ori_ori_n539_));
  NO2        o517(.A(ori_ori_n539_), .B(ori_ori_n388_), .Y(ori_ori_n540_));
  AOI220     o518(.A0(ori_ori_n540_), .A1(ori_ori_n36_), .B0(ori_ori_n537_), .B1(ori_ori_n45_), .Y(ori_ori_n541_));
  NA4        o519(.A(ori_ori_n541_), .B(ori_ori_n534_), .C(ori_ori_n518_), .D(ori_ori_n508_), .Y(ori6));
  NA4        o520(.A(ori_ori_n261_), .B(ori_ori_n316_), .C(ori_ori_n64_), .D(ori_ori_n90_), .Y(ori_ori_n543_));
  INV        o521(.A(ori_ori_n543_), .Y(ori_ori_n544_));
  NO2        o522(.A(ori_ori_n165_), .B(ori_ori_n319_), .Y(ori_ori_n545_));
  NO2        o523(.A(i_11_), .B(i_9_), .Y(ori_ori_n546_));
  NO2        o524(.A(ori_ori_n544_), .B(ori_ori_n216_), .Y(ori_ori_n547_));
  OR2        o525(.A(ori_ori_n547_), .B(i_12_), .Y(ori_ori_n548_));
  NA2        o526(.A(ori_ori_n373_), .B(ori_ori_n58_), .Y(ori_ori_n549_));
  BUFFER     o527(.A(ori_ori_n412_), .Y(ori_ori_n550_));
  NA2        o528(.A(ori_ori_n550_), .B(ori_ori_n549_), .Y(ori_ori_n551_));
  INV        o529(.A(ori_ori_n150_), .Y(ori_ori_n552_));
  AOI220     o530(.A0(ori_ori_n552_), .A1(ori_ori_n546_), .B0(ori_ori_n551_), .B1(ori_ori_n66_), .Y(ori_ori_n553_));
  INV        o531(.A(ori_ori_n215_), .Y(ori_ori_n554_));
  NA2        o532(.A(ori_ori_n68_), .B(ori_ori_n117_), .Y(ori_ori_n555_));
  INV        o533(.A(ori_ori_n110_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n556_), .B(ori_ori_n45_), .Y(ori_ori_n557_));
  AOI210     o535(.A0(ori_ori_n557_), .A1(ori_ori_n555_), .B0(ori_ori_n554_), .Y(ori_ori_n558_));
  NO2        o536(.A(ori_ori_n181_), .B(i_9_), .Y(ori_ori_n559_));
  NA2        o537(.A(ori_ori_n559_), .B(ori_ori_n538_), .Y(ori_ori_n560_));
  AOI210     o538(.A0(ori_ori_n560_), .A1(ori_ori_n336_), .B0(ori_ori_n144_), .Y(ori_ori_n561_));
  NO2        o539(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n562_));
  NAi32      o540(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n563_));
  NO2        o541(.A(ori_ori_n485_), .B(ori_ori_n563_), .Y(ori_ori_n564_));
  OR3        o542(.A(ori_ori_n564_), .B(ori_ori_n561_), .C(ori_ori_n558_), .Y(ori_ori_n565_));
  NO2        o543(.A(ori_ori_n466_), .B(i_2_), .Y(ori_ori_n566_));
  NA3        o544(.A(ori_ori_n288_), .B(ori_ori_n129_), .C(ori_ori_n62_), .Y(ori_ori_n567_));
  OR2        o545(.A(ori_ori_n505_), .B(ori_ori_n36_), .Y(ori_ori_n568_));
  NA2        o546(.A(ori_ori_n568_), .B(ori_ori_n567_), .Y(ori_ori_n569_));
  OAI210     o547(.A0(i_6_), .A1(i_11_), .B0(ori_ori_n76_), .Y(ori_ori_n570_));
  AOI220     o548(.A0(ori_ori_n570_), .A1(ori_ori_n364_), .B0(ori_ori_n545_), .B1(ori_ori_n479_), .Y(ori_ori_n571_));
  NA3        o549(.A(ori_ori_n250_), .B(ori_ori_n174_), .C(ori_ori_n129_), .Y(ori_ori_n572_));
  NA3        o550(.A(ori_ori_n572_), .B(ori_ori_n571_), .C(ori_ori_n394_), .Y(ori_ori_n573_));
  AO210      o551(.A0(ori_ori_n338_), .A1(ori_ori_n45_), .B0(ori_ori_n77_), .Y(ori_ori_n574_));
  NA3        o552(.A(ori_ori_n574_), .B(ori_ori_n317_), .C(ori_ori_n164_), .Y(ori_ori_n575_));
  NA2        o553(.A(ori_ori_n288_), .B(ori_ori_n286_), .Y(ori_ori_n576_));
  NO2        o554(.A(ori_ori_n401_), .B(ori_ori_n91_), .Y(ori_ori_n577_));
  OAI210     o555(.A0(ori_ori_n577_), .A1(ori_ori_n99_), .B0(ori_ori_n270_), .Y(ori_ori_n578_));
  NA3        o556(.A(ori_ori_n578_), .B(ori_ori_n576_), .C(ori_ori_n575_), .Y(ori_ori_n579_));
  NO4        o557(.A(ori_ori_n579_), .B(ori_ori_n573_), .C(ori_ori_n569_), .D(ori_ori_n565_), .Y(ori_ori_n580_));
  NA4        o558(.A(ori_ori_n580_), .B(ori_ori_n553_), .C(ori_ori_n548_), .D(ori_ori_n256_), .Y(ori3));
  NA2        o559(.A(i_12_), .B(i_10_), .Y(ori_ori_n582_));
  NA2        o560(.A(ori_ori_n572_), .B(ori_ori_n394_), .Y(ori_ori_n583_));
  NA2        o561(.A(ori_ori_n583_), .B(ori_ori_n39_), .Y(ori_ori_n584_));
  NOi21      o562(.An(ori_ori_n87_), .B(ori_ori_n514_), .Y(ori_ori_n585_));
  NO3        o563(.A(ori_ori_n417_), .B(ori_ori_n296_), .C(ori_ori_n117_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n271_), .B(ori_ori_n44_), .Y(ori_ori_n587_));
  AN2        o565(.A(ori_ori_n294_), .B(ori_ori_n53_), .Y(ori_ori_n588_));
  NO3        o566(.A(ori_ori_n588_), .B(ori_ori_n586_), .C(ori_ori_n585_), .Y(ori_ori_n589_));
  AOI210     o567(.A0(ori_ori_n589_), .A1(ori_ori_n584_), .B0(ori_ori_n47_), .Y(ori_ori_n590_));
  NO3        o568(.A(ori_ori_n258_), .B(ori_ori_n38_), .C(i_0_), .Y(ori_ori_n591_));
  NA2        o569(.A(ori_ori_n144_), .B(ori_ori_n365_), .Y(ori_ori_n592_));
  NOi21      o570(.An(ori_ori_n592_), .B(ori_ori_n591_), .Y(ori_ori_n593_));
  NO2        o571(.A(ori_ori_n593_), .B(ori_ori_n58_), .Y(ori_ori_n594_));
  NOi21      o572(.An(i_5_), .B(i_9_), .Y(ori_ori_n595_));
  NA2        o573(.A(ori_ori_n595_), .B(ori_ori_n285_), .Y(ori_ori_n596_));
  BUFFER     o574(.A(ori_ori_n193_), .Y(ori_ori_n597_));
  AOI210     o575(.A0(ori_ori_n597_), .A1(ori_ori_n314_), .B0(ori_ori_n458_), .Y(ori_ori_n598_));
  NO2        o576(.A(ori_ori_n598_), .B(ori_ori_n596_), .Y(ori_ori_n599_));
  NO3        o577(.A(ori_ori_n599_), .B(ori_ori_n594_), .C(ori_ori_n590_), .Y(ori_ori_n600_));
  NA2        o578(.A(ori_ori_n144_), .B(ori_ori_n24_), .Y(ori_ori_n601_));
  NO2        o579(.A(ori_ori_n450_), .B(ori_ori_n385_), .Y(ori_ori_n602_));
  NO2        o580(.A(ori_ori_n602_), .B(ori_ori_n601_), .Y(ori_ori_n603_));
  INV        o581(.A(ori_ori_n603_), .Y(ori_ori_n604_));
  NA2        o582(.A(ori_ori_n366_), .B(i_0_), .Y(ori_ori_n605_));
  NO3        o583(.A(ori_ori_n605_), .B(ori_ori_n259_), .C(ori_ori_n78_), .Y(ori_ori_n606_));
  NO4        o584(.A(ori_ori_n377_), .B(i_12_), .C(ori_ori_n273_), .D(i_6_), .Y(ori_ori_n607_));
  AOI210     o585(.A0(ori_ori_n607_), .A1(i_11_), .B0(ori_ori_n606_), .Y(ori_ori_n608_));
  NA2        o586(.A(ori_ori_n503_), .B(ori_ori_n216_), .Y(ori_ori_n609_));
  AOI210     o587(.A0(ori_ori_n317_), .A1(ori_ori_n78_), .B0(ori_ori_n55_), .Y(ori_ori_n610_));
  NO2        o588(.A(ori_ori_n610_), .B(ori_ori_n609_), .Y(ori_ori_n611_));
  NO2        o589(.A(ori_ori_n183_), .B(ori_ori_n131_), .Y(ori_ori_n612_));
  INV        o590(.A(ori_ori_n348_), .Y(ori_ori_n613_));
  NO4        o591(.A(ori_ori_n100_), .B(ori_ori_n55_), .C(ori_ori_n709_), .D(i_5_), .Y(ori_ori_n614_));
  AO220      o592(.A0(ori_ori_n614_), .A1(ori_ori_n613_), .B0(ori_ori_n612_), .B1(i_6_), .Y(ori_ori_n615_));
  NO2        o593(.A(ori_ori_n615_), .B(ori_ori_n611_), .Y(ori_ori_n616_));
  NA3        o594(.A(ori_ori_n616_), .B(ori_ori_n608_), .C(ori_ori_n604_), .Y(ori_ori_n617_));
  NO2        o595(.A(ori_ori_n92_), .B(ori_ori_n37_), .Y(ori_ori_n618_));
  NA2        o596(.A(i_11_), .B(i_9_), .Y(ori_ori_n619_));
  NO3        o597(.A(i_12_), .B(ori_ori_n619_), .C(ori_ori_n393_), .Y(ori_ori_n620_));
  AN2        o598(.A(ori_ori_n620_), .B(ori_ori_n618_), .Y(ori_ori_n621_));
  NA2        o599(.A(ori_ori_n262_), .B(ori_ori_n143_), .Y(ori_ori_n622_));
  INV        o600(.A(ori_ori_n622_), .Y(ori_ori_n623_));
  NO2        o601(.A(ori_ori_n619_), .B(ori_ori_n66_), .Y(ori_ori_n624_));
  NO2        o602(.A(ori_ori_n623_), .B(ori_ori_n621_), .Y(ori_ori_n625_));
  NA2        o603(.A(ori_ori_n138_), .B(ori_ori_n92_), .Y(ori_ori_n626_));
  NA2        o604(.A(ori_ori_n395_), .B(ori_ori_n216_), .Y(ori_ori_n627_));
  NO2        o605(.A(ori_ori_n627_), .B(ori_ori_n587_), .Y(ori_ori_n628_));
  INV        o606(.A(ori_ori_n628_), .Y(ori_ori_n629_));
  INV        o607(.A(ori_ori_n214_), .Y(ori_ori_n630_));
  NA2        o608(.A(ori_ori_n629_), .B(ori_ori_n625_), .Y(ori_ori_n631_));
  NO2        o609(.A(ori_ori_n582_), .B(ori_ori_n213_), .Y(ori_ori_n632_));
  OA210      o610(.A0(ori_ori_n313_), .A1(ori_ori_n168_), .B0(ori_ori_n312_), .Y(ori_ori_n633_));
  NA2        o611(.A(ori_ori_n632_), .B(ori_ori_n624_), .Y(ori_ori_n634_));
  NA2        o612(.A(ori_ori_n624_), .B(ori_ori_n208_), .Y(ori_ori_n635_));
  INV        o613(.A(ori_ori_n635_), .Y(ori_ori_n636_));
  NA2        o614(.A(ori_ori_n636_), .B(ori_ori_n313_), .Y(ori_ori_n637_));
  NO3        o615(.A(ori_ori_n377_), .B(ori_ori_n234_), .C(ori_ori_n24_), .Y(ori_ori_n638_));
  NO2        o616(.A(ori_ori_n351_), .B(ori_ori_n638_), .Y(ori_ori_n639_));
  NAi21      o617(.An(i_9_), .B(i_5_), .Y(ori_ori_n640_));
  NO2        o618(.A(ori_ori_n640_), .B(ori_ori_n267_), .Y(ori_ori_n641_));
  NA2        o619(.A(ori_ori_n641_), .B(ori_ori_n407_), .Y(ori_ori_n642_));
  OAI220     o620(.A0(ori_ori_n642_), .A1(ori_ori_n75_), .B0(ori_ori_n639_), .B1(ori_ori_n139_), .Y(ori_ori_n643_));
  NO2        o621(.A(ori_ori_n643_), .B(ori_ori_n340_), .Y(ori_ori_n644_));
  NA3        o622(.A(ori_ori_n644_), .B(ori_ori_n637_), .C(ori_ori_n634_), .Y(ori_ori_n645_));
  NO3        o623(.A(ori_ori_n645_), .B(ori_ori_n631_), .C(ori_ori_n617_), .Y(ori_ori_n646_));
  NO2        o624(.A(i_0_), .B(ori_ori_n489_), .Y(ori_ori_n647_));
  AOI210     o625(.A0(ori_ori_n549_), .A1(ori_ori_n457_), .B0(ori_ori_n626_), .Y(ori_ori_n648_));
  INV        o626(.A(ori_ori_n648_), .Y(ori_ori_n649_));
  NA2        o627(.A(ori_ori_n178_), .B(ori_ori_n171_), .Y(ori_ori_n650_));
  AOI210     o628(.A0(ori_ori_n650_), .A1(ori_ori_n605_), .B0(ori_ori_n131_), .Y(ori_ori_n651_));
  INV        o629(.A(ori_ori_n651_), .Y(ori_ori_n652_));
  NA2        o630(.A(ori_ori_n652_), .B(ori_ori_n649_), .Y(ori_ori_n653_));
  NO3        o631(.A(ori_ori_n159_), .B(ori_ori_n258_), .C(i_0_), .Y(ori_ori_n654_));
  OAI210     o632(.A0(ori_ori_n654_), .A1(ori_ori_n69_), .B0(i_13_), .Y(ori_ori_n655_));
  INV        o633(.A(ori_ori_n655_), .Y(ori_ori_n656_));
  INV        o634(.A(ori_ori_n84_), .Y(ori_ori_n657_));
  AOI210     o635(.A0(ori_ori_n657_), .A1(ori_ori_n647_), .B0(ori_ori_n97_), .Y(ori_ori_n658_));
  OR2        o636(.A(ori_ori_n658_), .B(i_5_), .Y(ori_ori_n659_));
  AOI210     o637(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n141_), .Y(ori_ori_n660_));
  NA2        o638(.A(ori_ori_n660_), .B(ori_ori_n633_), .Y(ori_ori_n661_));
  NO3        o639(.A(ori_ori_n587_), .B(ori_ori_n52_), .C(ori_ori_n47_), .Y(ori_ori_n662_));
  NA2        o640(.A(ori_ori_n322_), .B(ori_ori_n318_), .Y(ori_ori_n663_));
  NO3        o641(.A(ori_ori_n663_), .B(ori_ori_n662_), .C(ori_ori_n706_), .Y(ori_ori_n664_));
  NA3        o642(.A(ori_ori_n261_), .B(ori_ori_n138_), .C(ori_ori_n137_), .Y(ori_ori_n665_));
  NA3        o643(.A(i_5_), .B(ori_ori_n205_), .C(ori_ori_n171_), .Y(ori_ori_n666_));
  NA2        o644(.A(ori_ori_n666_), .B(ori_ori_n665_), .Y(ori_ori_n667_));
  NO3        o645(.A(ori_ori_n619_), .B(ori_ori_n164_), .C(ori_ori_n147_), .Y(ori_ori_n668_));
  NO2        o646(.A(ori_ori_n668_), .B(ori_ori_n667_), .Y(ori_ori_n669_));
  NA4        o647(.A(ori_ori_n669_), .B(ori_ori_n664_), .C(ori_ori_n661_), .D(ori_ori_n659_), .Y(ori_ori_n670_));
  BUFFER     o648(.A(ori_ori_n176_), .Y(ori_ori_n671_));
  NO3        o649(.A(ori_ori_n175_), .B(i_0_), .C(i_12_), .Y(ori_ori_n672_));
  AOI220     o650(.A0(ori_ori_n672_), .A1(ori_ori_n671_), .B0(ori_ori_n544_), .B1(ori_ori_n142_), .Y(ori_ori_n673_));
  INV        o651(.A(ori_ori_n673_), .Y(ori_ori_n674_));
  NO4        o652(.A(ori_ori_n674_), .B(ori_ori_n670_), .C(ori_ori_n656_), .D(ori_ori_n653_), .Y(ori_ori_n675_));
  OAI210     o653(.A0(ori_ori_n566_), .A1(ori_ori_n562_), .B0(ori_ori_n37_), .Y(ori_ori_n676_));
  NA2        o654(.A(ori_ori_n676_), .B(ori_ori_n400_), .Y(ori_ori_n677_));
  NA2        o655(.A(ori_ori_n677_), .B(ori_ori_n157_), .Y(ori_ori_n678_));
  BUFFER     o656(.A(ori_ori_n466_), .Y(ori_ori_n679_));
  NA2        o657(.A(ori_ori_n145_), .B(ori_ori_n146_), .Y(ori_ori_n680_));
  AO210      o658(.A0(ori_ori_n679_), .A1(ori_ori_n33_), .B0(ori_ori_n680_), .Y(ori_ori_n681_));
  NAi31      o659(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n682_));
  NO2        o660(.A(ori_ori_n63_), .B(ori_ori_n682_), .Y(ori_ori_n683_));
  NO2        o661(.A(ori_ori_n683_), .B(ori_ori_n430_), .Y(ori_ori_n684_));
  NA2        o662(.A(ori_ori_n684_), .B(ori_ori_n681_), .Y(ori_ori_n685_));
  NO2        o663(.A(ori_ori_n304_), .B(ori_ori_n193_), .Y(ori_ori_n686_));
  AOI210     o664(.A0(ori_ori_n685_), .A1(ori_ori_n47_), .B0(ori_ori_n686_), .Y(ori_ori_n687_));
  AOI210     o665(.A0(ori_ori_n687_), .A1(ori_ori_n678_), .B0(ori_ori_n66_), .Y(ori_ori_n688_));
  INV        o666(.A(ori_ori_n255_), .Y(ori_ori_n689_));
  NO2        o667(.A(ori_ori_n689_), .B(ori_ori_n509_), .Y(ori_ori_n690_));
  OAI210     o668(.A0(ori_ori_n195_), .A1(ori_ori_n133_), .B0(ori_ori_n78_), .Y(ori_ori_n691_));
  NO2        o669(.A(ori_ori_n691_), .B(i_11_), .Y(ori_ori_n692_));
  NO3        o670(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(i_4_), .Y(ori_ori_n693_));
  OAI210     o671(.A0(ori_ori_n630_), .A1(ori_ori_n209_), .B0(ori_ori_n693_), .Y(ori_ori_n694_));
  NO2        o672(.A(ori_ori_n694_), .B(ori_ori_n489_), .Y(ori_ori_n695_));
  NO4        o673(.A(ori_ori_n640_), .B(i_11_), .C(ori_ori_n182_), .D(ori_ori_n181_), .Y(ori_ori_n696_));
  NO2        o674(.A(ori_ori_n696_), .B(ori_ori_n363_), .Y(ori_ori_n697_));
  INV        o675(.A(ori_ori_n240_), .Y(ori_ori_n698_));
  AOI210     o676(.A0(ori_ori_n698_), .A1(ori_ori_n697_), .B0(ori_ori_n40_), .Y(ori_ori_n699_));
  NO3        o677(.A(ori_ori_n699_), .B(ori_ori_n695_), .C(ori_ori_n692_), .Y(ori_ori_n700_));
  INV        o678(.A(ori_ori_n700_), .Y(ori_ori_n701_));
  NO3        o679(.A(ori_ori_n701_), .B(ori_ori_n690_), .C(ori_ori_n688_), .Y(ori_ori_n702_));
  NA4        o680(.A(ori_ori_n702_), .B(ori_ori_n675_), .C(ori_ori_n646_), .D(ori_ori_n600_), .Y(ori4));
  INV        o681(.A(ori_ori_n350_), .Y(ori_ori_n706_));
  INV        o682(.A(i_6_), .Y(ori_ori_n707_));
  INV        o683(.A(ori_ori_n269_), .Y(ori_ori_n708_));
  INV        o684(.A(i_3_), .Y(ori_ori_n709_));
  INV        o685(.A(i_2_), .Y(ori_ori_n710_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_0_), .B(i_2_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_7_), .B(i_9_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NA3        m031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n54_));
  NO2        m032(.A(i_1_), .B(i_6_), .Y(mai_mai_n55_));
  NA2        m033(.A(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  OAI210     m034(.A0(mai_mai_n56_), .A1(mai_mai_n55_), .B0(mai_mai_n54_), .Y(mai_mai_n57_));
  NA2        m035(.A(mai_mai_n57_), .B(i_12_), .Y(mai_mai_n58_));
  NAi21      m036(.An(i_2_), .B(i_7_), .Y(mai_mai_n59_));
  INV        m037(.A(i_1_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n61_));
  NA3        m039(.A(mai_mai_n61_), .B(mai_mai_n59_), .C(mai_mai_n31_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_1_), .B(i_10_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NAi31      m042(.An(mai_mai_n64_), .B(mai_mai_n62_), .C(mai_mai_n58_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n67_));
  NA2        m045(.A(i_1_), .B(i_6_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n25_), .Y(mai_mai_n69_));
  INV        m047(.A(i_0_), .Y(mai_mai_n70_));
  NAi21      m048(.An(i_5_), .B(i_10_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_5_), .B(i_9_), .Y(mai_mai_n72_));
  AOI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n71_), .B0(mai_mai_n70_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n69_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n74_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n65_), .B0(i_0_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_12_), .B(i_5_), .Y(mai_mai_n77_));
  NA2        m055(.A(i_2_), .B(i_8_), .Y(mai_mai_n78_));
  NO2        m056(.A(i_3_), .B(i_9_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_3_), .B(i_7_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n80_), .B(mai_mai_n79_), .C(mai_mai_n60_), .Y(mai_mai_n81_));
  INV        m059(.A(i_6_), .Y(mai_mai_n82_));
  NO2        m060(.A(i_2_), .B(i_7_), .Y(mai_mai_n83_));
  INV        m061(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  NA2        m062(.A(mai_mai_n81_), .B(mai_mai_n84_), .Y(mai_mai_n85_));
  NAi21      m063(.An(i_6_), .B(i_10_), .Y(mai_mai_n86_));
  NA2        m064(.A(i_6_), .B(i_9_), .Y(mai_mai_n87_));
  AOI210     m065(.A0(mai_mai_n87_), .A1(mai_mai_n86_), .B0(mai_mai_n60_), .Y(mai_mai_n88_));
  NA2        m066(.A(i_2_), .B(i_6_), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n49_), .C(mai_mai_n25_), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n90_), .B(mai_mai_n88_), .Y(mai_mai_n91_));
  AOI210     m069(.A0(mai_mai_n91_), .A1(mai_mai_n85_), .B0(mai_mai_n77_), .Y(mai_mai_n92_));
  AN3        m070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n93_));
  NAi21      m071(.An(i_6_), .B(i_11_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_5_), .B(i_8_), .Y(mai_mai_n95_));
  NOi21      m073(.An(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  AOI220     m074(.A0(mai_mai_n96_), .A1(mai_mai_n59_), .B0(mai_mai_n93_), .B1(mai_mai_n32_), .Y(mai_mai_n97_));
  INV        m075(.A(i_7_), .Y(mai_mai_n98_));
  NA2        m076(.A(mai_mai_n46_), .B(mai_mai_n98_), .Y(mai_mai_n99_));
  NO2        m077(.A(i_0_), .B(i_5_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n82_), .Y(mai_mai_n101_));
  NA2        m079(.A(i_12_), .B(i_3_), .Y(mai_mai_n102_));
  INV        m080(.A(mai_mai_n102_), .Y(mai_mai_n103_));
  NA3        m081(.A(mai_mai_n103_), .B(mai_mai_n101_), .C(mai_mai_n99_), .Y(mai_mai_n104_));
  NAi21      m082(.An(i_7_), .B(i_11_), .Y(mai_mai_n105_));
  NO3        m083(.A(mai_mai_n105_), .B(mai_mai_n86_), .C(mai_mai_n51_), .Y(mai_mai_n106_));
  AN2        m084(.A(i_2_), .B(i_10_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(i_7_), .Y(mai_mai_n108_));
  OR2        m086(.A(mai_mai_n77_), .B(mai_mai_n55_), .Y(mai_mai_n109_));
  NO2        m087(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n110_));
  NO3        m088(.A(mai_mai_n110_), .B(mai_mai_n109_), .C(mai_mai_n108_), .Y(mai_mai_n111_));
  NA2        m089(.A(i_12_), .B(i_7_), .Y(mai_mai_n112_));
  NA2        m090(.A(i_11_), .B(i_12_), .Y(mai_mai_n113_));
  INV        m091(.A(mai_mai_n113_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n114_), .B(mai_mai_n111_), .Y(mai_mai_n115_));
  NAi41      m093(.An(mai_mai_n106_), .B(mai_mai_n115_), .C(mai_mai_n104_), .D(mai_mai_n97_), .Y(mai_mai_n116_));
  NOi21      m094(.An(i_1_), .B(i_5_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(i_11_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n98_), .B(mai_mai_n37_), .Y(mai_mai_n119_));
  NA2        m097(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n120_), .B(mai_mai_n119_), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n121_), .B(mai_mai_n46_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n123_));
  NAi21      m101(.An(i_3_), .B(i_8_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(mai_mai_n59_), .Y(mai_mai_n125_));
  NOi31      m103(.An(mai_mai_n125_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n126_));
  NO2        m104(.A(i_1_), .B(mai_mai_n82_), .Y(mai_mai_n127_));
  NO2        m105(.A(i_6_), .B(i_5_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(i_3_), .Y(mai_mai_n129_));
  OAI220     m107(.A0(mai_mai_n129_), .A1(mai_mai_n105_), .B0(mai_mai_n126_), .B1(mai_mai_n118_), .Y(mai_mai_n130_));
  NO3        m108(.A(mai_mai_n130_), .B(mai_mai_n116_), .C(mai_mai_n92_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(mai_mai_n76_), .Y(mai2));
  NO2        m110(.A(mai_mai_n60_), .B(mai_mai_n37_), .Y(mai_mai_n133_));
  NA2        m111(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n135_));
  NA4        m113(.A(mai_mai_n135_), .B(mai_mai_n74_), .C(mai_mai_n66_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m114(.A(i_8_), .B(i_7_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n137_), .B(i_6_), .Y(mai_mai_n138_));
  NO2        m116(.A(i_12_), .B(i_13_), .Y(mai_mai_n139_));
  NAi21      m117(.An(i_5_), .B(i_11_), .Y(mai_mai_n140_));
  NOi21      m118(.An(mai_mai_n139_), .B(mai_mai_n140_), .Y(mai_mai_n141_));
  NO2        m119(.A(i_0_), .B(i_1_), .Y(mai_mai_n142_));
  NA2        m120(.A(i_2_), .B(i_3_), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n143_), .B(i_4_), .Y(mai_mai_n144_));
  NA3        m122(.A(mai_mai_n144_), .B(mai_mai_n142_), .C(mai_mai_n141_), .Y(mai_mai_n145_));
  AN2        m123(.A(mai_mai_n139_), .B(mai_mai_n79_), .Y(mai_mai_n146_));
  NA2        m124(.A(i_1_), .B(i_5_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n70_), .B(mai_mai_n46_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(i_13_), .Y(mai_mai_n150_));
  OR2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n77_), .C(i_13_), .Y(mai_mai_n152_));
  NAi32      m130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n153_));
  NAi21      m131(.An(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m132(.An(i_4_), .B(i_10_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NO3        m134(.A(mai_mai_n70_), .B(i_2_), .C(i_1_), .Y(mai_mai_n157_));
  INV        m135(.A(mai_mai_n157_), .Y(mai_mai_n158_));
  OAI210     m136(.A0(mai_mai_n158_), .A1(mai_mai_n156_), .B0(mai_mai_n154_), .Y(mai_mai_n159_));
  NO2        m137(.A(mai_mai_n159_), .B(mai_mai_n150_), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n160_), .A1(mai_mai_n145_), .B0(mai_mai_n138_), .Y(mai_mai_n161_));
  INV        m139(.A(i_1_), .Y(mai_mai_n162_));
  NA2        m140(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n163_));
  NOi21      m141(.An(i_4_), .B(i_9_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_11_), .B(i_13_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  OR2        m144(.A(mai_mai_n166_), .B(mai_mai_n163_), .Y(mai_mai_n167_));
  NO2        m145(.A(i_4_), .B(i_5_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_12_), .B(i_11_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(i_13_), .Y(mai_mai_n170_));
  NA3        m148(.A(mai_mai_n170_), .B(mai_mai_n168_), .C(mai_mai_n79_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n167_), .B0(mai_mai_n162_), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n70_), .B(mai_mai_n60_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(mai_mai_n46_), .Y(mai_mai_n174_));
  NAi31      m152(.An(mai_mai_n959_), .B(mai_mai_n146_), .C(i_11_), .Y(mai_mai_n175_));
  NA2        m153(.A(i_3_), .B(i_5_), .Y(mai_mai_n176_));
  AOI210     m154(.A0(mai_mai_n166_), .A1(mai_mai_n175_), .B0(mai_mai_n174_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n178_));
  NO2        m156(.A(i_13_), .B(i_10_), .Y(mai_mai_n179_));
  NA3        m157(.A(mai_mai_n179_), .B(mai_mai_n178_), .C(mai_mai_n44_), .Y(mai_mai_n180_));
  NO2        m158(.A(i_2_), .B(i_1_), .Y(mai_mai_n181_));
  NA2        m159(.A(mai_mai_n181_), .B(i_3_), .Y(mai_mai_n182_));
  NAi21      m160(.An(i_4_), .B(i_12_), .Y(mai_mai_n183_));
  NO3        m161(.A(mai_mai_n183_), .B(mai_mai_n182_), .C(mai_mai_n180_), .Y(mai_mai_n184_));
  NO3        m162(.A(mai_mai_n184_), .B(mai_mai_n177_), .C(mai_mai_n172_), .Y(mai_mai_n185_));
  INV        m163(.A(i_8_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n961_), .B(i_6_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_3_), .B(mai_mai_n82_), .C(mai_mai_n48_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(mai_mai_n110_), .Y(mai_mai_n189_));
  NO3        m167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n190_));
  NA3        m168(.A(mai_mai_n190_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n191_));
  NO3        m169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n192_));
  OAI210     m170(.A0(mai_mai_n93_), .A1(i_12_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  AOI210     m171(.A0(mai_mai_n193_), .A1(mai_mai_n191_), .B0(mai_mai_n189_), .Y(mai_mai_n194_));
  NO2        m172(.A(i_3_), .B(i_8_), .Y(mai_mai_n195_));
  NO3        m173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n196_));
  NO2        m174(.A(i_13_), .B(i_9_), .Y(mai_mai_n197_));
  NA3        m175(.A(mai_mai_n197_), .B(i_6_), .C(mai_mai_n186_), .Y(mai_mai_n198_));
  NAi21      m176(.An(i_12_), .B(i_3_), .Y(mai_mai_n199_));
  BUFFER     m177(.A(mai_mai_n198_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n201_));
  NO3        m179(.A(i_0_), .B(i_2_), .C(mai_mai_n60_), .Y(mai_mai_n202_));
  NA3        m180(.A(mai_mai_n202_), .B(mai_mai_n201_), .C(i_10_), .Y(mai_mai_n203_));
  NO2        m181(.A(mai_mai_n203_), .B(mai_mai_n200_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(mai_mai_n194_), .Y(mai_mai_n205_));
  OAI220     m183(.A0(mai_mai_n205_), .A1(i_4_), .B0(mai_mai_n187_), .B1(mai_mai_n185_), .Y(mai_mai_n206_));
  NAi21      m184(.An(i_12_), .B(i_7_), .Y(mai_mai_n207_));
  NA3        m185(.A(i_13_), .B(mai_mai_n186_), .C(i_10_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n209_));
  NA2        m187(.A(i_0_), .B(i_5_), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n210_), .B(mai_mai_n101_), .Y(mai_mai_n211_));
  OAI220     m189(.A0(mai_mai_n211_), .A1(mai_mai_n182_), .B0(mai_mai_n174_), .B1(mai_mai_n129_), .Y(mai_mai_n212_));
  NAi31      m190(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n70_), .B(mai_mai_n26_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n46_), .B(mai_mai_n60_), .Y(mai_mai_n216_));
  NA3        m194(.A(mai_mai_n216_), .B(mai_mai_n215_), .C(mai_mai_n214_), .Y(mai_mai_n217_));
  INV        m195(.A(i_13_), .Y(mai_mai_n218_));
  NO2        m196(.A(i_12_), .B(mai_mai_n218_), .Y(mai_mai_n219_));
  NA3        m197(.A(mai_mai_n219_), .B(mai_mai_n190_), .C(mai_mai_n188_), .Y(mai_mai_n220_));
  OAI210     m198(.A0(mai_mai_n217_), .A1(mai_mai_n213_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  AOI220     m199(.A0(mai_mai_n221_), .A1(mai_mai_n137_), .B0(mai_mai_n212_), .B1(mai_mai_n209_), .Y(mai_mai_n222_));
  NO2        m200(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n176_), .B(i_4_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n225_));
  OR2        m203(.A(i_8_), .B(i_7_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n226_), .B(mai_mai_n82_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n51_), .B(i_1_), .Y(mai_mai_n228_));
  NA2        m206(.A(mai_mai_n228_), .B(mai_mai_n227_), .Y(mai_mai_n229_));
  INV        m207(.A(i_12_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n44_), .B(mai_mai_n230_), .Y(mai_mai_n231_));
  NO3        m209(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n232_));
  NA2        m210(.A(i_2_), .B(i_1_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n229_), .B(mai_mai_n225_), .Y(mai_mai_n234_));
  NO3        m212(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n235_));
  NAi21      m213(.An(i_4_), .B(i_3_), .Y(mai_mai_n236_));
  INV        m214(.A(mai_mai_n72_), .Y(mai_mai_n237_));
  NO2        m215(.A(i_0_), .B(i_6_), .Y(mai_mai_n238_));
  NOi41      m216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n239_));
  NA2        m217(.A(mai_mai_n239_), .B(mai_mai_n238_), .Y(mai_mai_n240_));
  INV        m218(.A(mai_mai_n234_), .Y(mai_mai_n241_));
  NO2        m219(.A(i_11_), .B(mai_mai_n218_), .Y(mai_mai_n242_));
  NOi21      m220(.An(i_1_), .B(i_6_), .Y(mai_mai_n243_));
  NAi21      m221(.An(i_3_), .B(i_7_), .Y(mai_mai_n244_));
  NA2        m222(.A(mai_mai_n230_), .B(i_9_), .Y(mai_mai_n245_));
  OR4        m223(.A(mai_mai_n245_), .B(mai_mai_n244_), .C(mai_mai_n243_), .D(mai_mai_n178_), .Y(mai_mai_n246_));
  NO2        m224(.A(i_12_), .B(i_3_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n248_));
  NA2        m226(.A(i_3_), .B(i_9_), .Y(mai_mai_n249_));
  NAi21      m227(.An(i_7_), .B(i_10_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n250_), .B(mai_mai_n249_), .Y(mai_mai_n251_));
  NA3        m229(.A(mai_mai_n251_), .B(mai_mai_n248_), .C(mai_mai_n61_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n252_), .B(mai_mai_n246_), .Y(mai_mai_n253_));
  NA3        m231(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n254_));
  INV        m232(.A(mai_mai_n138_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n230_), .B(i_13_), .Y(mai_mai_n256_));
  NO2        m234(.A(mai_mai_n256_), .B(mai_mai_n72_), .Y(mai_mai_n257_));
  AOI220     m235(.A0(mai_mai_n257_), .A1(mai_mai_n255_), .B0(mai_mai_n253_), .B1(mai_mai_n242_), .Y(mai_mai_n258_));
  NO2        m236(.A(mai_mai_n226_), .B(mai_mai_n37_), .Y(mai_mai_n259_));
  NA2        m237(.A(i_12_), .B(i_6_), .Y(mai_mai_n260_));
  OR2        m238(.A(i_13_), .B(i_9_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n236_), .B(i_2_), .Y(mai_mai_n262_));
  NA2        m240(.A(mai_mai_n242_), .B(i_9_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n148_), .B(mai_mai_n60_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n244_), .B(i_8_), .Y(mai_mai_n265_));
  NO2        m243(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n266_));
  NA3        m244(.A(mai_mai_n266_), .B(mai_mai_n265_), .C(i_13_), .Y(mai_mai_n267_));
  NA3        m245(.A(i_6_), .B(mai_mai_n259_), .C(mai_mai_n219_), .Y(mai_mai_n268_));
  AOI210     m246(.A0(mai_mai_n268_), .A1(mai_mai_n267_), .B0(mai_mai_n264_), .Y(mai_mai_n269_));
  INV        m247(.A(mai_mai_n269_), .Y(mai_mai_n270_));
  NA4        m248(.A(mai_mai_n270_), .B(mai_mai_n258_), .C(mai_mai_n241_), .D(mai_mai_n222_), .Y(mai_mai_n271_));
  NO3        m249(.A(i_12_), .B(mai_mai_n218_), .C(mai_mai_n37_), .Y(mai_mai_n272_));
  INV        m250(.A(mai_mai_n272_), .Y(mai_mai_n273_));
  NA2        m251(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n274_));
  NO3        m252(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n275_));
  AOI220     m253(.A0(mai_mai_n275_), .A1(mai_mai_n188_), .B0(i_6_), .B1(mai_mai_n228_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(mai_mai_n274_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n233_), .B(i_0_), .Y(mai_mai_n278_));
  AOI220     m256(.A0(mai_mai_n278_), .A1(mai_mai_n961_), .B0(i_1_), .B1(mai_mai_n137_), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n266_), .B(mai_mai_n26_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n280_), .B(mai_mai_n279_), .Y(mai_mai_n281_));
  NA2        m259(.A(i_0_), .B(i_1_), .Y(mai_mai_n282_));
  NO2        m260(.A(mai_mai_n282_), .B(i_2_), .Y(mai_mai_n283_));
  NO2        m261(.A(mai_mai_n56_), .B(i_6_), .Y(mai_mai_n284_));
  NA2        m262(.A(mai_mai_n284_), .B(mai_mai_n283_), .Y(mai_mai_n285_));
  OAI210     m263(.A0(mai_mai_n158_), .A1(mai_mai_n138_), .B0(mai_mai_n285_), .Y(mai_mai_n286_));
  NO3        m264(.A(mai_mai_n286_), .B(mai_mai_n281_), .C(mai_mai_n277_), .Y(mai_mai_n287_));
  NO2        m265(.A(i_3_), .B(i_10_), .Y(mai_mai_n288_));
  NA3        m266(.A(mai_mai_n288_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n289_));
  NO2        m267(.A(i_2_), .B(mai_mai_n98_), .Y(mai_mai_n290_));
  NA2        m268(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n291_), .B(i_8_), .Y(mai_mai_n292_));
  NA2        m270(.A(mai_mai_n292_), .B(mai_mai_n290_), .Y(mai_mai_n293_));
  AN2        m271(.A(i_3_), .B(i_10_), .Y(mai_mai_n294_));
  NA3        m272(.A(mai_mai_n294_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n295_));
  NO2        m273(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n296_));
  NO2        m274(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n297_));
  OR2        m275(.A(mai_mai_n293_), .B(mai_mai_n289_), .Y(mai_mai_n298_));
  OAI220     m276(.A0(mai_mai_n298_), .A1(i_6_), .B0(mai_mai_n287_), .B1(mai_mai_n273_), .Y(mai_mai_n299_));
  NO4        m277(.A(mai_mai_n299_), .B(mai_mai_n271_), .C(mai_mai_n206_), .D(mai_mai_n161_), .Y(mai_mai_n300_));
  NO3        m278(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n301_));
  NO3        m279(.A(i_6_), .B(mai_mai_n186_), .C(i_7_), .Y(mai_mai_n302_));
  AOI210     m280(.A0(mai_mai_n186_), .A1(mai_mai_n233_), .B0(mai_mai_n163_), .Y(mai_mai_n303_));
  NO2        m281(.A(i_2_), .B(i_3_), .Y(mai_mai_n304_));
  OR2        m282(.A(i_0_), .B(i_5_), .Y(mai_mai_n305_));
  NA2        m283(.A(mai_mai_n210_), .B(mai_mai_n305_), .Y(mai_mai_n306_));
  NA4        m284(.A(mai_mai_n306_), .B(mai_mai_n227_), .C(mai_mai_n304_), .D(i_1_), .Y(mai_mai_n307_));
  NA3        m285(.A(mai_mai_n278_), .B(i_6_), .C(mai_mai_n110_), .Y(mai_mai_n308_));
  NAi21      m286(.An(i_8_), .B(i_7_), .Y(mai_mai_n309_));
  NO2        m287(.A(mai_mai_n309_), .B(i_6_), .Y(mai_mai_n310_));
  NO2        m288(.A(mai_mai_n151_), .B(mai_mai_n46_), .Y(mai_mai_n311_));
  NA2        m289(.A(mai_mai_n311_), .B(mai_mai_n310_), .Y(mai_mai_n312_));
  NA3        m290(.A(mai_mai_n312_), .B(mai_mai_n308_), .C(mai_mai_n307_), .Y(mai_mai_n313_));
  OAI210     m291(.A0(mai_mai_n313_), .A1(mai_mai_n303_), .B0(i_4_), .Y(mai_mai_n314_));
  NO2        m292(.A(i_12_), .B(i_10_), .Y(mai_mai_n315_));
  NOi21      m293(.An(i_5_), .B(i_0_), .Y(mai_mai_n316_));
  NA4        m294(.A(mai_mai_n80_), .B(mai_mai_n36_), .C(mai_mai_n82_), .D(i_8_), .Y(mai_mai_n317_));
  NO2        m295(.A(i_6_), .B(i_8_), .Y(mai_mai_n318_));
  NOi21      m296(.An(i_0_), .B(i_2_), .Y(mai_mai_n319_));
  AN2        m297(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n320_));
  NO2        m298(.A(i_1_), .B(i_7_), .Y(mai_mai_n321_));
  AO220      m299(.A0(mai_mai_n321_), .A1(mai_mai_n320_), .B0(mai_mai_n310_), .B1(mai_mai_n228_), .Y(mai_mai_n322_));
  NA3        m300(.A(mai_mai_n322_), .B(i_4_), .C(i_5_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n323_), .B(mai_mai_n314_), .Y(mai_mai_n324_));
  INV        m302(.A(i_6_), .Y(mai_mai_n325_));
  INV        m303(.A(mai_mai_n306_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n100_), .B(mai_mai_n120_), .Y(mai_mai_n327_));
  OAI210     m305(.A0(mai_mai_n327_), .A1(mai_mai_n326_), .B0(i_3_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n282_), .B(mai_mai_n78_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(mai_mai_n128_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n89_), .B(mai_mai_n186_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n331_), .B(mai_mai_n60_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n332_), .A1(mai_mai_n330_), .B0(i_7_), .Y(mai_mai_n333_));
  NO2        m311(.A(mai_mai_n186_), .B(i_9_), .Y(mai_mai_n334_));
  NO3        m312(.A(mai_mai_n334_), .B(mai_mai_n333_), .C(mai_mai_n281_), .Y(mai_mai_n335_));
  AOI210     m313(.A0(mai_mai_n335_), .A1(mai_mai_n328_), .B0(mai_mai_n156_), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n324_), .A1(mai_mai_n301_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  NOi32      m315(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n338_));
  INV        m316(.A(mai_mai_n338_), .Y(mai_mai_n339_));
  NAi21      m317(.An(i_0_), .B(i_6_), .Y(mai_mai_n340_));
  NAi21      m318(.An(i_1_), .B(i_5_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n342_));
  NA2        m320(.A(mai_mai_n342_), .B(mai_mai_n25_), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n153_), .B0(mai_mai_n240_), .Y(mai_mai_n344_));
  NAi41      m322(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n345_));
  NO2        m323(.A(mai_mai_n153_), .B(mai_mai_n151_), .Y(mai_mai_n346_));
  NOi32      m324(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n347_));
  NO2        m325(.A(i_1_), .B(mai_mai_n98_), .Y(mai_mai_n348_));
  NAi21      m326(.An(i_3_), .B(i_4_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n349_), .B(i_9_), .Y(mai_mai_n350_));
  AN2        m328(.A(i_6_), .B(i_7_), .Y(mai_mai_n351_));
  OAI210     m329(.A0(mai_mai_n351_), .A1(mai_mai_n348_), .B0(mai_mai_n350_), .Y(mai_mai_n352_));
  NA2        m330(.A(i_2_), .B(i_7_), .Y(mai_mai_n353_));
  NO2        m331(.A(mai_mai_n349_), .B(i_10_), .Y(mai_mai_n354_));
  NA3        m332(.A(mai_mai_n354_), .B(mai_mai_n353_), .C(mai_mai_n238_), .Y(mai_mai_n355_));
  AOI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n352_), .B0(mai_mai_n178_), .Y(mai_mai_n356_));
  AOI210     m334(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n357_));
  OAI210     m335(.A0(mai_mai_n357_), .A1(mai_mai_n181_), .B0(mai_mai_n354_), .Y(mai_mai_n358_));
  NO2        m336(.A(mai_mai_n358_), .B(i_5_), .Y(mai_mai_n359_));
  NO4        m337(.A(mai_mai_n359_), .B(mai_mai_n356_), .C(mai_mai_n346_), .D(mai_mai_n344_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n360_), .B(mai_mai_n339_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n56_), .B(mai_mai_n25_), .Y(mai_mai_n362_));
  AN2        m340(.A(i_12_), .B(i_5_), .Y(mai_mai_n363_));
  NO2        m341(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n364_));
  NA2        m342(.A(mai_mai_n364_), .B(mai_mai_n363_), .Y(mai_mai_n365_));
  NO2        m343(.A(i_11_), .B(i_6_), .Y(mai_mai_n366_));
  NA3        m344(.A(mai_mai_n366_), .B(mai_mai_n311_), .C(mai_mai_n218_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n367_), .B(mai_mai_n365_), .Y(mai_mai_n368_));
  NO2        m346(.A(mai_mai_n236_), .B(i_5_), .Y(mai_mai_n369_));
  NO2        m347(.A(i_5_), .B(i_10_), .Y(mai_mai_n370_));
  NA2        m348(.A(mai_mai_n139_), .B(mai_mai_n45_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n371_), .B(mai_mai_n236_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n372_), .B(mai_mai_n362_), .Y(mai_mai_n373_));
  NO2        m351(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n374_));
  INV        m352(.A(mai_mai_n368_), .Y(mai_mai_n375_));
  NO3        m353(.A(mai_mai_n82_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n376_));
  NO2        m354(.A(i_11_), .B(i_12_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n370_), .B(mai_mai_n230_), .Y(mai_mai_n378_));
  NA3        m356(.A(mai_mai_n110_), .B(i_4_), .C(i_11_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(mai_mai_n213_), .Y(mai_mai_n380_));
  NAi21      m358(.An(i_13_), .B(i_0_), .Y(mai_mai_n381_));
  INV        m359(.A(mai_mai_n381_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n380_), .B(mai_mai_n382_), .Y(mai_mai_n383_));
  NA3        m361(.A(mai_mai_n383_), .B(mai_mai_n375_), .C(mai_mai_n373_), .Y(mai_mai_n384_));
  NO3        m362(.A(i_1_), .B(i_12_), .C(mai_mai_n82_), .Y(mai_mai_n385_));
  NO2        m363(.A(i_0_), .B(i_11_), .Y(mai_mai_n386_));
  INV        m364(.A(i_5_), .Y(mai_mai_n387_));
  AN2        m365(.A(i_1_), .B(i_6_), .Y(mai_mai_n388_));
  NOi21      m366(.An(i_2_), .B(i_12_), .Y(mai_mai_n389_));
  NA2        m367(.A(mai_mai_n389_), .B(mai_mai_n388_), .Y(mai_mai_n390_));
  NO2        m368(.A(mai_mai_n390_), .B(mai_mai_n387_), .Y(mai_mai_n391_));
  NA2        m369(.A(mai_mai_n137_), .B(i_9_), .Y(mai_mai_n392_));
  NO2        m370(.A(mai_mai_n392_), .B(i_4_), .Y(mai_mai_n393_));
  NA2        m371(.A(mai_mai_n391_), .B(mai_mai_n393_), .Y(mai_mai_n394_));
  NAi21      m372(.An(i_9_), .B(i_4_), .Y(mai_mai_n395_));
  OR2        m373(.A(i_13_), .B(i_10_), .Y(mai_mai_n396_));
  NO3        m374(.A(mai_mai_n396_), .B(mai_mai_n113_), .C(mai_mai_n395_), .Y(mai_mai_n397_));
  OR2        m375(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n398_));
  NO2        m376(.A(mai_mai_n98_), .B(mai_mai_n25_), .Y(mai_mai_n399_));
  NA2        m377(.A(mai_mai_n272_), .B(mai_mai_n399_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n266_), .B(mai_mai_n202_), .Y(mai_mai_n401_));
  OAI220     m379(.A0(mai_mai_n401_), .A1(mai_mai_n398_), .B0(mai_mai_n400_), .B1(mai_mai_n100_), .Y(mai_mai_n402_));
  INV        m380(.A(mai_mai_n402_), .Y(mai_mai_n403_));
  AOI210     m381(.A0(mai_mai_n403_), .A1(mai_mai_n394_), .B0(mai_mai_n26_), .Y(mai_mai_n404_));
  NA2        m382(.A(mai_mai_n308_), .B(mai_mai_n307_), .Y(mai_mai_n405_));
  AOI220     m383(.A0(mai_mai_n284_), .A1(mai_mai_n275_), .B0(mai_mai_n278_), .B1(i_6_), .Y(mai_mai_n406_));
  NO2        m384(.A(mai_mai_n406_), .B(mai_mai_n163_), .Y(mai_mai_n407_));
  NO2        m385(.A(mai_mai_n176_), .B(mai_mai_n82_), .Y(mai_mai_n408_));
  AOI220     m386(.A0(mai_mai_n408_), .A1(mai_mai_n283_), .B0(i_6_), .B1(mai_mai_n202_), .Y(mai_mai_n409_));
  NO2        m387(.A(mai_mai_n409_), .B(mai_mai_n274_), .Y(mai_mai_n410_));
  NO3        m388(.A(mai_mai_n410_), .B(mai_mai_n407_), .C(mai_mai_n405_), .Y(mai_mai_n411_));
  NA2        m389(.A(mai_mai_n188_), .B(mai_mai_n93_), .Y(mai_mai_n412_));
  NA2        m390(.A(mai_mai_n311_), .B(mai_mai_n82_), .Y(mai_mai_n413_));
  AOI210     m391(.A0(mai_mai_n413_), .A1(mai_mai_n412_), .B0(mai_mai_n309_), .Y(mai_mai_n414_));
  NA2        m392(.A(mai_mai_n186_), .B(i_10_), .Y(mai_mai_n415_));
  NA3        m393(.A(mai_mai_n248_), .B(mai_mai_n61_), .C(i_2_), .Y(mai_mai_n416_));
  NA2        m394(.A(mai_mai_n284_), .B(mai_mai_n228_), .Y(mai_mai_n417_));
  OAI220     m395(.A0(mai_mai_n417_), .A1(mai_mai_n176_), .B0(mai_mai_n416_), .B1(mai_mai_n415_), .Y(mai_mai_n418_));
  NA3        m396(.A(mai_mai_n321_), .B(mai_mai_n320_), .C(i_5_), .Y(mai_mai_n419_));
  INV        m397(.A(mai_mai_n302_), .Y(mai_mai_n420_));
  OAI210     m398(.A0(mai_mai_n420_), .A1(mai_mai_n182_), .B0(mai_mai_n419_), .Y(mai_mai_n421_));
  NO3        m399(.A(mai_mai_n421_), .B(mai_mai_n418_), .C(mai_mai_n414_), .Y(mai_mai_n422_));
  AOI210     m400(.A0(mai_mai_n422_), .A1(mai_mai_n411_), .B0(mai_mai_n263_), .Y(mai_mai_n423_));
  NO4        m401(.A(mai_mai_n423_), .B(mai_mai_n404_), .C(mai_mai_n384_), .D(mai_mai_n361_), .Y(mai_mai_n424_));
  NO2        m402(.A(mai_mai_n60_), .B(i_4_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n70_), .B(i_13_), .Y(mai_mai_n426_));
  NO2        m404(.A(i_10_), .B(i_9_), .Y(mai_mai_n427_));
  NAi21      m405(.An(i_12_), .B(i_8_), .Y(mai_mai_n428_));
  NO2        m406(.A(mai_mai_n428_), .B(i_3_), .Y(mai_mai_n429_));
  INV        m407(.A(i_0_), .Y(mai_mai_n430_));
  NA2        m408(.A(mai_mai_n260_), .B(mai_mai_n94_), .Y(mai_mai_n431_));
  NA2        m409(.A(i_8_), .B(i_9_), .Y(mai_mai_n432_));
  NO3        m410(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n433_));
  NA3        m411(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n434_));
  OR2        m412(.A(mai_mai_n282_), .B(mai_mai_n198_), .Y(mai_mai_n435_));
  BUFFER     m413(.A(mai_mai_n285_), .Y(mai_mai_n436_));
  OA220      m414(.A0(mai_mai_n436_), .A1(mai_mai_n156_), .B0(mai_mai_n435_), .B1(mai_mai_n225_), .Y(mai_mai_n437_));
  NA2        m415(.A(mai_mai_n93_), .B(i_13_), .Y(mai_mai_n438_));
  NA2        m416(.A(mai_mai_n408_), .B(mai_mai_n362_), .Y(mai_mai_n439_));
  NO2        m417(.A(i_2_), .B(i_13_), .Y(mai_mai_n440_));
  NA3        m418(.A(mai_mai_n440_), .B(mai_mai_n155_), .C(mai_mai_n96_), .Y(mai_mai_n441_));
  OAI220     m419(.A0(mai_mai_n441_), .A1(mai_mai_n230_), .B0(mai_mai_n439_), .B1(mai_mai_n438_), .Y(mai_mai_n442_));
  NO3        m420(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n443_));
  NO2        m421(.A(i_6_), .B(i_7_), .Y(mai_mai_n444_));
  NA2        m422(.A(mai_mai_n444_), .B(mai_mai_n443_), .Y(mai_mai_n445_));
  NO2        m423(.A(mai_mai_n70_), .B(i_3_), .Y(mai_mai_n446_));
  NOi21      m424(.An(i_2_), .B(i_7_), .Y(mai_mai_n447_));
  NAi31      m425(.An(i_11_), .B(mai_mai_n447_), .C(mai_mai_n446_), .Y(mai_mai_n448_));
  INV        m426(.A(mai_mai_n396_), .Y(mai_mai_n449_));
  NA3        m427(.A(mai_mai_n449_), .B(mai_mai_n425_), .C(mai_mai_n72_), .Y(mai_mai_n450_));
  NO2        m428(.A(mai_mai_n450_), .B(mai_mai_n448_), .Y(mai_mai_n451_));
  NO2        m429(.A(i_6_), .B(i_10_), .Y(mai_mai_n452_));
  NA4        m430(.A(mai_mai_n452_), .B(mai_mai_n301_), .C(i_8_), .D(mai_mai_n230_), .Y(mai_mai_n453_));
  NO2        m431(.A(mai_mai_n453_), .B(mai_mai_n149_), .Y(mai_mai_n454_));
  NA3        m432(.A(mai_mai_n239_), .B(mai_mai_n165_), .C(mai_mai_n128_), .Y(mai_mai_n455_));
  NA2        m433(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n456_));
  NO2        m434(.A(mai_mai_n151_), .B(i_3_), .Y(mai_mai_n457_));
  NAi31      m435(.An(mai_mai_n456_), .B(mai_mai_n457_), .C(mai_mai_n219_), .Y(mai_mai_n458_));
  NA3        m436(.A(mai_mai_n374_), .B(mai_mai_n173_), .C(mai_mai_n144_), .Y(mai_mai_n459_));
  NA3        m437(.A(mai_mai_n459_), .B(mai_mai_n458_), .C(mai_mai_n455_), .Y(mai_mai_n460_));
  NO4        m438(.A(mai_mai_n460_), .B(mai_mai_n454_), .C(mai_mai_n451_), .D(mai_mai_n442_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n433_), .B(mai_mai_n370_), .Y(mai_mai_n462_));
  NO2        m440(.A(mai_mai_n462_), .B(mai_mai_n217_), .Y(mai_mai_n463_));
  NAi21      m441(.An(mai_mai_n208_), .B(mai_mai_n377_), .Y(mai_mai_n464_));
  NO2        m442(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n465_));
  NO2        m443(.A(i_0_), .B(mai_mai_n82_), .Y(mai_mai_n466_));
  NA3        m444(.A(mai_mai_n466_), .B(mai_mai_n465_), .C(mai_mai_n137_), .Y(mai_mai_n467_));
  OR3        m445(.A(mai_mai_n291_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n468_));
  NO2        m446(.A(mai_mai_n468_), .B(mai_mai_n467_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n470_));
  NA2        m448(.A(mai_mai_n301_), .B(mai_mai_n232_), .Y(mai_mai_n471_));
  OAI220     m449(.A0(mai_mai_n471_), .A1(mai_mai_n416_), .B0(mai_mai_n470_), .B1(mai_mai_n438_), .Y(mai_mai_n472_));
  NA4        m450(.A(mai_mai_n294_), .B(mai_mai_n216_), .C(mai_mai_n70_), .D(mai_mai_n230_), .Y(mai_mai_n473_));
  NO2        m451(.A(mai_mai_n473_), .B(mai_mai_n445_), .Y(mai_mai_n474_));
  NO4        m452(.A(mai_mai_n474_), .B(mai_mai_n472_), .C(mai_mai_n469_), .D(mai_mai_n463_), .Y(mai_mai_n475_));
  NA3        m453(.A(mai_mai_n475_), .B(mai_mai_n461_), .C(mai_mai_n437_), .Y(mai_mai_n476_));
  NA3        m454(.A(mai_mai_n294_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n477_));
  INV        m455(.A(mai_mai_n477_), .Y(mai_mai_n478_));
  BUFFER     m456(.A(mai_mai_n275_), .Y(mai_mai_n479_));
  NA2        m457(.A(mai_mai_n479_), .B(mai_mai_n478_), .Y(mai_mai_n480_));
  INV        m458(.A(mai_mai_n157_), .Y(mai_mai_n481_));
  OAI210     m459(.A0(mai_mai_n481_), .A1(mai_mai_n225_), .B0(mai_mai_n295_), .Y(mai_mai_n482_));
  NA2        m460(.A(mai_mai_n482_), .B(mai_mai_n310_), .Y(mai_mai_n483_));
  NA2        m461(.A(mai_mai_n363_), .B(mai_mai_n218_), .Y(mai_mai_n484_));
  NA2        m462(.A(mai_mai_n351_), .B(mai_mai_n347_), .Y(mai_mai_n485_));
  OR2        m463(.A(mai_mai_n484_), .B(mai_mai_n485_), .Y(mai_mai_n486_));
  NO2        m464(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n487_));
  AOI210     m465(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n397_), .Y(mai_mai_n488_));
  NA2        m466(.A(mai_mai_n488_), .B(mai_mai_n486_), .Y(mai_mai_n489_));
  INV        m467(.A(mai_mai_n489_), .Y(mai_mai_n490_));
  NO2        m468(.A(i_7_), .B(mai_mai_n191_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n176_), .B(mai_mai_n82_), .Y(mai_mai_n492_));
  NA2        m470(.A(mai_mai_n492_), .B(mai_mai_n491_), .Y(mai_mai_n493_));
  NA4        m471(.A(mai_mai_n493_), .B(mai_mai_n490_), .C(mai_mai_n483_), .D(mai_mai_n480_), .Y(mai_mai_n494_));
  NA2        m472(.A(mai_mai_n369_), .B(mai_mai_n283_), .Y(mai_mai_n495_));
  OAI210     m473(.A0(mai_mai_n365_), .A1(mai_mai_n162_), .B0(mai_mai_n495_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n958_), .B(mai_mai_n218_), .Y(mai_mai_n497_));
  NA2        m475(.A(mai_mai_n452_), .B(mai_mai_n27_), .Y(mai_mai_n498_));
  NO2        m476(.A(mai_mai_n498_), .B(mai_mai_n497_), .Y(mai_mai_n499_));
  NOi31      m477(.An(mai_mai_n302_), .B(mai_mai_n396_), .C(mai_mai_n38_), .Y(mai_mai_n500_));
  OAI210     m478(.A0(mai_mai_n500_), .A1(mai_mai_n499_), .B0(mai_mai_n496_), .Y(mai_mai_n501_));
  NO2        m479(.A(i_8_), .B(i_7_), .Y(mai_mai_n502_));
  OAI210     m480(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n503_));
  NA2        m481(.A(mai_mai_n503_), .B(mai_mai_n216_), .Y(mai_mai_n504_));
  NA2        m482(.A(mai_mai_n228_), .B(mai_mai_n197_), .Y(mai_mai_n505_));
  OAI220     m483(.A0(mai_mai_n505_), .A1(mai_mai_n176_), .B0(mai_mai_n504_), .B1(mai_mai_n236_), .Y(mai_mai_n506_));
  NA2        m484(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n507_));
  NO2        m485(.A(mai_mai_n507_), .B(i_6_), .Y(mai_mai_n508_));
  NA3        m486(.A(mai_mai_n508_), .B(mai_mai_n506_), .C(mai_mai_n502_), .Y(mai_mai_n509_));
  AOI220     m487(.A0(mai_mai_n408_), .A1(mai_mai_n311_), .B0(i_2_), .B1(mai_mai_n238_), .Y(mai_mai_n510_));
  OAI220     m488(.A0(mai_mai_n510_), .A1(mai_mai_n256_), .B0(mai_mai_n438_), .B1(mai_mai_n129_), .Y(mai_mai_n511_));
  NA2        m489(.A(mai_mai_n511_), .B(mai_mai_n259_), .Y(mai_mai_n512_));
  NOi31      m490(.An(mai_mai_n278_), .B(mai_mai_n289_), .C(mai_mai_n959_), .Y(mai_mai_n513_));
  NO2        m491(.A(mai_mai_n214_), .B(mai_mai_n44_), .Y(mai_mai_n514_));
  NO2        m492(.A(mai_mai_n151_), .B(i_5_), .Y(mai_mai_n515_));
  NA2        m493(.A(mai_mai_n515_), .B(mai_mai_n304_), .Y(mai_mai_n516_));
  NO2        m494(.A(mai_mai_n516_), .B(mai_mai_n514_), .Y(mai_mai_n517_));
  OAI210     m495(.A0(mai_mai_n517_), .A1(mai_mai_n513_), .B0(mai_mai_n433_), .Y(mai_mai_n518_));
  NA4        m496(.A(mai_mai_n518_), .B(mai_mai_n512_), .C(mai_mai_n509_), .D(mai_mai_n501_), .Y(mai_mai_n519_));
  NA3        m497(.A(mai_mai_n210_), .B(mai_mai_n68_), .C(mai_mai_n44_), .Y(mai_mai_n520_));
  NA2        m498(.A(mai_mai_n272_), .B(mai_mai_n80_), .Y(mai_mai_n521_));
  AOI210     m499(.A0(mai_mai_n520_), .A1(mai_mai_n330_), .B0(mai_mai_n521_), .Y(mai_mai_n522_));
  NO2        m500(.A(mai_mai_n56_), .B(mai_mai_n167_), .Y(mai_mai_n523_));
  NA2        m501(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n524_));
  NA2        m502(.A(mai_mai_n427_), .B(mai_mai_n214_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n524_), .B(mai_mai_n525_), .Y(mai_mai_n526_));
  NO3        m504(.A(mai_mai_n526_), .B(mai_mai_n523_), .C(mai_mai_n522_), .Y(mai_mai_n527_));
  NO4        m505(.A(mai_mai_n243_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n528_));
  NO3        m506(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n529_));
  NO2        m507(.A(mai_mai_n226_), .B(mai_mai_n36_), .Y(mai_mai_n530_));
  AN2        m508(.A(mai_mai_n530_), .B(mai_mai_n529_), .Y(mai_mai_n531_));
  OA210      m509(.A0(mai_mai_n531_), .A1(mai_mai_n528_), .B0(mai_mai_n338_), .Y(mai_mai_n532_));
  NO2        m510(.A(mai_mai_n396_), .B(i_1_), .Y(mai_mai_n533_));
  NOi31      m511(.An(mai_mai_n533_), .B(mai_mai_n431_), .C(mai_mai_n70_), .Y(mai_mai_n534_));
  AN3        m512(.A(mai_mai_n534_), .B(mai_mai_n393_), .C(i_2_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n406_), .B(mai_mai_n171_), .Y(mai_mai_n536_));
  NO3        m514(.A(mai_mai_n536_), .B(mai_mai_n535_), .C(mai_mai_n532_), .Y(mai_mai_n537_));
  NOi21      m515(.An(i_10_), .B(i_6_), .Y(mai_mai_n538_));
  NO2        m516(.A(mai_mai_n112_), .B(mai_mai_n23_), .Y(mai_mai_n539_));
  NA2        m517(.A(mai_mai_n302_), .B(mai_mai_n157_), .Y(mai_mai_n540_));
  AOI220     m518(.A0(mai_mai_n540_), .A1(mai_mai_n417_), .B0(mai_mai_n166_), .B1(mai_mai_n175_), .Y(mai_mai_n541_));
  NO2        m519(.A(mai_mai_n190_), .B(mai_mai_n37_), .Y(mai_mai_n542_));
  NOi31      m520(.An(mai_mai_n141_), .B(mai_mai_n542_), .C(mai_mai_n317_), .Y(mai_mai_n543_));
  NO2        m521(.A(mai_mai_n543_), .B(mai_mai_n541_), .Y(mai_mai_n544_));
  INV        m522(.A(mai_mai_n304_), .Y(mai_mai_n545_));
  NO2        m523(.A(i_12_), .B(mai_mai_n82_), .Y(mai_mai_n546_));
  NO3        m524(.A(i_4_), .B(mai_mai_n325_), .C(mai_mai_n289_), .Y(mai_mai_n547_));
  OR2        m525(.A(i_2_), .B(i_5_), .Y(mai_mai_n548_));
  OR2        m526(.A(mai_mai_n548_), .B(mai_mai_n388_), .Y(mai_mai_n549_));
  NA2        m527(.A(mai_mai_n353_), .B(mai_mai_n238_), .Y(mai_mai_n550_));
  AOI210     m528(.A0(mai_mai_n550_), .A1(mai_mai_n549_), .B0(mai_mai_n464_), .Y(mai_mai_n551_));
  NO2        m529(.A(mai_mai_n551_), .B(mai_mai_n547_), .Y(mai_mai_n552_));
  NA4        m530(.A(mai_mai_n552_), .B(mai_mai_n544_), .C(mai_mai_n537_), .D(mai_mai_n527_), .Y(mai_mai_n553_));
  NO4        m531(.A(mai_mai_n553_), .B(mai_mai_n519_), .C(mai_mai_n494_), .D(mai_mai_n476_), .Y(mai_mai_n554_));
  NA4        m532(.A(mai_mai_n554_), .B(mai_mai_n424_), .C(mai_mai_n337_), .D(mai_mai_n300_), .Y(mai7));
  NO2        m533(.A(mai_mai_n89_), .B(mai_mai_n52_), .Y(mai_mai_n556_));
  NA2        m534(.A(mai_mai_n452_), .B(mai_mai_n80_), .Y(mai_mai_n557_));
  NA2        m535(.A(i_11_), .B(mai_mai_n186_), .Y(mai_mai_n558_));
  NA3        m536(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n559_));
  NO2        m537(.A(mai_mai_n230_), .B(i_4_), .Y(mai_mai_n560_));
  NA2        m538(.A(mai_mai_n560_), .B(i_8_), .Y(mai_mai_n561_));
  NO2        m539(.A(mai_mai_n102_), .B(mai_mai_n559_), .Y(mai_mai_n562_));
  NA2        m540(.A(i_2_), .B(mai_mai_n82_), .Y(mai_mai_n563_));
  OAI210     m541(.A0(mai_mai_n83_), .A1(mai_mai_n195_), .B0(mai_mai_n196_), .Y(mai_mai_n564_));
  NO2        m542(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n565_));
  NA2        m543(.A(i_4_), .B(i_8_), .Y(mai_mai_n566_));
  AOI210     m544(.A0(mai_mai_n566_), .A1(mai_mai_n294_), .B0(mai_mai_n565_), .Y(mai_mai_n567_));
  OAI220     m545(.A0(mai_mai_n567_), .A1(mai_mai_n563_), .B0(mai_mai_n564_), .B1(i_13_), .Y(mai_mai_n568_));
  NO3        m546(.A(mai_mai_n568_), .B(mai_mai_n562_), .C(mai_mai_n556_), .Y(mai_mai_n569_));
  AOI210     m547(.A0(mai_mai_n124_), .A1(mai_mai_n59_), .B0(i_10_), .Y(mai_mai_n570_));
  AOI210     m548(.A0(mai_mai_n570_), .A1(mai_mai_n230_), .B0(mai_mai_n155_), .Y(mai_mai_n571_));
  OR2        m549(.A(i_6_), .B(i_10_), .Y(mai_mai_n572_));
  NO2        m550(.A(mai_mai_n572_), .B(mai_mai_n23_), .Y(mai_mai_n573_));
  OR3        m551(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n574_));
  NO3        m552(.A(mai_mai_n574_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n575_));
  INV        m553(.A(mai_mai_n192_), .Y(mai_mai_n576_));
  NO2        m554(.A(mai_mai_n575_), .B(mai_mai_n573_), .Y(mai_mai_n577_));
  OA220      m555(.A0(mai_mai_n577_), .A1(mai_mai_n545_), .B0(mai_mai_n571_), .B1(mai_mai_n261_), .Y(mai_mai_n578_));
  AOI210     m556(.A0(mai_mai_n578_), .A1(mai_mai_n569_), .B0(mai_mai_n60_), .Y(mai_mai_n579_));
  NOi21      m557(.An(i_11_), .B(i_7_), .Y(mai_mai_n580_));
  AO210      m558(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n581_));
  NO2        m559(.A(mai_mai_n581_), .B(mai_mai_n580_), .Y(mai_mai_n582_));
  NA3        m560(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n583_));
  NO3        m561(.A(mai_mai_n250_), .B(mai_mai_n199_), .C(mai_mai_n558_), .Y(mai_mai_n584_));
  OAI210     m562(.A0(mai_mai_n584_), .A1(mai_mai_n219_), .B0(mai_mai_n60_), .Y(mai_mai_n585_));
  NO2        m563(.A(mai_mai_n60_), .B(i_9_), .Y(mai_mai_n586_));
  NO2        m564(.A(i_1_), .B(i_12_), .Y(mai_mai_n587_));
  INV        m565(.A(mai_mai_n585_), .Y(mai_mai_n588_));
  NA2        m566(.A(mai_mai_n588_), .B(i_6_), .Y(mai_mai_n589_));
  NO2        m567(.A(mai_mai_n583_), .B(mai_mai_n105_), .Y(mai_mai_n590_));
  NA2        m568(.A(mai_mai_n590_), .B(mai_mai_n546_), .Y(mai_mai_n591_));
  NO2        m569(.A(i_6_), .B(i_11_), .Y(mai_mai_n592_));
  INV        m570(.A(mai_mai_n591_), .Y(mai_mai_n593_));
  NO4        m571(.A(mai_mai_n207_), .B(mai_mai_n124_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n594_));
  NA2        m572(.A(mai_mai_n594_), .B(mai_mai_n586_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n230_), .B(i_6_), .Y(mai_mai_n596_));
  NO3        m574(.A(mai_mai_n572_), .B(mai_mai_n226_), .C(mai_mai_n23_), .Y(mai_mai_n597_));
  AOI210     m575(.A0(i_1_), .A1(mai_mai_n251_), .B0(mai_mai_n597_), .Y(mai_mai_n598_));
  OAI210     m576(.A0(mai_mai_n598_), .A1(mai_mai_n44_), .B0(mai_mai_n595_), .Y(mai_mai_n599_));
  NA3        m577(.A(mai_mai_n502_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n600_));
  NA2        m578(.A(mai_mai_n133_), .B(i_9_), .Y(mai_mai_n601_));
  NA3        m579(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n603_));
  NA3        m581(.A(mai_mai_n603_), .B(mai_mai_n260_), .C(mai_mai_n44_), .Y(mai_mai_n604_));
  OAI220     m582(.A0(mai_mai_n604_), .A1(mai_mai_n602_), .B0(mai_mai_n601_), .B1(mai_mai_n956_), .Y(mai_mai_n605_));
  NA3        m583(.A(mai_mai_n586_), .B(mai_mai_n304_), .C(i_6_), .Y(mai_mai_n606_));
  NO2        m584(.A(mai_mai_n606_), .B(mai_mai_n23_), .Y(mai_mai_n607_));
  NAi21      m585(.An(mai_mai_n600_), .B(mai_mai_n88_), .Y(mai_mai_n608_));
  NA2        m586(.A(mai_mai_n603_), .B(mai_mai_n260_), .Y(mai_mai_n609_));
  NO2        m587(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n610_));
  NA2        m588(.A(mai_mai_n610_), .B(mai_mai_n24_), .Y(mai_mai_n611_));
  OAI210     m589(.A0(mai_mai_n611_), .A1(mai_mai_n609_), .B0(mai_mai_n608_), .Y(mai_mai_n612_));
  OR3        m590(.A(mai_mai_n612_), .B(mai_mai_n607_), .C(mai_mai_n605_), .Y(mai_mai_n613_));
  NO3        m591(.A(mai_mai_n613_), .B(mai_mai_n599_), .C(mai_mai_n593_), .Y(mai_mai_n614_));
  NO2        m592(.A(mai_mai_n230_), .B(mai_mai_n98_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n615_), .B(mai_mai_n580_), .Y(mai_mai_n616_));
  NA2        m594(.A(mai_mai_n616_), .B(i_1_), .Y(mai_mai_n617_));
  NO2        m595(.A(mai_mai_n617_), .B(mai_mai_n574_), .Y(mai_mai_n618_));
  NO2        m596(.A(mai_mai_n395_), .B(mai_mai_n82_), .Y(mai_mai_n619_));
  NA2        m597(.A(mai_mai_n618_), .B(mai_mai_n46_), .Y(mai_mai_n620_));
  NO2        m598(.A(i_8_), .B(mai_mai_n112_), .Y(mai_mai_n621_));
  AN2        m599(.A(mai_mai_n621_), .B(mai_mai_n508_), .Y(mai_mai_n622_));
  NO2        m600(.A(mai_mai_n226_), .B(mai_mai_n44_), .Y(mai_mai_n623_));
  NO3        m601(.A(mai_mai_n623_), .B(mai_mai_n297_), .C(mai_mai_n231_), .Y(mai_mai_n624_));
  NO2        m602(.A(mai_mai_n113_), .B(mai_mai_n37_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n625_), .B(i_6_), .Y(mai_mai_n626_));
  NO2        m604(.A(mai_mai_n82_), .B(i_9_), .Y(mai_mai_n627_));
  NO2        m605(.A(mai_mai_n627_), .B(mai_mai_n60_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n628_), .B(mai_mai_n587_), .Y(mai_mai_n629_));
  NO4        m607(.A(mai_mai_n629_), .B(mai_mai_n626_), .C(mai_mai_n624_), .D(i_4_), .Y(mai_mai_n630_));
  NA2        m608(.A(i_1_), .B(i_3_), .Y(mai_mai_n631_));
  NO2        m609(.A(mai_mai_n432_), .B(mai_mai_n89_), .Y(mai_mai_n632_));
  AOI210     m610(.A0(mai_mai_n623_), .A1(mai_mai_n538_), .B0(mai_mai_n632_), .Y(mai_mai_n633_));
  NO2        m611(.A(mai_mai_n633_), .B(mai_mai_n631_), .Y(mai_mai_n634_));
  NO3        m612(.A(mai_mai_n634_), .B(mai_mai_n630_), .C(mai_mai_n622_), .Y(mai_mai_n635_));
  NA4        m613(.A(mai_mai_n635_), .B(mai_mai_n620_), .C(mai_mai_n614_), .D(mai_mai_n589_), .Y(mai_mai_n636_));
  NO3        m614(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n637_));
  NOi21      m615(.An(mai_mai_n637_), .B(i_10_), .Y(mai_mai_n638_));
  OA210      m616(.A0(mai_mai_n638_), .A1(mai_mai_n239_), .B0(mai_mai_n82_), .Y(mai_mai_n639_));
  NA2        m617(.A(mai_mai_n351_), .B(mai_mai_n350_), .Y(mai_mai_n640_));
  NA3        m618(.A(mai_mai_n452_), .B(mai_mai_n487_), .C(mai_mai_n46_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n641_), .B(mai_mai_n640_), .Y(mai_mai_n642_));
  OAI210     m620(.A0(mai_mai_n642_), .A1(mai_mai_n639_), .B0(i_1_), .Y(mai_mai_n643_));
  AOI210     m621(.A0(mai_mai_n260_), .A1(mai_mai_n94_), .B0(i_1_), .Y(mai_mai_n644_));
  NO2        m622(.A(mai_mai_n349_), .B(i_2_), .Y(mai_mai_n645_));
  NA2        m623(.A(mai_mai_n645_), .B(mai_mai_n644_), .Y(mai_mai_n646_));
  OAI210     m624(.A0(mai_mai_n606_), .A1(mai_mai_n428_), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  INV        m625(.A(mai_mai_n647_), .Y(mai_mai_n648_));
  AOI210     m626(.A0(mai_mai_n648_), .A1(mai_mai_n643_), .B0(i_13_), .Y(mai_mai_n649_));
  OR2        m627(.A(i_11_), .B(i_7_), .Y(mai_mai_n650_));
  NO2        m628(.A(mai_mai_n52_), .B(i_12_), .Y(mai_mai_n651_));
  AOI220     m629(.A0(i_7_), .A1(mai_mai_n619_), .B0(mai_mai_n239_), .B1(mai_mai_n127_), .Y(mai_mai_n652_));
  OAI220     m630(.A0(mai_mai_n652_), .A1(mai_mai_n41_), .B0(mai_mai_n955_), .B1(mai_mai_n89_), .Y(mai_mai_n653_));
  INV        m631(.A(mai_mai_n653_), .Y(mai_mai_n654_));
  AOI210     m632(.A0(mai_mai_n428_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n655_));
  NOi31      m633(.An(mai_mai_n655_), .B(mai_mai_n557_), .C(mai_mai_n44_), .Y(mai_mai_n656_));
  NA2        m634(.A(mai_mai_n123_), .B(i_13_), .Y(mai_mai_n657_));
  NO2        m635(.A(mai_mai_n602_), .B(mai_mai_n112_), .Y(mai_mai_n658_));
  INV        m636(.A(mai_mai_n658_), .Y(mai_mai_n659_));
  OAI220     m637(.A0(mai_mai_n659_), .A1(mai_mai_n68_), .B0(mai_mai_n657_), .B1(mai_mai_n644_), .Y(mai_mai_n660_));
  NA2        m638(.A(mai_mai_n26_), .B(mai_mai_n186_), .Y(mai_mai_n661_));
  NA2        m639(.A(mai_mai_n661_), .B(i_7_), .Y(mai_mai_n662_));
  NO3        m640(.A(mai_mai_n447_), .B(mai_mai_n230_), .C(mai_mai_n82_), .Y(mai_mai_n663_));
  NA2        m641(.A(mai_mai_n663_), .B(mai_mai_n662_), .Y(mai_mai_n664_));
  AOI220     m642(.A0(mai_mai_n366_), .A1(mai_mai_n603_), .B0(mai_mai_n88_), .B1(mai_mai_n99_), .Y(mai_mai_n665_));
  OAI220     m643(.A0(mai_mai_n665_), .A1(mai_mai_n561_), .B0(mai_mai_n664_), .B1(mai_mai_n576_), .Y(mai_mai_n666_));
  NO3        m644(.A(mai_mai_n666_), .B(mai_mai_n660_), .C(mai_mai_n656_), .Y(mai_mai_n667_));
  OR2        m645(.A(i_11_), .B(i_6_), .Y(mai_mai_n668_));
  NA3        m646(.A(mai_mai_n560_), .B(mai_mai_n661_), .C(i_7_), .Y(mai_mai_n669_));
  AOI210     m647(.A0(mai_mai_n669_), .A1(mai_mai_n659_), .B0(mai_mai_n668_), .Y(mai_mai_n670_));
  NA3        m648(.A(mai_mai_n389_), .B(mai_mai_n565_), .C(mai_mai_n94_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n592_), .B(i_13_), .Y(mai_mai_n672_));
  NAi21      m650(.An(i_11_), .B(i_12_), .Y(mai_mai_n673_));
  NOi41      m651(.An(mai_mai_n108_), .B(mai_mai_n673_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n674_));
  INV        m652(.A(mai_mai_n674_), .Y(mai_mai_n675_));
  NA3        m653(.A(mai_mai_n675_), .B(mai_mai_n672_), .C(mai_mai_n671_), .Y(mai_mai_n676_));
  OAI210     m654(.A0(mai_mai_n676_), .A1(mai_mai_n670_), .B0(mai_mai_n60_), .Y(mai_mai_n677_));
  NO2        m655(.A(i_2_), .B(i_12_), .Y(mai_mai_n678_));
  NA2        m656(.A(mai_mai_n348_), .B(mai_mai_n678_), .Y(mai_mai_n679_));
  NO3        m657(.A(i_9_), .B(mai_mai_n364_), .C(mai_mai_n560_), .Y(mai_mai_n680_));
  NA2        m658(.A(mai_mai_n680_), .B(mai_mai_n348_), .Y(mai_mai_n681_));
  NO2        m659(.A(mai_mai_n124_), .B(i_2_), .Y(mai_mai_n682_));
  NA2        m660(.A(mai_mai_n682_), .B(mai_mai_n587_), .Y(mai_mai_n683_));
  NA3        m661(.A(mai_mai_n683_), .B(mai_mai_n681_), .C(mai_mai_n679_), .Y(mai_mai_n684_));
  NA3        m662(.A(mai_mai_n684_), .B(mai_mai_n45_), .C(mai_mai_n218_), .Y(mai_mai_n685_));
  NA4        m663(.A(mai_mai_n685_), .B(mai_mai_n677_), .C(mai_mai_n667_), .D(mai_mai_n654_), .Y(mai_mai_n686_));
  OR4        m664(.A(mai_mai_n686_), .B(mai_mai_n649_), .C(mai_mai_n636_), .D(mai_mai_n579_), .Y(mai5));
  NA2        m665(.A(mai_mai_n616_), .B(mai_mai_n262_), .Y(mai_mai_n688_));
  AN2        m666(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n689_));
  NA3        m667(.A(mai_mai_n689_), .B(mai_mai_n678_), .C(mai_mai_n105_), .Y(mai_mai_n690_));
  NO2        m668(.A(mai_mai_n561_), .B(i_11_), .Y(mai_mai_n691_));
  NA2        m669(.A(mai_mai_n83_), .B(mai_mai_n691_), .Y(mai_mai_n692_));
  NA3        m670(.A(mai_mai_n692_), .B(mai_mai_n690_), .C(mai_mai_n688_), .Y(mai_mai_n693_));
  NO3        m671(.A(i_11_), .B(mai_mai_n230_), .C(i_13_), .Y(mai_mai_n694_));
  NO2        m672(.A(mai_mai_n120_), .B(mai_mai_n23_), .Y(mai_mai_n695_));
  NA2        m673(.A(i_12_), .B(i_8_), .Y(mai_mai_n696_));
  INV        m674(.A(mai_mai_n427_), .Y(mai_mai_n697_));
  AOI220     m675(.A0(mai_mai_n304_), .A1(mai_mai_n539_), .B0(i_12_), .B1(mai_mai_n695_), .Y(mai_mai_n698_));
  INV        m676(.A(mai_mai_n698_), .Y(mai_mai_n699_));
  NO2        m677(.A(mai_mai_n699_), .B(mai_mai_n693_), .Y(mai_mai_n700_));
  INV        m678(.A(mai_mai_n165_), .Y(mai_mai_n701_));
  INV        m679(.A(mai_mai_n239_), .Y(mai_mai_n702_));
  OAI210     m680(.A0(mai_mai_n645_), .A1(mai_mai_n429_), .B0(mai_mai_n108_), .Y(mai_mai_n703_));
  AOI210     m681(.A0(mai_mai_n703_), .A1(mai_mai_n702_), .B0(mai_mai_n701_), .Y(mai_mai_n704_));
  INV        m682(.A(mai_mai_n399_), .Y(mai_mai_n705_));
  NA2        m683(.A(mai_mai_n705_), .B(i_2_), .Y(mai_mai_n706_));
  INV        m684(.A(mai_mai_n706_), .Y(mai_mai_n707_));
  AOI210     m685(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n396_), .Y(mai_mai_n708_));
  AOI210     m686(.A0(mai_mai_n708_), .A1(mai_mai_n707_), .B0(mai_mai_n704_), .Y(mai_mai_n709_));
  NO2        m687(.A(mai_mai_n183_), .B(mai_mai_n121_), .Y(mai_mai_n710_));
  OAI210     m688(.A0(mai_mai_n710_), .A1(mai_mai_n695_), .B0(i_2_), .Y(mai_mai_n711_));
  INV        m689(.A(mai_mai_n166_), .Y(mai_mai_n712_));
  NO3        m690(.A(mai_mai_n581_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n713_));
  AOI210     m691(.A0(mai_mai_n712_), .A1(mai_mai_n83_), .B0(mai_mai_n713_), .Y(mai_mai_n714_));
  AOI210     m692(.A0(mai_mai_n714_), .A1(mai_mai_n711_), .B0(mai_mai_n186_), .Y(mai_mai_n715_));
  OA210      m693(.A0(mai_mai_n582_), .A1(mai_mai_n122_), .B0(i_13_), .Y(mai_mai_n716_));
  INV        m694(.A(mai_mai_n146_), .Y(mai_mai_n717_));
  NO2        m695(.A(mai_mai_n717_), .B(mai_mai_n353_), .Y(mai_mai_n718_));
  AOI210     m696(.A0(mai_mai_n199_), .A1(mai_mai_n143_), .B0(mai_mai_n487_), .Y(mai_mai_n719_));
  NA2        m697(.A(mai_mai_n719_), .B(mai_mai_n399_), .Y(mai_mai_n720_));
  NO2        m698(.A(mai_mai_n99_), .B(mai_mai_n44_), .Y(mai_mai_n721_));
  INV        m699(.A(mai_mai_n290_), .Y(mai_mai_n722_));
  NA4        m700(.A(mai_mai_n722_), .B(mai_mai_n294_), .C(mai_mai_n120_), .D(mai_mai_n42_), .Y(mai_mai_n723_));
  OAI210     m701(.A0(mai_mai_n723_), .A1(mai_mai_n721_), .B0(mai_mai_n720_), .Y(mai_mai_n724_));
  NO4        m702(.A(mai_mai_n724_), .B(mai_mai_n718_), .C(mai_mai_n716_), .D(mai_mai_n715_), .Y(mai_mai_n725_));
  NO2        m703(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n726_), .B(mai_mai_n122_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n727_), .B(mai_mai_n558_), .Y(mai_mai_n728_));
  NA2        m706(.A(mai_mai_n728_), .B(mai_mai_n36_), .Y(mai_mai_n729_));
  NA4        m707(.A(mai_mai_n729_), .B(mai_mai_n725_), .C(mai_mai_n709_), .D(mai_mai_n700_), .Y(mai6));
  NO3        m708(.A(i_9_), .B(mai_mai_n296_), .C(i_1_), .Y(mai_mai_n731_));
  NO2        m709(.A(mai_mai_n178_), .B(mai_mai_n134_), .Y(mai_mai_n732_));
  OAI210     m710(.A0(mai_mai_n732_), .A1(mai_mai_n731_), .B0(mai_mai_n682_), .Y(mai_mai_n733_));
  NO2        m711(.A(mai_mai_n213_), .B(mai_mai_n456_), .Y(mai_mai_n734_));
  INV        m712(.A(mai_mai_n316_), .Y(mai_mai_n735_));
  AO210      m713(.A0(mai_mai_n735_), .A1(mai_mai_n733_), .B0(i_12_), .Y(mai_mai_n736_));
  NA2        m714(.A(mai_mai_n354_), .B(mai_mai_n321_), .Y(mai_mai_n737_));
  NA2        m715(.A(mai_mai_n546_), .B(mai_mai_n60_), .Y(mai_mai_n738_));
  NA2        m716(.A(mai_mai_n638_), .B(mai_mai_n68_), .Y(mai_mai_n739_));
  NA3        m717(.A(mai_mai_n739_), .B(mai_mai_n738_), .C(mai_mai_n737_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n740_), .B(mai_mai_n70_), .Y(mai_mai_n741_));
  INV        m719(.A(mai_mai_n315_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n72_), .B(mai_mai_n127_), .Y(mai_mai_n743_));
  INV        m721(.A(mai_mai_n120_), .Y(mai_mai_n744_));
  NA2        m722(.A(mai_mai_n744_), .B(mai_mai_n46_), .Y(mai_mai_n745_));
  AOI210     m723(.A0(mai_mai_n745_), .A1(mai_mai_n743_), .B0(mai_mai_n742_), .Y(mai_mai_n746_));
  NO2        m724(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n747_));
  NA3        m725(.A(mai_mai_n747_), .B(mai_mai_n444_), .C(mai_mai_n370_), .Y(mai_mai_n748_));
  OAI210     m726(.A0(mai_mai_n637_), .A1(mai_mai_n530_), .B0(mai_mai_n529_), .Y(mai_mai_n749_));
  NA2        m727(.A(mai_mai_n749_), .B(mai_mai_n748_), .Y(mai_mai_n750_));
  OR2        m728(.A(mai_mai_n750_), .B(mai_mai_n746_), .Y(mai_mai_n751_));
  NO2        m729(.A(mai_mai_n650_), .B(i_2_), .Y(mai_mai_n752_));
  NA2        m730(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n753_));
  NO2        m731(.A(mai_mai_n753_), .B(mai_mai_n388_), .Y(mai_mai_n754_));
  NA2        m732(.A(mai_mai_n754_), .B(mai_mai_n752_), .Y(mai_mai_n755_));
  AO210      m733(.A0(mai_mai_n342_), .A1(mai_mai_n334_), .B0(mai_mai_n376_), .Y(mai_mai_n756_));
  NA3        m734(.A(mai_mai_n756_), .B(mai_mai_n247_), .C(i_7_), .Y(mai_mai_n757_));
  OR2        m735(.A(mai_mai_n582_), .B(mai_mai_n429_), .Y(mai_mai_n758_));
  NA2        m736(.A(mai_mai_n758_), .B(mai_mai_n142_), .Y(mai_mai_n759_));
  AO210      m737(.A0(mai_mai_n462_), .A1(mai_mai_n697_), .B0(mai_mai_n36_), .Y(mai_mai_n760_));
  NA4        m738(.A(mai_mai_n760_), .B(mai_mai_n759_), .C(mai_mai_n757_), .D(mai_mai_n755_), .Y(mai_mai_n761_));
  NO2        m739(.A(i_6_), .B(i_11_), .Y(mai_mai_n762_));
  AOI220     m740(.A0(mai_mai_n762_), .A1(mai_mai_n529_), .B0(mai_mai_n734_), .B1(mai_mai_n662_), .Y(mai_mai_n763_));
  NA3        m741(.A(mai_mai_n353_), .B(mai_mai_n232_), .C(mai_mai_n142_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n376_), .B(mai_mai_n67_), .Y(mai_mai_n765_));
  NA4        m743(.A(mai_mai_n765_), .B(mai_mai_n764_), .C(mai_mai_n763_), .D(mai_mai_n564_), .Y(mai_mai_n766_));
  AOI210     m744(.A0(mai_mai_n429_), .A1(mai_mai_n427_), .B0(mai_mai_n528_), .Y(mai_mai_n767_));
  NO2        m745(.A(mai_mai_n572_), .B(mai_mai_n99_), .Y(mai_mai_n768_));
  OAI210     m746(.A0(mai_mai_n768_), .A1(mai_mai_n109_), .B0(mai_mai_n386_), .Y(mai_mai_n769_));
  INV        m747(.A(mai_mai_n549_), .Y(mai_mai_n770_));
  NA3        m748(.A(mai_mai_n770_), .B(mai_mai_n315_), .C(i_7_), .Y(mai_mai_n771_));
  NA3        m749(.A(mai_mai_n771_), .B(mai_mai_n769_), .C(mai_mai_n767_), .Y(mai_mai_n772_));
  NO4        m750(.A(mai_mai_n772_), .B(mai_mai_n766_), .C(mai_mai_n761_), .D(mai_mai_n751_), .Y(mai_mai_n773_));
  NA4        m751(.A(mai_mai_n773_), .B(mai_mai_n741_), .C(mai_mai_n736_), .D(mai_mai_n360_), .Y(mai3));
  NA2        m752(.A(i_6_), .B(i_7_), .Y(mai_mai_n775_));
  NO2        m753(.A(mai_mai_n775_), .B(i_0_), .Y(mai_mai_n776_));
  NO2        m754(.A(i_11_), .B(mai_mai_n230_), .Y(mai_mai_n777_));
  NA2        m755(.A(mai_mai_n278_), .B(mai_mai_n777_), .Y(mai_mai_n778_));
  NO2        m756(.A(mai_mai_n778_), .B(mai_mai_n186_), .Y(mai_mai_n779_));
  NO3        m757(.A(mai_mai_n430_), .B(mai_mai_n86_), .C(mai_mai_n44_), .Y(mai_mai_n780_));
  OA210      m758(.A0(mai_mai_n780_), .A1(mai_mai_n779_), .B0(mai_mai_n168_), .Y(mai_mai_n781_));
  NA2        m759(.A(mai_mai_n764_), .B(mai_mai_n352_), .Y(mai_mai_n782_));
  NA2        m760(.A(mai_mai_n782_), .B(mai_mai_n40_), .Y(mai_mai_n783_));
  AN2        m761(.A(mai_mai_n431_), .B(mai_mai_n53_), .Y(mai_mai_n784_));
  AOI210     m762(.A0(mai_mai_n957_), .A1(mai_mai_n783_), .B0(mai_mai_n48_), .Y(mai_mai_n785_));
  NO4        m763(.A(mai_mai_n357_), .B(mai_mai_n363_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n786_));
  INV        m764(.A(mai_mai_n786_), .Y(mai_mai_n787_));
  NA2        m765(.A(mai_mai_n655_), .B(mai_mai_n627_), .Y(mai_mai_n788_));
  NA2        m766(.A(mai_mai_n319_), .B(i_5_), .Y(mai_mai_n789_));
  OAI220     m767(.A0(mai_mai_n789_), .A1(mai_mai_n788_), .B0(mai_mai_n787_), .B1(mai_mai_n60_), .Y(mai_mai_n790_));
  NOi21      m768(.An(i_5_), .B(i_9_), .Y(mai_mai_n791_));
  NA2        m769(.A(mai_mai_n791_), .B(mai_mai_n426_), .Y(mai_mai_n792_));
  NO3        m770(.A(mai_mai_n392_), .B(mai_mai_n260_), .C(mai_mai_n70_), .Y(mai_mai_n793_));
  NO2        m771(.A(mai_mai_n169_), .B(mai_mai_n143_), .Y(mai_mai_n794_));
  AOI210     m772(.A0(mai_mai_n794_), .A1(mai_mai_n238_), .B0(mai_mai_n793_), .Y(mai_mai_n795_));
  NO2        m773(.A(mai_mai_n795_), .B(mai_mai_n959_), .Y(mai_mai_n796_));
  NO4        m774(.A(mai_mai_n796_), .B(mai_mai_n790_), .C(mai_mai_n785_), .D(mai_mai_n781_), .Y(mai_mai_n797_));
  NA2        m775(.A(mai_mai_n178_), .B(mai_mai_n24_), .Y(mai_mai_n798_));
  NA2        m776(.A(mai_mai_n301_), .B(mai_mai_n125_), .Y(mai_mai_n799_));
  NAi21      m777(.An(mai_mai_n156_), .B(i_5_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n799_), .B(mai_mai_n378_), .Y(mai_mai_n801_));
  INV        m779(.A(mai_mai_n801_), .Y(mai_mai_n802_));
  NO2        m780(.A(mai_mai_n370_), .B(mai_mai_n282_), .Y(mai_mai_n803_));
  NA2        m781(.A(mai_mai_n803_), .B(mai_mai_n658_), .Y(mai_mai_n804_));
  NO4        m782(.A(mai_mai_n548_), .B(mai_mai_n207_), .C(mai_mai_n396_), .D(mai_mai_n388_), .Y(mai_mai_n805_));
  AN2        m783(.A(mai_mai_n93_), .B(mai_mai_n237_), .Y(mai_mai_n806_));
  NA2        m784(.A(mai_mai_n694_), .B(mai_mai_n316_), .Y(mai_mai_n807_));
  AOI210     m785(.A0(mai_mai_n452_), .A1(mai_mai_n83_), .B0(mai_mai_n55_), .Y(mai_mai_n808_));
  OAI220     m786(.A0(mai_mai_n808_), .A1(mai_mai_n807_), .B0(mai_mai_n611_), .B1(mai_mai_n504_), .Y(mai_mai_n809_));
  NO2        m787(.A(mai_mai_n245_), .B(mai_mai_n147_), .Y(mai_mai_n810_));
  NA2        m788(.A(i_0_), .B(i_10_), .Y(mai_mai_n811_));
  AN2        m789(.A(mai_mai_n810_), .B(i_6_), .Y(mai_mai_n812_));
  AOI220     m790(.A0(mai_mai_n319_), .A1(mai_mai_n95_), .B0(mai_mai_n178_), .B1(mai_mai_n80_), .Y(mai_mai_n813_));
  NA2        m791(.A(mai_mai_n533_), .B(i_4_), .Y(mai_mai_n814_));
  NA2        m792(.A(mai_mai_n181_), .B(mai_mai_n195_), .Y(mai_mai_n815_));
  OAI220     m793(.A0(mai_mai_n815_), .A1(mai_mai_n807_), .B0(mai_mai_n814_), .B1(mai_mai_n813_), .Y(mai_mai_n816_));
  NO4        m794(.A(mai_mai_n816_), .B(mai_mai_n812_), .C(mai_mai_n809_), .D(mai_mai_n806_), .Y(mai_mai_n817_));
  NA3        m795(.A(mai_mai_n817_), .B(mai_mai_n804_), .C(mai_mai_n802_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n819_));
  NA2        m797(.A(mai_mai_n374_), .B(mai_mai_n173_), .Y(mai_mai_n820_));
  NA2        m798(.A(mai_mai_n820_), .B(mai_mai_n154_), .Y(mai_mai_n821_));
  NO2        m799(.A(mai_mai_n169_), .B(i_0_), .Y(mai_mai_n822_));
  INV        m800(.A(mai_mai_n822_), .Y(mai_mai_n823_));
  NA2        m801(.A(mai_mai_n444_), .B(mai_mai_n224_), .Y(mai_mai_n824_));
  INV        m802(.A(mai_mai_n385_), .Y(mai_mai_n825_));
  OAI220     m803(.A0(mai_mai_n825_), .A1(mai_mai_n792_), .B0(mai_mai_n824_), .B1(mai_mai_n823_), .Y(mai_mai_n826_));
  NO2        m804(.A(mai_mai_n826_), .B(mai_mai_n821_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n610_), .B(mai_mai_n117_), .Y(mai_mai_n828_));
  NO2        m806(.A(i_6_), .B(mai_mai_n828_), .Y(mai_mai_n829_));
  AOI210     m807(.A0(mai_mai_n428_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n830_));
  NA2        m808(.A(mai_mai_n165_), .B(mai_mai_n100_), .Y(mai_mai_n831_));
  NOi32      m809(.An(mai_mai_n830_), .Bn(mai_mai_n181_), .C(mai_mai_n831_), .Y(mai_mai_n832_));
  NO2        m810(.A(mai_mai_n832_), .B(mai_mai_n829_), .Y(mai_mai_n833_));
  NOi21      m811(.An(i_7_), .B(i_5_), .Y(mai_mai_n834_));
  NOi31      m812(.An(mai_mai_n834_), .B(i_0_), .C(mai_mai_n673_), .Y(mai_mai_n835_));
  NA3        m813(.A(mai_mai_n835_), .B(mai_mai_n364_), .C(i_6_), .Y(mai_mai_n836_));
  OA210      m814(.A0(mai_mai_n831_), .A1(mai_mai_n485_), .B0(mai_mai_n836_), .Y(mai_mai_n837_));
  NO3        m815(.A(mai_mai_n381_), .B(mai_mai_n345_), .C(mai_mai_n341_), .Y(mai_mai_n838_));
  NO2        m816(.A(mai_mai_n254_), .B(mai_mai_n305_), .Y(mai_mai_n839_));
  NO2        m817(.A(mai_mai_n673_), .B(mai_mai_n249_), .Y(mai_mai_n840_));
  AOI210     m818(.A0(mai_mai_n840_), .A1(mai_mai_n839_), .B0(mai_mai_n838_), .Y(mai_mai_n841_));
  NA4        m819(.A(mai_mai_n841_), .B(mai_mai_n837_), .C(mai_mai_n833_), .D(mai_mai_n827_), .Y(mai_mai_n842_));
  NO2        m820(.A(mai_mai_n798_), .B(mai_mai_n233_), .Y(mai_mai_n843_));
  AN2        m821(.A(mai_mai_n318_), .B(mai_mai_n316_), .Y(mai_mai_n844_));
  NA2        m822(.A(mai_mai_n843_), .B(i_10_), .Y(mai_mai_n845_));
  OA210      m823(.A0(mai_mai_n444_), .A1(mai_mai_n216_), .B0(mai_mai_n443_), .Y(mai_mai_n846_));
  NA3        m824(.A(mai_mai_n443_), .B(mai_mai_n389_), .C(mai_mai_n45_), .Y(mai_mai_n847_));
  OAI210     m825(.A0(mai_mai_n800_), .A1(i_6_), .B0(mai_mai_n847_), .Y(mai_mai_n848_));
  INV        m826(.A(mai_mai_n180_), .Y(mai_mai_n849_));
  AOI220     m827(.A0(mai_mai_n849_), .A1(mai_mai_n444_), .B0(mai_mai_n848_), .B1(mai_mai_n70_), .Y(mai_mai_n850_));
  NA2        m828(.A(mai_mai_n89_), .B(mai_mai_n44_), .Y(mai_mai_n851_));
  NO2        m829(.A(mai_mai_n72_), .B(mai_mai_n696_), .Y(mai_mai_n852_));
  NA2        m830(.A(mai_mai_n852_), .B(mai_mai_n851_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n853_), .B(mai_mai_n47_), .Y(mai_mai_n854_));
  NO2        m832(.A(mai_mai_n559_), .B(mai_mai_n102_), .Y(mai_mai_n855_));
  NA2        m833(.A(mai_mai_n855_), .B(i_0_), .Y(mai_mai_n856_));
  NO2        m834(.A(mai_mai_n856_), .B(mai_mai_n82_), .Y(mai_mai_n857_));
  NO3        m835(.A(mai_mai_n857_), .B(mai_mai_n854_), .C(mai_mai_n489_), .Y(mai_mai_n858_));
  NA3        m836(.A(mai_mai_n858_), .B(mai_mai_n850_), .C(mai_mai_n845_), .Y(mai_mai_n859_));
  NO3        m837(.A(mai_mai_n859_), .B(mai_mai_n842_), .C(mai_mai_n818_), .Y(mai_mai_n860_));
  NO2        m838(.A(i_0_), .B(mai_mai_n673_), .Y(mai_mai_n861_));
  NA2        m839(.A(mai_mai_n70_), .B(mai_mai_n44_), .Y(mai_mai_n862_));
  INV        m840(.A(mai_mai_n862_), .Y(mai_mai_n863_));
  NO3        m841(.A(mai_mai_n102_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n864_));
  AO220      m842(.A0(mai_mai_n864_), .A1(mai_mai_n863_), .B0(mai_mai_n861_), .B1(mai_mai_n168_), .Y(mai_mai_n865_));
  AOI210     m843(.A0(mai_mai_n738_), .A1(mai_mai_n640_), .B0(mai_mai_n831_), .Y(mai_mai_n866_));
  AOI210     m844(.A0(mai_mai_n865_), .A1(mai_mai_n331_), .B0(mai_mai_n866_), .Y(mai_mai_n867_));
  NA3        m845(.A(mai_mai_n141_), .B(mai_mai_n627_), .C(mai_mai_n70_), .Y(mai_mai_n868_));
  NO2        m846(.A(mai_mai_n749_), .B(mai_mai_n381_), .Y(mai_mai_n869_));
  NA3        m847(.A(mai_mai_n776_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n870_));
  NA2        m848(.A(mai_mai_n777_), .B(i_9_), .Y(mai_mai_n871_));
  AOI210     m849(.A0(mai_mai_n870_), .A1(mai_mai_n467_), .B0(mai_mai_n871_), .Y(mai_mai_n872_));
  NA2        m850(.A(mai_mai_n238_), .B(mai_mai_n223_), .Y(mai_mai_n873_));
  NO2        m851(.A(mai_mai_n873_), .B(mai_mai_n147_), .Y(mai_mai_n874_));
  NO3        m852(.A(mai_mai_n874_), .B(mai_mai_n872_), .C(mai_mai_n869_), .Y(mai_mai_n875_));
  NA3        m853(.A(mai_mai_n875_), .B(mai_mai_n868_), .C(mai_mai_n867_), .Y(mai_mai_n876_));
  NA2        m854(.A(mai_mai_n844_), .B(mai_mai_n353_), .Y(mai_mai_n877_));
  AOI210     m855(.A0(mai_mai_n289_), .A1(mai_mai_n156_), .B0(mai_mai_n877_), .Y(mai_mai_n878_));
  NA2        m856(.A(mai_mai_n40_), .B(mai_mai_n44_), .Y(mai_mai_n879_));
  NA2        m857(.A(mai_mai_n819_), .B(mai_mai_n457_), .Y(mai_mai_n880_));
  AOI210     m858(.A0(mai_mai_n879_), .A1(mai_mai_n156_), .B0(mai_mai_n880_), .Y(mai_mai_n881_));
  NO2        m859(.A(mai_mai_n881_), .B(mai_mai_n878_), .Y(mai_mai_n882_));
  NO3        m860(.A(mai_mai_n811_), .B(mai_mai_n791_), .C(mai_mai_n183_), .Y(mai_mai_n883_));
  AOI220     m861(.A0(mai_mai_n883_), .A1(i_11_), .B0(mai_mai_n534_), .B1(mai_mai_n72_), .Y(mai_mai_n884_));
  NO3        m862(.A(mai_mai_n201_), .B(mai_mai_n363_), .C(i_0_), .Y(mai_mai_n885_));
  OAI210     m863(.A0(mai_mai_n885_), .A1(mai_mai_n73_), .B0(i_13_), .Y(mai_mai_n886_));
  INV        m864(.A(mai_mai_n210_), .Y(mai_mai_n887_));
  OAI220     m865(.A0(mai_mai_n497_), .A1(mai_mai_n134_), .B0(mai_mai_n596_), .B1(mai_mai_n576_), .Y(mai_mai_n888_));
  NA3        m866(.A(mai_mai_n888_), .B(i_7_), .C(mai_mai_n887_), .Y(mai_mai_n889_));
  NA4        m867(.A(mai_mai_n889_), .B(mai_mai_n886_), .C(mai_mai_n884_), .D(mai_mai_n882_), .Y(mai_mai_n890_));
  INV        m868(.A(mai_mai_n106_), .Y(mai_mai_n891_));
  NA2        m869(.A(mai_mai_n834_), .B(mai_mai_n457_), .Y(mai_mai_n892_));
  INV        m870(.A(mai_mai_n170_), .Y(mai_mai_n893_));
  OA220      m871(.A0(mai_mai_n893_), .A1(mai_mai_n892_), .B0(mai_mai_n891_), .B1(i_5_), .Y(mai_mai_n894_));
  AOI210     m872(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n169_), .Y(mai_mai_n895_));
  NA2        m873(.A(mai_mai_n895_), .B(mai_mai_n846_), .Y(mai_mai_n896_));
  NA3        m874(.A(mai_mai_n370_), .B(mai_mai_n320_), .C(mai_mai_n214_), .Y(mai_mai_n897_));
  INV        m875(.A(mai_mai_n897_), .Y(mai_mai_n898_));
  NOi31      m876(.An(mai_mai_n369_), .B(mai_mai_n862_), .C(mai_mai_n233_), .Y(mai_mai_n899_));
  NO2        m877(.A(mai_mai_n899_), .B(mai_mai_n898_), .Y(mai_mai_n900_));
  NA4        m878(.A(mai_mai_n900_), .B(mai_mai_n441_), .C(mai_mai_n896_), .D(mai_mai_n894_), .Y(mai_mai_n901_));
  NA3        m879(.A(mai_mai_n294_), .B(i_5_), .C(mai_mai_n186_), .Y(mai_mai_n902_));
  NAi31      m880(.An(mai_mai_n235_), .B(mai_mai_n902_), .C(mai_mai_n236_), .Y(mai_mai_n903_));
  NO4        m881(.A(mai_mai_n233_), .B(mai_mai_n201_), .C(i_0_), .D(i_12_), .Y(mai_mai_n904_));
  NA2        m882(.A(mai_mai_n904_), .B(mai_mai_n903_), .Y(mai_mai_n905_));
  AN2        m883(.A(mai_mai_n811_), .B(mai_mai_n147_), .Y(mai_mai_n906_));
  NO4        m884(.A(mai_mai_n906_), .B(i_12_), .C(mai_mai_n600_), .D(mai_mai_n127_), .Y(mai_mai_n907_));
  NA2        m885(.A(mai_mai_n907_), .B(mai_mai_n210_), .Y(mai_mai_n908_));
  NA3        m886(.A(mai_mai_n95_), .B(mai_mai_n538_), .C(i_11_), .Y(mai_mai_n909_));
  NA2        m887(.A(mai_mai_n834_), .B(mai_mai_n440_), .Y(mai_mai_n910_));
  NA2        m888(.A(mai_mai_n61_), .B(mai_mai_n98_), .Y(mai_mai_n911_));
  OAI220     m889(.A0(mai_mai_n911_), .A1(mai_mai_n902_), .B0(mai_mai_n910_), .B1(mai_mai_n628_), .Y(mai_mai_n912_));
  NA2        m890(.A(mai_mai_n912_), .B(mai_mai_n822_), .Y(mai_mai_n913_));
  NA3        m891(.A(mai_mai_n913_), .B(mai_mai_n908_), .C(mai_mai_n905_), .Y(mai_mai_n914_));
  NO4        m892(.A(mai_mai_n914_), .B(mai_mai_n901_), .C(mai_mai_n890_), .D(mai_mai_n876_), .Y(mai_mai_n915_));
  OAI210     m893(.A0(mai_mai_n752_), .A1(mai_mai_n747_), .B0(mai_mai_n37_), .Y(mai_mai_n916_));
  NA3        m894(.A(mai_mai_n830_), .B(mai_mai_n348_), .C(i_5_), .Y(mai_mai_n917_));
  NA3        m895(.A(mai_mai_n917_), .B(mai_mai_n916_), .C(mai_mai_n571_), .Y(mai_mai_n918_));
  NA2        m896(.A(mai_mai_n918_), .B(mai_mai_n197_), .Y(mai_mai_n919_));
  BUFFER     m897(.A(mai_mai_n349_), .Y(mai_mai_n920_));
  NA2        m898(.A(mai_mai_n179_), .B(mai_mai_n181_), .Y(mai_mai_n921_));
  AO210      m899(.A0(mai_mai_n920_), .A1(mai_mai_n33_), .B0(mai_mai_n921_), .Y(mai_mai_n922_));
  OAI210     m900(.A0(mai_mai_n575_), .A1(mai_mai_n573_), .B0(mai_mai_n304_), .Y(mai_mai_n923_));
  NAi31      m901(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n924_));
  NO2        m902(.A(mai_mai_n67_), .B(mai_mai_n924_), .Y(mai_mai_n925_));
  NO2        m903(.A(mai_mai_n925_), .B(mai_mai_n597_), .Y(mai_mai_n926_));
  NA3        m904(.A(mai_mai_n926_), .B(mai_mai_n923_), .C(mai_mai_n922_), .Y(mai_mai_n927_));
  NO2        m905(.A(mai_mai_n434_), .B(mai_mai_n260_), .Y(mai_mai_n928_));
  NO4        m906(.A(mai_mai_n226_), .B(mai_mai_n140_), .C(mai_mai_n631_), .D(mai_mai_n37_), .Y(mai_mai_n929_));
  NO3        m907(.A(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n805_), .Y(mai_mai_n930_));
  OAI210     m908(.A0(mai_mai_n909_), .A1(mai_mai_n143_), .B0(mai_mai_n930_), .Y(mai_mai_n931_));
  AOI210     m909(.A0(mai_mai_n927_), .A1(mai_mai_n48_), .B0(mai_mai_n931_), .Y(mai_mai_n932_));
  AOI210     m910(.A0(mai_mai_n932_), .A1(mai_mai_n919_), .B0(mai_mai_n70_), .Y(mai_mai_n933_));
  NO2        m911(.A(mai_mai_n531_), .B(mai_mai_n359_), .Y(mai_mai_n934_));
  NO2        m912(.A(mai_mai_n934_), .B(mai_mai_n701_), .Y(mai_mai_n935_));
  OAI210     m913(.A0(mai_mai_n77_), .A1(mai_mai_n52_), .B0(mai_mai_n105_), .Y(mai_mai_n936_));
  NA2        m914(.A(mai_mai_n936_), .B(mai_mai_n73_), .Y(mai_mai_n937_));
  AOI210     m915(.A0(mai_mai_n895_), .A1(mai_mai_n819_), .B0(mai_mai_n835_), .Y(mai_mai_n938_));
  AOI210     m916(.A0(mai_mai_n938_), .A1(mai_mai_n937_), .B0(mai_mai_n631_), .Y(mai_mai_n939_));
  NA2        m917(.A(mai_mai_n254_), .B(mai_mai_n54_), .Y(mai_mai_n940_));
  NA2        m918(.A(mai_mai_n940_), .B(mai_mai_n73_), .Y(mai_mai_n941_));
  NO2        m919(.A(mai_mai_n941_), .B(mai_mai_n230_), .Y(mai_mai_n942_));
  NA3        m920(.A(mai_mai_n93_), .B(mai_mai_n296_), .C(mai_mai_n31_), .Y(mai_mai_n943_));
  INV        m921(.A(mai_mai_n943_), .Y(mai_mai_n944_));
  NO3        m922(.A(mai_mai_n944_), .B(mai_mai_n942_), .C(mai_mai_n939_), .Y(mai_mai_n945_));
  OAI210     m923(.A0(mai_mai_n960_), .A1(mai_mai_n830_), .B0(mai_mai_n197_), .Y(mai_mai_n946_));
  NA2        m924(.A(mai_mai_n157_), .B(i_5_), .Y(mai_mai_n947_));
  NO2        m925(.A(mai_mai_n946_), .B(mai_mai_n947_), .Y(mai_mai_n948_));
  INV        m926(.A(mai_mai_n948_), .Y(mai_mai_n949_));
  OAI210     m927(.A0(mai_mai_n945_), .A1(i_4_), .B0(mai_mai_n949_), .Y(mai_mai_n950_));
  NO3        m928(.A(mai_mai_n950_), .B(mai_mai_n935_), .C(mai_mai_n933_), .Y(mai_mai_n951_));
  NA4        m929(.A(mai_mai_n951_), .B(mai_mai_n915_), .C(mai_mai_n860_), .D(mai_mai_n797_), .Y(mai4));
  INV        m930(.A(mai_mai_n651_), .Y(mai_mai_n955_));
  INV        m931(.A(i_2_), .Y(mai_mai_n956_));
  INV        m932(.A(mai_mai_n784_), .Y(mai_mai_n957_));
  INV        m933(.A(i_12_), .Y(mai_mai_n958_));
  INV        m934(.A(i_5_), .Y(mai_mai_n959_));
  INV        m935(.A(i_12_), .Y(mai_mai_n960_));
  INV        m936(.A(i_7_), .Y(mai_mai_n961_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(i_1_), .B(i_10_), .Y(men_men_n64_));
  NO2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NAi21      u0043(.An(men_men_n65_), .B(men_men_n61_), .Y(men_men_n66_));
  NA2        u0044(.A(men_men_n51_), .B(i_2_), .Y(men_men_n67_));
  AOI210     u0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n68_));
  NA2        u0046(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO2        u0047(.A(men_men_n69_), .B(men_men_n25_), .Y(men_men_n70_));
  INV        u0048(.A(i_0_), .Y(men_men_n71_));
  NAi21      u0049(.An(i_5_), .B(i_10_), .Y(men_men_n72_));
  NA2        u0050(.A(i_5_), .B(i_9_), .Y(men_men_n73_));
  AOI210     u0051(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n71_), .Y(men_men_n74_));
  NO2        u0052(.A(men_men_n74_), .B(men_men_n70_), .Y(men_men_n75_));
  INV        u0053(.A(men_men_n75_), .Y(men_men_n76_));
  OAI210     u0054(.A0(men_men_n76_), .A1(men_men_n66_), .B0(i_0_), .Y(men_men_n77_));
  NA2        u0055(.A(i_12_), .B(i_5_), .Y(men_men_n78_));
  NA2        u0056(.A(i_2_), .B(i_8_), .Y(men_men_n79_));
  NO2        u0057(.A(men_men_n79_), .B(men_men_n58_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_9_), .Y(men_men_n81_));
  NO2        u0059(.A(i_3_), .B(i_7_), .Y(men_men_n82_));
  INV        u0060(.A(i_6_), .Y(men_men_n83_));
  OR4        u0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n84_));
  NO2        u0062(.A(i_2_), .B(i_7_), .Y(men_men_n85_));
  NAi21      u0063(.An(i_6_), .B(i_10_), .Y(men_men_n86_));
  NA2        u0064(.A(i_6_), .B(i_9_), .Y(men_men_n87_));
  NA2        u0065(.A(i_2_), .B(i_6_), .Y(men_men_n88_));
  NO2        u0066(.A(men_men_n1019_), .B(men_men_n78_), .Y(men_men_n89_));
  AN3        u0067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n90_));
  NAi21      u0068(.An(i_6_), .B(i_11_), .Y(men_men_n91_));
  NO2        u0069(.A(i_5_), .B(i_8_), .Y(men_men_n92_));
  NOi21      u0070(.An(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  AOI220     u0071(.A0(men_men_n93_), .A1(men_men_n62_), .B0(men_men_n90_), .B1(men_men_n32_), .Y(men_men_n94_));
  INV        u0072(.A(i_7_), .Y(men_men_n95_));
  NA2        u0073(.A(men_men_n47_), .B(men_men_n95_), .Y(men_men_n96_));
  NO2        u0074(.A(i_0_), .B(i_5_), .Y(men_men_n97_));
  NO2        u0075(.A(men_men_n97_), .B(men_men_n83_), .Y(men_men_n98_));
  NA2        u0076(.A(i_12_), .B(i_3_), .Y(men_men_n99_));
  INV        u0077(.A(men_men_n99_), .Y(men_men_n100_));
  NA3        u0078(.A(men_men_n100_), .B(men_men_n98_), .C(men_men_n96_), .Y(men_men_n101_));
  NAi21      u0079(.An(i_7_), .B(i_11_), .Y(men_men_n102_));
  AN2        u0080(.A(i_2_), .B(i_10_), .Y(men_men_n103_));
  NO2        u0081(.A(men_men_n103_), .B(i_7_), .Y(men_men_n104_));
  OR2        u0082(.A(men_men_n78_), .B(men_men_n58_), .Y(men_men_n105_));
  NO2        u0083(.A(i_8_), .B(men_men_n95_), .Y(men_men_n106_));
  NO3        u0084(.A(men_men_n106_), .B(men_men_n105_), .C(men_men_n104_), .Y(men_men_n107_));
  NA2        u0085(.A(i_12_), .B(i_7_), .Y(men_men_n108_));
  NO2        u0086(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n109_));
  NA2        u0087(.A(men_men_n109_), .B(i_0_), .Y(men_men_n110_));
  NA2        u0088(.A(i_11_), .B(i_12_), .Y(men_men_n111_));
  OAI210     u0089(.A0(men_men_n110_), .A1(men_men_n108_), .B0(men_men_n111_), .Y(men_men_n112_));
  NO2        u0090(.A(men_men_n112_), .B(men_men_n107_), .Y(men_men_n113_));
  NA3        u0091(.A(men_men_n113_), .B(men_men_n101_), .C(men_men_n94_), .Y(men_men_n114_));
  NOi21      u0092(.An(i_1_), .B(i_5_), .Y(men_men_n115_));
  NA2        u0093(.A(men_men_n115_), .B(i_11_), .Y(men_men_n116_));
  NA2        u0094(.A(men_men_n95_), .B(men_men_n37_), .Y(men_men_n117_));
  NA2        u0095(.A(i_7_), .B(men_men_n25_), .Y(men_men_n118_));
  NA2        u0096(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NO2        u0097(.A(men_men_n119_), .B(men_men_n47_), .Y(men_men_n120_));
  NA2        u0098(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n121_));
  NAi21      u0099(.An(i_3_), .B(i_8_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n122_), .B(men_men_n62_), .Y(men_men_n123_));
  NOi21      u0101(.An(men_men_n123_), .B(men_men_n121_), .Y(men_men_n124_));
  NO2        u0102(.A(i_1_), .B(men_men_n83_), .Y(men_men_n125_));
  NO2        u0103(.A(i_6_), .B(i_5_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n126_), .B(i_3_), .Y(men_men_n127_));
  AO210      u0105(.A0(men_men_n127_), .A1(men_men_n48_), .B0(men_men_n125_), .Y(men_men_n128_));
  OAI220     u0106(.A0(men_men_n128_), .A1(men_men_n102_), .B0(men_men_n124_), .B1(men_men_n116_), .Y(men_men_n129_));
  NO3        u0107(.A(men_men_n129_), .B(men_men_n114_), .C(men_men_n89_), .Y(men_men_n130_));
  NA3        u0108(.A(men_men_n130_), .B(men_men_n77_), .C(men_men_n56_), .Y(men2));
  NO2        u0109(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n132_));
  INV        u0110(.A(i_6_), .Y(men_men_n133_));
  NA2        u0111(.A(men_men_n133_), .B(men_men_n132_), .Y(men_men_n134_));
  NA4        u0112(.A(men_men_n134_), .B(men_men_n75_), .C(men_men_n67_), .D(men_men_n30_), .Y(men0));
  AN2        u0113(.A(i_8_), .B(i_7_), .Y(men_men_n136_));
  NA2        u0114(.A(men_men_n136_), .B(i_6_), .Y(men_men_n137_));
  NO2        u0115(.A(i_12_), .B(i_13_), .Y(men_men_n138_));
  NAi21      u0116(.An(i_5_), .B(i_11_), .Y(men_men_n139_));
  NOi21      u0117(.An(men_men_n138_), .B(men_men_n139_), .Y(men_men_n140_));
  NO2        u0118(.A(i_0_), .B(i_1_), .Y(men_men_n141_));
  NA2        u0119(.A(i_2_), .B(i_3_), .Y(men_men_n142_));
  NO2        u0120(.A(men_men_n142_), .B(i_4_), .Y(men_men_n143_));
  NA3        u0121(.A(men_men_n143_), .B(men_men_n141_), .C(men_men_n140_), .Y(men_men_n144_));
  OR2        u0122(.A(men_men_n144_), .B(men_men_n25_), .Y(men_men_n145_));
  AN2        u0123(.A(men_men_n138_), .B(men_men_n81_), .Y(men_men_n146_));
  NO2        u0124(.A(men_men_n146_), .B(men_men_n27_), .Y(men_men_n147_));
  NA2        u0125(.A(i_1_), .B(i_5_), .Y(men_men_n148_));
  NO2        u0126(.A(men_men_n71_), .B(men_men_n47_), .Y(men_men_n149_));
  NA2        u0127(.A(men_men_n149_), .B(men_men_n36_), .Y(men_men_n150_));
  NO3        u0128(.A(men_men_n150_), .B(men_men_n148_), .C(men_men_n147_), .Y(men_men_n151_));
  OR2        u0129(.A(i_0_), .B(i_1_), .Y(men_men_n152_));
  NO3        u0130(.A(men_men_n152_), .B(men_men_n78_), .C(i_13_), .Y(men_men_n153_));
  NAi32      u0131(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n154_));
  NAi21      u0132(.An(men_men_n154_), .B(men_men_n153_), .Y(men_men_n155_));
  NOi21      u0133(.An(i_4_), .B(i_10_), .Y(men_men_n156_));
  NA2        u0134(.A(men_men_n156_), .B(men_men_n40_), .Y(men_men_n157_));
  NO2        u0135(.A(i_3_), .B(i_5_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n71_), .B(i_2_), .C(i_1_), .Y(men_men_n159_));
  NA2        u0137(.A(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  OAI210     u0138(.A0(men_men_n160_), .A1(men_men_n157_), .B0(men_men_n155_), .Y(men_men_n161_));
  NO2        u0139(.A(men_men_n161_), .B(men_men_n151_), .Y(men_men_n162_));
  AOI210     u0140(.A0(men_men_n162_), .A1(men_men_n145_), .B0(men_men_n137_), .Y(men_men_n163_));
  NA3        u0141(.A(men_men_n71_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n164_));
  NOi21      u0142(.An(i_4_), .B(i_9_), .Y(men_men_n165_));
  NOi21      u0143(.An(i_11_), .B(i_13_), .Y(men_men_n166_));
  NA2        u0144(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  NO2        u0145(.A(i_4_), .B(i_5_), .Y(men_men_n168_));
  NAi21      u0146(.An(i_12_), .B(i_11_), .Y(men_men_n169_));
  NO2        u0147(.A(men_men_n169_), .B(i_13_), .Y(men_men_n170_));
  NA3        u0148(.A(men_men_n170_), .B(men_men_n168_), .C(men_men_n81_), .Y(men_men_n171_));
  AOI210     u0149(.A0(men_men_n171_), .A1(men_men_n167_), .B0(men_men_n164_), .Y(men_men_n172_));
  NO2        u0150(.A(men_men_n71_), .B(men_men_n63_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n36_), .B(i_5_), .Y(men_men_n174_));
  NAi31      u0152(.An(men_men_n174_), .B(men_men_n146_), .C(i_11_), .Y(men_men_n175_));
  NA2        u0153(.A(i_3_), .B(i_5_), .Y(men_men_n176_));
  OR2        u0154(.A(men_men_n176_), .B(men_men_n167_), .Y(men_men_n177_));
  AOI210     u0155(.A0(men_men_n177_), .A1(men_men_n175_), .B0(men_men_n63_), .Y(men_men_n178_));
  NO2        u0156(.A(men_men_n71_), .B(i_5_), .Y(men_men_n179_));
  NO2        u0157(.A(i_13_), .B(i_10_), .Y(men_men_n180_));
  NA3        u0158(.A(men_men_n180_), .B(men_men_n179_), .C(men_men_n45_), .Y(men_men_n181_));
  NO2        u0159(.A(i_2_), .B(i_1_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n182_), .B(i_3_), .Y(men_men_n183_));
  NAi21      u0161(.An(i_4_), .B(i_12_), .Y(men_men_n184_));
  NO4        u0162(.A(men_men_n184_), .B(men_men_n183_), .C(men_men_n181_), .D(men_men_n25_), .Y(men_men_n185_));
  NO3        u0163(.A(men_men_n185_), .B(men_men_n178_), .C(men_men_n172_), .Y(men_men_n186_));
  INV        u0164(.A(i_8_), .Y(men_men_n187_));
  NO2        u0165(.A(men_men_n187_), .B(i_7_), .Y(men_men_n188_));
  NA2        u0166(.A(men_men_n188_), .B(i_6_), .Y(men_men_n189_));
  NO3        u0167(.A(i_3_), .B(men_men_n83_), .C(men_men_n49_), .Y(men_men_n190_));
  NA2        u0168(.A(men_men_n190_), .B(men_men_n106_), .Y(men_men_n191_));
  NO3        u0169(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n192_));
  NA3        u0170(.A(men_men_n192_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n193_));
  NO3        u0171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n194_));
  OAI210     u0172(.A0(men_men_n90_), .A1(i_12_), .B0(men_men_n194_), .Y(men_men_n195_));
  AOI210     u0173(.A0(men_men_n195_), .A1(men_men_n193_), .B0(men_men_n191_), .Y(men_men_n196_));
  NO2        u0174(.A(i_3_), .B(i_8_), .Y(men_men_n197_));
  NO3        u0175(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n198_));
  NA3        u0176(.A(men_men_n198_), .B(men_men_n197_), .C(men_men_n40_), .Y(men_men_n199_));
  NO2        u0177(.A(men_men_n97_), .B(men_men_n58_), .Y(men_men_n200_));
  NO2        u0178(.A(i_13_), .B(i_9_), .Y(men_men_n201_));
  NA3        u0179(.A(men_men_n201_), .B(i_6_), .C(men_men_n187_), .Y(men_men_n202_));
  NAi21      u0180(.An(i_12_), .B(i_3_), .Y(men_men_n203_));
  OR2        u0181(.A(men_men_n203_), .B(men_men_n202_), .Y(men_men_n204_));
  NO2        u0182(.A(men_men_n45_), .B(i_5_), .Y(men_men_n205_));
  NO3        u0183(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n206_));
  INV        u0184(.A(men_men_n206_), .Y(men_men_n207_));
  OAI220     u0185(.A0(men_men_n207_), .A1(men_men_n204_), .B0(men_men_n97_), .B1(men_men_n199_), .Y(men_men_n208_));
  AOI210     u0186(.A0(men_men_n208_), .A1(i_7_), .B0(men_men_n196_), .Y(men_men_n209_));
  OAI220     u0187(.A0(men_men_n209_), .A1(i_4_), .B0(men_men_n189_), .B1(men_men_n186_), .Y(men_men_n210_));
  NAi21      u0188(.An(i_12_), .B(i_7_), .Y(men_men_n211_));
  NA3        u0189(.A(i_13_), .B(men_men_n187_), .C(i_10_), .Y(men_men_n212_));
  NO2        u0190(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  NA2        u0191(.A(i_0_), .B(i_5_), .Y(men_men_n214_));
  OAI220     u0192(.A0(men_men_n83_), .A1(men_men_n183_), .B0(men_men_n63_), .B1(men_men_n127_), .Y(men_men_n215_));
  NAi31      u0193(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n216_));
  NO2        u0194(.A(men_men_n36_), .B(i_13_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n47_), .B(men_men_n63_), .Y(men_men_n218_));
  NA3        u0196(.A(men_men_n218_), .B(i_0_), .C(men_men_n217_), .Y(men_men_n219_));
  INV        u0197(.A(i_13_), .Y(men_men_n220_));
  NO2        u0198(.A(i_12_), .B(men_men_n220_), .Y(men_men_n221_));
  NA3        u0199(.A(men_men_n221_), .B(men_men_n192_), .C(men_men_n190_), .Y(men_men_n222_));
  OAI210     u0200(.A0(men_men_n219_), .A1(men_men_n216_), .B0(men_men_n222_), .Y(men_men_n223_));
  AOI220     u0201(.A0(men_men_n223_), .A1(men_men_n136_), .B0(men_men_n215_), .B1(men_men_n213_), .Y(men_men_n224_));
  NO2        u0202(.A(i_12_), .B(men_men_n37_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n176_), .B(i_4_), .Y(men_men_n226_));
  NA2        u0204(.A(men_men_n226_), .B(men_men_n225_), .Y(men_men_n227_));
  OR2        u0205(.A(i_8_), .B(i_7_), .Y(men_men_n228_));
  NO2        u0206(.A(men_men_n228_), .B(men_men_n83_), .Y(men_men_n229_));
  NO2        u0207(.A(men_men_n54_), .B(i_1_), .Y(men_men_n230_));
  NA2        u0208(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n231_));
  INV        u0209(.A(i_12_), .Y(men_men_n232_));
  NO3        u0210(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n233_));
  NA2        u0211(.A(i_2_), .B(i_1_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n231_), .B(men_men_n227_), .Y(men_men_n235_));
  NO3        u0213(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n236_));
  NAi21      u0214(.An(i_4_), .B(i_3_), .Y(men_men_n237_));
  NO2        u0215(.A(i_0_), .B(i_6_), .Y(men_men_n238_));
  NOi41      u0216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n234_), .B(men_men_n176_), .Y(men_men_n241_));
  NAi21      u0219(.An(men_men_n240_), .B(men_men_n241_), .Y(men_men_n242_));
  INV        u0220(.A(men_men_n242_), .Y(men_men_n243_));
  AOI220     u0221(.A0(men_men_n243_), .A1(men_men_n40_), .B0(men_men_n235_), .B1(men_men_n201_), .Y(men_men_n244_));
  NO2        u0222(.A(i_11_), .B(men_men_n220_), .Y(men_men_n245_));
  NOi21      u0223(.An(i_1_), .B(i_6_), .Y(men_men_n246_));
  NAi21      u0224(.An(i_3_), .B(i_7_), .Y(men_men_n247_));
  NO2        u0225(.A(i_12_), .B(i_3_), .Y(men_men_n248_));
  NA2        u0226(.A(i_3_), .B(i_9_), .Y(men_men_n249_));
  NA3        u0227(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n250_));
  INV        u0228(.A(men_men_n137_), .Y(men_men_n251_));
  NA2        u0229(.A(men_men_n232_), .B(i_13_), .Y(men_men_n252_));
  NO2        u0230(.A(men_men_n252_), .B(men_men_n73_), .Y(men_men_n253_));
  NA2        u0231(.A(men_men_n253_), .B(men_men_n251_), .Y(men_men_n254_));
  NO2        u0232(.A(men_men_n228_), .B(men_men_n37_), .Y(men_men_n255_));
  NA2        u0233(.A(i_12_), .B(i_6_), .Y(men_men_n256_));
  OR2        u0234(.A(i_13_), .B(i_9_), .Y(men_men_n257_));
  NO3        u0235(.A(men_men_n257_), .B(men_men_n256_), .C(men_men_n49_), .Y(men_men_n258_));
  NO2        u0236(.A(men_men_n237_), .B(i_2_), .Y(men_men_n259_));
  NA3        u0237(.A(men_men_n259_), .B(men_men_n258_), .C(men_men_n45_), .Y(men_men_n260_));
  NA2        u0238(.A(men_men_n245_), .B(i_9_), .Y(men_men_n261_));
  OAI210     u0239(.A0(men_men_n63_), .A1(men_men_n261_), .B0(men_men_n260_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n149_), .B(men_men_n63_), .Y(men_men_n263_));
  NO3        u0241(.A(i_11_), .B(men_men_n220_), .C(men_men_n25_), .Y(men_men_n264_));
  NO2        u0242(.A(men_men_n247_), .B(i_8_), .Y(men_men_n265_));
  NO2        u0243(.A(i_6_), .B(men_men_n49_), .Y(men_men_n266_));
  NA2        u0244(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n267_));
  NO3        u0245(.A(men_men_n26_), .B(men_men_n83_), .C(i_5_), .Y(men_men_n268_));
  NA3        u0246(.A(men_men_n268_), .B(men_men_n255_), .C(men_men_n221_), .Y(men_men_n269_));
  AOI210     u0247(.A0(men_men_n269_), .A1(men_men_n267_), .B0(men_men_n263_), .Y(men_men_n270_));
  AOI210     u0248(.A0(men_men_n262_), .A1(men_men_n255_), .B0(men_men_n270_), .Y(men_men_n271_));
  NA4        u0249(.A(men_men_n271_), .B(men_men_n254_), .C(men_men_n244_), .D(men_men_n224_), .Y(men_men_n272_));
  NO3        u0250(.A(i_12_), .B(men_men_n220_), .C(men_men_n37_), .Y(men_men_n273_));
  INV        u0251(.A(men_men_n273_), .Y(men_men_n274_));
  NO3        u0252(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n275_));
  AOI220     u0253(.A0(men_men_n275_), .A1(men_men_n190_), .B0(men_men_n158_), .B1(men_men_n230_), .Y(men_men_n276_));
  NO2        u0254(.A(men_men_n276_), .B(men_men_n1025_), .Y(men_men_n277_));
  NO3        u0255(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n278_));
  NO2        u0256(.A(men_men_n234_), .B(i_0_), .Y(men_men_n279_));
  AOI220     u0257(.A0(men_men_n279_), .A1(men_men_n188_), .B0(men_men_n278_), .B1(men_men_n136_), .Y(men_men_n280_));
  NA2        u0258(.A(men_men_n266_), .B(men_men_n26_), .Y(men_men_n281_));
  NO2        u0259(.A(men_men_n281_), .B(men_men_n280_), .Y(men_men_n282_));
  NA2        u0260(.A(i_0_), .B(i_1_), .Y(men_men_n283_));
  NO2        u0261(.A(men_men_n283_), .B(i_2_), .Y(men_men_n284_));
  NO2        u0262(.A(men_men_n59_), .B(i_6_), .Y(men_men_n285_));
  NA3        u0263(.A(men_men_n285_), .B(men_men_n284_), .C(men_men_n158_), .Y(men_men_n286_));
  OAI210     u0264(.A0(men_men_n160_), .A1(men_men_n137_), .B0(men_men_n286_), .Y(men_men_n287_));
  NO3        u0265(.A(men_men_n287_), .B(men_men_n282_), .C(men_men_n277_), .Y(men_men_n288_));
  NO2        u0266(.A(i_3_), .B(i_10_), .Y(men_men_n289_));
  NA3        u0267(.A(men_men_n289_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n290_));
  NO2        u0268(.A(i_2_), .B(men_men_n95_), .Y(men_men_n291_));
  NA2        u0269(.A(i_1_), .B(men_men_n36_), .Y(men_men_n292_));
  NOi21      u0270(.An(men_men_n214_), .B(men_men_n97_), .Y(men_men_n293_));
  NA3        u0271(.A(men_men_n293_), .B(i_1_), .C(men_men_n291_), .Y(men_men_n294_));
  AN2        u0272(.A(i_3_), .B(i_10_), .Y(men_men_n295_));
  NA4        u0273(.A(men_men_n295_), .B(men_men_n192_), .C(men_men_n170_), .D(men_men_n168_), .Y(men_men_n296_));
  NO2        u0274(.A(i_5_), .B(men_men_n37_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n298_));
  OR2        u0276(.A(men_men_n294_), .B(men_men_n290_), .Y(men_men_n299_));
  OAI220     u0277(.A0(men_men_n299_), .A1(i_6_), .B0(men_men_n288_), .B1(men_men_n274_), .Y(men_men_n300_));
  NO4        u0278(.A(men_men_n300_), .B(men_men_n272_), .C(men_men_n210_), .D(men_men_n163_), .Y(men_men_n301_));
  NO3        u0279(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n59_), .B(men_men_n83_), .Y(men_men_n303_));
  NA2        u0281(.A(men_men_n279_), .B(men_men_n303_), .Y(men_men_n304_));
  NO3        u0282(.A(i_6_), .B(men_men_n187_), .C(i_7_), .Y(men_men_n305_));
  NA2        u0283(.A(men_men_n305_), .B(men_men_n192_), .Y(men_men_n306_));
  AOI210     u0284(.A0(men_men_n306_), .A1(men_men_n304_), .B0(i_5_), .Y(men_men_n307_));
  NO2        u0285(.A(i_2_), .B(i_3_), .Y(men_men_n308_));
  OR2        u0286(.A(i_0_), .B(i_5_), .Y(men_men_n309_));
  NA2        u0287(.A(men_men_n214_), .B(men_men_n309_), .Y(men_men_n310_));
  NA4        u0288(.A(men_men_n310_), .B(men_men_n229_), .C(men_men_n308_), .D(i_1_), .Y(men_men_n311_));
  NA3        u0289(.A(men_men_n279_), .B(men_men_n158_), .C(men_men_n106_), .Y(men_men_n312_));
  NAi21      u0290(.An(i_8_), .B(i_7_), .Y(men_men_n313_));
  NO2        u0291(.A(men_men_n152_), .B(men_men_n47_), .Y(men_men_n314_));
  NA3        u0292(.A(men_men_n314_), .B(i_7_), .C(men_men_n158_), .Y(men_men_n315_));
  NA3        u0293(.A(men_men_n315_), .B(men_men_n312_), .C(men_men_n311_), .Y(men_men_n316_));
  OAI210     u0294(.A0(men_men_n316_), .A1(men_men_n307_), .B0(i_4_), .Y(men_men_n317_));
  NO2        u0295(.A(i_12_), .B(i_10_), .Y(men_men_n318_));
  NOi21      u0296(.An(i_5_), .B(i_0_), .Y(men_men_n319_));
  NO2        u0297(.A(men_men_n292_), .B(men_men_n122_), .Y(men_men_n320_));
  NA4        u0298(.A(men_men_n82_), .B(men_men_n36_), .C(men_men_n83_), .D(i_8_), .Y(men_men_n321_));
  NA2        u0299(.A(men_men_n320_), .B(men_men_n318_), .Y(men_men_n322_));
  NO2        u0300(.A(i_6_), .B(i_8_), .Y(men_men_n323_));
  AN2        u0301(.A(i_0_), .B(men_men_n323_), .Y(men_men_n324_));
  NO2        u0302(.A(i_1_), .B(i_7_), .Y(men_men_n325_));
  NA2        u0303(.A(men_men_n324_), .B(men_men_n42_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n326_), .B(men_men_n322_), .C(men_men_n317_), .Y(men_men_n327_));
  NO3        u0305(.A(men_men_n228_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n328_));
  NO3        u0306(.A(men_men_n313_), .B(i_2_), .C(i_1_), .Y(men_men_n329_));
  OAI210     u0307(.A0(men_men_n329_), .A1(men_men_n328_), .B0(i_6_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n246_), .B(men_men_n291_), .C(men_men_n187_), .Y(men_men_n331_));
  NA2        u0309(.A(men_men_n331_), .B(men_men_n330_), .Y(men_men_n332_));
  NA2        u0310(.A(men_men_n332_), .B(i_3_), .Y(men_men_n333_));
  NO2        u0311(.A(men_men_n283_), .B(men_men_n79_), .Y(men_men_n334_));
  NA2        u0312(.A(men_men_n334_), .B(men_men_n126_), .Y(men_men_n335_));
  NO2        u0313(.A(men_men_n88_), .B(men_men_n187_), .Y(men_men_n336_));
  NA2        u0314(.A(men_men_n293_), .B(men_men_n336_), .Y(men_men_n337_));
  AOI210     u0315(.A0(men_men_n337_), .A1(men_men_n335_), .B0(i_3_), .Y(men_men_n338_));
  NO2        u0316(.A(men_men_n187_), .B(i_9_), .Y(men_men_n339_));
  NA2        u0317(.A(men_men_n339_), .B(men_men_n200_), .Y(men_men_n340_));
  NO2        u0318(.A(men_men_n338_), .B(men_men_n282_), .Y(men_men_n341_));
  AOI210     u0319(.A0(men_men_n341_), .A1(men_men_n333_), .B0(men_men_n157_), .Y(men_men_n342_));
  AOI210     u0320(.A0(men_men_n327_), .A1(men_men_n302_), .B0(men_men_n342_), .Y(men_men_n343_));
  NOi32      u0321(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n344_));
  INV        u0322(.A(men_men_n344_), .Y(men_men_n345_));
  NAi21      u0323(.An(i_1_), .B(i_5_), .Y(men_men_n346_));
  INV        u0324(.A(men_men_n240_), .Y(men_men_n347_));
  NAi41      u0325(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n348_));
  OAI220     u0326(.A0(men_men_n348_), .A1(men_men_n346_), .B0(men_men_n216_), .B1(men_men_n154_), .Y(men_men_n349_));
  AOI210     u0327(.A0(men_men_n348_), .A1(men_men_n154_), .B0(men_men_n152_), .Y(men_men_n350_));
  NOi32      u0328(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n351_));
  NAi21      u0329(.An(i_6_), .B(i_1_), .Y(men_men_n352_));
  NA3        u0330(.A(men_men_n352_), .B(men_men_n351_), .C(men_men_n47_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n353_), .B(i_0_), .Y(men_men_n354_));
  OR3        u0332(.A(men_men_n354_), .B(men_men_n350_), .C(men_men_n349_), .Y(men_men_n355_));
  NO2        u0333(.A(i_1_), .B(men_men_n95_), .Y(men_men_n356_));
  NAi21      u0334(.An(i_3_), .B(i_4_), .Y(men_men_n357_));
  NO2        u0335(.A(men_men_n357_), .B(i_9_), .Y(men_men_n358_));
  AN2        u0336(.A(i_6_), .B(i_7_), .Y(men_men_n359_));
  OAI210     u0337(.A0(men_men_n359_), .A1(men_men_n356_), .B0(men_men_n358_), .Y(men_men_n360_));
  NA2        u0338(.A(i_2_), .B(i_7_), .Y(men_men_n361_));
  NO2        u0339(.A(men_men_n357_), .B(i_10_), .Y(men_men_n362_));
  NA3        u0340(.A(men_men_n362_), .B(men_men_n361_), .C(men_men_n238_), .Y(men_men_n363_));
  AOI210     u0341(.A0(men_men_n363_), .A1(men_men_n360_), .B0(men_men_n179_), .Y(men_men_n364_));
  AOI220     u0342(.A0(men_men_n362_), .A1(men_men_n325_), .B0(men_men_n233_), .B1(men_men_n182_), .Y(men_men_n365_));
  NO2        u0343(.A(men_men_n365_), .B(i_5_), .Y(men_men_n366_));
  NO4        u0344(.A(men_men_n366_), .B(men_men_n364_), .C(men_men_n355_), .D(men_men_n347_), .Y(men_men_n367_));
  NO2        u0345(.A(men_men_n367_), .B(men_men_n345_), .Y(men_men_n368_));
  NO2        u0346(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n369_));
  AN2        u0347(.A(i_12_), .B(i_5_), .Y(men_men_n370_));
  NO2        u0348(.A(i_4_), .B(men_men_n26_), .Y(men_men_n371_));
  NA2        u0349(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  NO2        u0350(.A(i_11_), .B(i_6_), .Y(men_men_n373_));
  NA3        u0351(.A(men_men_n373_), .B(men_men_n314_), .C(men_men_n220_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n374_), .B(men_men_n372_), .Y(men_men_n375_));
  NO2        u0353(.A(men_men_n237_), .B(i_5_), .Y(men_men_n376_));
  NO2        u0354(.A(i_5_), .B(i_10_), .Y(men_men_n377_));
  AOI220     u0355(.A0(men_men_n377_), .A1(men_men_n259_), .B0(men_men_n376_), .B1(men_men_n192_), .Y(men_men_n378_));
  NO2        u0356(.A(men_men_n1020_), .B(men_men_n378_), .Y(men_men_n379_));
  OAI210     u0357(.A0(men_men_n379_), .A1(men_men_n375_), .B0(men_men_n369_), .Y(men_men_n380_));
  NO2        u0358(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n144_), .B(men_men_n83_), .Y(men_men_n382_));
  OAI210     u0360(.A0(men_men_n382_), .A1(men_men_n375_), .B0(men_men_n381_), .Y(men_men_n383_));
  NO3        u0361(.A(men_men_n83_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n384_));
  NA2        u0362(.A(men_men_n289_), .B(men_men_n87_), .Y(men_men_n385_));
  NO2        u0363(.A(i_11_), .B(i_12_), .Y(men_men_n386_));
  NA2        u0364(.A(men_men_n386_), .B(men_men_n36_), .Y(men_men_n387_));
  NO2        u0365(.A(men_men_n385_), .B(men_men_n387_), .Y(men_men_n388_));
  NA2        u0366(.A(men_men_n377_), .B(men_men_n232_), .Y(men_men_n389_));
  INV        u0367(.A(men_men_n42_), .Y(men_men_n390_));
  NO2        u0368(.A(men_men_n390_), .B(men_men_n216_), .Y(men_men_n391_));
  NAi21      u0369(.An(i_13_), .B(i_0_), .Y(men_men_n392_));
  NO2        u0370(.A(men_men_n392_), .B(men_men_n234_), .Y(men_men_n393_));
  OAI210     u0371(.A0(men_men_n391_), .A1(men_men_n388_), .B0(men_men_n393_), .Y(men_men_n394_));
  NA3        u0372(.A(men_men_n394_), .B(men_men_n383_), .C(men_men_n380_), .Y(men_men_n395_));
  NA2        u0373(.A(men_men_n45_), .B(men_men_n220_), .Y(men_men_n396_));
  NO3        u0374(.A(i_1_), .B(i_12_), .C(men_men_n83_), .Y(men_men_n397_));
  NO2        u0375(.A(i_0_), .B(i_11_), .Y(men_men_n398_));
  AN2        u0376(.A(i_1_), .B(i_6_), .Y(men_men_n399_));
  NOi21      u0377(.An(i_2_), .B(i_12_), .Y(men_men_n400_));
  NA2        u0378(.A(men_men_n400_), .B(men_men_n399_), .Y(men_men_n401_));
  INV        u0379(.A(men_men_n401_), .Y(men_men_n402_));
  NA2        u0380(.A(men_men_n136_), .B(i_9_), .Y(men_men_n403_));
  NO2        u0381(.A(men_men_n403_), .B(i_4_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n402_), .B(men_men_n404_), .Y(men_men_n405_));
  NAi21      u0383(.An(i_9_), .B(i_4_), .Y(men_men_n406_));
  OR2        u0384(.A(i_13_), .B(i_10_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n167_), .B(men_men_n117_), .Y(men_men_n408_));
  BUFFER     u0386(.A(men_men_n212_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n95_), .B(men_men_n25_), .Y(men_men_n410_));
  NA2        u0388(.A(men_men_n266_), .B(men_men_n206_), .Y(men_men_n411_));
  NO2        u0389(.A(men_men_n411_), .B(men_men_n409_), .Y(men_men_n412_));
  INV        u0390(.A(men_men_n412_), .Y(men_men_n413_));
  AOI210     u0391(.A0(men_men_n413_), .A1(men_men_n405_), .B0(men_men_n26_), .Y(men_men_n414_));
  NA2        u0392(.A(men_men_n312_), .B(men_men_n311_), .Y(men_men_n415_));
  AOI220     u0393(.A0(men_men_n285_), .A1(men_men_n275_), .B0(men_men_n279_), .B1(men_men_n303_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n416_), .B(i_5_), .Y(men_men_n417_));
  NO2        u0395(.A(men_men_n176_), .B(men_men_n83_), .Y(men_men_n418_));
  AOI220     u0396(.A0(men_men_n418_), .A1(men_men_n284_), .B0(men_men_n268_), .B1(men_men_n206_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n419_), .B(men_men_n1025_), .Y(men_men_n420_));
  NO3        u0398(.A(men_men_n420_), .B(men_men_n417_), .C(men_men_n415_), .Y(men_men_n421_));
  INV        u0399(.A(men_men_n90_), .Y(men_men_n422_));
  NA3        u0400(.A(men_men_n314_), .B(men_men_n158_), .C(men_men_n83_), .Y(men_men_n423_));
  AOI210     u0401(.A0(men_men_n423_), .A1(men_men_n422_), .B0(men_men_n313_), .Y(men_men_n424_));
  NA2        u0402(.A(men_men_n285_), .B(men_men_n230_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n425_), .B(men_men_n176_), .Y(men_men_n426_));
  NO2        u0404(.A(i_3_), .B(men_men_n49_), .Y(men_men_n427_));
  NA3        u0405(.A(men_men_n325_), .B(men_men_n324_), .C(men_men_n427_), .Y(men_men_n428_));
  NA2        u0406(.A(men_men_n305_), .B(men_men_n310_), .Y(men_men_n429_));
  OAI210     u0407(.A0(men_men_n429_), .A1(men_men_n183_), .B0(men_men_n428_), .Y(men_men_n430_));
  NO3        u0408(.A(men_men_n430_), .B(men_men_n426_), .C(men_men_n424_), .Y(men_men_n431_));
  AOI210     u0409(.A0(men_men_n431_), .A1(men_men_n421_), .B0(men_men_n261_), .Y(men_men_n432_));
  NO4        u0410(.A(men_men_n432_), .B(men_men_n414_), .C(men_men_n395_), .D(men_men_n368_), .Y(men_men_n433_));
  NO2        u0411(.A(men_men_n71_), .B(i_13_), .Y(men_men_n434_));
  NO2        u0412(.A(i_10_), .B(i_9_), .Y(men_men_n435_));
  NAi21      u0413(.An(i_12_), .B(i_8_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(i_3_), .Y(men_men_n437_));
  NA2        u0415(.A(i_2_), .B(men_men_n98_), .Y(men_men_n438_));
  NO2        u0416(.A(men_men_n438_), .B(men_men_n199_), .Y(men_men_n439_));
  NA2        u0417(.A(men_men_n298_), .B(i_0_), .Y(men_men_n440_));
  NO3        u0418(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n441_));
  NA2        u0419(.A(men_men_n256_), .B(men_men_n91_), .Y(men_men_n442_));
  NA2        u0420(.A(men_men_n442_), .B(men_men_n441_), .Y(men_men_n443_));
  NA2        u0421(.A(i_8_), .B(i_9_), .Y(men_men_n444_));
  NA2        u0422(.A(men_men_n273_), .B(men_men_n200_), .Y(men_men_n445_));
  OAI220     u0423(.A0(men_men_n445_), .A1(men_men_n444_), .B0(men_men_n443_), .B1(men_men_n440_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n245_), .B(men_men_n297_), .Y(men_men_n447_));
  NO3        u0425(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n448_));
  INV        u0426(.A(men_men_n448_), .Y(men_men_n449_));
  NA3        u0427(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n450_));
  NA4        u0428(.A(men_men_n139_), .B(men_men_n109_), .C(men_men_n78_), .D(men_men_n23_), .Y(men_men_n451_));
  OAI220     u0429(.A0(men_men_n451_), .A1(men_men_n450_), .B0(men_men_n449_), .B1(men_men_n447_), .Y(men_men_n452_));
  NO3        u0430(.A(men_men_n452_), .B(men_men_n446_), .C(men_men_n439_), .Y(men_men_n453_));
  NA2        u0431(.A(men_men_n284_), .B(men_men_n102_), .Y(men_men_n454_));
  OR2        u0432(.A(men_men_n454_), .B(men_men_n202_), .Y(men_men_n455_));
  OR2        u0433(.A(men_men_n340_), .B(men_men_n95_), .Y(men_men_n456_));
  OA220      u0434(.A0(men_men_n456_), .A1(men_men_n157_), .B0(men_men_n455_), .B1(men_men_n227_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n90_), .B(i_13_), .Y(men_men_n458_));
  NA2        u0436(.A(men_men_n418_), .B(men_men_n369_), .Y(men_men_n459_));
  NO2        u0437(.A(i_2_), .B(i_13_), .Y(men_men_n460_));
  NA3        u0438(.A(men_men_n460_), .B(men_men_n156_), .C(men_men_n93_), .Y(men_men_n461_));
  NO2        u0439(.A(men_men_n459_), .B(men_men_n458_), .Y(men_men_n462_));
  NO3        u0440(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n463_));
  NO2        u0441(.A(i_6_), .B(i_7_), .Y(men_men_n464_));
  NA2        u0442(.A(men_men_n464_), .B(men_men_n463_), .Y(men_men_n465_));
  NO2        u0443(.A(i_11_), .B(i_1_), .Y(men_men_n466_));
  OR2        u0444(.A(i_11_), .B(i_8_), .Y(men_men_n467_));
  NOi21      u0445(.An(i_2_), .B(i_7_), .Y(men_men_n468_));
  NAi31      u0446(.An(men_men_n467_), .B(men_men_n468_), .C(i_0_), .Y(men_men_n469_));
  NO2        u0447(.A(men_men_n407_), .B(i_6_), .Y(men_men_n470_));
  NA2        u0448(.A(men_men_n470_), .B(i_1_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n471_), .B(men_men_n469_), .Y(men_men_n472_));
  NO2        u0450(.A(i_3_), .B(men_men_n187_), .Y(men_men_n473_));
  NO2        u0451(.A(i_6_), .B(i_10_), .Y(men_men_n474_));
  NA3        u0452(.A(men_men_n474_), .B(men_men_n302_), .C(men_men_n473_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n475_), .B(men_men_n150_), .Y(men_men_n476_));
  NA3        u0454(.A(men_men_n239_), .B(men_men_n166_), .C(men_men_n126_), .Y(men_men_n477_));
  NO2        u0455(.A(men_men_n152_), .B(i_3_), .Y(men_men_n478_));
  NA3        u0456(.A(men_men_n381_), .B(men_men_n173_), .C(men_men_n143_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n479_), .B(men_men_n477_), .Y(men_men_n480_));
  NO4        u0458(.A(men_men_n480_), .B(men_men_n476_), .C(men_men_n472_), .D(men_men_n462_), .Y(men_men_n481_));
  NA2        u0459(.A(men_men_n441_), .B(men_men_n370_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n448_), .B(men_men_n377_), .Y(men_men_n483_));
  NO2        u0461(.A(men_men_n483_), .B(men_men_n219_), .Y(men_men_n484_));
  NAi21      u0462(.An(men_men_n212_), .B(men_men_n386_), .Y(men_men_n485_));
  NA2        u0463(.A(men_men_n325_), .B(men_men_n214_), .Y(men_men_n486_));
  NO2        u0464(.A(men_men_n26_), .B(i_5_), .Y(men_men_n487_));
  NA3        u0465(.A(i_6_), .B(men_men_n487_), .C(men_men_n136_), .Y(men_men_n488_));
  OR3        u0466(.A(men_men_n292_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n489_));
  OAI220     u0467(.A0(men_men_n489_), .A1(men_men_n488_), .B0(men_men_n486_), .B1(men_men_n485_), .Y(men_men_n490_));
  NA3        u0468(.A(men_men_n295_), .B(men_men_n218_), .C(men_men_n71_), .Y(men_men_n491_));
  NO2        u0469(.A(men_men_n491_), .B(men_men_n465_), .Y(men_men_n492_));
  NO3        u0470(.A(men_men_n492_), .B(men_men_n490_), .C(men_men_n484_), .Y(men_men_n493_));
  NA4        u0471(.A(men_men_n493_), .B(men_men_n481_), .C(men_men_n457_), .D(men_men_n453_), .Y(men_men_n494_));
  NA3        u0472(.A(men_men_n295_), .B(men_men_n170_), .C(men_men_n168_), .Y(men_men_n495_));
  OAI210     u0473(.A0(men_men_n290_), .A1(men_men_n174_), .B0(men_men_n495_), .Y(men_men_n496_));
  AN2        u0474(.A(men_men_n275_), .B(men_men_n229_), .Y(men_men_n497_));
  NA2        u0475(.A(men_men_n497_), .B(men_men_n496_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n116_), .B(men_men_n105_), .Y(men_men_n499_));
  AN2        u0477(.A(men_men_n499_), .B(men_men_n441_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n302_), .B(men_men_n159_), .Y(men_men_n501_));
  OAI210     u0479(.A0(men_men_n501_), .A1(men_men_n227_), .B0(men_men_n296_), .Y(men_men_n502_));
  AOI220     u0480(.A0(men_men_n502_), .A1(i_7_), .B0(men_men_n500_), .B1(men_men_n298_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n344_), .B(men_men_n71_), .Y(men_men_n504_));
  NA2        u0482(.A(men_men_n359_), .B(men_men_n351_), .Y(men_men_n505_));
  NO2        u0483(.A(men_men_n36_), .B(i_8_), .Y(men_men_n506_));
  NA2        u0484(.A(men_men_n39_), .B(i_13_), .Y(men_men_n507_));
  OAI210     u0485(.A0(i_8_), .A1(men_men_n63_), .B0(men_men_n128_), .Y(men_men_n508_));
  AOI210     u0486(.A0(men_men_n188_), .A1(i_9_), .B0(men_men_n255_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n509_), .B(men_men_n193_), .Y(men_men_n510_));
  OR2        u0488(.A(men_men_n176_), .B(i_4_), .Y(men_men_n511_));
  INV        u0489(.A(men_men_n511_), .Y(men_men_n512_));
  AOI220     u0490(.A0(men_men_n512_), .A1(men_men_n510_), .B0(men_men_n508_), .B1(men_men_n408_), .Y(men_men_n513_));
  NA4        u0491(.A(men_men_n513_), .B(men_men_n507_), .C(men_men_n503_), .D(men_men_n498_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n376_), .B(men_men_n284_), .Y(men_men_n515_));
  OAI210     u0493(.A0(men_men_n372_), .A1(men_men_n164_), .B0(men_men_n515_), .Y(men_men_n516_));
  NO2        u0494(.A(i_12_), .B(men_men_n187_), .Y(men_men_n517_));
  NOi31      u0495(.An(men_men_n305_), .B(men_men_n407_), .C(men_men_n38_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n518_), .B(men_men_n516_), .Y(men_men_n519_));
  NO2        u0497(.A(i_8_), .B(i_7_), .Y(men_men_n520_));
  OAI210     u0498(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n521_));
  NA2        u0499(.A(men_men_n521_), .B(men_men_n218_), .Y(men_men_n522_));
  NA2        u0500(.A(men_men_n45_), .B(i_10_), .Y(men_men_n523_));
  NO2        u0501(.A(men_men_n523_), .B(i_6_), .Y(men_men_n524_));
  NA3        u0502(.A(men_men_n524_), .B(men_men_n1024_), .C(men_men_n520_), .Y(men_men_n525_));
  AOI220     u0503(.A0(men_men_n418_), .A1(men_men_n314_), .B0(men_men_n241_), .B1(men_men_n238_), .Y(men_men_n526_));
  OAI220     u0504(.A0(men_men_n526_), .A1(men_men_n252_), .B0(men_men_n458_), .B1(men_men_n127_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n527_), .B(men_men_n255_), .Y(men_men_n528_));
  NO2        u0506(.A(men_men_n290_), .B(men_men_n174_), .Y(men_men_n529_));
  NA3        u0507(.A(men_men_n295_), .B(men_men_n168_), .C(men_men_n90_), .Y(men_men_n530_));
  NO2        u0508(.A(men_men_n152_), .B(i_5_), .Y(men_men_n531_));
  NA3        u0509(.A(men_men_n531_), .B(men_men_n396_), .C(men_men_n308_), .Y(men_men_n532_));
  NA2        u0510(.A(men_men_n532_), .B(men_men_n530_), .Y(men_men_n533_));
  OAI210     u0511(.A0(men_men_n533_), .A1(men_men_n529_), .B0(men_men_n448_), .Y(men_men_n534_));
  NA4        u0512(.A(men_men_n534_), .B(men_men_n528_), .C(men_men_n525_), .D(men_men_n519_), .Y(men_men_n535_));
  NA3        u0513(.A(men_men_n214_), .B(men_men_n69_), .C(men_men_n45_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n273_), .B(men_men_n82_), .Y(men_men_n537_));
  AOI210     u0515(.A0(men_men_n536_), .A1(men_men_n335_), .B0(men_men_n537_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n285_), .B(men_men_n275_), .Y(men_men_n539_));
  NO2        u0517(.A(men_men_n539_), .B(men_men_n167_), .Y(men_men_n540_));
  NA2        u0518(.A(i_0_), .B(men_men_n49_), .Y(men_men_n541_));
  NA3        u0519(.A(men_men_n517_), .B(men_men_n264_), .C(men_men_n541_), .Y(men_men_n542_));
  NO2        u0520(.A(i_1_), .B(men_men_n542_), .Y(men_men_n543_));
  NO3        u0521(.A(men_men_n543_), .B(men_men_n540_), .C(men_men_n538_), .Y(men_men_n544_));
  NO4        u0522(.A(men_men_n246_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n545_));
  NO3        u0523(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n546_));
  NO2        u0524(.A(men_men_n228_), .B(men_men_n36_), .Y(men_men_n547_));
  AN2        u0525(.A(men_men_n547_), .B(men_men_n546_), .Y(men_men_n548_));
  OA210      u0526(.A0(men_men_n548_), .A1(men_men_n545_), .B0(men_men_n344_), .Y(men_men_n549_));
  NO2        u0527(.A(men_men_n407_), .B(i_1_), .Y(men_men_n550_));
  NOi31      u0528(.An(men_men_n550_), .B(men_men_n442_), .C(men_men_n71_), .Y(men_men_n551_));
  AN3        u0529(.A(men_men_n551_), .B(men_men_n404_), .C(men_men_n487_), .Y(men_men_n552_));
  NO2        u0530(.A(men_men_n416_), .B(men_men_n171_), .Y(men_men_n553_));
  NO3        u0531(.A(men_men_n553_), .B(men_men_n552_), .C(men_men_n549_), .Y(men_men_n554_));
  NOi21      u0532(.An(i_10_), .B(i_6_), .Y(men_men_n555_));
  NO2        u0533(.A(men_men_n83_), .B(men_men_n25_), .Y(men_men_n556_));
  AOI220     u0534(.A0(men_men_n273_), .A1(men_men_n556_), .B0(men_men_n264_), .B1(men_men_n555_), .Y(men_men_n557_));
  NO2        u0535(.A(men_men_n557_), .B(men_men_n440_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n108_), .B(men_men_n23_), .Y(men_men_n559_));
  NA2        u0537(.A(men_men_n305_), .B(men_men_n159_), .Y(men_men_n560_));
  AOI220     u0538(.A0(men_men_n560_), .A1(men_men_n425_), .B0(men_men_n177_), .B1(men_men_n175_), .Y(men_men_n561_));
  NOi21      u0539(.An(men_men_n140_), .B(men_men_n321_), .Y(men_men_n562_));
  NO3        u0540(.A(men_men_n562_), .B(men_men_n561_), .C(men_men_n558_), .Y(men_men_n563_));
  NO2        u0541(.A(men_men_n504_), .B(men_men_n365_), .Y(men_men_n564_));
  INV        u0542(.A(men_men_n308_), .Y(men_men_n565_));
  NO2        u0543(.A(i_12_), .B(men_men_n83_), .Y(men_men_n566_));
  NA3        u0544(.A(men_men_n566_), .B(men_men_n264_), .C(men_men_n541_), .Y(men_men_n567_));
  NA3        u0545(.A(men_men_n373_), .B(men_men_n273_), .C(men_men_n214_), .Y(men_men_n568_));
  AOI210     u0546(.A0(men_men_n568_), .A1(men_men_n567_), .B0(men_men_n565_), .Y(men_men_n569_));
  NA2        u0547(.A(men_men_n168_), .B(i_0_), .Y(men_men_n570_));
  NO3        u0548(.A(men_men_n570_), .B(men_men_n330_), .C(men_men_n290_), .Y(men_men_n571_));
  OR2        u0549(.A(i_2_), .B(i_5_), .Y(men_men_n572_));
  OR2        u0550(.A(men_men_n572_), .B(men_men_n399_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n573_), .B(men_men_n485_), .Y(men_men_n574_));
  NO4        u0552(.A(men_men_n574_), .B(men_men_n571_), .C(men_men_n569_), .D(men_men_n564_), .Y(men_men_n575_));
  NA4        u0553(.A(men_men_n575_), .B(men_men_n563_), .C(men_men_n554_), .D(men_men_n544_), .Y(men_men_n576_));
  NO4        u0554(.A(men_men_n576_), .B(men_men_n535_), .C(men_men_n514_), .D(men_men_n494_), .Y(men_men_n577_));
  NA4        u0555(.A(men_men_n577_), .B(men_men_n433_), .C(men_men_n343_), .D(men_men_n301_), .Y(men7));
  NO2        u0556(.A(men_men_n102_), .B(men_men_n86_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n371_), .B(men_men_n579_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n474_), .B(men_men_n82_), .Y(men_men_n581_));
  NA2        u0559(.A(i_11_), .B(men_men_n187_), .Y(men_men_n582_));
  OAI210     u0560(.A0(men_men_n1023_), .A1(men_men_n581_), .B0(men_men_n580_), .Y(men_men_n583_));
  NA3        u0561(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n232_), .B(i_4_), .Y(men_men_n585_));
  NO2        u0563(.A(men_men_n99_), .B(men_men_n584_), .Y(men_men_n586_));
  NA2        u0564(.A(i_2_), .B(men_men_n83_), .Y(men_men_n587_));
  OAI210     u0565(.A0(men_men_n85_), .A1(men_men_n197_), .B0(men_men_n198_), .Y(men_men_n588_));
  NO2        u0566(.A(i_7_), .B(men_men_n37_), .Y(men_men_n589_));
  NA2        u0567(.A(i_4_), .B(i_8_), .Y(men_men_n590_));
  AOI210     u0568(.A0(men_men_n590_), .A1(men_men_n295_), .B0(men_men_n589_), .Y(men_men_n591_));
  NO2        u0569(.A(men_men_n591_), .B(men_men_n587_), .Y(men_men_n592_));
  NO3        u0570(.A(men_men_n592_), .B(men_men_n586_), .C(men_men_n583_), .Y(men_men_n593_));
  INV        u0571(.A(men_men_n156_), .Y(men_men_n594_));
  OR2        u0572(.A(i_6_), .B(i_10_), .Y(men_men_n595_));
  NO2        u0573(.A(men_men_n595_), .B(men_men_n23_), .Y(men_men_n596_));
  OR3        u0574(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n597_));
  NO3        u0575(.A(men_men_n597_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n598_));
  INV        u0576(.A(men_men_n194_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n598_), .B(men_men_n596_), .Y(men_men_n600_));
  OA220      u0578(.A0(men_men_n600_), .A1(men_men_n565_), .B0(men_men_n594_), .B1(men_men_n257_), .Y(men_men_n601_));
  AOI210     u0579(.A0(men_men_n601_), .A1(men_men_n593_), .B0(men_men_n63_), .Y(men_men_n602_));
  NOi21      u0580(.An(i_11_), .B(i_7_), .Y(men_men_n603_));
  AO210      u0581(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n604_), .B(men_men_n603_), .Y(men_men_n605_));
  NA2        u0583(.A(men_men_n605_), .B(men_men_n201_), .Y(men_men_n606_));
  NA3        u0584(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n607_));
  AOI210     u0585(.A0(men_men_n607_), .A1(men_men_n606_), .B0(men_men_n63_), .Y(men_men_n608_));
  AO210      u0586(.A0(men_men_n84_), .A1(men_men_n365_), .B0(men_men_n41_), .Y(men_men_n609_));
  NA2        u0587(.A(men_men_n221_), .B(men_men_n63_), .Y(men_men_n610_));
  NA2        u0588(.A(men_men_n400_), .B(men_men_n31_), .Y(men_men_n611_));
  OR2        u0589(.A(men_men_n203_), .B(men_men_n102_), .Y(men_men_n612_));
  NA2        u0590(.A(men_men_n612_), .B(men_men_n611_), .Y(men_men_n613_));
  NO2        u0591(.A(men_men_n63_), .B(i_9_), .Y(men_men_n614_));
  NO2        u0592(.A(men_men_n614_), .B(i_4_), .Y(men_men_n615_));
  NA2        u0593(.A(men_men_n615_), .B(men_men_n613_), .Y(men_men_n616_));
  NO2        u0594(.A(i_1_), .B(i_12_), .Y(men_men_n617_));
  NA3        u0595(.A(men_men_n617_), .B(men_men_n103_), .C(men_men_n24_), .Y(men_men_n618_));
  NA4        u0596(.A(men_men_n618_), .B(men_men_n616_), .C(men_men_n610_), .D(men_men_n609_), .Y(men_men_n619_));
  OAI210     u0597(.A0(men_men_n619_), .A1(men_men_n608_), .B0(i_6_), .Y(men_men_n620_));
  NO2        u0598(.A(i_6_), .B(i_11_), .Y(men_men_n621_));
  INV        u0599(.A(men_men_n443_), .Y(men_men_n622_));
  NO4        u0600(.A(men_men_n211_), .B(men_men_n122_), .C(i_13_), .D(men_men_n83_), .Y(men_men_n623_));
  NA2        u0601(.A(men_men_n623_), .B(men_men_n614_), .Y(men_men_n624_));
  INV        u0602(.A(men_men_n624_), .Y(men_men_n625_));
  NA3        u0603(.A(men_men_n520_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n626_));
  NA2        u0604(.A(men_men_n132_), .B(i_9_), .Y(men_men_n627_));
  NO2        u0605(.A(men_men_n47_), .B(i_1_), .Y(men_men_n628_));
  NO2        u0606(.A(men_men_n627_), .B(men_men_n1016_), .Y(men_men_n629_));
  NA3        u0607(.A(men_men_n614_), .B(men_men_n308_), .C(i_6_), .Y(men_men_n630_));
  NO2        u0608(.A(men_men_n630_), .B(men_men_n23_), .Y(men_men_n631_));
  AOI210     u0609(.A0(men_men_n466_), .A1(men_men_n410_), .B0(men_men_n236_), .Y(men_men_n632_));
  NO2        u0610(.A(men_men_n632_), .B(men_men_n587_), .Y(men_men_n633_));
  NA2        u0611(.A(men_men_n628_), .B(men_men_n256_), .Y(men_men_n634_));
  NO2        u0612(.A(i_11_), .B(men_men_n37_), .Y(men_men_n635_));
  NA2        u0613(.A(men_men_n635_), .B(men_men_n24_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n636_), .B(men_men_n634_), .Y(men_men_n637_));
  OR4        u0615(.A(men_men_n637_), .B(men_men_n633_), .C(men_men_n631_), .D(men_men_n629_), .Y(men_men_n638_));
  NO3        u0616(.A(men_men_n638_), .B(men_men_n625_), .C(men_men_n622_), .Y(men_men_n639_));
  NO2        u0617(.A(men_men_n232_), .B(men_men_n95_), .Y(men_men_n640_));
  NO2        u0618(.A(men_men_n640_), .B(men_men_n603_), .Y(men_men_n641_));
  NA2        u0619(.A(men_men_n641_), .B(i_1_), .Y(men_men_n642_));
  NO2        u0620(.A(men_men_n642_), .B(men_men_n597_), .Y(men_men_n643_));
  NO2        u0621(.A(men_men_n406_), .B(men_men_n83_), .Y(men_men_n644_));
  NA2        u0622(.A(men_men_n643_), .B(men_men_n47_), .Y(men_men_n645_));
  NA2        u0623(.A(i_3_), .B(men_men_n187_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n228_), .B(men_men_n45_), .Y(men_men_n647_));
  NO3        u0625(.A(men_men_n647_), .B(men_men_n298_), .C(i_12_), .Y(men_men_n648_));
  NO2        u0626(.A(men_men_n111_), .B(men_men_n37_), .Y(men_men_n649_));
  NO2        u0627(.A(men_men_n649_), .B(i_6_), .Y(men_men_n650_));
  NO2        u0628(.A(men_men_n83_), .B(i_9_), .Y(men_men_n651_));
  NO2        u0629(.A(men_men_n651_), .B(men_men_n63_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n652_), .B(men_men_n617_), .Y(men_men_n653_));
  NO4        u0631(.A(men_men_n653_), .B(men_men_n650_), .C(men_men_n648_), .D(i_4_), .Y(men_men_n654_));
  NA2        u0632(.A(i_1_), .B(i_3_), .Y(men_men_n655_));
  INV        u0633(.A(men_men_n654_), .Y(men_men_n656_));
  NA4        u0634(.A(men_men_n656_), .B(men_men_n645_), .C(men_men_n639_), .D(men_men_n620_), .Y(men_men_n657_));
  NO3        u0635(.A(men_men_n467_), .B(i_3_), .C(i_7_), .Y(men_men_n658_));
  NOi21      u0636(.An(men_men_n658_), .B(i_10_), .Y(men_men_n659_));
  OA210      u0637(.A0(men_men_n659_), .A1(men_men_n239_), .B0(men_men_n83_), .Y(men_men_n660_));
  NA3        u0638(.A(men_men_n474_), .B(men_men_n506_), .C(men_men_n47_), .Y(men_men_n661_));
  NO3        u0639(.A(men_men_n468_), .B(men_men_n590_), .C(men_men_n83_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(men_men_n25_), .Y(men_men_n663_));
  NA3        u0641(.A(men_men_n156_), .B(men_men_n82_), .C(men_men_n83_), .Y(men_men_n664_));
  NA3        u0642(.A(men_men_n664_), .B(men_men_n663_), .C(men_men_n661_), .Y(men_men_n665_));
  OAI210     u0643(.A0(men_men_n665_), .A1(men_men_n660_), .B0(i_1_), .Y(men_men_n666_));
  AOI210     u0644(.A0(men_men_n256_), .A1(men_men_n91_), .B0(i_1_), .Y(men_men_n667_));
  NO2        u0645(.A(men_men_n357_), .B(i_2_), .Y(men_men_n668_));
  NA2        u0646(.A(men_men_n668_), .B(men_men_n667_), .Y(men_men_n669_));
  OAI210     u0647(.A0(men_men_n630_), .A1(men_men_n436_), .B0(men_men_n669_), .Y(men_men_n670_));
  INV        u0648(.A(men_men_n670_), .Y(men_men_n671_));
  AOI210     u0649(.A0(men_men_n671_), .A1(men_men_n666_), .B0(i_13_), .Y(men_men_n672_));
  NA3        u0650(.A(i_11_), .B(men_men_n100_), .C(men_men_n132_), .Y(men_men_n673_));
  AOI220     u0651(.A0(men_men_n460_), .A1(men_men_n156_), .B0(i_2_), .B1(men_men_n132_), .Y(men_men_n674_));
  OAI210     u0652(.A0(men_men_n674_), .A1(men_men_n45_), .B0(men_men_n673_), .Y(men_men_n675_));
  NO2        u0653(.A(men_men_n55_), .B(i_12_), .Y(men_men_n676_));
  NO2        u0654(.A(men_men_n468_), .B(men_men_n24_), .Y(men_men_n677_));
  AOI220     u0655(.A0(men_men_n677_), .A1(men_men_n644_), .B0(men_men_n239_), .B1(men_men_n125_), .Y(men_men_n678_));
  OAI220     u0656(.A0(men_men_n678_), .A1(men_men_n41_), .B0(men_men_n1015_), .B1(men_men_n88_), .Y(men_men_n679_));
  AOI210     u0657(.A0(men_men_n675_), .A1(men_men_n323_), .B0(men_men_n679_), .Y(men_men_n680_));
  AOI220     u0658(.A0(i_12_), .A1(men_men_n70_), .B0(men_men_n373_), .B1(men_men_n628_), .Y(men_men_n681_));
  NO2        u0659(.A(men_men_n681_), .B(men_men_n237_), .Y(men_men_n682_));
  AOI210     u0660(.A0(men_men_n436_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n683_));
  NOi31      u0661(.An(men_men_n683_), .B(men_men_n581_), .C(men_men_n45_), .Y(men_men_n684_));
  NA2        u0662(.A(men_men_n121_), .B(i_13_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n685_), .B(men_men_n667_), .Y(men_men_n686_));
  NO3        u0664(.A(men_men_n69_), .B(men_men_n32_), .C(men_men_n95_), .Y(men_men_n687_));
  NA2        u0665(.A(men_men_n26_), .B(men_men_n187_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n1017_), .B(men_men_n599_), .Y(men_men_n689_));
  NO4        u0667(.A(men_men_n689_), .B(men_men_n686_), .C(men_men_n684_), .D(men_men_n682_), .Y(men_men_n690_));
  OR2        u0668(.A(i_11_), .B(i_6_), .Y(men_men_n691_));
  NA3        u0669(.A(men_men_n585_), .B(men_men_n688_), .C(i_7_), .Y(men_men_n692_));
  NO2        u0670(.A(men_men_n692_), .B(men_men_n691_), .Y(men_men_n693_));
  NA3        u0671(.A(men_men_n400_), .B(men_men_n589_), .C(men_men_n91_), .Y(men_men_n694_));
  NA2        u0672(.A(men_men_n621_), .B(i_13_), .Y(men_men_n695_));
  NA2        u0673(.A(men_men_n96_), .B(men_men_n688_), .Y(men_men_n696_));
  NAi21      u0674(.An(i_11_), .B(i_12_), .Y(men_men_n697_));
  NOi41      u0675(.An(men_men_n104_), .B(men_men_n697_), .C(i_13_), .D(men_men_n83_), .Y(men_men_n698_));
  NO3        u0676(.A(men_men_n468_), .B(men_men_n566_), .C(men_men_n590_), .Y(men_men_n699_));
  AOI220     u0677(.A0(men_men_n699_), .A1(men_men_n302_), .B0(men_men_n698_), .B1(men_men_n696_), .Y(men_men_n700_));
  NA3        u0678(.A(men_men_n700_), .B(men_men_n695_), .C(men_men_n694_), .Y(men_men_n701_));
  OAI210     u0679(.A0(men_men_n701_), .A1(men_men_n693_), .B0(men_men_n63_), .Y(men_men_n702_));
  NO2        u0680(.A(i_2_), .B(i_12_), .Y(men_men_n703_));
  NA2        u0681(.A(men_men_n356_), .B(men_men_n703_), .Y(men_men_n704_));
  NA2        u0682(.A(i_8_), .B(men_men_n25_), .Y(men_men_n705_));
  NO3        u0683(.A(men_men_n705_), .B(men_men_n371_), .C(men_men_n585_), .Y(men_men_n706_));
  OAI210     u0684(.A0(men_men_n706_), .A1(men_men_n358_), .B0(men_men_n356_), .Y(men_men_n707_));
  NO2        u0685(.A(men_men_n122_), .B(i_2_), .Y(men_men_n708_));
  NA2        u0686(.A(men_men_n707_), .B(men_men_n704_), .Y(men_men_n709_));
  NA3        u0687(.A(men_men_n709_), .B(men_men_n46_), .C(men_men_n220_), .Y(men_men_n710_));
  NA4        u0688(.A(men_men_n710_), .B(men_men_n702_), .C(men_men_n690_), .D(men_men_n680_), .Y(men_men_n711_));
  OR4        u0689(.A(men_men_n711_), .B(men_men_n672_), .C(men_men_n657_), .D(men_men_n602_), .Y(men5));
  AOI210     u0690(.A0(men_men_n641_), .A1(men_men_n259_), .B0(men_men_n408_), .Y(men_men_n713_));
  AN2        u0691(.A(men_men_n24_), .B(i_10_), .Y(men_men_n714_));
  NA3        u0692(.A(men_men_n714_), .B(men_men_n703_), .C(men_men_n102_), .Y(men_men_n715_));
  NA2        u0693(.A(men_men_n715_), .B(men_men_n713_), .Y(men_men_n716_));
  NO3        u0694(.A(i_11_), .B(men_men_n232_), .C(i_13_), .Y(men_men_n717_));
  NO2        u0695(.A(men_men_n118_), .B(men_men_n23_), .Y(men_men_n718_));
  NA2        u0696(.A(i_12_), .B(i_8_), .Y(men_men_n719_));
  OAI210     u0697(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n719_), .Y(men_men_n720_));
  INV        u0698(.A(men_men_n435_), .Y(men_men_n721_));
  AOI220     u0699(.A0(men_men_n308_), .A1(men_men_n559_), .B0(men_men_n720_), .B1(men_men_n718_), .Y(men_men_n722_));
  INV        u0700(.A(men_men_n722_), .Y(men_men_n723_));
  NO2        u0701(.A(men_men_n723_), .B(men_men_n716_), .Y(men_men_n724_));
  INV        u0702(.A(men_men_n166_), .Y(men_men_n725_));
  INV        u0703(.A(men_men_n239_), .Y(men_men_n726_));
  OAI210     u0704(.A0(men_men_n668_), .A1(men_men_n437_), .B0(men_men_n104_), .Y(men_men_n727_));
  AOI210     u0705(.A0(men_men_n727_), .A1(men_men_n726_), .B0(men_men_n725_), .Y(men_men_n728_));
  NO2        u0706(.A(men_men_n444_), .B(men_men_n26_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n729_), .B(men_men_n410_), .Y(men_men_n730_));
  NA2        u0708(.A(men_men_n730_), .B(i_2_), .Y(men_men_n731_));
  INV        u0709(.A(men_men_n731_), .Y(men_men_n732_));
  AOI210     u0710(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n407_), .Y(men_men_n733_));
  AOI210     u0711(.A0(men_men_n733_), .A1(men_men_n732_), .B0(men_men_n728_), .Y(men_men_n734_));
  NO2        u0712(.A(men_men_n184_), .B(men_men_n119_), .Y(men_men_n735_));
  OAI210     u0713(.A0(men_men_n735_), .A1(men_men_n718_), .B0(i_2_), .Y(men_men_n736_));
  NO2        u0714(.A(men_men_n736_), .B(men_men_n187_), .Y(men_men_n737_));
  OA210      u0715(.A0(men_men_n605_), .A1(men_men_n120_), .B0(i_13_), .Y(men_men_n738_));
  NA2        u0716(.A(men_men_n194_), .B(men_men_n197_), .Y(men_men_n739_));
  NA2        u0717(.A(men_men_n146_), .B(men_men_n582_), .Y(men_men_n740_));
  AOI210     u0718(.A0(men_men_n740_), .A1(men_men_n739_), .B0(men_men_n361_), .Y(men_men_n741_));
  AOI210     u0719(.A0(men_men_n203_), .A1(men_men_n142_), .B0(men_men_n506_), .Y(men_men_n742_));
  NA2        u0720(.A(men_men_n742_), .B(men_men_n410_), .Y(men_men_n743_));
  NO2        u0721(.A(men_men_n96_), .B(men_men_n45_), .Y(men_men_n744_));
  INV        u0722(.A(men_men_n291_), .Y(men_men_n745_));
  NA4        u0723(.A(men_men_n745_), .B(men_men_n295_), .C(men_men_n118_), .D(men_men_n43_), .Y(men_men_n746_));
  OAI210     u0724(.A0(men_men_n746_), .A1(men_men_n744_), .B0(men_men_n743_), .Y(men_men_n747_));
  NO4        u0725(.A(men_men_n747_), .B(men_men_n741_), .C(men_men_n738_), .D(men_men_n737_), .Y(men_men_n748_));
  NA2        u0726(.A(men_men_n559_), .B(men_men_n28_), .Y(men_men_n749_));
  NA2        u0727(.A(men_men_n717_), .B(men_men_n265_), .Y(men_men_n750_));
  NA2        u0728(.A(men_men_n750_), .B(men_men_n749_), .Y(men_men_n751_));
  NO2        u0729(.A(men_men_n62_), .B(i_12_), .Y(men_men_n752_));
  NO2        u0730(.A(men_men_n752_), .B(men_men_n120_), .Y(men_men_n753_));
  NO2        u0731(.A(men_men_n753_), .B(men_men_n582_), .Y(men_men_n754_));
  AOI220     u0732(.A0(men_men_n754_), .A1(men_men_n36_), .B0(men_men_n751_), .B1(men_men_n47_), .Y(men_men_n755_));
  NA4        u0733(.A(men_men_n755_), .B(men_men_n748_), .C(men_men_n734_), .D(men_men_n724_), .Y(men6));
  NA2        u0734(.A(men_men_n25_), .B(men_men_n708_), .Y(men_men_n757_));
  NA4        u0735(.A(men_men_n377_), .B(men_men_n473_), .C(men_men_n69_), .D(men_men_n95_), .Y(men_men_n758_));
  INV        u0736(.A(men_men_n758_), .Y(men_men_n759_));
  NO2        u0737(.A(i_11_), .B(i_9_), .Y(men_men_n760_));
  NO2        u0738(.A(men_men_n759_), .B(men_men_n319_), .Y(men_men_n761_));
  AO210      u0739(.A0(men_men_n761_), .A1(men_men_n757_), .B0(i_12_), .Y(men_men_n762_));
  NA2        u0740(.A(men_men_n362_), .B(men_men_n325_), .Y(men_men_n763_));
  NA2        u0741(.A(men_men_n566_), .B(men_men_n63_), .Y(men_men_n764_));
  INV        u0742(.A(men_men_n659_), .Y(men_men_n765_));
  NA4        u0743(.A(men_men_n84_), .B(men_men_n765_), .C(men_men_n764_), .D(men_men_n763_), .Y(men_men_n766_));
  INV        u0744(.A(men_men_n191_), .Y(men_men_n767_));
  AOI220     u0745(.A0(men_men_n767_), .A1(men_men_n760_), .B0(men_men_n766_), .B1(men_men_n71_), .Y(men_men_n768_));
  NO2        u0746(.A(men_men_n246_), .B(i_9_), .Y(men_men_n769_));
  NA2        u0747(.A(men_men_n769_), .B(men_men_n752_), .Y(men_men_n770_));
  AOI210     u0748(.A0(men_men_n770_), .A1(men_men_n505_), .B0(men_men_n179_), .Y(men_men_n771_));
  NA3        u0749(.A(men_men_n1022_), .B(men_men_n464_), .C(men_men_n377_), .Y(men_men_n772_));
  NAi32      u0750(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n773_));
  AOI210     u0751(.A0(men_men_n691_), .A1(men_men_n84_), .B0(men_men_n773_), .Y(men_men_n774_));
  OAI210     u0752(.A0(men_men_n658_), .A1(men_men_n547_), .B0(men_men_n546_), .Y(men_men_n775_));
  NAi31      u0753(.An(men_men_n774_), .B(men_men_n775_), .C(men_men_n772_), .Y(men_men_n776_));
  OR2        u0754(.A(men_men_n776_), .B(men_men_n771_), .Y(men_men_n777_));
  NO2        u0755(.A(i_11_), .B(i_2_), .Y(men_men_n778_));
  NA2        u0756(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n779_));
  NO2        u0757(.A(men_men_n779_), .B(men_men_n399_), .Y(men_men_n780_));
  NA2        u0758(.A(men_men_n780_), .B(men_men_n778_), .Y(men_men_n781_));
  NA3        u0759(.A(men_men_n339_), .B(men_men_n248_), .C(i_7_), .Y(men_men_n782_));
  BUFFER     u0760(.A(men_men_n605_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(men_men_n141_), .Y(men_men_n784_));
  OR2        u0762(.A(men_men_n721_), .B(men_men_n36_), .Y(men_men_n785_));
  NA4        u0763(.A(men_men_n785_), .B(men_men_n784_), .C(men_men_n782_), .D(men_men_n781_), .Y(men_men_n786_));
  NA2        u0764(.A(men_men_n384_), .B(men_men_n68_), .Y(men_men_n787_));
  NA2        u0765(.A(men_men_n787_), .B(men_men_n588_), .Y(men_men_n788_));
  NA3        u0766(.A(men_men_n506_), .B(men_men_n474_), .C(men_men_n214_), .Y(men_men_n789_));
  INV        u0767(.A(men_men_n545_), .Y(men_men_n790_));
  NA2        u0768(.A(men_men_n105_), .B(men_men_n398_), .Y(men_men_n791_));
  NA2        u0769(.A(men_men_n238_), .B(men_men_n47_), .Y(men_men_n792_));
  INV        u0770(.A(men_men_n573_), .Y(men_men_n793_));
  NA3        u0771(.A(men_men_n793_), .B(men_men_n318_), .C(i_7_), .Y(men_men_n794_));
  NA4        u0772(.A(men_men_n794_), .B(men_men_n791_), .C(men_men_n790_), .D(men_men_n789_), .Y(men_men_n795_));
  NO4        u0773(.A(men_men_n795_), .B(men_men_n788_), .C(men_men_n786_), .D(men_men_n777_), .Y(men_men_n796_));
  NA4        u0774(.A(men_men_n796_), .B(men_men_n768_), .C(men_men_n762_), .D(men_men_n367_), .Y(men3));
  NA2        u0775(.A(i_12_), .B(i_10_), .Y(men_men_n798_));
  NA2        u0776(.A(i_6_), .B(i_7_), .Y(men_men_n799_));
  NO2        u0777(.A(men_men_n799_), .B(i_0_), .Y(men_men_n800_));
  NO2        u0778(.A(i_11_), .B(men_men_n232_), .Y(men_men_n801_));
  OAI210     u0779(.A0(men_men_n800_), .A1(men_men_n279_), .B0(men_men_n801_), .Y(men_men_n802_));
  NO2        u0780(.A(men_men_n802_), .B(men_men_n187_), .Y(men_men_n803_));
  NO3        u0781(.A(men_men_n440_), .B(men_men_n86_), .C(men_men_n45_), .Y(men_men_n804_));
  OA210      u0782(.A0(men_men_n804_), .A1(men_men_n803_), .B0(men_men_n168_), .Y(men_men_n805_));
  NA2        u0783(.A(men_men_n588_), .B(men_men_n360_), .Y(men_men_n806_));
  NA2        u0784(.A(men_men_n806_), .B(men_men_n40_), .Y(men_men_n807_));
  NO3        u0785(.A(men_men_n612_), .B(men_men_n444_), .C(men_men_n125_), .Y(men_men_n808_));
  NA2        u0786(.A(men_men_n400_), .B(men_men_n46_), .Y(men_men_n809_));
  AOI210     u0787(.A0(men_men_n1018_), .A1(men_men_n807_), .B0(men_men_n49_), .Y(men_men_n810_));
  NA2        u0788(.A(men_men_n179_), .B(men_men_n555_), .Y(men_men_n811_));
  NA2        u0789(.A(men_men_n683_), .B(men_men_n651_), .Y(men_men_n812_));
  NA2        u0790(.A(i_0_), .B(men_men_n427_), .Y(men_men_n813_));
  OAI220     u0791(.A0(men_men_n813_), .A1(men_men_n812_), .B0(men_men_n811_), .B1(men_men_n63_), .Y(men_men_n814_));
  NOi21      u0792(.An(i_5_), .B(i_9_), .Y(men_men_n815_));
  NA2        u0793(.A(men_men_n815_), .B(men_men_n434_), .Y(men_men_n816_));
  AOI210     u0794(.A0(men_men_n256_), .A1(men_men_n466_), .B0(men_men_n662_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n169_), .B(men_men_n142_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n818_), .B(men_men_n238_), .Y(men_men_n819_));
  OAI220     u0797(.A0(men_men_n819_), .A1(men_men_n174_), .B0(men_men_n817_), .B1(men_men_n816_), .Y(men_men_n820_));
  NO4        u0798(.A(men_men_n820_), .B(men_men_n814_), .C(men_men_n810_), .D(men_men_n805_), .Y(men_men_n821_));
  NA2        u0799(.A(men_men_n179_), .B(men_men_n24_), .Y(men_men_n822_));
  NO2        u0800(.A(men_men_n649_), .B(men_men_n579_), .Y(men_men_n823_));
  NO2        u0801(.A(men_men_n823_), .B(men_men_n822_), .Y(men_men_n824_));
  NA2        u0802(.A(men_men_n302_), .B(men_men_n123_), .Y(men_men_n825_));
  NAi21      u0803(.An(men_men_n157_), .B(men_men_n427_), .Y(men_men_n826_));
  OAI220     u0804(.A0(men_men_n826_), .A1(men_men_n792_), .B0(men_men_n825_), .B1(men_men_n389_), .Y(men_men_n827_));
  NO2        u0805(.A(men_men_n827_), .B(men_men_n824_), .Y(men_men_n828_));
  NA2        u0806(.A(men_men_n556_), .B(i_0_), .Y(men_men_n829_));
  NO2        u0807(.A(men_men_n829_), .B(men_men_n372_), .Y(men_men_n830_));
  NO4        u0808(.A(men_men_n572_), .B(men_men_n211_), .C(men_men_n407_), .D(men_men_n399_), .Y(men_men_n831_));
  AOI210     u0809(.A0(men_men_n831_), .A1(i_11_), .B0(men_men_n830_), .Y(men_men_n832_));
  NA2        u0810(.A(men_men_n717_), .B(men_men_n319_), .Y(men_men_n833_));
  INV        u0811(.A(men_men_n58_), .Y(men_men_n834_));
  OAI220     u0812(.A0(men_men_n834_), .A1(men_men_n833_), .B0(men_men_n636_), .B1(men_men_n522_), .Y(men_men_n835_));
  NA2        u0813(.A(i_0_), .B(i_10_), .Y(men_men_n836_));
  OAI210     u0814(.A0(men_men_n836_), .A1(men_men_n83_), .B0(men_men_n523_), .Y(men_men_n837_));
  NO4        u0815(.A(men_men_n108_), .B(men_men_n58_), .C(men_men_n646_), .D(i_5_), .Y(men_men_n838_));
  AN2        u0816(.A(men_men_n838_), .B(men_men_n837_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n179_), .B(men_men_n82_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n550_), .B(i_4_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n182_), .B(men_men_n197_), .Y(men_men_n842_));
  OAI220     u0820(.A0(men_men_n842_), .A1(men_men_n833_), .B0(men_men_n841_), .B1(men_men_n840_), .Y(men_men_n843_));
  NO3        u0821(.A(men_men_n843_), .B(men_men_n839_), .C(men_men_n835_), .Y(men_men_n844_));
  NA3        u0822(.A(men_men_n844_), .B(men_men_n832_), .C(men_men_n828_), .Y(men_men_n845_));
  NO2        u0823(.A(men_men_n97_), .B(men_men_n37_), .Y(men_men_n846_));
  NA2        u0824(.A(i_11_), .B(i_9_), .Y(men_men_n847_));
  NO3        u0825(.A(i_12_), .B(men_men_n847_), .C(men_men_n587_), .Y(men_men_n848_));
  AN2        u0826(.A(men_men_n848_), .B(men_men_n846_), .Y(men_men_n849_));
  NO2        u0827(.A(men_men_n49_), .B(i_7_), .Y(men_men_n850_));
  NA2        u0828(.A(men_men_n381_), .B(men_men_n173_), .Y(men_men_n851_));
  NA2        u0829(.A(men_men_n851_), .B(men_men_n155_), .Y(men_men_n852_));
  NO2        u0830(.A(men_men_n847_), .B(men_men_n71_), .Y(men_men_n853_));
  NO2        u0831(.A(men_men_n169_), .B(i_0_), .Y(men_men_n854_));
  INV        u0832(.A(men_men_n854_), .Y(men_men_n855_));
  NA2        u0833(.A(men_men_n464_), .B(men_men_n226_), .Y(men_men_n856_));
  AOI210     u0834(.A0(men_men_n359_), .A1(men_men_n42_), .B0(men_men_n397_), .Y(men_men_n857_));
  OAI220     u0835(.A0(men_men_n857_), .A1(men_men_n816_), .B0(men_men_n856_), .B1(men_men_n855_), .Y(men_men_n858_));
  NO3        u0836(.A(men_men_n858_), .B(men_men_n852_), .C(men_men_n849_), .Y(men_men_n859_));
  NA2        u0837(.A(men_men_n635_), .B(men_men_n115_), .Y(men_men_n860_));
  NO2        u0838(.A(i_6_), .B(men_men_n860_), .Y(men_men_n861_));
  AOI210     u0839(.A0(men_men_n436_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n862_));
  NA2        u0840(.A(men_men_n166_), .B(men_men_n97_), .Y(men_men_n863_));
  NOi32      u0841(.An(men_men_n862_), .Bn(men_men_n182_), .C(men_men_n863_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n589_), .B(men_men_n319_), .Y(men_men_n865_));
  NO2        u0843(.A(men_men_n865_), .B(men_men_n809_), .Y(men_men_n866_));
  NO3        u0844(.A(men_men_n866_), .B(men_men_n864_), .C(men_men_n861_), .Y(men_men_n867_));
  NOi21      u0845(.An(i_7_), .B(i_5_), .Y(men_men_n868_));
  NOi31      u0846(.An(men_men_n868_), .B(i_0_), .C(men_men_n697_), .Y(men_men_n869_));
  NA3        u0847(.A(men_men_n869_), .B(men_men_n371_), .C(i_6_), .Y(men_men_n870_));
  OA210      u0848(.A0(men_men_n863_), .A1(men_men_n505_), .B0(men_men_n870_), .Y(men_men_n871_));
  NO3        u0849(.A(men_men_n392_), .B(men_men_n348_), .C(men_men_n346_), .Y(men_men_n872_));
  NO2        u0850(.A(men_men_n250_), .B(men_men_n309_), .Y(men_men_n873_));
  NO2        u0851(.A(men_men_n697_), .B(men_men_n249_), .Y(men_men_n874_));
  AOI210     u0852(.A0(men_men_n874_), .A1(men_men_n873_), .B0(men_men_n872_), .Y(men_men_n875_));
  NA4        u0853(.A(men_men_n875_), .B(men_men_n871_), .C(men_men_n867_), .D(men_men_n859_), .Y(men_men_n876_));
  NO2        u0854(.A(men_men_n822_), .B(men_men_n234_), .Y(men_men_n877_));
  AN2        u0855(.A(men_men_n323_), .B(men_men_n319_), .Y(men_men_n878_));
  AN2        u0856(.A(men_men_n878_), .B(men_men_n818_), .Y(men_men_n879_));
  OAI210     u0857(.A0(men_men_n879_), .A1(men_men_n877_), .B0(i_10_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n798_), .B(men_men_n308_), .Y(men_men_n881_));
  NA2        u0859(.A(men_men_n881_), .B(men_men_n853_), .Y(men_men_n882_));
  NA3        u0860(.A(men_men_n463_), .B(men_men_n400_), .C(men_men_n46_), .Y(men_men_n883_));
  OAI210     u0861(.A0(men_men_n826_), .A1(i_7_), .B0(men_men_n883_), .Y(men_men_n884_));
  NO2        u0862(.A(men_men_n248_), .B(men_men_n47_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n853_), .B(men_men_n295_), .Y(men_men_n886_));
  OAI210     u0864(.A0(men_men_n885_), .A1(men_men_n181_), .B0(men_men_n886_), .Y(men_men_n887_));
  AOI220     u0865(.A0(men_men_n887_), .A1(men_men_n464_), .B0(men_men_n884_), .B1(men_men_n71_), .Y(men_men_n888_));
  NO2        u0866(.A(men_men_n73_), .B(men_men_n719_), .Y(men_men_n889_));
  AOI210     u0867(.A0(men_men_n168_), .A1(men_men_n579_), .B0(men_men_n889_), .Y(men_men_n890_));
  NO2        u0868(.A(men_men_n890_), .B(men_men_n48_), .Y(men_men_n891_));
  NO3        u0869(.A(men_men_n572_), .B(i_0_), .C(men_men_n24_), .Y(men_men_n892_));
  AOI210     u0870(.A0(men_men_n677_), .A1(men_men_n531_), .B0(men_men_n892_), .Y(men_men_n893_));
  NAi21      u0871(.An(i_9_), .B(i_5_), .Y(men_men_n894_));
  NO2        u0872(.A(men_men_n894_), .B(men_men_n392_), .Y(men_men_n895_));
  NO2        u0873(.A(men_men_n584_), .B(men_men_n99_), .Y(men_men_n896_));
  AOI220     u0874(.A0(men_men_n896_), .A1(i_0_), .B0(men_men_n895_), .B1(men_men_n605_), .Y(men_men_n897_));
  OAI220     u0875(.A0(men_men_n897_), .A1(men_men_n83_), .B0(men_men_n893_), .B1(men_men_n167_), .Y(men_men_n898_));
  NO2        u0876(.A(men_men_n898_), .B(men_men_n891_), .Y(men_men_n899_));
  NA4        u0877(.A(men_men_n899_), .B(men_men_n888_), .C(men_men_n882_), .D(men_men_n880_), .Y(men_men_n900_));
  NO3        u0878(.A(men_men_n900_), .B(men_men_n876_), .C(men_men_n845_), .Y(men_men_n901_));
  NO2        u0879(.A(i_0_), .B(men_men_n697_), .Y(men_men_n902_));
  NA2        u0880(.A(men_men_n71_), .B(men_men_n45_), .Y(men_men_n903_));
  NO3        u0881(.A(men_men_n99_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n904_));
  AO220      u0882(.A0(men_men_n904_), .A1(men_men_n45_), .B0(men_men_n902_), .B1(men_men_n168_), .Y(men_men_n905_));
  NO2        u0883(.A(men_men_n764_), .B(men_men_n863_), .Y(men_men_n906_));
  AOI210     u0884(.A0(men_men_n905_), .A1(men_men_n336_), .B0(men_men_n906_), .Y(men_men_n907_));
  NA2        u0885(.A(men_men_n708_), .B(men_men_n140_), .Y(men_men_n908_));
  INV        u0886(.A(men_men_n908_), .Y(men_men_n909_));
  NA2        u0887(.A(men_men_n909_), .B(men_men_n651_), .Y(men_men_n910_));
  NO2        u0888(.A(men_men_n775_), .B(men_men_n392_), .Y(men_men_n911_));
  NA3        u0889(.A(men_men_n800_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n912_));
  NA2        u0890(.A(men_men_n801_), .B(i_9_), .Y(men_men_n913_));
  AOI210     u0891(.A0(men_men_n912_), .A1(men_men_n488_), .B0(men_men_n913_), .Y(men_men_n914_));
  OAI210     u0892(.A0(men_men_n238_), .A1(i_9_), .B0(men_men_n225_), .Y(men_men_n915_));
  AOI210     u0893(.A0(men_men_n915_), .A1(men_men_n829_), .B0(men_men_n148_), .Y(men_men_n916_));
  NO3        u0894(.A(men_men_n916_), .B(men_men_n914_), .C(men_men_n911_), .Y(men_men_n917_));
  NA3        u0895(.A(men_men_n917_), .B(men_men_n910_), .C(men_men_n907_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n878_), .B(men_men_n361_), .Y(men_men_n919_));
  AOI210     u0897(.A0(men_men_n290_), .A1(men_men_n157_), .B0(men_men_n919_), .Y(men_men_n920_));
  NA3        u0898(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n921_));
  NA2        u0899(.A(men_men_n850_), .B(men_men_n478_), .Y(men_men_n922_));
  AOI210     u0900(.A0(men_men_n921_), .A1(men_men_n157_), .B0(men_men_n922_), .Y(men_men_n923_));
  NO2        u0901(.A(men_men_n923_), .B(men_men_n920_), .Y(men_men_n924_));
  NO3        u0902(.A(men_men_n836_), .B(men_men_n815_), .C(men_men_n184_), .Y(men_men_n925_));
  AOI220     u0903(.A0(men_men_n925_), .A1(i_11_), .B0(men_men_n551_), .B1(men_men_n73_), .Y(men_men_n926_));
  NO3        u0904(.A(men_men_n205_), .B(men_men_n370_), .C(i_0_), .Y(men_men_n927_));
  OAI210     u0905(.A0(men_men_n927_), .A1(men_men_n74_), .B0(i_13_), .Y(men_men_n928_));
  INV        u0906(.A(men_men_n214_), .Y(men_men_n929_));
  NO2        u0907(.A(i_12_), .B(men_men_n599_), .Y(men_men_n930_));
  NA3        u0908(.A(men_men_n930_), .B(men_men_n1021_), .C(men_men_n929_), .Y(men_men_n931_));
  NA4        u0909(.A(men_men_n931_), .B(men_men_n928_), .C(men_men_n926_), .D(men_men_n924_), .Y(men_men_n932_));
  NO2        u0910(.A(men_men_n237_), .B(men_men_n88_), .Y(men_men_n933_));
  NA2        u0911(.A(men_men_n933_), .B(men_men_n902_), .Y(men_men_n934_));
  AOI220     u0912(.A0(men_men_n868_), .A1(men_men_n478_), .B0(men_men_n800_), .B1(men_men_n158_), .Y(men_men_n935_));
  NA2        u0913(.A(men_men_n339_), .B(men_men_n170_), .Y(men_men_n936_));
  OA220      u0914(.A0(men_men_n936_), .A1(men_men_n935_), .B0(men_men_n934_), .B1(i_5_), .Y(men_men_n937_));
  AOI210     u0915(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n169_), .Y(men_men_n938_));
  NA3        u0916(.A(men_men_n596_), .B(men_men_n179_), .C(men_men_n82_), .Y(men_men_n939_));
  NA2        u0917(.A(men_men_n939_), .B(men_men_n530_), .Y(men_men_n940_));
  NO3        u0918(.A(men_men_n809_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n941_));
  NA3        u0919(.A(men_men_n482_), .B(men_men_n477_), .C(men_men_n461_), .Y(men_men_n942_));
  NO3        u0920(.A(men_men_n942_), .B(men_men_n941_), .C(men_men_n940_), .Y(men_men_n943_));
  NA3        u0921(.A(men_men_n377_), .B(men_men_n166_), .C(men_men_n165_), .Y(men_men_n944_));
  NA3        u0922(.A(men_men_n850_), .B(men_men_n279_), .C(men_men_n225_), .Y(men_men_n945_));
  NA2        u0923(.A(men_men_n945_), .B(men_men_n944_), .Y(men_men_n946_));
  NA3        u0924(.A(men_men_n377_), .B(men_men_n324_), .C(men_men_n217_), .Y(men_men_n947_));
  INV        u0925(.A(men_men_n947_), .Y(men_men_n948_));
  NOi31      u0926(.An(men_men_n376_), .B(men_men_n903_), .C(men_men_n234_), .Y(men_men_n949_));
  NO3        u0927(.A(men_men_n847_), .B(men_men_n214_), .C(men_men_n184_), .Y(men_men_n950_));
  NO4        u0928(.A(men_men_n950_), .B(men_men_n949_), .C(men_men_n948_), .D(men_men_n946_), .Y(men_men_n951_));
  NA3        u0929(.A(men_men_n951_), .B(men_men_n943_), .C(men_men_n937_), .Y(men_men_n952_));
  INV        u0930(.A(men_men_n598_), .Y(men_men_n953_));
  NO3        u0931(.A(men_men_n953_), .B(men_men_n541_), .C(i_3_), .Y(men_men_n954_));
  NO2        u0932(.A(men_men_n83_), .B(i_5_), .Y(men_men_n955_));
  NA3        u0933(.A(men_men_n801_), .B(men_men_n103_), .C(men_men_n118_), .Y(men_men_n956_));
  INV        u0934(.A(men_men_n956_), .Y(men_men_n957_));
  AOI210     u0935(.A0(men_men_n957_), .A1(men_men_n955_), .B0(men_men_n954_), .Y(men_men_n958_));
  NA3        u0936(.A(men_men_n295_), .B(i_5_), .C(men_men_n187_), .Y(men_men_n959_));
  NA2        u0937(.A(men_men_n959_), .B(men_men_n237_), .Y(men_men_n960_));
  NO4        u0938(.A(men_men_n234_), .B(men_men_n205_), .C(i_0_), .D(i_12_), .Y(men_men_n961_));
  AOI220     u0939(.A0(men_men_n961_), .A1(men_men_n960_), .B0(men_men_n759_), .B1(men_men_n170_), .Y(men_men_n962_));
  AN2        u0940(.A(men_men_n836_), .B(men_men_n148_), .Y(men_men_n963_));
  NO4        u0941(.A(men_men_n963_), .B(i_12_), .C(men_men_n626_), .D(men_men_n125_), .Y(men_men_n964_));
  NA2        u0942(.A(men_men_n964_), .B(men_men_n214_), .Y(men_men_n965_));
  NA3        u0943(.A(men_men_n92_), .B(men_men_n555_), .C(i_11_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n966_), .B(men_men_n150_), .Y(men_men_n967_));
  NA2        u0945(.A(men_men_n868_), .B(men_men_n460_), .Y(men_men_n968_));
  OAI220     u0946(.A0(i_7_), .A1(men_men_n959_), .B0(men_men_n968_), .B1(men_men_n652_), .Y(men_men_n969_));
  AOI210     u0947(.A0(men_men_n969_), .A1(men_men_n854_), .B0(men_men_n967_), .Y(men_men_n970_));
  NA4        u0948(.A(men_men_n970_), .B(men_men_n965_), .C(men_men_n962_), .D(men_men_n958_), .Y(men_men_n971_));
  NO4        u0949(.A(men_men_n971_), .B(men_men_n952_), .C(men_men_n932_), .D(men_men_n918_), .Y(men_men_n972_));
  NA3        u0950(.A(men_men_n862_), .B(men_men_n356_), .C(i_5_), .Y(men_men_n973_));
  NA2        u0951(.A(men_men_n973_), .B(men_men_n594_), .Y(men_men_n974_));
  NA2        u0952(.A(men_men_n974_), .B(men_men_n201_), .Y(men_men_n975_));
  NA2        u0953(.A(men_men_n180_), .B(men_men_n182_), .Y(men_men_n976_));
  AO210      u0954(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n976_), .Y(men_men_n977_));
  OAI210     u0955(.A0(men_men_n598_), .A1(men_men_n596_), .B0(men_men_n308_), .Y(men_men_n978_));
  NA2        u0956(.A(men_men_n978_), .B(men_men_n977_), .Y(men_men_n979_));
  NO4        u0957(.A(men_men_n228_), .B(men_men_n139_), .C(men_men_n655_), .D(men_men_n37_), .Y(men_men_n980_));
  NO2        u0958(.A(men_men_n980_), .B(men_men_n831_), .Y(men_men_n981_));
  OAI210     u0959(.A0(men_men_n966_), .A1(men_men_n142_), .B0(men_men_n981_), .Y(men_men_n982_));
  AOI210     u0960(.A0(men_men_n979_), .A1(men_men_n49_), .B0(men_men_n982_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n983_), .A1(men_men_n975_), .B0(men_men_n71_), .Y(men_men_n984_));
  NO2        u0962(.A(men_men_n548_), .B(men_men_n366_), .Y(men_men_n985_));
  NO2        u0963(.A(men_men_n985_), .B(men_men_n725_), .Y(men_men_n986_));
  INV        u0964(.A(men_men_n74_), .Y(men_men_n987_));
  AOI210     u0965(.A0(men_men_n938_), .A1(men_men_n850_), .B0(men_men_n869_), .Y(men_men_n988_));
  AOI210     u0966(.A0(men_men_n988_), .A1(men_men_n987_), .B0(men_men_n655_), .Y(men_men_n989_));
  NA2        u0967(.A(i_8_), .B(men_men_n74_), .Y(men_men_n990_));
  NO2        u0968(.A(men_men_n990_), .B(men_men_n232_), .Y(men_men_n991_));
  NA3        u0969(.A(men_men_n90_), .B(men_men_n297_), .C(men_men_n31_), .Y(men_men_n992_));
  INV        u0970(.A(men_men_n992_), .Y(men_men_n993_));
  NO3        u0971(.A(men_men_n993_), .B(men_men_n991_), .C(men_men_n989_), .Y(men_men_n994_));
  OAI210     u0972(.A0(men_men_n258_), .A1(men_men_n153_), .B0(men_men_n85_), .Y(men_men_n995_));
  NA3        u0973(.A(men_men_n729_), .B(men_men_n279_), .C(men_men_n78_), .Y(men_men_n996_));
  AOI210     u0974(.A0(men_men_n996_), .A1(men_men_n995_), .B0(i_11_), .Y(men_men_n997_));
  NA2        u0975(.A(men_men_n590_), .B(men_men_n211_), .Y(men_men_n998_));
  OAI210     u0976(.A0(men_men_n998_), .A1(men_men_n862_), .B0(men_men_n201_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n159_), .B(i_5_), .Y(men_men_n1000_));
  NO2        u0978(.A(men_men_n999_), .B(men_men_n1000_), .Y(men_men_n1001_));
  NO3        u0979(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1002_));
  OAI210     u0980(.A0(men_men_n873_), .A1(men_men_n297_), .B0(men_men_n1002_), .Y(men_men_n1003_));
  NO2        u0981(.A(men_men_n1003_), .B(men_men_n697_), .Y(men_men_n1004_));
  NO3        u0982(.A(men_men_n894_), .B(men_men_n467_), .C(men_men_n247_), .Y(men_men_n1005_));
  NO2        u0983(.A(men_men_n1005_), .B(men_men_n545_), .Y(men_men_n1006_));
  INV        u0984(.A(men_men_n349_), .Y(men_men_n1007_));
  AOI210     u0985(.A0(men_men_n1007_), .A1(men_men_n1006_), .B0(men_men_n41_), .Y(men_men_n1008_));
  NO4        u0986(.A(men_men_n1008_), .B(men_men_n1004_), .C(men_men_n1001_), .D(men_men_n997_), .Y(men_men_n1009_));
  OAI210     u0987(.A0(men_men_n994_), .A1(i_4_), .B0(men_men_n1009_), .Y(men_men_n1010_));
  NO3        u0988(.A(men_men_n1010_), .B(men_men_n986_), .C(men_men_n984_), .Y(men_men_n1011_));
  NA4        u0989(.A(men_men_n1011_), .B(men_men_n972_), .C(men_men_n901_), .D(men_men_n821_), .Y(men4));
  INV        u0990(.A(men_men_n676_), .Y(men_men_n1015_));
  INV        u0991(.A(i_2_), .Y(men_men_n1016_));
  INV        u0992(.A(men_men_n687_), .Y(men_men_n1017_));
  INV        u0993(.A(men_men_n808_), .Y(men_men_n1018_));
  INV        u0994(.A(men_men_n80_), .Y(men_men_n1019_));
  INV        u0995(.A(men_men_n138_), .Y(men_men_n1020_));
  INV        u0996(.A(i_3_), .Y(men_men_n1021_));
  INV        u0997(.A(i_11_), .Y(men_men_n1022_));
  INV        u0998(.A(men_men_n138_), .Y(men_men_n1023_));
  INV        u0999(.A(men_men_n237_), .Y(men_men_n1024_));
  INV        u1000(.A(i_8_), .Y(men_men_n1025_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule