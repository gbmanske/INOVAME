//Benchmark atmr_max1024_476_0.0156

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n62_), .B(ori_ori_n36_), .Y(ori_ori_n63_));
  INV        o047(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NO3        o048(.A(ori_ori_n64_), .B(ori_ori_n61_), .C(ori_ori_n60_), .Y(ori_ori_n65_));
  NO2        o049(.A(x7), .B(x6), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n67_));
  NO2        o051(.A(x8), .B(x2), .Y(ori_ori_n68_));
  INV        o052(.A(ori_ori_n68_), .Y(ori_ori_n69_));
  NO2        o053(.A(ori_ori_n69_), .B(x1), .Y(ori_ori_n70_));
  OA210      o054(.A0(ori_ori_n70_), .A1(ori_ori_n67_), .B0(ori_ori_n66_), .Y(ori_ori_n71_));
  OAI210     o055(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n72_));
  OAI210     o056(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n72_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n71_), .Y(ori_ori_n74_));
  OAI210     o058(.A0(ori_ori_n74_), .A1(ori_ori_n65_), .B0(x4), .Y(ori_ori_n75_));
  NA2        o059(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n76_));
  OAI210     o060(.A0(ori_ori_n76_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n77_));
  NA2        o061(.A(x5), .B(x3), .Y(ori_ori_n78_));
  NO2        o062(.A(x8), .B(x6), .Y(ori_ori_n79_));
  NO4        o063(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(ori_ori_n66_), .D(ori_ori_n54_), .Y(ori_ori_n80_));
  NAi21      o064(.An(x4), .B(x3), .Y(ori_ori_n81_));
  INV        o065(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n82_), .B(ori_ori_n22_), .Y(ori_ori_n83_));
  NO2        o067(.A(x4), .B(x2), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n84_), .B(x3), .Y(ori_ori_n85_));
  NO3        o069(.A(ori_ori_n85_), .B(ori_ori_n83_), .C(ori_ori_n18_), .Y(ori_ori_n86_));
  NO3        o070(.A(ori_ori_n86_), .B(ori_ori_n80_), .C(ori_ori_n77_), .Y(ori_ori_n87_));
  NA2        o071(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n88_), .B(ori_ori_n25_), .Y(ori_ori_n89_));
  INV        o073(.A(x8), .Y(ori_ori_n90_));
  NA2        o074(.A(x2), .B(x1), .Y(ori_ori_n91_));
  NO2        o075(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n92_));
  NO2        o076(.A(ori_ori_n92_), .B(ori_ori_n89_), .Y(ori_ori_n93_));
  NO2        o077(.A(ori_ori_n93_), .B(ori_ori_n26_), .Y(ori_ori_n94_));
  AOI210     o078(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n96_));
  NO3        o080(.A(ori_ori_n96_), .B(ori_ori_n95_), .C(ori_ori_n94_), .Y(ori_ori_n97_));
  NA2        o081(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n98_));
  NO2        o082(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n99_));
  OAI210     o083(.A0(ori_ori_n99_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n100_));
  AOI210     o084(.A0(ori_ori_n98_), .A1(ori_ori_n52_), .B0(ori_ori_n100_), .Y(ori_ori_n101_));
  NO2        o085(.A(x3), .B(x2), .Y(ori_ori_n102_));
  NA3        o086(.A(ori_ori_n102_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n103_));
  AOI210     o087(.A0(x8), .A1(x6), .B0(ori_ori_n103_), .Y(ori_ori_n104_));
  NA2        o088(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n105_));
  OAI210     o089(.A0(ori_ori_n105_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n106_));
  NO4        o090(.A(ori_ori_n106_), .B(ori_ori_n104_), .C(ori_ori_n101_), .D(ori_ori_n97_), .Y(ori_ori_n107_));
  AO210      o091(.A0(ori_ori_n87_), .A1(ori_ori_n75_), .B0(ori_ori_n107_), .Y(ori02));
  NO2        o092(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n109_));
  NO2        o093(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n110_));
  NA2        o094(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n111_));
  NA2        o095(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n112_));
  INV        o096(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  AOI220     o097(.A0(ori_ori_n113_), .A1(ori_ori_n110_), .B0(ori_ori_n109_), .B1(x4), .Y(ori_ori_n114_));
  NO3        o098(.A(ori_ori_n114_), .B(x7), .C(x5), .Y(ori_ori_n115_));
  NA2        o099(.A(x9), .B(x2), .Y(ori_ori_n116_));
  OR2        o100(.A(x8), .B(x0), .Y(ori_ori_n117_));
  INV        o101(.A(ori_ori_n117_), .Y(ori_ori_n118_));
  NAi21      o102(.An(x2), .B(x8), .Y(ori_ori_n119_));
  INV        o103(.A(ori_ori_n119_), .Y(ori_ori_n120_));
  NO2        o104(.A(x4), .B(x1), .Y(ori_ori_n121_));
  NA3        o105(.A(ori_ori_n121_), .B(x2), .C(ori_ori_n60_), .Y(ori_ori_n122_));
  NOi21      o106(.An(x0), .B(x1), .Y(ori_ori_n123_));
  NO3        o107(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n124_));
  NOi21      o108(.An(x0), .B(x4), .Y(ori_ori_n125_));
  NAi21      o109(.An(x8), .B(x7), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n126_), .B(ori_ori_n62_), .Y(ori_ori_n127_));
  AOI220     o111(.A0(ori_ori_n127_), .A1(ori_ori_n125_), .B0(ori_ori_n124_), .B1(ori_ori_n123_), .Y(ori_ori_n128_));
  AOI210     o112(.A0(ori_ori_n128_), .A1(ori_ori_n122_), .B0(ori_ori_n78_), .Y(ori_ori_n129_));
  NO2        o113(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n130_));
  NA2        o114(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n131_));
  AOI210     o115(.A0(ori_ori_n131_), .A1(ori_ori_n105_), .B0(ori_ori_n112_), .Y(ori_ori_n132_));
  OAI210     o116(.A0(ori_ori_n132_), .A1(ori_ori_n35_), .B0(ori_ori_n130_), .Y(ori_ori_n133_));
  NAi21      o117(.An(x0), .B(x4), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n134_), .B(x1), .Y(ori_ori_n135_));
  NO2        o119(.A(x7), .B(x0), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n84_), .B(ori_ori_n99_), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n137_), .B(x3), .Y(ori_ori_n138_));
  OAI210     o122(.A0(ori_ori_n136_), .A1(ori_ori_n135_), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n140_));
  NA2        o124(.A(x5), .B(x0), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n142_));
  NA3        o126(.A(ori_ori_n142_), .B(ori_ori_n141_), .C(ori_ori_n140_), .Y(ori_ori_n143_));
  NA4        o127(.A(ori_ori_n143_), .B(ori_ori_n139_), .C(ori_ori_n133_), .D(ori_ori_n36_), .Y(ori_ori_n144_));
  NO3        o128(.A(ori_ori_n144_), .B(ori_ori_n129_), .C(ori_ori_n115_), .Y(ori_ori_n145_));
  NO3        o129(.A(ori_ori_n78_), .B(ori_ori_n76_), .C(ori_ori_n24_), .Y(ori_ori_n146_));
  NO2        o130(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n147_));
  AOI220     o131(.A0(ori_ori_n123_), .A1(ori_ori_n147_), .B0(ori_ori_n67_), .B1(ori_ori_n17_), .Y(ori_ori_n148_));
  NO3        o132(.A(ori_ori_n148_), .B(ori_ori_n60_), .C(ori_ori_n62_), .Y(ori_ori_n149_));
  NA2        o133(.A(x7), .B(x3), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n98_), .B(x5), .Y(ori_ori_n151_));
  NO2        o135(.A(x9), .B(x7), .Y(ori_ori_n152_));
  NOi21      o136(.An(x8), .B(x0), .Y(ori_ori_n153_));
  OA210      o137(.A0(ori_ori_n152_), .A1(x1), .B0(ori_ori_n153_), .Y(ori_ori_n154_));
  NO2        o138(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n155_));
  INV        o139(.A(x7), .Y(ori_ori_n156_));
  NA2        o140(.A(ori_ori_n156_), .B(ori_ori_n18_), .Y(ori_ori_n157_));
  AOI220     o141(.A0(ori_ori_n157_), .A1(ori_ori_n155_), .B0(ori_ori_n109_), .B1(ori_ori_n38_), .Y(ori_ori_n158_));
  NO2        o142(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n159_), .B(ori_ori_n125_), .Y(ori_ori_n160_));
  NO2        o144(.A(ori_ori_n160_), .B(ori_ori_n158_), .Y(ori_ori_n161_));
  AOI210     o145(.A0(ori_ori_n154_), .A1(ori_ori_n151_), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  OAI210     o146(.A0(ori_ori_n150_), .A1(ori_ori_n50_), .B0(ori_ori_n162_), .Y(ori_ori_n163_));
  NA2        o147(.A(x5), .B(x1), .Y(ori_ori_n164_));
  INV        o148(.A(ori_ori_n164_), .Y(ori_ori_n165_));
  AOI210     o149(.A0(ori_ori_n165_), .A1(ori_ori_n125_), .B0(ori_ori_n36_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n62_), .B(ori_ori_n90_), .Y(ori_ori_n167_));
  NAi21      o151(.An(x2), .B(x7), .Y(ori_ori_n168_));
  NO3        o152(.A(ori_ori_n168_), .B(ori_ori_n167_), .C(ori_ori_n48_), .Y(ori_ori_n169_));
  NA2        o153(.A(ori_ori_n169_), .B(ori_ori_n67_), .Y(ori_ori_n170_));
  NAi31      o154(.An(ori_ori_n78_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n171_));
  NA3        o155(.A(ori_ori_n171_), .B(ori_ori_n170_), .C(ori_ori_n166_), .Y(ori_ori_n172_));
  NO4        o156(.A(ori_ori_n172_), .B(ori_ori_n163_), .C(ori_ori_n149_), .D(ori_ori_n146_), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n173_), .B(ori_ori_n145_), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n141_), .B(ori_ori_n137_), .Y(ori_ori_n175_));
  NA2        o159(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n176_));
  NA2        o160(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n177_));
  NA3        o161(.A(ori_ori_n177_), .B(ori_ori_n176_), .C(ori_ori_n24_), .Y(ori_ori_n178_));
  AN2        o162(.A(ori_ori_n178_), .B(ori_ori_n142_), .Y(ori_ori_n179_));
  NA2        o163(.A(x8), .B(x0), .Y(ori_ori_n180_));
  NO2        o164(.A(ori_ori_n156_), .B(ori_ori_n25_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n123_), .B(x4), .Y(ori_ori_n182_));
  NA2        o166(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n183_));
  AOI210     o167(.A0(ori_ori_n180_), .A1(ori_ori_n131_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  NA2        o168(.A(x2), .B(x0), .Y(ori_ori_n185_));
  NA2        o169(.A(x4), .B(x1), .Y(ori_ori_n186_));
  NAi21      o170(.An(ori_ori_n121_), .B(ori_ori_n186_), .Y(ori_ori_n187_));
  NOi31      o171(.An(ori_ori_n187_), .B(ori_ori_n159_), .C(ori_ori_n185_), .Y(ori_ori_n188_));
  NO4        o172(.A(ori_ori_n188_), .B(ori_ori_n184_), .C(ori_ori_n179_), .D(ori_ori_n175_), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n189_), .B(ori_ori_n43_), .Y(ori_ori_n190_));
  NO2        o174(.A(ori_ori_n178_), .B(ori_ori_n76_), .Y(ori_ori_n191_));
  INV        o175(.A(ori_ori_n130_), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n105_), .B(ori_ori_n17_), .Y(ori_ori_n193_));
  AOI210     o177(.A0(ori_ori_n35_), .A1(ori_ori_n90_), .B0(ori_ori_n193_), .Y(ori_ori_n194_));
  NO3        o178(.A(ori_ori_n194_), .B(ori_ori_n192_), .C(x7), .Y(ori_ori_n195_));
  NA3        o179(.A(ori_ori_n187_), .B(ori_ori_n192_), .C(ori_ori_n42_), .Y(ori_ori_n196_));
  OAI210     o180(.A0(ori_ori_n177_), .A1(ori_ori_n137_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  NO3        o181(.A(ori_ori_n197_), .B(ori_ori_n195_), .C(ori_ori_n191_), .Y(ori_ori_n198_));
  NO2        o182(.A(ori_ori_n198_), .B(x3), .Y(ori_ori_n199_));
  NO3        o183(.A(ori_ori_n199_), .B(ori_ori_n190_), .C(ori_ori_n174_), .Y(ori03));
  NO2        o184(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n201_));
  NO2        o185(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n202_));
  INV        o186(.A(ori_ori_n202_), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n204_));
  OAI210     o188(.A0(ori_ori_n204_), .A1(ori_ori_n25_), .B0(ori_ori_n63_), .Y(ori_ori_n205_));
  OAI220     o189(.A0(ori_ori_n205_), .A1(ori_ori_n17_), .B0(ori_ori_n203_), .B1(ori_ori_n105_), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n206_), .B(ori_ori_n201_), .Y(ori_ori_n207_));
  NO2        o191(.A(ori_ori_n78_), .B(x6), .Y(ori_ori_n208_));
  NA2        o192(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n209_));
  NO2        o193(.A(ori_ori_n209_), .B(x4), .Y(ori_ori_n210_));
  NO2        o194(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n211_));
  AN2        o195(.A(ori_ori_n208_), .B(ori_ori_n55_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n212_), .B(ori_ori_n62_), .Y(ori_ori_n213_));
  NA2        o197(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n214_));
  NO2        o198(.A(ori_ori_n214_), .B(ori_ori_n209_), .Y(ori_ori_n215_));
  NA2        o199(.A(x9), .B(ori_ori_n54_), .Y(ori_ori_n216_));
  NA2        o200(.A(ori_ori_n216_), .B(x4), .Y(ori_ori_n217_));
  NA2        o201(.A(ori_ori_n209_), .B(ori_ori_n81_), .Y(ori_ori_n218_));
  AOI210     o202(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n185_), .Y(ori_ori_n219_));
  AOI220     o203(.A0(ori_ori_n219_), .A1(ori_ori_n218_), .B0(ori_ori_n217_), .B1(ori_ori_n215_), .Y(ori_ori_n220_));
  NO3        o204(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n221_));
  NO2        o205(.A(x5), .B(x1), .Y(ori_ori_n222_));
  NO2        o206(.A(ori_ori_n214_), .B(ori_ori_n176_), .Y(ori_ori_n223_));
  NO3        o207(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n224_));
  NO2        o208(.A(ori_ori_n224_), .B(ori_ori_n223_), .Y(ori_ori_n225_));
  INV        o209(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NA2        o210(.A(ori_ori_n226_), .B(ori_ori_n48_), .Y(ori_ori_n227_));
  NA4        o211(.A(ori_ori_n227_), .B(ori_ori_n220_), .C(ori_ori_n213_), .D(ori_ori_n207_), .Y(ori_ori_n228_));
  NO2        o212(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n229_));
  NA2        o213(.A(ori_ori_n229_), .B(ori_ori_n19_), .Y(ori_ori_n230_));
  NO2        o214(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n231_));
  NO2        o215(.A(ori_ori_n231_), .B(x6), .Y(ori_ori_n232_));
  NOi21      o216(.An(ori_ori_n84_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NA2        o217(.A(ori_ori_n62_), .B(ori_ori_n90_), .Y(ori_ori_n234_));
  NA3        o218(.A(ori_ori_n234_), .B(ori_ori_n231_), .C(x6), .Y(ori_ori_n235_));
  AOI210     o219(.A0(ori_ori_n235_), .A1(ori_ori_n233_), .B0(ori_ori_n156_), .Y(ori_ori_n236_));
  AO210      o220(.A0(ori_ori_n236_), .A1(ori_ori_n230_), .B0(ori_ori_n181_), .Y(ori_ori_n237_));
  NA2        o221(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n238_));
  OAI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n25_), .B0(ori_ori_n177_), .Y(ori_ori_n239_));
  NO3        o223(.A(ori_ori_n186_), .B(ori_ori_n62_), .C(x6), .Y(ori_ori_n240_));
  AOI220     o224(.A0(ori_ori_n240_), .A1(ori_ori_n239_), .B0(ori_ori_n142_), .B1(ori_ori_n89_), .Y(ori_ori_n241_));
  NA2        o225(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n242_));
  OAI210     o226(.A0(ori_ori_n118_), .A1(ori_ori_n79_), .B0(x4), .Y(ori_ori_n243_));
  AOI210     o227(.A0(ori_ori_n243_), .A1(ori_ori_n242_), .B0(ori_ori_n78_), .Y(ori_ori_n244_));
  NO2        o228(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n245_));
  NO2        o229(.A(ori_ori_n164_), .B(ori_ori_n43_), .Y(ori_ori_n246_));
  OAI210     o230(.A0(ori_ori_n246_), .A1(ori_ori_n223_), .B0(ori_ori_n245_), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n202_), .B(ori_ori_n135_), .Y(ori_ori_n248_));
  NA3        o232(.A(ori_ori_n214_), .B(ori_ori_n130_), .C(x6), .Y(ori_ori_n249_));
  OAI210     o233(.A0(ori_ori_n90_), .A1(ori_ori_n36_), .B0(ori_ori_n67_), .Y(ori_ori_n250_));
  NA4        o234(.A(ori_ori_n250_), .B(ori_ori_n249_), .C(ori_ori_n248_), .D(ori_ori_n247_), .Y(ori_ori_n251_));
  OAI210     o235(.A0(ori_ori_n251_), .A1(ori_ori_n244_), .B0(x2), .Y(ori_ori_n252_));
  NA3        o236(.A(ori_ori_n252_), .B(ori_ori_n241_), .C(ori_ori_n237_), .Y(ori_ori_n253_));
  AOI210     o237(.A0(ori_ori_n228_), .A1(x8), .B0(ori_ori_n253_), .Y(ori_ori_n254_));
  NO2        o238(.A(ori_ori_n90_), .B(x3), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n255_), .B(ori_ori_n210_), .Y(ori_ori_n256_));
  NO3        o240(.A(ori_ori_n88_), .B(ori_ori_n79_), .C(ori_ori_n25_), .Y(ori_ori_n257_));
  AOI210     o241(.A0(ori_ori_n232_), .A1(ori_ori_n159_), .B0(ori_ori_n257_), .Y(ori_ori_n258_));
  AOI210     o242(.A0(ori_ori_n258_), .A1(ori_ori_n256_), .B0(x2), .Y(ori_ori_n259_));
  NO2        o243(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n260_));
  AOI220     o244(.A0(ori_ori_n210_), .A1(ori_ori_n193_), .B0(ori_ori_n260_), .B1(ori_ori_n67_), .Y(ori_ori_n261_));
  NA2        o245(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n262_));
  NA3        o246(.A(ori_ori_n25_), .B(x3), .C(x2), .Y(ori_ori_n263_));
  AOI210     o247(.A0(ori_ori_n263_), .A1(ori_ori_n141_), .B0(ori_ori_n262_), .Y(ori_ori_n264_));
  NA2        o248(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n265_));
  NO2        o249(.A(ori_ori_n265_), .B(ori_ori_n25_), .Y(ori_ori_n266_));
  OAI210     o250(.A0(ori_ori_n266_), .A1(ori_ori_n264_), .B0(ori_ori_n121_), .Y(ori_ori_n267_));
  NA2        o251(.A(ori_ori_n214_), .B(x6), .Y(ori_ori_n268_));
  NO2        o252(.A(ori_ori_n214_), .B(x6), .Y(ori_ori_n269_));
  NAi21      o253(.An(ori_ori_n167_), .B(ori_ori_n269_), .Y(ori_ori_n270_));
  NA3        o254(.A(ori_ori_n270_), .B(ori_ori_n268_), .C(ori_ori_n147_), .Y(ori_ori_n271_));
  NA4        o255(.A(ori_ori_n271_), .B(ori_ori_n267_), .C(ori_ori_n261_), .D(ori_ori_n156_), .Y(ori_ori_n272_));
  NA2        o256(.A(ori_ori_n202_), .B(ori_ori_n231_), .Y(ori_ori_n273_));
  NO2        o257(.A(x9), .B(x6), .Y(ori_ori_n274_));
  NO2        o258(.A(ori_ori_n141_), .B(ori_ori_n18_), .Y(ori_ori_n275_));
  NAi21      o259(.An(ori_ori_n275_), .B(ori_ori_n263_), .Y(ori_ori_n276_));
  NAi21      o260(.An(x1), .B(x4), .Y(ori_ori_n277_));
  AOI210     o261(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n278_));
  OAI210     o262(.A0(ori_ori_n141_), .A1(x3), .B0(ori_ori_n278_), .Y(ori_ori_n279_));
  AOI220     o263(.A0(ori_ori_n279_), .A1(ori_ori_n277_), .B0(ori_ori_n276_), .B1(ori_ori_n274_), .Y(ori_ori_n280_));
  NA2        o264(.A(ori_ori_n280_), .B(ori_ori_n273_), .Y(ori_ori_n281_));
  NA2        o265(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n282_));
  NO2        o266(.A(ori_ori_n282_), .B(ori_ori_n273_), .Y(ori_ori_n283_));
  NA2        o267(.A(x6), .B(x2), .Y(ori_ori_n284_));
  NO2        o268(.A(ori_ori_n182_), .B(ori_ori_n46_), .Y(ori_ori_n285_));
  OAI210     o269(.A0(ori_ori_n285_), .A1(ori_ori_n283_), .B0(ori_ori_n281_), .Y(ori_ori_n286_));
  NA2        o270(.A(x9), .B(ori_ori_n43_), .Y(ori_ori_n287_));
  NO2        o271(.A(ori_ori_n287_), .B(ori_ori_n209_), .Y(ori_ori_n288_));
  OR3        o272(.A(ori_ori_n288_), .B(ori_ori_n208_), .C(ori_ori_n151_), .Y(ori_ori_n289_));
  NA2        o273(.A(x4), .B(x0), .Y(ori_ori_n290_));
  NA2        o274(.A(ori_ori_n289_), .B(ori_ori_n42_), .Y(ori_ori_n291_));
  AOI210     o275(.A0(ori_ori_n291_), .A1(ori_ori_n286_), .B0(x8), .Y(ori_ori_n292_));
  INV        o276(.A(ori_ori_n262_), .Y(ori_ori_n293_));
  OAI210     o277(.A0(ori_ori_n275_), .A1(ori_ori_n222_), .B0(ori_ori_n293_), .Y(ori_ori_n294_));
  INV        o278(.A(ori_ori_n180_), .Y(ori_ori_n295_));
  OAI210     o279(.A0(ori_ori_n295_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n296_));
  AOI210     o280(.A0(ori_ori_n296_), .A1(ori_ori_n294_), .B0(ori_ori_n238_), .Y(ori_ori_n297_));
  NO4        o281(.A(ori_ori_n297_), .B(ori_ori_n292_), .C(ori_ori_n272_), .D(ori_ori_n259_), .Y(ori_ori_n298_));
  NO2        o282(.A(ori_ori_n167_), .B(x1), .Y(ori_ori_n299_));
  NO3        o283(.A(ori_ori_n299_), .B(x3), .C(ori_ori_n36_), .Y(ori_ori_n300_));
  OAI210     o284(.A0(ori_ori_n300_), .A1(ori_ori_n269_), .B0(x2), .Y(ori_ori_n301_));
  OAI210     o285(.A0(ori_ori_n295_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n302_));
  AOI210     o286(.A0(ori_ori_n302_), .A1(ori_ori_n301_), .B0(ori_ori_n192_), .Y(ori_ori_n303_));
  NOi21      o287(.An(ori_ori_n284_), .B(ori_ori_n17_), .Y(ori_ori_n304_));
  NA3        o288(.A(ori_ori_n304_), .B(ori_ori_n222_), .C(ori_ori_n40_), .Y(ori_ori_n305_));
  AOI210     o289(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n306_));
  NA3        o290(.A(ori_ori_n306_), .B(ori_ori_n165_), .C(ori_ori_n32_), .Y(ori_ori_n307_));
  NA2        o291(.A(x3), .B(x2), .Y(ori_ori_n308_));
  AOI220     o292(.A0(ori_ori_n308_), .A1(ori_ori_n238_), .B0(ori_ori_n307_), .B1(ori_ori_n305_), .Y(ori_ori_n309_));
  NAi21      o293(.An(x4), .B(x0), .Y(ori_ori_n310_));
  NO3        o294(.A(ori_ori_n310_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n311_));
  OAI210     o295(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n311_), .Y(ori_ori_n312_));
  OAI220     o296(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n313_));
  NO2        o297(.A(x9), .B(x8), .Y(ori_ori_n314_));
  NA3        o298(.A(ori_ori_n314_), .B(ori_ori_n36_), .C(ori_ori_n54_), .Y(ori_ori_n315_));
  OAI210     o299(.A0(ori_ori_n306_), .A1(ori_ori_n304_), .B0(ori_ori_n315_), .Y(ori_ori_n316_));
  AOI220     o300(.A0(ori_ori_n316_), .A1(ori_ori_n82_), .B0(ori_ori_n313_), .B1(ori_ori_n31_), .Y(ori_ori_n317_));
  AOI210     o301(.A0(ori_ori_n317_), .A1(ori_ori_n312_), .B0(ori_ori_n25_), .Y(ori_ori_n318_));
  NA3        o302(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n319_));
  OAI210     o303(.A0(ori_ori_n306_), .A1(ori_ori_n304_), .B0(ori_ori_n319_), .Y(ori_ori_n320_));
  INV        o304(.A(ori_ori_n223_), .Y(ori_ori_n321_));
  NA2        o305(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n322_));
  OR2        o306(.A(ori_ori_n322_), .B(ori_ori_n290_), .Y(ori_ori_n323_));
  OAI220     o307(.A0(ori_ori_n323_), .A1(ori_ori_n164_), .B0(ori_ori_n242_), .B1(ori_ori_n321_), .Y(ori_ori_n324_));
  AO210      o308(.A0(ori_ori_n320_), .A1(ori_ori_n151_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  NO4        o309(.A(ori_ori_n325_), .B(ori_ori_n318_), .C(ori_ori_n309_), .D(ori_ori_n303_), .Y(ori_ori_n326_));
  OAI210     o310(.A0(ori_ori_n298_), .A1(ori_ori_n254_), .B0(ori_ori_n326_), .Y(ori04));
  NO2        o311(.A(x2), .B(x1), .Y(ori_ori_n328_));
  OAI210     o312(.A0(ori_ori_n265_), .A1(ori_ori_n328_), .B0(ori_ori_n36_), .Y(ori_ori_n329_));
  NO2        o313(.A(ori_ori_n328_), .B(ori_ori_n310_), .Y(ori_ori_n330_));
  AOI210     o314(.A0(ori_ori_n62_), .A1(x4), .B0(ori_ori_n111_), .Y(ori_ori_n331_));
  OAI210     o315(.A0(ori_ori_n331_), .A1(ori_ori_n330_), .B0(ori_ori_n255_), .Y(ori_ori_n332_));
  NO2        o316(.A(ori_ori_n282_), .B(ori_ori_n88_), .Y(ori_ori_n333_));
  NO2        o317(.A(ori_ori_n333_), .B(ori_ori_n36_), .Y(ori_ori_n334_));
  NO2        o318(.A(ori_ori_n308_), .B(ori_ori_n211_), .Y(ori_ori_n335_));
  NA2        o319(.A(ori_ori_n335_), .B(ori_ori_n90_), .Y(ori_ori_n336_));
  NA3        o320(.A(ori_ori_n336_), .B(ori_ori_n334_), .C(ori_ori_n332_), .Y(ori_ori_n337_));
  NA2        o321(.A(ori_ori_n337_), .B(ori_ori_n329_), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n216_), .B(ori_ori_n112_), .Y(ori_ori_n339_));
  NO3        o323(.A(ori_ori_n262_), .B(ori_ori_n119_), .C(ori_ori_n18_), .Y(ori_ori_n340_));
  NO2        o324(.A(ori_ori_n340_), .B(ori_ori_n339_), .Y(ori_ori_n341_));
  OAI210     o325(.A0(ori_ori_n117_), .A1(ori_ori_n105_), .B0(ori_ori_n180_), .Y(ori_ori_n342_));
  NA3        o326(.A(ori_ori_n342_), .B(x6), .C(x3), .Y(ori_ori_n343_));
  NOi21      o327(.An(ori_ori_n153_), .B(ori_ori_n131_), .Y(ori_ori_n344_));
  AOI210     o328(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n345_));
  OAI220     o329(.A0(ori_ori_n345_), .A1(ori_ori_n322_), .B0(ori_ori_n282_), .B1(ori_ori_n319_), .Y(ori_ori_n346_));
  AOI210     o330(.A0(ori_ori_n344_), .A1(ori_ori_n63_), .B0(ori_ori_n346_), .Y(ori_ori_n347_));
  NA2        o331(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n348_));
  OAI210     o332(.A0(ori_ori_n105_), .A1(ori_ori_n17_), .B0(ori_ori_n348_), .Y(ori_ori_n349_));
  AOI220     o333(.A0(ori_ori_n349_), .A1(ori_ori_n79_), .B0(ori_ori_n333_), .B1(ori_ori_n90_), .Y(ori_ori_n350_));
  NA4        o334(.A(ori_ori_n350_), .B(ori_ori_n347_), .C(ori_ori_n343_), .D(ori_ori_n341_), .Y(ori_ori_n351_));
  OAI210     o335(.A0(ori_ori_n110_), .A1(x3), .B0(ori_ori_n311_), .Y(ori_ori_n352_));
  NA2        o336(.A(ori_ori_n221_), .B(ori_ori_n84_), .Y(ori_ori_n353_));
  NA3        o337(.A(ori_ori_n353_), .B(ori_ori_n352_), .C(ori_ori_n156_), .Y(ori_ori_n354_));
  AOI210     o338(.A0(ori_ori_n351_), .A1(x4), .B0(ori_ori_n354_), .Y(ori_ori_n355_));
  NA3        o339(.A(ori_ori_n330_), .B(ori_ori_n216_), .C(ori_ori_n90_), .Y(ori_ori_n356_));
  NOi21      o340(.An(x4), .B(x0), .Y(ori_ori_n357_));
  XO2        o341(.A(x4), .B(x0), .Y(ori_ori_n358_));
  OAI210     o342(.A0(ori_ori_n358_), .A1(ori_ori_n116_), .B0(ori_ori_n277_), .Y(ori_ori_n359_));
  AOI220     o343(.A0(ori_ori_n359_), .A1(x8), .B0(ori_ori_n357_), .B1(ori_ori_n91_), .Y(ori_ori_n360_));
  AOI210     o344(.A0(ori_ori_n360_), .A1(ori_ori_n356_), .B0(x3), .Y(ori_ori_n361_));
  INV        o345(.A(ori_ori_n91_), .Y(ori_ori_n362_));
  NO2        o346(.A(ori_ori_n90_), .B(x4), .Y(ori_ori_n363_));
  AOI220     o347(.A0(ori_ori_n363_), .A1(ori_ori_n44_), .B0(ori_ori_n125_), .B1(ori_ori_n362_), .Y(ori_ori_n364_));
  NO3        o348(.A(ori_ori_n358_), .B(ori_ori_n167_), .C(x2), .Y(ori_ori_n365_));
  NO3        o349(.A(ori_ori_n234_), .B(ori_ori_n28_), .C(ori_ori_n24_), .Y(ori_ori_n366_));
  NO2        o350(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n367_));
  NA4        o351(.A(ori_ori_n367_), .B(ori_ori_n364_), .C(ori_ori_n230_), .D(x6), .Y(ori_ori_n368_));
  OAI220     o352(.A0(ori_ori_n310_), .A1(ori_ori_n88_), .B0(ori_ori_n185_), .B1(ori_ori_n90_), .Y(ori_ori_n369_));
  NO2        o353(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n370_));
  OR2        o354(.A(ori_ori_n363_), .B(ori_ori_n370_), .Y(ori_ori_n371_));
  NO2        o355(.A(ori_ori_n153_), .B(ori_ori_n105_), .Y(ori_ori_n372_));
  AOI220     o356(.A0(ori_ori_n372_), .A1(ori_ori_n371_), .B0(ori_ori_n369_), .B1(ori_ori_n61_), .Y(ori_ori_n373_));
  NO2        o357(.A(ori_ori_n153_), .B(ori_ori_n81_), .Y(ori_ori_n374_));
  NO2        o358(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n375_));
  NOi21      o359(.An(ori_ori_n121_), .B(ori_ori_n27_), .Y(ori_ori_n376_));
  AOI210     o360(.A0(ori_ori_n375_), .A1(ori_ori_n374_), .B0(ori_ori_n376_), .Y(ori_ori_n377_));
  OAI210     o361(.A0(ori_ori_n373_), .A1(ori_ori_n62_), .B0(ori_ori_n377_), .Y(ori_ori_n378_));
  OAI220     o362(.A0(ori_ori_n378_), .A1(x6), .B0(ori_ori_n368_), .B1(ori_ori_n361_), .Y(ori_ori_n379_));
  OAI210     o363(.A0(ori_ori_n63_), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n380_));
  OAI210     o364(.A0(ori_ori_n380_), .A1(ori_ori_n90_), .B0(ori_ori_n323_), .Y(ori_ori_n381_));
  AOI210     o365(.A0(ori_ori_n381_), .A1(ori_ori_n18_), .B0(ori_ori_n156_), .Y(ori_ori_n382_));
  AO220      o366(.A0(ori_ori_n382_), .A1(ori_ori_n379_), .B0(ori_ori_n355_), .B1(ori_ori_n338_), .Y(ori_ori_n383_));
  NA2        o367(.A(ori_ori_n375_), .B(x6), .Y(ori_ori_n384_));
  AOI210     o368(.A0(x6), .A1(x1), .B0(ori_ori_n155_), .Y(ori_ori_n385_));
  NA2        o369(.A(ori_ori_n363_), .B(x0), .Y(ori_ori_n386_));
  NA2        o370(.A(ori_ori_n84_), .B(x6), .Y(ori_ori_n387_));
  OAI210     o371(.A0(ori_ori_n386_), .A1(ori_ori_n385_), .B0(ori_ori_n387_), .Y(ori_ori_n388_));
  AOI220     o372(.A0(ori_ori_n388_), .A1(ori_ori_n384_), .B0(ori_ori_n224_), .B1(ori_ori_n49_), .Y(ori_ori_n389_));
  NA2        o373(.A(ori_ori_n389_), .B(ori_ori_n383_), .Y(ori_ori_n390_));
  AOI210     o374(.A0(ori_ori_n204_), .A1(x8), .B0(ori_ori_n110_), .Y(ori_ori_n391_));
  NA2        o375(.A(ori_ori_n391_), .B(ori_ori_n348_), .Y(ori_ori_n392_));
  NA3        o376(.A(ori_ori_n392_), .B(ori_ori_n201_), .C(ori_ori_n156_), .Y(ori_ori_n393_));
  OAI210     o377(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n238_), .Y(ori_ori_n394_));
  AO220      o378(.A0(ori_ori_n394_), .A1(ori_ori_n152_), .B0(ori_ori_n109_), .B1(x4), .Y(ori_ori_n395_));
  NA3        o379(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n396_));
  NA2        o380(.A(ori_ori_n229_), .B(x0), .Y(ori_ori_n397_));
  OAI220     o381(.A0(ori_ori_n397_), .A1(ori_ori_n216_), .B0(ori_ori_n396_), .B1(ori_ori_n362_), .Y(ori_ori_n398_));
  AOI210     o382(.A0(ori_ori_n395_), .A1(ori_ori_n118_), .B0(ori_ori_n398_), .Y(ori_ori_n399_));
  AOI210     o383(.A0(ori_ori_n399_), .A1(ori_ori_n393_), .B0(ori_ori_n25_), .Y(ori_ori_n400_));
  NA3        o384(.A(ori_ori_n120_), .B(ori_ori_n229_), .C(x0), .Y(ori_ori_n401_));
  OAI210     o385(.A0(ori_ori_n201_), .A1(ori_ori_n68_), .B0(ori_ori_n211_), .Y(ori_ori_n402_));
  NA3        o386(.A(ori_ori_n204_), .B(ori_ori_n231_), .C(x8), .Y(ori_ori_n403_));
  AOI210     o387(.A0(ori_ori_n403_), .A1(ori_ori_n402_), .B0(ori_ori_n25_), .Y(ori_ori_n404_));
  AOI210     o388(.A0(ori_ori_n119_), .A1(ori_ori_n117_), .B0(ori_ori_n42_), .Y(ori_ori_n405_));
  NOi31      o389(.An(ori_ori_n405_), .B(ori_ori_n370_), .C(ori_ori_n186_), .Y(ori_ori_n406_));
  OAI210     o390(.A0(ori_ori_n406_), .A1(ori_ori_n404_), .B0(ori_ori_n152_), .Y(ori_ori_n407_));
  NAi31      o391(.An(ori_ori_n50_), .B(ori_ori_n299_), .C(ori_ori_n181_), .Y(ori_ori_n408_));
  NA3        o392(.A(ori_ori_n408_), .B(ori_ori_n407_), .C(ori_ori_n401_), .Y(ori_ori_n409_));
  OAI210     o393(.A0(ori_ori_n409_), .A1(ori_ori_n400_), .B0(x6), .Y(ori_ori_n410_));
  OAI210     o394(.A0(ori_ori_n167_), .A1(ori_ori_n48_), .B0(ori_ori_n136_), .Y(ori_ori_n411_));
  NA3        o395(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n412_));
  AOI220     o396(.A0(ori_ori_n412_), .A1(ori_ori_n411_), .B0(ori_ori_n40_), .B1(ori_ori_n32_), .Y(ori_ori_n413_));
  NO2        o397(.A(ori_ori_n156_), .B(x0), .Y(ori_ori_n414_));
  AOI220     o398(.A0(ori_ori_n414_), .A1(ori_ori_n229_), .B0(ori_ori_n201_), .B1(ori_ori_n156_), .Y(ori_ori_n415_));
  AOI210     o399(.A0(ori_ori_n127_), .A1(ori_ori_n260_), .B0(x1), .Y(ori_ori_n416_));
  OAI210     o400(.A0(ori_ori_n415_), .A1(x8), .B0(ori_ori_n416_), .Y(ori_ori_n417_));
  NAi31      o401(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n418_));
  OAI210     o402(.A0(ori_ori_n418_), .A1(x4), .B0(ori_ori_n168_), .Y(ori_ori_n419_));
  NA3        o403(.A(ori_ori_n419_), .B(ori_ori_n150_), .C(x9), .Y(ori_ori_n420_));
  NO4        o404(.A(ori_ori_n126_), .B(ori_ori_n310_), .C(x9), .D(x2), .Y(ori_ori_n421_));
  NOi21      o405(.An(ori_ori_n124_), .B(ori_ori_n185_), .Y(ori_ori_n422_));
  NO3        o406(.A(ori_ori_n422_), .B(ori_ori_n421_), .C(ori_ori_n18_), .Y(ori_ori_n423_));
  NO3        o407(.A(x9), .B(ori_ori_n156_), .C(x0), .Y(ori_ori_n424_));
  AOI220     o408(.A0(ori_ori_n424_), .A1(ori_ori_n255_), .B0(ori_ori_n374_), .B1(ori_ori_n156_), .Y(ori_ori_n425_));
  NA4        o409(.A(ori_ori_n425_), .B(ori_ori_n423_), .C(ori_ori_n420_), .D(ori_ori_n50_), .Y(ori_ori_n426_));
  OAI210     o410(.A0(ori_ori_n417_), .A1(ori_ori_n413_), .B0(ori_ori_n426_), .Y(ori_ori_n427_));
  NOi31      o411(.An(ori_ori_n414_), .B(ori_ori_n32_), .C(x8), .Y(ori_ori_n428_));
  AOI210     o412(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n134_), .Y(ori_ori_n429_));
  NO3        o413(.A(ori_ori_n429_), .B(ori_ori_n124_), .C(ori_ori_n43_), .Y(ori_ori_n430_));
  NOi31      o414(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n431_));
  AOI220     o415(.A0(ori_ori_n431_), .A1(ori_ori_n357_), .B0(ori_ori_n125_), .B1(x3), .Y(ori_ori_n432_));
  AOI210     o416(.A0(ori_ori_n277_), .A1(ori_ori_n60_), .B0(ori_ori_n123_), .Y(ori_ori_n433_));
  OAI210     o417(.A0(ori_ori_n433_), .A1(x3), .B0(ori_ori_n432_), .Y(ori_ori_n434_));
  NO3        o418(.A(ori_ori_n434_), .B(ori_ori_n430_), .C(x2), .Y(ori_ori_n435_));
  OAI220     o419(.A0(ori_ori_n358_), .A1(ori_ori_n314_), .B0(ori_ori_n310_), .B1(ori_ori_n43_), .Y(ori_ori_n436_));
  AOI210     o420(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n396_), .Y(ori_ori_n437_));
  AOI220     o421(.A0(ori_ori_n437_), .A1(ori_ori_n90_), .B0(ori_ori_n436_), .B1(ori_ori_n156_), .Y(ori_ori_n438_));
  NO2        o422(.A(ori_ori_n438_), .B(ori_ori_n54_), .Y(ori_ori_n439_));
  NO3        o423(.A(ori_ori_n439_), .B(ori_ori_n435_), .C(ori_ori_n428_), .Y(ori_ori_n440_));
  AOI210     o424(.A0(ori_ori_n440_), .A1(ori_ori_n427_), .B0(ori_ori_n25_), .Y(ori_ori_n441_));
  NA4        o425(.A(ori_ori_n31_), .B(ori_ori_n90_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n442_));
  NO3        o426(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n443_));
  NO3        o427(.A(ori_ori_n68_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n444_));
  AOI220     o428(.A0(ori_ori_n444_), .A1(ori_ori_n278_), .B0(ori_ori_n443_), .B1(ori_ori_n405_), .Y(ori_ori_n445_));
  NO2        o429(.A(ori_ori_n445_), .B(ori_ori_n102_), .Y(ori_ori_n446_));
  NO3        o430(.A(ori_ori_n282_), .B(ori_ori_n180_), .C(ori_ori_n40_), .Y(ori_ori_n447_));
  OAI210     o431(.A0(ori_ori_n447_), .A1(ori_ori_n446_), .B0(x7), .Y(ori_ori_n448_));
  NA2        o432(.A(ori_ori_n234_), .B(x7), .Y(ori_ori_n449_));
  NA3        o433(.A(ori_ori_n449_), .B(ori_ori_n155_), .C(ori_ori_n135_), .Y(ori_ori_n450_));
  NA3        o434(.A(ori_ori_n450_), .B(ori_ori_n448_), .C(ori_ori_n442_), .Y(ori_ori_n451_));
  OAI210     o435(.A0(ori_ori_n451_), .A1(ori_ori_n441_), .B0(ori_ori_n36_), .Y(ori_ori_n452_));
  NO2        o436(.A(ori_ori_n424_), .B(ori_ori_n211_), .Y(ori_ori_n453_));
  NO4        o437(.A(ori_ori_n453_), .B(ori_ori_n78_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n454_));
  NA2        o438(.A(ori_ori_n265_), .B(ori_ori_n21_), .Y(ori_ori_n455_));
  NO2        o439(.A(ori_ori_n164_), .B(ori_ori_n136_), .Y(ori_ori_n456_));
  NA2        o440(.A(ori_ori_n456_), .B(ori_ori_n455_), .Y(ori_ori_n457_));
  AOI210     o441(.A0(ori_ori_n457_), .A1(ori_ori_n171_), .B0(ori_ori_n28_), .Y(ori_ori_n458_));
  AOI220     o442(.A0(ori_ori_n370_), .A1(ori_ori_n90_), .B0(ori_ori_n153_), .B1(ori_ori_n204_), .Y(ori_ori_n459_));
  NA3        o443(.A(ori_ori_n459_), .B(ori_ori_n418_), .C(ori_ori_n88_), .Y(ori_ori_n460_));
  NA2        o444(.A(ori_ori_n460_), .B(ori_ori_n181_), .Y(ori_ori_n461_));
  OAI220     o445(.A0(ori_ori_n287_), .A1(ori_ori_n69_), .B0(ori_ori_n164_), .B1(ori_ori_n43_), .Y(ori_ori_n462_));
  NA2        o446(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n463_));
  OAI210     o447(.A0(ori_ori_n152_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n464_));
  NO3        o448(.A(ori_ori_n431_), .B(x3), .C(ori_ori_n54_), .Y(ori_ori_n465_));
  NA2        o449(.A(ori_ori_n465_), .B(ori_ori_n464_), .Y(ori_ori_n466_));
  OAI210     o450(.A0(ori_ori_n157_), .A1(ori_ori_n463_), .B0(ori_ori_n466_), .Y(ori_ori_n467_));
  AOI220     o451(.A0(ori_ori_n467_), .A1(x0), .B0(ori_ori_n462_), .B1(ori_ori_n136_), .Y(ori_ori_n468_));
  AOI210     o452(.A0(ori_ori_n468_), .A1(ori_ori_n461_), .B0(ori_ori_n242_), .Y(ori_ori_n469_));
  NO3        o453(.A(ori_ori_n469_), .B(ori_ori_n458_), .C(ori_ori_n454_), .Y(ori_ori_n470_));
  NA3        o454(.A(ori_ori_n470_), .B(ori_ori_n452_), .C(ori_ori_n410_), .Y(ori_ori_n471_));
  AOI210     o455(.A0(ori_ori_n390_), .A1(ori_ori_n25_), .B0(ori_ori_n471_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  INV        m047(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  NO2        m048(.A(x7), .B(x6), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(x8), .B(x2), .Y(mai_mai_n67_));
  INV        m051(.A(mai_mai_n67_), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n68_), .B(x1), .Y(mai_mai_n69_));
  OA210      m053(.A0(mai_mai_n69_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  NAi31      m056(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n73_));
  OAI220     m057(.A0(mai_mai_n73_), .A1(mai_mai_n43_), .B0(mai_mai_n72_), .B1(mai_mai_n70_), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n74_), .B(x4), .Y(mai_mai_n75_));
  NA2        m059(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n76_));
  OAI210     m060(.A0(mai_mai_n76_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n77_));
  NA2        m061(.A(x5), .B(x3), .Y(mai_mai_n78_));
  NO2        m062(.A(x8), .B(x6), .Y(mai_mai_n79_));
  NO4        m063(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(mai_mai_n65_), .D(mai_mai_n54_), .Y(mai_mai_n80_));
  NAi21      m064(.An(x4), .B(x3), .Y(mai_mai_n81_));
  INV        m065(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(mai_mai_n22_), .Y(mai_mai_n83_));
  NO2        m067(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(x3), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n83_), .C(mai_mai_n18_), .Y(mai_mai_n86_));
  NO3        m070(.A(mai_mai_n86_), .B(mai_mai_n80_), .C(mai_mai_n77_), .Y(mai_mai_n87_));
  NO4        m071(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n43_), .D(x1), .Y(mai_mai_n88_));
  NA2        m072(.A(mai_mai_n62_), .B(mai_mai_n48_), .Y(mai_mai_n89_));
  INV        m073(.A(mai_mai_n89_), .Y(mai_mai_n90_));
  NA2        m074(.A(mai_mai_n88_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  NA2        m075(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n25_), .Y(mai_mai_n93_));
  INV        m077(.A(x8), .Y(mai_mai_n94_));
  NA2        m078(.A(x2), .B(x1), .Y(mai_mai_n95_));
  INV        m079(.A(mai_mai_n93_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n96_), .B(mai_mai_n26_), .Y(mai_mai_n97_));
  AOI210     m081(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n98_));
  OAI210     m082(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n99_));
  NO3        m083(.A(mai_mai_n99_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n100_));
  NA2        m084(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n101_));
  NO2        m085(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n102_));
  OAI210     m086(.A0(mai_mai_n102_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n103_));
  AOI210     m087(.A0(mai_mai_n101_), .A1(mai_mai_n52_), .B0(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m088(.A(x3), .B(x2), .Y(mai_mai_n105_));
  NA3        m089(.A(mai_mai_n105_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n106_));
  AOI210     m090(.A0(x8), .A1(x6), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  NA2        m091(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n108_));
  OAI210     m092(.A0(mai_mai_n108_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n109_));
  NO4        m093(.A(mai_mai_n109_), .B(mai_mai_n107_), .C(mai_mai_n104_), .D(mai_mai_n100_), .Y(mai_mai_n110_));
  AO220      m094(.A0(mai_mai_n110_), .A1(mai_mai_n91_), .B0(mai_mai_n87_), .B1(mai_mai_n75_), .Y(mai02));
  NO2        m095(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n112_));
  NO2        m096(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n113_));
  NA2        m097(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n114_));
  NA2        m098(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n115_));
  OAI210     m099(.A0(mai_mai_n89_), .A1(mai_mai_n114_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  AOI220     m100(.A0(mai_mai_n116_), .A1(mai_mai_n113_), .B0(mai_mai_n112_), .B1(x4), .Y(mai_mai_n117_));
  NO3        m101(.A(mai_mai_n117_), .B(x7), .C(x5), .Y(mai_mai_n118_));
  NA2        m102(.A(x9), .B(x2), .Y(mai_mai_n119_));
  OR2        m103(.A(x8), .B(x0), .Y(mai_mai_n120_));
  INV        m104(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NAi21      m105(.An(x2), .B(x8), .Y(mai_mai_n122_));
  INV        m106(.A(mai_mai_n122_), .Y(mai_mai_n123_));
  OAI220     m107(.A0(mai_mai_n123_), .A1(mai_mai_n121_), .B0(mai_mai_n119_), .B1(x7), .Y(mai_mai_n124_));
  NO2        m108(.A(x4), .B(x1), .Y(mai_mai_n125_));
  NA3        m109(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(mai_mai_n60_), .Y(mai_mai_n126_));
  NOi21      m110(.An(x0), .B(x1), .Y(mai_mai_n127_));
  NO3        m111(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n128_));
  NOi21      m112(.An(x0), .B(x4), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n126_), .B(mai_mai_n78_), .Y(mai_mai_n130_));
  NO2        m114(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n131_));
  NA2        m115(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n132_));
  AOI210     m116(.A0(mai_mai_n132_), .A1(mai_mai_n108_), .B0(mai_mai_n115_), .Y(mai_mai_n133_));
  OAI210     m117(.A0(mai_mai_n133_), .A1(mai_mai_n35_), .B0(mai_mai_n131_), .Y(mai_mai_n134_));
  NAi21      m118(.An(x0), .B(x4), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n135_), .B(x1), .Y(mai_mai_n136_));
  NO2        m120(.A(x7), .B(x0), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n84_), .B(mai_mai_n102_), .Y(mai_mai_n138_));
  NO2        m122(.A(mai_mai_n138_), .B(x3), .Y(mai_mai_n139_));
  OAI210     m123(.A0(mai_mai_n137_), .A1(mai_mai_n136_), .B0(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n141_));
  NA2        m125(.A(x5), .B(x0), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n143_));
  NA3        m127(.A(mai_mai_n143_), .B(mai_mai_n142_), .C(mai_mai_n141_), .Y(mai_mai_n144_));
  NA4        m128(.A(mai_mai_n144_), .B(mai_mai_n140_), .C(mai_mai_n134_), .D(mai_mai_n36_), .Y(mai_mai_n145_));
  NO3        m129(.A(mai_mai_n145_), .B(mai_mai_n130_), .C(mai_mai_n118_), .Y(mai_mai_n146_));
  NO3        m130(.A(mai_mai_n78_), .B(mai_mai_n76_), .C(mai_mai_n24_), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n148_));
  NA2        m132(.A(x7), .B(x3), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n101_), .B(x5), .Y(mai_mai_n150_));
  NO2        m134(.A(x9), .B(x7), .Y(mai_mai_n151_));
  NOi21      m135(.An(x8), .B(x0), .Y(mai_mai_n152_));
  OA210      m136(.A0(mai_mai_n151_), .A1(x1), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n154_));
  INV        m138(.A(x7), .Y(mai_mai_n155_));
  NA2        m139(.A(mai_mai_n155_), .B(mai_mai_n18_), .Y(mai_mai_n156_));
  AOI220     m140(.A0(mai_mai_n156_), .A1(mai_mai_n154_), .B0(mai_mai_n112_), .B1(mai_mai_n38_), .Y(mai_mai_n157_));
  NO2        m141(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n158_));
  NO2        m142(.A(mai_mai_n158_), .B(mai_mai_n129_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n159_), .B(mai_mai_n157_), .Y(mai_mai_n160_));
  AOI210     m144(.A0(mai_mai_n153_), .A1(mai_mai_n150_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  OAI210     m145(.A0(mai_mai_n149_), .A1(mai_mai_n50_), .B0(mai_mai_n161_), .Y(mai_mai_n162_));
  NA2        m146(.A(x5), .B(x1), .Y(mai_mai_n163_));
  INV        m147(.A(mai_mai_n163_), .Y(mai_mai_n164_));
  AOI210     m148(.A0(mai_mai_n164_), .A1(mai_mai_n129_), .B0(mai_mai_n36_), .Y(mai_mai_n165_));
  NO2        m149(.A(mai_mai_n62_), .B(mai_mai_n94_), .Y(mai_mai_n166_));
  NAi21      m150(.An(x2), .B(x7), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n167_), .B(mai_mai_n48_), .Y(mai_mai_n168_));
  NA2        m152(.A(mai_mai_n168_), .B(mai_mai_n66_), .Y(mai_mai_n169_));
  NAi31      m153(.An(mai_mai_n78_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n170_));
  NA3        m154(.A(mai_mai_n170_), .B(mai_mai_n169_), .C(mai_mai_n165_), .Y(mai_mai_n171_));
  NO3        m155(.A(mai_mai_n171_), .B(mai_mai_n162_), .C(mai_mai_n147_), .Y(mai_mai_n172_));
  NO2        m156(.A(mai_mai_n172_), .B(mai_mai_n146_), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n142_), .B(mai_mai_n138_), .Y(mai_mai_n174_));
  NA2        m158(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n175_));
  NA2        m159(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n176_));
  NA3        m160(.A(mai_mai_n176_), .B(mai_mai_n175_), .C(mai_mai_n24_), .Y(mai_mai_n177_));
  AN2        m161(.A(mai_mai_n177_), .B(mai_mai_n143_), .Y(mai_mai_n178_));
  NA2        m162(.A(x8), .B(x0), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n155_), .B(mai_mai_n25_), .Y(mai_mai_n180_));
  NO2        m164(.A(mai_mai_n127_), .B(x4), .Y(mai_mai_n181_));
  NA2        m165(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  AOI210     m166(.A0(mai_mai_n179_), .A1(mai_mai_n132_), .B0(mai_mai_n182_), .Y(mai_mai_n183_));
  NA2        m167(.A(x2), .B(x0), .Y(mai_mai_n184_));
  NA2        m168(.A(x4), .B(x1), .Y(mai_mai_n185_));
  NAi21      m169(.An(mai_mai_n125_), .B(mai_mai_n185_), .Y(mai_mai_n186_));
  NOi31      m170(.An(mai_mai_n186_), .B(mai_mai_n158_), .C(mai_mai_n184_), .Y(mai_mai_n187_));
  NO4        m171(.A(mai_mai_n187_), .B(mai_mai_n183_), .C(mai_mai_n178_), .D(mai_mai_n174_), .Y(mai_mai_n188_));
  NO2        m172(.A(mai_mai_n188_), .B(mai_mai_n43_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n177_), .B(mai_mai_n76_), .Y(mai_mai_n190_));
  INV        m174(.A(mai_mai_n131_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n108_), .B(mai_mai_n17_), .Y(mai_mai_n192_));
  AOI210     m176(.A0(mai_mai_n35_), .A1(mai_mai_n94_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  NO3        m177(.A(mai_mai_n193_), .B(mai_mai_n191_), .C(x7), .Y(mai_mai_n194_));
  NA3        m178(.A(mai_mai_n186_), .B(mai_mai_n191_), .C(mai_mai_n42_), .Y(mai_mai_n195_));
  OAI210     m179(.A0(mai_mai_n176_), .A1(mai_mai_n138_), .B0(mai_mai_n195_), .Y(mai_mai_n196_));
  NO3        m180(.A(mai_mai_n196_), .B(mai_mai_n194_), .C(mai_mai_n190_), .Y(mai_mai_n197_));
  NO2        m181(.A(mai_mai_n197_), .B(x3), .Y(mai_mai_n198_));
  NO3        m182(.A(mai_mai_n198_), .B(mai_mai_n189_), .C(mai_mai_n173_), .Y(mai03));
  NO2        m183(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n200_));
  NO2        m184(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n78_), .B(x6), .Y(mai_mai_n203_));
  NA2        m187(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n204_));
  NO2        m188(.A(mai_mai_n204_), .B(x4), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n206_));
  AO220      m190(.A0(mai_mai_n206_), .A1(mai_mai_n205_), .B0(mai_mai_n203_), .B1(mai_mai_n55_), .Y(mai_mai_n207_));
  INV        m191(.A(mai_mai_n207_), .Y(mai_mai_n208_));
  NA2        m192(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n209_));
  NA2        m193(.A(x9), .B(mai_mai_n54_), .Y(mai_mai_n210_));
  NA2        m194(.A(mai_mai_n204_), .B(mai_mai_n81_), .Y(mai_mai_n211_));
  AOI210     m195(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n184_), .Y(mai_mai_n212_));
  NA2        m196(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n213_));
  NO3        m197(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n214_));
  NO2        m198(.A(x5), .B(x1), .Y(mai_mai_n215_));
  AOI220     m199(.A0(mai_mai_n215_), .A1(mai_mai_n17_), .B0(mai_mai_n105_), .B1(x5), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n209_), .B(mai_mai_n175_), .Y(mai_mai_n217_));
  NO3        m201(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n218_));
  NO2        m202(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n219_));
  OAI210     m203(.A0(mai_mai_n216_), .A1(mai_mai_n64_), .B0(mai_mai_n219_), .Y(mai_mai_n220_));
  AOI220     m204(.A0(mai_mai_n220_), .A1(mai_mai_n48_), .B0(mai_mai_n214_), .B1(mai_mai_n131_), .Y(mai_mai_n221_));
  NA3        m205(.A(mai_mai_n221_), .B(mai_mai_n213_), .C(mai_mai_n208_), .Y(mai_mai_n222_));
  NO2        m206(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n223_), .B(mai_mai_n19_), .Y(mai_mai_n224_));
  NO2        m208(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n225_));
  NO2        m209(.A(mai_mai_n225_), .B(x6), .Y(mai_mai_n226_));
  NOi21      m210(.An(mai_mai_n84_), .B(mai_mai_n226_), .Y(mai_mai_n227_));
  NA2        m211(.A(mai_mai_n62_), .B(mai_mai_n94_), .Y(mai_mai_n228_));
  NA3        m212(.A(mai_mai_n228_), .B(mai_mai_n225_), .C(x6), .Y(mai_mai_n229_));
  AOI210     m213(.A0(mai_mai_n229_), .A1(mai_mai_n227_), .B0(mai_mai_n155_), .Y(mai_mai_n230_));
  AO210      m214(.A0(mai_mai_n230_), .A1(mai_mai_n224_), .B0(mai_mai_n180_), .Y(mai_mai_n231_));
  NA2        m215(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n232_));
  OAI210     m216(.A0(mai_mai_n232_), .A1(mai_mai_n25_), .B0(mai_mai_n176_), .Y(mai_mai_n233_));
  NO3        m217(.A(mai_mai_n185_), .B(mai_mai_n62_), .C(x6), .Y(mai_mai_n234_));
  AOI220     m218(.A0(mai_mai_n234_), .A1(mai_mai_n233_), .B0(mai_mai_n143_), .B1(mai_mai_n93_), .Y(mai_mai_n235_));
  NA2        m219(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n236_));
  OAI210     m220(.A0(mai_mai_n121_), .A1(mai_mai_n79_), .B0(x4), .Y(mai_mai_n237_));
  AOI210     m221(.A0(mai_mai_n237_), .A1(mai_mai_n236_), .B0(mai_mai_n78_), .Y(mai_mai_n238_));
  NA2        m222(.A(mai_mai_n201_), .B(mai_mai_n136_), .Y(mai_mai_n239_));
  NA3        m223(.A(mai_mai_n209_), .B(mai_mai_n131_), .C(x6), .Y(mai_mai_n240_));
  OAI210     m224(.A0(mai_mai_n94_), .A1(mai_mai_n36_), .B0(mai_mai_n66_), .Y(mai_mai_n241_));
  NA3        m225(.A(mai_mai_n241_), .B(mai_mai_n240_), .C(mai_mai_n239_), .Y(mai_mai_n242_));
  OAI210     m226(.A0(mai_mai_n242_), .A1(mai_mai_n238_), .B0(x2), .Y(mai_mai_n243_));
  NA3        m227(.A(mai_mai_n243_), .B(mai_mai_n235_), .C(mai_mai_n231_), .Y(mai_mai_n244_));
  AOI210     m228(.A0(mai_mai_n222_), .A1(x8), .B0(mai_mai_n244_), .Y(mai_mai_n245_));
  NO2        m229(.A(mai_mai_n94_), .B(x3), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n246_), .B(mai_mai_n205_), .Y(mai_mai_n247_));
  NO3        m231(.A(mai_mai_n92_), .B(mai_mai_n79_), .C(mai_mai_n25_), .Y(mai_mai_n248_));
  AOI210     m232(.A0(mai_mai_n226_), .A1(mai_mai_n158_), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  AOI210     m233(.A0(mai_mai_n249_), .A1(mai_mai_n247_), .B0(x2), .Y(mai_mai_n250_));
  NO2        m234(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n251_));
  AOI220     m235(.A0(mai_mai_n205_), .A1(mai_mai_n192_), .B0(mai_mai_n251_), .B1(mai_mai_n66_), .Y(mai_mai_n252_));
  NA2        m236(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n253_));
  NA3        m237(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n254_));
  AOI210     m238(.A0(mai_mai_n254_), .A1(mai_mai_n142_), .B0(mai_mai_n253_), .Y(mai_mai_n255_));
  NA2        m239(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n256_));
  NO2        m240(.A(mai_mai_n256_), .B(mai_mai_n25_), .Y(mai_mai_n257_));
  OAI210     m241(.A0(mai_mai_n257_), .A1(mai_mai_n255_), .B0(mai_mai_n125_), .Y(mai_mai_n258_));
  NA2        m242(.A(mai_mai_n209_), .B(x6), .Y(mai_mai_n259_));
  NO2        m243(.A(mai_mai_n209_), .B(x6), .Y(mai_mai_n260_));
  NAi21      m244(.An(mai_mai_n166_), .B(mai_mai_n260_), .Y(mai_mai_n261_));
  NA3        m245(.A(mai_mai_n261_), .B(mai_mai_n259_), .C(mai_mai_n148_), .Y(mai_mai_n262_));
  NA4        m246(.A(mai_mai_n262_), .B(mai_mai_n258_), .C(mai_mai_n252_), .D(mai_mai_n155_), .Y(mai_mai_n263_));
  NA2        m247(.A(mai_mai_n201_), .B(mai_mai_n225_), .Y(mai_mai_n264_));
  NO2        m248(.A(x9), .B(x6), .Y(mai_mai_n265_));
  NO2        m249(.A(mai_mai_n142_), .B(mai_mai_n18_), .Y(mai_mai_n266_));
  NAi21      m250(.An(mai_mai_n266_), .B(mai_mai_n254_), .Y(mai_mai_n267_));
  NAi21      m251(.An(x1), .B(x4), .Y(mai_mai_n268_));
  AOI210     m252(.A0(x3), .A1(x2), .B0(mai_mai_n48_), .Y(mai_mai_n269_));
  OAI210     m253(.A0(mai_mai_n142_), .A1(x3), .B0(mai_mai_n269_), .Y(mai_mai_n270_));
  AOI220     m254(.A0(mai_mai_n270_), .A1(mai_mai_n268_), .B0(mai_mai_n267_), .B1(mai_mai_n265_), .Y(mai_mai_n271_));
  NA2        m255(.A(mai_mai_n271_), .B(mai_mai_n264_), .Y(mai_mai_n272_));
  NA2        m256(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n273_));
  NO3        m257(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n274_));
  NA2        m258(.A(mai_mai_n108_), .B(mai_mai_n25_), .Y(mai_mai_n275_));
  NA2        m259(.A(x6), .B(x2), .Y(mai_mai_n276_));
  NO2        m260(.A(mai_mai_n276_), .B(mai_mai_n175_), .Y(mai_mai_n277_));
  AOI210     m261(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  OAI220     m262(.A0(mai_mai_n278_), .A1(mai_mai_n43_), .B0(mai_mai_n181_), .B1(mai_mai_n46_), .Y(mai_mai_n279_));
  NA2        m263(.A(mai_mai_n279_), .B(mai_mai_n272_), .Y(mai_mai_n280_));
  NA2        m264(.A(x9), .B(mai_mai_n43_), .Y(mai_mai_n281_));
  NO2        m265(.A(mai_mai_n281_), .B(mai_mai_n204_), .Y(mai_mai_n282_));
  OR3        m266(.A(mai_mai_n282_), .B(mai_mai_n203_), .C(mai_mai_n150_), .Y(mai_mai_n283_));
  NA2        m267(.A(x4), .B(x0), .Y(mai_mai_n284_));
  NO3        m268(.A(mai_mai_n73_), .B(mai_mai_n284_), .C(x6), .Y(mai_mai_n285_));
  AOI210     m269(.A0(mai_mai_n283_), .A1(mai_mai_n42_), .B0(mai_mai_n285_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n286_), .A1(mai_mai_n280_), .B0(x8), .Y(mai_mai_n287_));
  INV        m271(.A(mai_mai_n253_), .Y(mai_mai_n288_));
  OAI210     m272(.A0(mai_mai_n266_), .A1(mai_mai_n215_), .B0(mai_mai_n288_), .Y(mai_mai_n289_));
  INV        m273(.A(mai_mai_n179_), .Y(mai_mai_n290_));
  OAI210     m274(.A0(mai_mai_n290_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n291_));
  AOI210     m275(.A0(mai_mai_n291_), .A1(mai_mai_n289_), .B0(mai_mai_n232_), .Y(mai_mai_n292_));
  NO4        m276(.A(mai_mai_n292_), .B(mai_mai_n287_), .C(mai_mai_n263_), .D(mai_mai_n250_), .Y(mai_mai_n293_));
  NO2        m277(.A(mai_mai_n166_), .B(x1), .Y(mai_mai_n294_));
  NO3        m278(.A(mai_mai_n294_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n295_));
  OAI210     m279(.A0(mai_mai_n295_), .A1(mai_mai_n260_), .B0(x2), .Y(mai_mai_n296_));
  OAI210     m280(.A0(mai_mai_n290_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n297_), .A1(mai_mai_n296_), .B0(mai_mai_n191_), .Y(mai_mai_n298_));
  NOi21      m282(.An(mai_mai_n276_), .B(mai_mai_n17_), .Y(mai_mai_n299_));
  NA3        m283(.A(mai_mai_n299_), .B(mai_mai_n215_), .C(mai_mai_n40_), .Y(mai_mai_n300_));
  AOI210     m284(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n301_));
  NA3        m285(.A(mai_mai_n301_), .B(mai_mai_n164_), .C(mai_mai_n32_), .Y(mai_mai_n302_));
  NA2        m286(.A(x3), .B(x2), .Y(mai_mai_n303_));
  AOI220     m287(.A0(mai_mai_n303_), .A1(mai_mai_n232_), .B0(mai_mai_n302_), .B1(mai_mai_n300_), .Y(mai_mai_n304_));
  NAi21      m288(.An(x4), .B(x0), .Y(mai_mai_n305_));
  NO3        m289(.A(mai_mai_n305_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n306_));
  OAI210     m290(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  OAI220     m291(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n308_));
  NO2        m292(.A(x9), .B(x8), .Y(mai_mai_n309_));
  NO2        m293(.A(mai_mai_n301_), .B(mai_mai_n299_), .Y(mai_mai_n310_));
  AOI220     m294(.A0(mai_mai_n310_), .A1(mai_mai_n82_), .B0(mai_mai_n308_), .B1(mai_mai_n31_), .Y(mai_mai_n311_));
  AOI210     m295(.A0(mai_mai_n311_), .A1(mai_mai_n307_), .B0(mai_mai_n25_), .Y(mai_mai_n312_));
  NA3        m296(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n313_));
  OAI210     m297(.A0(mai_mai_n301_), .A1(mai_mai_n299_), .B0(mai_mai_n313_), .Y(mai_mai_n314_));
  INV        m298(.A(mai_mai_n217_), .Y(mai_mai_n315_));
  NA2        m299(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n316_));
  OR2        m300(.A(mai_mai_n316_), .B(mai_mai_n284_), .Y(mai_mai_n317_));
  OAI220     m301(.A0(mai_mai_n317_), .A1(mai_mai_n163_), .B0(mai_mai_n236_), .B1(mai_mai_n315_), .Y(mai_mai_n318_));
  AO210      m302(.A0(mai_mai_n314_), .A1(mai_mai_n150_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  NO4        m303(.A(mai_mai_n319_), .B(mai_mai_n312_), .C(mai_mai_n304_), .D(mai_mai_n298_), .Y(mai_mai_n320_));
  OAI210     m304(.A0(mai_mai_n293_), .A1(mai_mai_n245_), .B0(mai_mai_n320_), .Y(mai04));
  OAI210     m305(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n322_));
  NA3        m306(.A(mai_mai_n322_), .B(mai_mai_n274_), .C(mai_mai_n85_), .Y(mai_mai_n323_));
  NO2        m307(.A(x2), .B(x1), .Y(mai_mai_n324_));
  OAI210     m308(.A0(mai_mai_n256_), .A1(mai_mai_n324_), .B0(mai_mai_n36_), .Y(mai_mai_n325_));
  NO2        m309(.A(mai_mai_n324_), .B(mai_mai_n305_), .Y(mai_mai_n326_));
  AOI210     m310(.A0(mai_mai_n62_), .A1(x4), .B0(mai_mai_n114_), .Y(mai_mai_n327_));
  OAI210     m311(.A0(mai_mai_n327_), .A1(mai_mai_n326_), .B0(mai_mai_n246_), .Y(mai_mai_n328_));
  NO2        m312(.A(mai_mai_n273_), .B(mai_mai_n92_), .Y(mai_mai_n329_));
  NO2        m313(.A(mai_mai_n329_), .B(mai_mai_n36_), .Y(mai_mai_n330_));
  NO2        m314(.A(mai_mai_n303_), .B(mai_mai_n206_), .Y(mai_mai_n331_));
  NA2        m315(.A(x9), .B(x0), .Y(mai_mai_n332_));
  AOI210     m316(.A0(mai_mai_n92_), .A1(mai_mai_n76_), .B0(mai_mai_n332_), .Y(mai_mai_n333_));
  OAI210     m317(.A0(mai_mai_n333_), .A1(mai_mai_n331_), .B0(mai_mai_n94_), .Y(mai_mai_n334_));
  NA3        m318(.A(mai_mai_n334_), .B(mai_mai_n330_), .C(mai_mai_n328_), .Y(mai_mai_n335_));
  NA2        m319(.A(mai_mai_n335_), .B(mai_mai_n325_), .Y(mai_mai_n336_));
  NO2        m320(.A(mai_mai_n210_), .B(mai_mai_n115_), .Y(mai_mai_n337_));
  NO3        m321(.A(mai_mai_n253_), .B(mai_mai_n122_), .C(mai_mai_n18_), .Y(mai_mai_n338_));
  NO2        m322(.A(mai_mai_n338_), .B(mai_mai_n337_), .Y(mai_mai_n339_));
  OAI210     m323(.A0(mai_mai_n120_), .A1(mai_mai_n108_), .B0(mai_mai_n179_), .Y(mai_mai_n340_));
  NA3        m324(.A(mai_mai_n340_), .B(x6), .C(x3), .Y(mai_mai_n341_));
  NOi21      m325(.An(mai_mai_n152_), .B(mai_mai_n132_), .Y(mai_mai_n342_));
  AOI210     m326(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n343_));
  OAI220     m327(.A0(mai_mai_n343_), .A1(mai_mai_n316_), .B0(mai_mai_n273_), .B1(mai_mai_n313_), .Y(mai_mai_n344_));
  AOI210     m328(.A0(mai_mai_n342_), .A1(mai_mai_n63_), .B0(mai_mai_n344_), .Y(mai_mai_n345_));
  NA2        m329(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n346_));
  OAI210     m330(.A0(mai_mai_n108_), .A1(mai_mai_n17_), .B0(mai_mai_n346_), .Y(mai_mai_n347_));
  AOI220     m331(.A0(mai_mai_n347_), .A1(mai_mai_n79_), .B0(mai_mai_n329_), .B1(mai_mai_n94_), .Y(mai_mai_n348_));
  NA4        m332(.A(mai_mai_n348_), .B(mai_mai_n345_), .C(mai_mai_n341_), .D(mai_mai_n339_), .Y(mai_mai_n349_));
  OAI210     m333(.A0(mai_mai_n113_), .A1(x3), .B0(mai_mai_n306_), .Y(mai_mai_n350_));
  NA3        m334(.A(mai_mai_n228_), .B(mai_mai_n214_), .C(mai_mai_n84_), .Y(mai_mai_n351_));
  NA3        m335(.A(mai_mai_n351_), .B(mai_mai_n350_), .C(mai_mai_n155_), .Y(mai_mai_n352_));
  AOI210     m336(.A0(mai_mai_n349_), .A1(x4), .B0(mai_mai_n352_), .Y(mai_mai_n353_));
  NA3        m337(.A(mai_mai_n326_), .B(mai_mai_n210_), .C(mai_mai_n94_), .Y(mai_mai_n354_));
  NOi21      m338(.An(x4), .B(x0), .Y(mai_mai_n355_));
  XO2        m339(.A(x4), .B(x0), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n356_), .A1(mai_mai_n119_), .B0(mai_mai_n268_), .Y(mai_mai_n357_));
  AOI220     m341(.A0(mai_mai_n357_), .A1(x8), .B0(mai_mai_n355_), .B1(mai_mai_n95_), .Y(mai_mai_n358_));
  AOI210     m342(.A0(mai_mai_n358_), .A1(mai_mai_n354_), .B0(x3), .Y(mai_mai_n359_));
  INV        m343(.A(mai_mai_n95_), .Y(mai_mai_n360_));
  NO2        m344(.A(mai_mai_n94_), .B(x4), .Y(mai_mai_n361_));
  AOI220     m345(.A0(mai_mai_n361_), .A1(mai_mai_n44_), .B0(mai_mai_n129_), .B1(mai_mai_n360_), .Y(mai_mai_n362_));
  NO3        m346(.A(mai_mai_n356_), .B(mai_mai_n166_), .C(x2), .Y(mai_mai_n363_));
  INV        m347(.A(mai_mai_n363_), .Y(mai_mai_n364_));
  NA4        m348(.A(mai_mai_n364_), .B(mai_mai_n362_), .C(mai_mai_n224_), .D(x6), .Y(mai_mai_n365_));
  OAI220     m349(.A0(mai_mai_n305_), .A1(mai_mai_n92_), .B0(mai_mai_n184_), .B1(mai_mai_n94_), .Y(mai_mai_n366_));
  NO2        m350(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n367_));
  OR2        m351(.A(mai_mai_n361_), .B(mai_mai_n367_), .Y(mai_mai_n368_));
  NO2        m352(.A(mai_mai_n152_), .B(mai_mai_n108_), .Y(mai_mai_n369_));
  AOI220     m353(.A0(mai_mai_n369_), .A1(mai_mai_n368_), .B0(mai_mai_n366_), .B1(mai_mai_n61_), .Y(mai_mai_n370_));
  NO2        m354(.A(mai_mai_n152_), .B(mai_mai_n81_), .Y(mai_mai_n371_));
  NO2        m355(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n372_));
  NOi21      m356(.An(mai_mai_n125_), .B(mai_mai_n27_), .Y(mai_mai_n373_));
  AOI210     m357(.A0(mai_mai_n372_), .A1(mai_mai_n371_), .B0(mai_mai_n373_), .Y(mai_mai_n374_));
  OAI210     m358(.A0(mai_mai_n370_), .A1(mai_mai_n62_), .B0(mai_mai_n374_), .Y(mai_mai_n375_));
  OAI220     m359(.A0(mai_mai_n375_), .A1(x6), .B0(mai_mai_n365_), .B1(mai_mai_n359_), .Y(mai_mai_n376_));
  OAI210     m360(.A0(mai_mai_n63_), .A1(mai_mai_n48_), .B0(mai_mai_n42_), .Y(mai_mai_n377_));
  OAI210     m361(.A0(mai_mai_n377_), .A1(mai_mai_n94_), .B0(mai_mai_n317_), .Y(mai_mai_n378_));
  AOI210     m362(.A0(mai_mai_n378_), .A1(mai_mai_n18_), .B0(mai_mai_n155_), .Y(mai_mai_n379_));
  AO220      m363(.A0(mai_mai_n379_), .A1(mai_mai_n376_), .B0(mai_mai_n353_), .B1(mai_mai_n336_), .Y(mai_mai_n380_));
  NA2        m364(.A(mai_mai_n372_), .B(x6), .Y(mai_mai_n381_));
  AOI210     m365(.A0(x6), .A1(x1), .B0(mai_mai_n154_), .Y(mai_mai_n382_));
  NA2        m366(.A(mai_mai_n361_), .B(x0), .Y(mai_mai_n383_));
  NA2        m367(.A(mai_mai_n84_), .B(x6), .Y(mai_mai_n384_));
  OAI210     m368(.A0(mai_mai_n383_), .A1(mai_mai_n382_), .B0(mai_mai_n384_), .Y(mai_mai_n385_));
  AOI220     m369(.A0(mai_mai_n385_), .A1(mai_mai_n381_), .B0(mai_mai_n218_), .B1(mai_mai_n49_), .Y(mai_mai_n386_));
  NA3        m370(.A(mai_mai_n386_), .B(mai_mai_n380_), .C(mai_mai_n323_), .Y(mai_mai_n387_));
  AOI210     m371(.A0(mai_mai_n202_), .A1(x8), .B0(mai_mai_n113_), .Y(mai_mai_n388_));
  NA2        m372(.A(mai_mai_n388_), .B(mai_mai_n346_), .Y(mai_mai_n389_));
  NA3        m373(.A(mai_mai_n389_), .B(mai_mai_n200_), .C(mai_mai_n155_), .Y(mai_mai_n390_));
  OAI210     m374(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n232_), .Y(mai_mai_n391_));
  AO220      m375(.A0(mai_mai_n391_), .A1(mai_mai_n151_), .B0(mai_mai_n112_), .B1(x4), .Y(mai_mai_n392_));
  NA3        m376(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n393_));
  NA2        m377(.A(mai_mai_n223_), .B(x0), .Y(mai_mai_n394_));
  OAI220     m378(.A0(mai_mai_n394_), .A1(mai_mai_n210_), .B0(mai_mai_n393_), .B1(mai_mai_n360_), .Y(mai_mai_n395_));
  AOI210     m379(.A0(mai_mai_n392_), .A1(mai_mai_n121_), .B0(mai_mai_n395_), .Y(mai_mai_n396_));
  AOI210     m380(.A0(mai_mai_n396_), .A1(mai_mai_n390_), .B0(mai_mai_n25_), .Y(mai_mai_n397_));
  NA3        m381(.A(mai_mai_n123_), .B(mai_mai_n223_), .C(x0), .Y(mai_mai_n398_));
  OAI210     m382(.A0(mai_mai_n200_), .A1(mai_mai_n67_), .B0(mai_mai_n206_), .Y(mai_mai_n399_));
  NA3        m383(.A(mai_mai_n202_), .B(mai_mai_n225_), .C(x8), .Y(mai_mai_n400_));
  AOI210     m384(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n25_), .Y(mai_mai_n401_));
  AOI210     m385(.A0(mai_mai_n122_), .A1(mai_mai_n120_), .B0(mai_mai_n42_), .Y(mai_mai_n402_));
  NOi31      m386(.An(mai_mai_n402_), .B(mai_mai_n367_), .C(mai_mai_n185_), .Y(mai_mai_n403_));
  OAI210     m387(.A0(mai_mai_n403_), .A1(mai_mai_n401_), .B0(mai_mai_n151_), .Y(mai_mai_n404_));
  NAi31      m388(.An(mai_mai_n50_), .B(mai_mai_n294_), .C(mai_mai_n180_), .Y(mai_mai_n405_));
  NA3        m389(.A(mai_mai_n405_), .B(mai_mai_n404_), .C(mai_mai_n398_), .Y(mai_mai_n406_));
  OAI210     m390(.A0(mai_mai_n406_), .A1(mai_mai_n397_), .B0(x6), .Y(mai_mai_n407_));
  OAI210     m391(.A0(mai_mai_n166_), .A1(mai_mai_n48_), .B0(mai_mai_n137_), .Y(mai_mai_n408_));
  NA3        m392(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n409_));
  AOI220     m393(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n410_));
  NO2        m394(.A(mai_mai_n155_), .B(x0), .Y(mai_mai_n411_));
  AOI220     m395(.A0(mai_mai_n411_), .A1(mai_mai_n223_), .B0(mai_mai_n200_), .B1(mai_mai_n155_), .Y(mai_mai_n412_));
  INV        m396(.A(x1), .Y(mai_mai_n413_));
  OAI210     m397(.A0(mai_mai_n412_), .A1(x8), .B0(mai_mai_n413_), .Y(mai_mai_n414_));
  NAi31      m398(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n415_));
  OAI210     m399(.A0(mai_mai_n415_), .A1(x4), .B0(mai_mai_n167_), .Y(mai_mai_n416_));
  NA3        m400(.A(mai_mai_n416_), .B(mai_mai_n149_), .C(x9), .Y(mai_mai_n417_));
  NO3        m401(.A(x9), .B(mai_mai_n155_), .C(x0), .Y(mai_mai_n418_));
  AOI220     m402(.A0(mai_mai_n418_), .A1(mai_mai_n246_), .B0(mai_mai_n371_), .B1(mai_mai_n155_), .Y(mai_mai_n419_));
  NA4        m403(.A(mai_mai_n419_), .B(x1), .C(mai_mai_n417_), .D(mai_mai_n50_), .Y(mai_mai_n420_));
  OAI210     m404(.A0(mai_mai_n414_), .A1(mai_mai_n410_), .B0(mai_mai_n420_), .Y(mai_mai_n421_));
  NOi31      m405(.An(mai_mai_n411_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n422_));
  AOI210     m406(.A0(mai_mai_n38_), .A1(x9), .B0(mai_mai_n135_), .Y(mai_mai_n423_));
  NO3        m407(.A(mai_mai_n423_), .B(mai_mai_n128_), .C(mai_mai_n43_), .Y(mai_mai_n424_));
  NOi31      m408(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n425_));
  AOI220     m409(.A0(mai_mai_n425_), .A1(mai_mai_n355_), .B0(mai_mai_n129_), .B1(x3), .Y(mai_mai_n426_));
  AOI210     m410(.A0(mai_mai_n268_), .A1(mai_mai_n60_), .B0(mai_mai_n127_), .Y(mai_mai_n427_));
  OAI210     m411(.A0(mai_mai_n427_), .A1(x3), .B0(mai_mai_n426_), .Y(mai_mai_n428_));
  NO3        m412(.A(mai_mai_n428_), .B(mai_mai_n424_), .C(x2), .Y(mai_mai_n429_));
  OAI220     m413(.A0(mai_mai_n356_), .A1(mai_mai_n309_), .B0(mai_mai_n305_), .B1(mai_mai_n43_), .Y(mai_mai_n430_));
  AOI210     m414(.A0(x9), .A1(mai_mai_n48_), .B0(mai_mai_n393_), .Y(mai_mai_n431_));
  AOI220     m415(.A0(mai_mai_n431_), .A1(mai_mai_n94_), .B0(mai_mai_n430_), .B1(mai_mai_n155_), .Y(mai_mai_n432_));
  NO2        m416(.A(mai_mai_n432_), .B(mai_mai_n54_), .Y(mai_mai_n433_));
  NO3        m417(.A(mai_mai_n433_), .B(mai_mai_n429_), .C(mai_mai_n422_), .Y(mai_mai_n434_));
  AOI210     m418(.A0(mai_mai_n434_), .A1(mai_mai_n421_), .B0(mai_mai_n25_), .Y(mai_mai_n435_));
  NA4        m419(.A(mai_mai_n31_), .B(mai_mai_n94_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n436_));
  NO3        m420(.A(mai_mai_n62_), .B(x4), .C(x1), .Y(mai_mai_n437_));
  NO3        m421(.A(mai_mai_n67_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n438_));
  AOI220     m422(.A0(mai_mai_n438_), .A1(mai_mai_n269_), .B0(mai_mai_n437_), .B1(mai_mai_n402_), .Y(mai_mai_n439_));
  NO2        m423(.A(mai_mai_n439_), .B(mai_mai_n105_), .Y(mai_mai_n440_));
  NO3        m424(.A(mai_mai_n273_), .B(mai_mai_n179_), .C(mai_mai_n40_), .Y(mai_mai_n441_));
  OAI210     m425(.A0(mai_mai_n441_), .A1(mai_mai_n440_), .B0(x7), .Y(mai_mai_n442_));
  NA2        m426(.A(mai_mai_n228_), .B(x7), .Y(mai_mai_n443_));
  NA3        m427(.A(mai_mai_n443_), .B(mai_mai_n154_), .C(mai_mai_n136_), .Y(mai_mai_n444_));
  NA3        m428(.A(mai_mai_n444_), .B(mai_mai_n442_), .C(mai_mai_n436_), .Y(mai_mai_n445_));
  OAI210     m429(.A0(mai_mai_n445_), .A1(mai_mai_n435_), .B0(mai_mai_n36_), .Y(mai_mai_n446_));
  NO2        m430(.A(mai_mai_n418_), .B(mai_mai_n206_), .Y(mai_mai_n447_));
  NO4        m431(.A(mai_mai_n447_), .B(mai_mai_n78_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n448_));
  NA2        m432(.A(mai_mai_n256_), .B(mai_mai_n21_), .Y(mai_mai_n449_));
  NO2        m433(.A(mai_mai_n163_), .B(mai_mai_n137_), .Y(mai_mai_n450_));
  NA2        m434(.A(mai_mai_n450_), .B(mai_mai_n449_), .Y(mai_mai_n451_));
  AOI210     m435(.A0(mai_mai_n451_), .A1(mai_mai_n170_), .B0(mai_mai_n28_), .Y(mai_mai_n452_));
  AOI220     m436(.A0(mai_mai_n367_), .A1(mai_mai_n94_), .B0(mai_mai_n152_), .B1(mai_mai_n202_), .Y(mai_mai_n453_));
  NA3        m437(.A(mai_mai_n453_), .B(mai_mai_n415_), .C(mai_mai_n92_), .Y(mai_mai_n454_));
  NA2        m438(.A(mai_mai_n454_), .B(mai_mai_n180_), .Y(mai_mai_n455_));
  OAI220     m439(.A0(mai_mai_n281_), .A1(mai_mai_n68_), .B0(mai_mai_n163_), .B1(mai_mai_n43_), .Y(mai_mai_n456_));
  NA2        m440(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n457_));
  AOI210     m441(.A0(mai_mai_n167_), .A1(mai_mai_n27_), .B0(mai_mai_n73_), .Y(mai_mai_n458_));
  OAI210     m442(.A0(mai_mai_n151_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n459_));
  NO3        m443(.A(mai_mai_n425_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n460_));
  AOI210     m444(.A0(mai_mai_n460_), .A1(mai_mai_n459_), .B0(mai_mai_n458_), .Y(mai_mai_n461_));
  OAI210     m445(.A0(mai_mai_n156_), .A1(mai_mai_n457_), .B0(mai_mai_n461_), .Y(mai_mai_n462_));
  AOI220     m446(.A0(mai_mai_n462_), .A1(x0), .B0(mai_mai_n456_), .B1(mai_mai_n137_), .Y(mai_mai_n463_));
  AOI210     m447(.A0(mai_mai_n463_), .A1(mai_mai_n455_), .B0(mai_mai_n236_), .Y(mai_mai_n464_));
  NA2        m448(.A(x9), .B(x5), .Y(mai_mai_n465_));
  NO4        m449(.A(mai_mai_n108_), .B(mai_mai_n465_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n466_));
  NO4        m450(.A(mai_mai_n466_), .B(mai_mai_n464_), .C(mai_mai_n452_), .D(mai_mai_n448_), .Y(mai_mai_n467_));
  NA3        m451(.A(mai_mai_n467_), .B(mai_mai_n446_), .C(mai_mai_n407_), .Y(mai_mai_n468_));
  AOI210     m452(.A0(mai_mai_n387_), .A1(mai_mai_n25_), .B0(mai_mai_n468_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n63_));
  INV        u047(.A(men_men_n63_), .Y(men_men_n64_));
  NO3        u048(.A(men_men_n64_), .B(men_men_n61_), .C(men_men_n60_), .Y(men_men_n65_));
  NO2        u049(.A(x7), .B(x6), .Y(men_men_n66_));
  NO2        u050(.A(men_men_n61_), .B(x5), .Y(men_men_n67_));
  NO2        u051(.A(x8), .B(x2), .Y(men_men_n68_));
  INV        u052(.A(men_men_n68_), .Y(men_men_n69_));
  AN2        u053(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n71_), .Y(men_men_n72_));
  NAi31      u056(.An(x1), .B(x9), .C(x5), .Y(men_men_n73_));
  NO2        u057(.A(men_men_n72_), .B(men_men_n70_), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n65_), .B0(x4), .Y(men_men_n75_));
  NA2        u059(.A(men_men_n48_), .B(x2), .Y(men_men_n76_));
  OAI210     u060(.A0(men_men_n76_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n77_));
  NA2        u061(.A(x5), .B(x3), .Y(men_men_n78_));
  NO2        u062(.A(x8), .B(x6), .Y(men_men_n79_));
  NO4        u063(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n66_), .D(men_men_n54_), .Y(men_men_n80_));
  NAi21      u064(.An(x4), .B(x3), .Y(men_men_n81_));
  INV        u065(.A(men_men_n81_), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(men_men_n22_), .Y(men_men_n83_));
  NO2        u067(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u068(.A(men_men_n84_), .B(x3), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n83_), .C(men_men_n18_), .Y(men_men_n86_));
  NO3        u070(.A(men_men_n86_), .B(men_men_n80_), .C(men_men_n77_), .Y(men_men_n87_));
  NO4        u071(.A(men_men_n21_), .B(x6), .C(men_men_n43_), .D(x1), .Y(men_men_n88_));
  NA2        u072(.A(men_men_n62_), .B(men_men_n48_), .Y(men_men_n89_));
  INV        u073(.A(men_men_n89_), .Y(men_men_n90_));
  OAI210     u074(.A0(men_men_n88_), .A1(men_men_n67_), .B0(men_men_n90_), .Y(men_men_n91_));
  NA2        u075(.A(x3), .B(men_men_n18_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n25_), .Y(men_men_n93_));
  INV        u077(.A(x8), .Y(men_men_n94_));
  NA2        u078(.A(x2), .B(x1), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n94_), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n93_), .Y(men_men_n97_));
  NO2        u081(.A(men_men_n97_), .B(men_men_n26_), .Y(men_men_n98_));
  AOI210     u082(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n99_));
  OAI210     u083(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n100_));
  NO3        u084(.A(men_men_n100_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n101_));
  NA2        u085(.A(x4), .B(men_men_n43_), .Y(men_men_n102_));
  NO2        u086(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n103_));
  OAI210     u087(.A0(men_men_n103_), .A1(men_men_n43_), .B0(men_men_n18_), .Y(men_men_n104_));
  AOI210     u088(.A0(men_men_n102_), .A1(men_men_n52_), .B0(men_men_n104_), .Y(men_men_n105_));
  NO2        u089(.A(x3), .B(x2), .Y(men_men_n106_));
  NA3        u090(.A(men_men_n106_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n107_));
  AOI210     u091(.A0(x8), .A1(x6), .B0(men_men_n107_), .Y(men_men_n108_));
  NA2        u092(.A(men_men_n54_), .B(x1), .Y(men_men_n109_));
  OAI210     u093(.A0(men_men_n109_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n110_));
  NO4        u094(.A(men_men_n110_), .B(men_men_n108_), .C(men_men_n105_), .D(men_men_n101_), .Y(men_men_n111_));
  AO220      u095(.A0(men_men_n111_), .A1(men_men_n91_), .B0(men_men_n87_), .B1(men_men_n75_), .Y(men02));
  NO2        u096(.A(x3), .B(men_men_n54_), .Y(men_men_n113_));
  NO2        u097(.A(x8), .B(men_men_n18_), .Y(men_men_n114_));
  NA2        u098(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n115_));
  NA2        u099(.A(men_men_n43_), .B(x0), .Y(men_men_n116_));
  OAI210     u100(.A0(men_men_n89_), .A1(men_men_n115_), .B0(men_men_n116_), .Y(men_men_n117_));
  AOI220     u101(.A0(men_men_n117_), .A1(men_men_n114_), .B0(men_men_n113_), .B1(x4), .Y(men_men_n118_));
  NO3        u102(.A(men_men_n118_), .B(x7), .C(x5), .Y(men_men_n119_));
  NA2        u103(.A(x9), .B(x2), .Y(men_men_n120_));
  OR2        u104(.A(x8), .B(x0), .Y(men_men_n121_));
  INV        u105(.A(men_men_n121_), .Y(men_men_n122_));
  NAi21      u106(.An(x2), .B(x8), .Y(men_men_n123_));
  INV        u107(.A(men_men_n123_), .Y(men_men_n124_));
  NO2        u108(.A(men_men_n124_), .B(men_men_n122_), .Y(men_men_n125_));
  NO2        u109(.A(x4), .B(x1), .Y(men_men_n126_));
  NA3        u110(.A(men_men_n126_), .B(men_men_n125_), .C(men_men_n60_), .Y(men_men_n127_));
  NOi21      u111(.An(x0), .B(x1), .Y(men_men_n128_));
  NO3        u112(.A(x9), .B(x8), .C(x7), .Y(men_men_n129_));
  NOi21      u113(.An(x0), .B(x4), .Y(men_men_n130_));
  NAi21      u114(.An(x8), .B(x7), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n131_), .B(men_men_n62_), .Y(men_men_n132_));
  AOI220     u116(.A0(men_men_n132_), .A1(men_men_n130_), .B0(men_men_n129_), .B1(men_men_n128_), .Y(men_men_n133_));
  AOI210     u117(.A0(men_men_n133_), .A1(men_men_n127_), .B0(men_men_n78_), .Y(men_men_n134_));
  NO2        u118(.A(x5), .B(men_men_n48_), .Y(men_men_n135_));
  NA2        u119(.A(x2), .B(men_men_n18_), .Y(men_men_n136_));
  AOI210     u120(.A0(men_men_n136_), .A1(men_men_n109_), .B0(men_men_n116_), .Y(men_men_n137_));
  OAI210     u121(.A0(men_men_n137_), .A1(men_men_n35_), .B0(men_men_n135_), .Y(men_men_n138_));
  NAi21      u122(.An(x0), .B(x4), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n139_), .B(x1), .Y(men_men_n140_));
  NO2        u124(.A(x7), .B(x0), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n84_), .B(men_men_n103_), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n142_), .B(x3), .Y(men_men_n143_));
  OAI210     u127(.A0(men_men_n141_), .A1(men_men_n140_), .B0(men_men_n143_), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n21_), .B(men_men_n43_), .Y(men_men_n145_));
  NA2        u129(.A(x5), .B(x0), .Y(men_men_n146_));
  NO2        u130(.A(men_men_n48_), .B(x2), .Y(men_men_n147_));
  NA3        u131(.A(men_men_n147_), .B(men_men_n146_), .C(men_men_n145_), .Y(men_men_n148_));
  NA4        u132(.A(men_men_n148_), .B(men_men_n144_), .C(men_men_n138_), .D(men_men_n36_), .Y(men_men_n149_));
  NO3        u133(.A(men_men_n149_), .B(men_men_n134_), .C(men_men_n119_), .Y(men_men_n150_));
  NO3        u134(.A(men_men_n78_), .B(men_men_n76_), .C(men_men_n24_), .Y(men_men_n151_));
  NO2        u135(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n152_));
  AOI220     u136(.A0(men_men_n128_), .A1(men_men_n152_), .B0(men_men_n67_), .B1(men_men_n17_), .Y(men_men_n153_));
  NO3        u137(.A(men_men_n153_), .B(men_men_n60_), .C(men_men_n62_), .Y(men_men_n154_));
  NA2        u138(.A(x7), .B(x3), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n102_), .B(x5), .Y(men_men_n156_));
  NO2        u140(.A(x9), .B(x7), .Y(men_men_n157_));
  NOi21      u141(.An(x8), .B(x0), .Y(men_men_n158_));
  OA210      u142(.A0(men_men_n157_), .A1(x1), .B0(men_men_n158_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n43_), .B(x2), .Y(men_men_n160_));
  INV        u144(.A(x7), .Y(men_men_n161_));
  NA2        u145(.A(men_men_n161_), .B(men_men_n18_), .Y(men_men_n162_));
  AOI220     u146(.A0(men_men_n162_), .A1(men_men_n160_), .B0(men_men_n113_), .B1(men_men_n38_), .Y(men_men_n163_));
  NO2        u147(.A(men_men_n25_), .B(x4), .Y(men_men_n164_));
  NO2        u148(.A(men_men_n164_), .B(men_men_n130_), .Y(men_men_n165_));
  NO2        u149(.A(men_men_n165_), .B(men_men_n163_), .Y(men_men_n166_));
  AOI210     u150(.A0(men_men_n159_), .A1(men_men_n156_), .B0(men_men_n166_), .Y(men_men_n167_));
  OAI210     u151(.A0(men_men_n155_), .A1(men_men_n50_), .B0(men_men_n167_), .Y(men_men_n168_));
  NA2        u152(.A(x5), .B(x1), .Y(men_men_n169_));
  INV        u153(.A(men_men_n169_), .Y(men_men_n170_));
  AOI210     u154(.A0(men_men_n170_), .A1(men_men_n130_), .B0(men_men_n36_), .Y(men_men_n171_));
  NO2        u155(.A(men_men_n62_), .B(men_men_n94_), .Y(men_men_n172_));
  NAi21      u156(.An(x2), .B(x7), .Y(men_men_n173_));
  NO3        u157(.A(men_men_n173_), .B(men_men_n172_), .C(men_men_n48_), .Y(men_men_n174_));
  NA2        u158(.A(men_men_n174_), .B(men_men_n67_), .Y(men_men_n175_));
  NAi31      u159(.An(men_men_n78_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n176_));
  NA3        u160(.A(men_men_n176_), .B(men_men_n175_), .C(men_men_n171_), .Y(men_men_n177_));
  NO4        u161(.A(men_men_n177_), .B(men_men_n168_), .C(men_men_n154_), .D(men_men_n151_), .Y(men_men_n178_));
  NO2        u162(.A(men_men_n178_), .B(men_men_n150_), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n146_), .B(men_men_n142_), .Y(men_men_n180_));
  NA2        u164(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n181_));
  NA2        u165(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n182_));
  NA3        u166(.A(men_men_n182_), .B(men_men_n181_), .C(men_men_n24_), .Y(men_men_n183_));
  AN2        u167(.A(men_men_n183_), .B(men_men_n147_), .Y(men_men_n184_));
  NA2        u168(.A(x8), .B(x0), .Y(men_men_n185_));
  NO2        u169(.A(men_men_n161_), .B(men_men_n25_), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n128_), .B(x4), .Y(men_men_n187_));
  NA2        u171(.A(men_men_n187_), .B(men_men_n186_), .Y(men_men_n188_));
  AOI210     u172(.A0(men_men_n185_), .A1(men_men_n136_), .B0(men_men_n188_), .Y(men_men_n189_));
  NA2        u173(.A(x2), .B(x0), .Y(men_men_n190_));
  NA2        u174(.A(x4), .B(x1), .Y(men_men_n191_));
  NAi21      u175(.An(men_men_n126_), .B(men_men_n191_), .Y(men_men_n192_));
  NOi31      u176(.An(men_men_n192_), .B(men_men_n164_), .C(men_men_n190_), .Y(men_men_n193_));
  NO4        u177(.A(men_men_n193_), .B(men_men_n189_), .C(men_men_n184_), .D(men_men_n180_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n194_), .B(men_men_n43_), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n183_), .B(men_men_n76_), .Y(men_men_n196_));
  INV        u180(.A(men_men_n135_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n109_), .B(men_men_n17_), .Y(men_men_n198_));
  AOI210     u182(.A0(men_men_n35_), .A1(men_men_n94_), .B0(men_men_n198_), .Y(men_men_n199_));
  NO3        u183(.A(men_men_n199_), .B(men_men_n197_), .C(x7), .Y(men_men_n200_));
  NA3        u184(.A(men_men_n192_), .B(men_men_n197_), .C(men_men_n42_), .Y(men_men_n201_));
  OAI210     u185(.A0(men_men_n182_), .A1(men_men_n142_), .B0(men_men_n201_), .Y(men_men_n202_));
  NO3        u186(.A(men_men_n202_), .B(men_men_n200_), .C(men_men_n196_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n203_), .B(x3), .Y(men_men_n204_));
  NO3        u188(.A(men_men_n204_), .B(men_men_n195_), .C(men_men_n179_), .Y(men03));
  NO2        u189(.A(men_men_n48_), .B(x3), .Y(men_men_n206_));
  NO2        u190(.A(x6), .B(men_men_n25_), .Y(men_men_n207_));
  INV        u191(.A(men_men_n207_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n54_), .B(x1), .Y(men_men_n209_));
  OAI210     u193(.A0(men_men_n209_), .A1(men_men_n25_), .B0(men_men_n63_), .Y(men_men_n210_));
  OAI220     u194(.A0(men_men_n210_), .A1(men_men_n17_), .B0(men_men_n208_), .B1(men_men_n109_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n211_), .B(men_men_n206_), .Y(men_men_n212_));
  NO2        u196(.A(men_men_n78_), .B(x6), .Y(men_men_n213_));
  NA2        u197(.A(x6), .B(men_men_n25_), .Y(men_men_n214_));
  NO2        u198(.A(men_men_n214_), .B(x4), .Y(men_men_n215_));
  NO2        u199(.A(men_men_n18_), .B(x0), .Y(men_men_n216_));
  AO220      u200(.A0(men_men_n216_), .A1(men_men_n215_), .B0(men_men_n213_), .B1(men_men_n55_), .Y(men_men_n217_));
  NA2        u201(.A(men_men_n217_), .B(men_men_n62_), .Y(men_men_n218_));
  NA2        u202(.A(x3), .B(men_men_n17_), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n219_), .B(men_men_n214_), .Y(men_men_n220_));
  NA2        u204(.A(x9), .B(men_men_n54_), .Y(men_men_n221_));
  NA2        u205(.A(men_men_n221_), .B(x4), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n214_), .B(men_men_n81_), .Y(men_men_n223_));
  AOI210     u207(.A0(men_men_n25_), .A1(x3), .B0(men_men_n190_), .Y(men_men_n224_));
  AOI220     u208(.A0(men_men_n224_), .A1(men_men_n223_), .B0(men_men_n222_), .B1(men_men_n220_), .Y(men_men_n225_));
  NO3        u209(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n226_));
  NO2        u210(.A(x5), .B(x1), .Y(men_men_n227_));
  AOI220     u211(.A0(men_men_n227_), .A1(men_men_n17_), .B0(men_men_n106_), .B1(x5), .Y(men_men_n228_));
  NO2        u212(.A(men_men_n219_), .B(men_men_n181_), .Y(men_men_n229_));
  NO3        u213(.A(x3), .B(x2), .C(x1), .Y(men_men_n230_));
  NO2        u214(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n228_), .A1(men_men_n64_), .B0(men_men_n231_), .Y(men_men_n232_));
  AOI220     u216(.A0(men_men_n232_), .A1(men_men_n48_), .B0(men_men_n226_), .B1(men_men_n135_), .Y(men_men_n233_));
  NA4        u217(.A(men_men_n233_), .B(men_men_n225_), .C(men_men_n218_), .D(men_men_n212_), .Y(men_men_n234_));
  NO2        u218(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n235_), .B(men_men_n19_), .Y(men_men_n236_));
  NO2        u220(.A(x3), .B(men_men_n17_), .Y(men_men_n237_));
  NO2        u221(.A(men_men_n237_), .B(x6), .Y(men_men_n238_));
  NOi21      u222(.An(men_men_n84_), .B(men_men_n238_), .Y(men_men_n239_));
  NA2        u223(.A(men_men_n62_), .B(men_men_n94_), .Y(men_men_n240_));
  NA3        u224(.A(men_men_n240_), .B(men_men_n237_), .C(x6), .Y(men_men_n241_));
  AOI210     u225(.A0(men_men_n241_), .A1(men_men_n239_), .B0(men_men_n161_), .Y(men_men_n242_));
  AO210      u226(.A0(men_men_n242_), .A1(men_men_n236_), .B0(men_men_n186_), .Y(men_men_n243_));
  NA2        u227(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n244_));
  NA2        u228(.A(men_men_n147_), .B(men_men_n93_), .Y(men_men_n245_));
  NA2        u229(.A(x6), .B(men_men_n48_), .Y(men_men_n246_));
  OAI210     u230(.A0(men_men_n122_), .A1(men_men_n79_), .B0(x4), .Y(men_men_n247_));
  AOI210     u231(.A0(men_men_n247_), .A1(men_men_n246_), .B0(men_men_n78_), .Y(men_men_n248_));
  NO2        u232(.A(men_men_n62_), .B(x6), .Y(men_men_n249_));
  NO2        u233(.A(men_men_n169_), .B(men_men_n43_), .Y(men_men_n250_));
  OAI210     u234(.A0(men_men_n250_), .A1(men_men_n229_), .B0(men_men_n249_), .Y(men_men_n251_));
  NA2        u235(.A(men_men_n207_), .B(men_men_n140_), .Y(men_men_n252_));
  NA3        u236(.A(men_men_n219_), .B(men_men_n135_), .C(x6), .Y(men_men_n253_));
  OAI210     u237(.A0(men_men_n94_), .A1(men_men_n36_), .B0(men_men_n67_), .Y(men_men_n254_));
  NA4        u238(.A(men_men_n254_), .B(men_men_n253_), .C(men_men_n252_), .D(men_men_n251_), .Y(men_men_n255_));
  OAI210     u239(.A0(men_men_n255_), .A1(men_men_n248_), .B0(x2), .Y(men_men_n256_));
  NA3        u240(.A(men_men_n256_), .B(men_men_n245_), .C(men_men_n243_), .Y(men_men_n257_));
  AOI210     u241(.A0(men_men_n234_), .A1(x8), .B0(men_men_n257_), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n94_), .B(x3), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n259_), .B(men_men_n215_), .Y(men_men_n260_));
  NO3        u244(.A(men_men_n92_), .B(men_men_n79_), .C(men_men_n25_), .Y(men_men_n261_));
  AOI210     u245(.A0(men_men_n238_), .A1(men_men_n164_), .B0(men_men_n261_), .Y(men_men_n262_));
  AOI210     u246(.A0(men_men_n262_), .A1(men_men_n260_), .B0(x2), .Y(men_men_n263_));
  NO2        u247(.A(x4), .B(men_men_n54_), .Y(men_men_n264_));
  AOI220     u248(.A0(men_men_n215_), .A1(men_men_n198_), .B0(men_men_n264_), .B1(men_men_n67_), .Y(men_men_n265_));
  NA2        u249(.A(men_men_n62_), .B(x6), .Y(men_men_n266_));
  NA2        u250(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n267_));
  NO2        u251(.A(men_men_n267_), .B(men_men_n25_), .Y(men_men_n268_));
  NA2        u252(.A(men_men_n268_), .B(men_men_n126_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n219_), .B(x6), .Y(men_men_n270_));
  NO2        u254(.A(men_men_n219_), .B(x6), .Y(men_men_n271_));
  NAi21      u255(.An(men_men_n172_), .B(men_men_n271_), .Y(men_men_n272_));
  NA3        u256(.A(men_men_n272_), .B(men_men_n270_), .C(men_men_n152_), .Y(men_men_n273_));
  NA4        u257(.A(men_men_n273_), .B(men_men_n269_), .C(men_men_n265_), .D(men_men_n161_), .Y(men_men_n274_));
  NA2        u258(.A(men_men_n207_), .B(men_men_n237_), .Y(men_men_n275_));
  NAi21      u259(.An(x1), .B(x4), .Y(men_men_n276_));
  AOI210     u260(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n277_));
  OAI210     u261(.A0(men_men_n146_), .A1(x3), .B0(men_men_n277_), .Y(men_men_n278_));
  NA2        u262(.A(men_men_n278_), .B(men_men_n276_), .Y(men_men_n279_));
  NA2        u263(.A(men_men_n279_), .B(men_men_n275_), .Y(men_men_n280_));
  NA2        u264(.A(men_men_n62_), .B(x2), .Y(men_men_n281_));
  NO2        u265(.A(men_men_n281_), .B(men_men_n275_), .Y(men_men_n282_));
  NO3        u266(.A(x9), .B(x6), .C(x0), .Y(men_men_n283_));
  NA2        u267(.A(men_men_n109_), .B(men_men_n25_), .Y(men_men_n284_));
  NA2        u268(.A(x6), .B(x2), .Y(men_men_n285_));
  NO2        u269(.A(men_men_n285_), .B(men_men_n181_), .Y(men_men_n286_));
  AOI210     u270(.A0(men_men_n284_), .A1(men_men_n283_), .B0(men_men_n286_), .Y(men_men_n287_));
  OAI220     u271(.A0(men_men_n287_), .A1(men_men_n43_), .B0(men_men_n187_), .B1(men_men_n46_), .Y(men_men_n288_));
  OAI210     u272(.A0(men_men_n288_), .A1(men_men_n282_), .B0(men_men_n280_), .Y(men_men_n289_));
  NA2        u273(.A(x9), .B(men_men_n43_), .Y(men_men_n290_));
  NO2        u274(.A(men_men_n290_), .B(men_men_n214_), .Y(men_men_n291_));
  OR3        u275(.A(men_men_n291_), .B(men_men_n213_), .C(men_men_n156_), .Y(men_men_n292_));
  NA2        u276(.A(x4), .B(x0), .Y(men_men_n293_));
  NO3        u277(.A(men_men_n73_), .B(men_men_n293_), .C(x6), .Y(men_men_n294_));
  AOI210     u278(.A0(men_men_n292_), .A1(men_men_n42_), .B0(men_men_n294_), .Y(men_men_n295_));
  AOI210     u279(.A0(men_men_n295_), .A1(men_men_n289_), .B0(x8), .Y(men_men_n296_));
  INV        u280(.A(men_men_n266_), .Y(men_men_n297_));
  NA2        u281(.A(men_men_n227_), .B(men_men_n297_), .Y(men_men_n298_));
  INV        u282(.A(men_men_n185_), .Y(men_men_n299_));
  OAI210     u283(.A0(men_men_n299_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n300_), .A1(men_men_n298_), .B0(men_men_n244_), .Y(men_men_n301_));
  NO4        u285(.A(men_men_n301_), .B(men_men_n296_), .C(men_men_n274_), .D(men_men_n263_), .Y(men_men_n302_));
  NO2        u286(.A(men_men_n172_), .B(x1), .Y(men_men_n303_));
  NO3        u287(.A(men_men_n303_), .B(x3), .C(men_men_n36_), .Y(men_men_n304_));
  OAI210     u288(.A0(men_men_n304_), .A1(men_men_n271_), .B0(x2), .Y(men_men_n305_));
  OAI210     u289(.A0(men_men_n299_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n306_));
  AOI210     u290(.A0(men_men_n306_), .A1(men_men_n305_), .B0(men_men_n197_), .Y(men_men_n307_));
  NOi21      u291(.An(men_men_n285_), .B(men_men_n17_), .Y(men_men_n308_));
  NA3        u292(.A(men_men_n308_), .B(men_men_n227_), .C(men_men_n40_), .Y(men_men_n309_));
  AOI210     u293(.A0(men_men_n36_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n310_));
  NA3        u294(.A(men_men_n310_), .B(men_men_n170_), .C(men_men_n32_), .Y(men_men_n311_));
  NA2        u295(.A(x3), .B(x2), .Y(men_men_n312_));
  AOI220     u296(.A0(men_men_n312_), .A1(men_men_n244_), .B0(men_men_n311_), .B1(men_men_n309_), .Y(men_men_n313_));
  NAi21      u297(.An(x4), .B(x0), .Y(men_men_n314_));
  NO3        u298(.A(men_men_n314_), .B(men_men_n44_), .C(x2), .Y(men_men_n315_));
  OAI210     u299(.A0(x6), .A1(men_men_n18_), .B0(men_men_n315_), .Y(men_men_n316_));
  OAI220     u300(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n317_));
  NO2        u301(.A(x9), .B(x8), .Y(men_men_n318_));
  NA3        u302(.A(men_men_n318_), .B(men_men_n36_), .C(men_men_n54_), .Y(men_men_n319_));
  OAI210     u303(.A0(men_men_n310_), .A1(men_men_n308_), .B0(men_men_n319_), .Y(men_men_n320_));
  AOI220     u304(.A0(men_men_n320_), .A1(men_men_n82_), .B0(men_men_n317_), .B1(men_men_n31_), .Y(men_men_n321_));
  AOI210     u305(.A0(men_men_n321_), .A1(men_men_n316_), .B0(men_men_n25_), .Y(men_men_n322_));
  NA3        u306(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n323_));
  OAI210     u307(.A0(men_men_n310_), .A1(men_men_n308_), .B0(men_men_n323_), .Y(men_men_n324_));
  INV        u308(.A(men_men_n229_), .Y(men_men_n325_));
  NA2        u309(.A(men_men_n36_), .B(men_men_n43_), .Y(men_men_n326_));
  OR2        u310(.A(men_men_n326_), .B(men_men_n293_), .Y(men_men_n327_));
  OAI220     u311(.A0(men_men_n327_), .A1(men_men_n169_), .B0(men_men_n246_), .B1(men_men_n325_), .Y(men_men_n328_));
  AO210      u312(.A0(men_men_n324_), .A1(men_men_n156_), .B0(men_men_n328_), .Y(men_men_n329_));
  NO4        u313(.A(men_men_n329_), .B(men_men_n322_), .C(men_men_n313_), .D(men_men_n307_), .Y(men_men_n330_));
  OAI210     u314(.A0(men_men_n302_), .A1(men_men_n258_), .B0(men_men_n330_), .Y(men04));
  OAI210     u315(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n332_));
  NA3        u316(.A(men_men_n332_), .B(men_men_n283_), .C(men_men_n85_), .Y(men_men_n333_));
  NO2        u317(.A(x2), .B(x1), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n267_), .A1(men_men_n334_), .B0(men_men_n36_), .Y(men_men_n335_));
  NO2        u319(.A(men_men_n334_), .B(men_men_n314_), .Y(men_men_n336_));
  AOI210     u320(.A0(men_men_n62_), .A1(x4), .B0(men_men_n115_), .Y(men_men_n337_));
  OAI210     u321(.A0(men_men_n337_), .A1(men_men_n336_), .B0(men_men_n259_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n281_), .B(men_men_n92_), .Y(men_men_n339_));
  NO2        u323(.A(men_men_n339_), .B(men_men_n36_), .Y(men_men_n340_));
  NO2        u324(.A(men_men_n312_), .B(men_men_n216_), .Y(men_men_n341_));
  NA2        u325(.A(x9), .B(x0), .Y(men_men_n342_));
  AOI210     u326(.A0(men_men_n92_), .A1(men_men_n76_), .B0(men_men_n342_), .Y(men_men_n343_));
  OAI210     u327(.A0(men_men_n343_), .A1(men_men_n341_), .B0(men_men_n94_), .Y(men_men_n344_));
  NA3        u328(.A(men_men_n344_), .B(men_men_n340_), .C(men_men_n338_), .Y(men_men_n345_));
  NA2        u329(.A(men_men_n345_), .B(men_men_n335_), .Y(men_men_n346_));
  NO2        u330(.A(men_men_n221_), .B(men_men_n116_), .Y(men_men_n347_));
  NO3        u331(.A(men_men_n266_), .B(men_men_n123_), .C(men_men_n18_), .Y(men_men_n348_));
  NO2        u332(.A(men_men_n348_), .B(men_men_n347_), .Y(men_men_n349_));
  OAI210     u333(.A0(men_men_n121_), .A1(men_men_n109_), .B0(men_men_n185_), .Y(men_men_n350_));
  NA3        u334(.A(men_men_n350_), .B(x6), .C(x3), .Y(men_men_n351_));
  NOi21      u335(.An(men_men_n158_), .B(men_men_n136_), .Y(men_men_n352_));
  AOI210     u336(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n353_));
  OAI220     u337(.A0(men_men_n353_), .A1(men_men_n326_), .B0(men_men_n281_), .B1(men_men_n323_), .Y(men_men_n354_));
  AOI210     u338(.A0(men_men_n352_), .A1(men_men_n63_), .B0(men_men_n354_), .Y(men_men_n355_));
  NA2        u339(.A(x2), .B(men_men_n17_), .Y(men_men_n356_));
  OAI210     u340(.A0(men_men_n109_), .A1(men_men_n17_), .B0(men_men_n356_), .Y(men_men_n357_));
  NA2        u341(.A(men_men_n357_), .B(men_men_n79_), .Y(men_men_n358_));
  NA4        u342(.A(men_men_n358_), .B(men_men_n355_), .C(men_men_n351_), .D(men_men_n349_), .Y(men_men_n359_));
  OAI210     u343(.A0(men_men_n114_), .A1(x3), .B0(men_men_n315_), .Y(men_men_n360_));
  NA3        u344(.A(men_men_n240_), .B(men_men_n226_), .C(men_men_n84_), .Y(men_men_n361_));
  NA3        u345(.A(men_men_n361_), .B(men_men_n360_), .C(men_men_n161_), .Y(men_men_n362_));
  AOI210     u346(.A0(men_men_n359_), .A1(x4), .B0(men_men_n362_), .Y(men_men_n363_));
  NA3        u347(.A(men_men_n336_), .B(men_men_n221_), .C(men_men_n94_), .Y(men_men_n364_));
  NOi21      u348(.An(x4), .B(x0), .Y(men_men_n365_));
  XO2        u349(.A(x4), .B(x0), .Y(men_men_n366_));
  OAI210     u350(.A0(men_men_n366_), .A1(men_men_n120_), .B0(men_men_n276_), .Y(men_men_n367_));
  AOI220     u351(.A0(men_men_n367_), .A1(x8), .B0(men_men_n365_), .B1(men_men_n95_), .Y(men_men_n368_));
  AOI210     u352(.A0(men_men_n368_), .A1(men_men_n364_), .B0(x3), .Y(men_men_n369_));
  INV        u353(.A(men_men_n95_), .Y(men_men_n370_));
  NO2        u354(.A(men_men_n94_), .B(x4), .Y(men_men_n371_));
  AOI220     u355(.A0(men_men_n371_), .A1(men_men_n44_), .B0(men_men_n130_), .B1(men_men_n370_), .Y(men_men_n372_));
  NO3        u356(.A(men_men_n366_), .B(men_men_n172_), .C(x2), .Y(men_men_n373_));
  NO3        u357(.A(men_men_n240_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n374_));
  NO2        u358(.A(men_men_n374_), .B(men_men_n373_), .Y(men_men_n375_));
  NA4        u359(.A(men_men_n375_), .B(men_men_n372_), .C(men_men_n236_), .D(x6), .Y(men_men_n376_));
  OAI220     u360(.A0(men_men_n314_), .A1(men_men_n92_), .B0(men_men_n190_), .B1(men_men_n94_), .Y(men_men_n377_));
  NO2        u361(.A(men_men_n43_), .B(x0), .Y(men_men_n378_));
  NA2        u362(.A(men_men_n377_), .B(men_men_n61_), .Y(men_men_n379_));
  NO2        u363(.A(men_men_n158_), .B(men_men_n81_), .Y(men_men_n380_));
  NO2        u364(.A(men_men_n35_), .B(x2), .Y(men_men_n381_));
  NOi21      u365(.An(men_men_n126_), .B(men_men_n27_), .Y(men_men_n382_));
  AOI210     u366(.A0(men_men_n381_), .A1(men_men_n380_), .B0(men_men_n382_), .Y(men_men_n383_));
  OAI210     u367(.A0(men_men_n379_), .A1(men_men_n62_), .B0(men_men_n383_), .Y(men_men_n384_));
  OAI220     u368(.A0(men_men_n384_), .A1(x6), .B0(men_men_n376_), .B1(men_men_n369_), .Y(men_men_n385_));
  OAI210     u369(.A0(men_men_n63_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n386_));
  OAI210     u370(.A0(men_men_n386_), .A1(men_men_n94_), .B0(men_men_n327_), .Y(men_men_n387_));
  AOI210     u371(.A0(men_men_n387_), .A1(men_men_n18_), .B0(men_men_n161_), .Y(men_men_n388_));
  AO220      u372(.A0(men_men_n388_), .A1(men_men_n385_), .B0(men_men_n363_), .B1(men_men_n346_), .Y(men_men_n389_));
  NA2        u373(.A(men_men_n381_), .B(x6), .Y(men_men_n390_));
  AOI210     u374(.A0(x6), .A1(x1), .B0(men_men_n160_), .Y(men_men_n391_));
  NA2        u375(.A(men_men_n371_), .B(x0), .Y(men_men_n392_));
  NA2        u376(.A(men_men_n84_), .B(x6), .Y(men_men_n393_));
  OAI210     u377(.A0(men_men_n392_), .A1(men_men_n391_), .B0(men_men_n393_), .Y(men_men_n394_));
  AOI220     u378(.A0(men_men_n394_), .A1(men_men_n390_), .B0(men_men_n230_), .B1(men_men_n49_), .Y(men_men_n395_));
  NA3        u379(.A(men_men_n395_), .B(men_men_n389_), .C(men_men_n333_), .Y(men_men_n396_));
  AOI210     u380(.A0(men_men_n209_), .A1(x8), .B0(men_men_n114_), .Y(men_men_n397_));
  NA2        u381(.A(men_men_n397_), .B(men_men_n356_), .Y(men_men_n398_));
  NA3        u382(.A(men_men_n398_), .B(men_men_n206_), .C(men_men_n161_), .Y(men_men_n399_));
  OAI210     u383(.A0(men_men_n28_), .A1(x1), .B0(men_men_n244_), .Y(men_men_n400_));
  AO220      u384(.A0(men_men_n400_), .A1(men_men_n157_), .B0(men_men_n113_), .B1(x4), .Y(men_men_n401_));
  NA3        u385(.A(x7), .B(x3), .C(x0), .Y(men_men_n402_));
  NA2        u386(.A(men_men_n235_), .B(x0), .Y(men_men_n403_));
  OAI220     u387(.A0(men_men_n403_), .A1(men_men_n221_), .B0(men_men_n402_), .B1(men_men_n370_), .Y(men_men_n404_));
  AOI210     u388(.A0(men_men_n401_), .A1(men_men_n122_), .B0(men_men_n404_), .Y(men_men_n405_));
  AOI210     u389(.A0(men_men_n405_), .A1(men_men_n399_), .B0(men_men_n25_), .Y(men_men_n406_));
  NA3        u390(.A(men_men_n124_), .B(men_men_n235_), .C(x0), .Y(men_men_n407_));
  NAi31      u391(.An(men_men_n50_), .B(men_men_n303_), .C(men_men_n186_), .Y(men_men_n408_));
  NA2        u392(.A(men_men_n408_), .B(men_men_n407_), .Y(men_men_n409_));
  OAI210     u393(.A0(men_men_n409_), .A1(men_men_n406_), .B0(x6), .Y(men_men_n410_));
  OAI210     u394(.A0(men_men_n172_), .A1(men_men_n48_), .B0(men_men_n141_), .Y(men_men_n411_));
  NA3        u395(.A(men_men_n55_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n412_));
  AOI220     u396(.A0(men_men_n412_), .A1(men_men_n411_), .B0(men_men_n40_), .B1(men_men_n32_), .Y(men_men_n413_));
  NO2        u397(.A(men_men_n161_), .B(x0), .Y(men_men_n414_));
  AOI220     u398(.A0(men_men_n414_), .A1(men_men_n235_), .B0(men_men_n206_), .B1(men_men_n161_), .Y(men_men_n415_));
  AOI210     u399(.A0(men_men_n132_), .A1(men_men_n264_), .B0(x1), .Y(men_men_n416_));
  OAI210     u400(.A0(men_men_n415_), .A1(x8), .B0(men_men_n416_), .Y(men_men_n417_));
  NAi31      u401(.An(x2), .B(x8), .C(x0), .Y(men_men_n418_));
  OAI210     u402(.A0(men_men_n418_), .A1(x4), .B0(men_men_n173_), .Y(men_men_n419_));
  NA3        u403(.A(men_men_n419_), .B(men_men_n155_), .C(x9), .Y(men_men_n420_));
  NO4        u404(.A(men_men_n131_), .B(men_men_n314_), .C(x9), .D(x2), .Y(men_men_n421_));
  NOi21      u405(.An(men_men_n129_), .B(men_men_n190_), .Y(men_men_n422_));
  NO3        u406(.A(men_men_n422_), .B(men_men_n421_), .C(men_men_n18_), .Y(men_men_n423_));
  NO3        u407(.A(x9), .B(men_men_n161_), .C(x0), .Y(men_men_n424_));
  AOI220     u408(.A0(men_men_n424_), .A1(men_men_n259_), .B0(men_men_n380_), .B1(men_men_n161_), .Y(men_men_n425_));
  NA4        u409(.A(men_men_n425_), .B(men_men_n423_), .C(men_men_n420_), .D(men_men_n50_), .Y(men_men_n426_));
  OAI210     u410(.A0(men_men_n417_), .A1(men_men_n413_), .B0(men_men_n426_), .Y(men_men_n427_));
  NOi31      u411(.An(men_men_n414_), .B(men_men_n32_), .C(x8), .Y(men_men_n428_));
  AOI210     u412(.A0(men_men_n38_), .A1(x9), .B0(men_men_n139_), .Y(men_men_n429_));
  NO3        u413(.A(men_men_n429_), .B(men_men_n129_), .C(men_men_n43_), .Y(men_men_n430_));
  NOi31      u414(.An(x1), .B(x8), .C(x7), .Y(men_men_n431_));
  AOI220     u415(.A0(men_men_n431_), .A1(men_men_n365_), .B0(men_men_n130_), .B1(x3), .Y(men_men_n432_));
  AOI210     u416(.A0(men_men_n276_), .A1(men_men_n60_), .B0(men_men_n128_), .Y(men_men_n433_));
  OAI210     u417(.A0(men_men_n433_), .A1(x3), .B0(men_men_n432_), .Y(men_men_n434_));
  NO3        u418(.A(men_men_n434_), .B(men_men_n430_), .C(x2), .Y(men_men_n435_));
  OAI220     u419(.A0(men_men_n366_), .A1(men_men_n318_), .B0(men_men_n314_), .B1(men_men_n43_), .Y(men_men_n436_));
  AOI210     u420(.A0(x9), .A1(men_men_n48_), .B0(men_men_n402_), .Y(men_men_n437_));
  AOI220     u421(.A0(men_men_n437_), .A1(men_men_n94_), .B0(men_men_n436_), .B1(men_men_n161_), .Y(men_men_n438_));
  NO2        u422(.A(men_men_n438_), .B(men_men_n54_), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n439_), .B(men_men_n435_), .C(men_men_n428_), .Y(men_men_n440_));
  AOI210     u424(.A0(men_men_n440_), .A1(men_men_n427_), .B0(men_men_n25_), .Y(men_men_n441_));
  NA4        u425(.A(men_men_n31_), .B(men_men_n94_), .C(x2), .D(men_men_n17_), .Y(men_men_n442_));
  NO3        u426(.A(men_men_n68_), .B(men_men_n18_), .C(x0), .Y(men_men_n443_));
  NA2        u427(.A(men_men_n443_), .B(men_men_n277_), .Y(men_men_n444_));
  NO2        u428(.A(men_men_n444_), .B(men_men_n106_), .Y(men_men_n445_));
  NO3        u429(.A(men_men_n281_), .B(men_men_n185_), .C(men_men_n40_), .Y(men_men_n446_));
  OAI210     u430(.A0(men_men_n446_), .A1(men_men_n445_), .B0(x7), .Y(men_men_n447_));
  NA2        u431(.A(men_men_n240_), .B(x7), .Y(men_men_n448_));
  NA3        u432(.A(men_men_n448_), .B(men_men_n160_), .C(men_men_n140_), .Y(men_men_n449_));
  NA3        u433(.A(men_men_n449_), .B(men_men_n447_), .C(men_men_n442_), .Y(men_men_n450_));
  OAI210     u434(.A0(men_men_n450_), .A1(men_men_n441_), .B0(men_men_n36_), .Y(men_men_n451_));
  NO2        u435(.A(men_men_n424_), .B(men_men_n216_), .Y(men_men_n452_));
  NO4        u436(.A(men_men_n452_), .B(men_men_n78_), .C(x4), .D(men_men_n54_), .Y(men_men_n453_));
  NA2        u437(.A(men_men_n267_), .B(men_men_n21_), .Y(men_men_n454_));
  NO2        u438(.A(men_men_n169_), .B(men_men_n141_), .Y(men_men_n455_));
  NA2        u439(.A(men_men_n455_), .B(men_men_n454_), .Y(men_men_n456_));
  AOI210     u440(.A0(men_men_n456_), .A1(men_men_n176_), .B0(men_men_n28_), .Y(men_men_n457_));
  AOI220     u441(.A0(men_men_n378_), .A1(men_men_n94_), .B0(men_men_n158_), .B1(men_men_n209_), .Y(men_men_n458_));
  NA3        u442(.A(men_men_n458_), .B(men_men_n418_), .C(men_men_n92_), .Y(men_men_n459_));
  NA2        u443(.A(men_men_n459_), .B(men_men_n186_), .Y(men_men_n460_));
  OAI220     u444(.A0(men_men_n290_), .A1(men_men_n69_), .B0(men_men_n169_), .B1(men_men_n43_), .Y(men_men_n461_));
  NA2        u445(.A(x3), .B(men_men_n54_), .Y(men_men_n462_));
  AOI210     u446(.A0(men_men_n173_), .A1(men_men_n27_), .B0(men_men_n73_), .Y(men_men_n463_));
  OAI210     u447(.A0(men_men_n157_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n464_));
  NO3        u448(.A(men_men_n431_), .B(x3), .C(men_men_n54_), .Y(men_men_n465_));
  AOI210     u449(.A0(men_men_n465_), .A1(men_men_n464_), .B0(men_men_n463_), .Y(men_men_n466_));
  OAI210     u450(.A0(men_men_n162_), .A1(men_men_n462_), .B0(men_men_n466_), .Y(men_men_n467_));
  AOI220     u451(.A0(men_men_n467_), .A1(x0), .B0(men_men_n461_), .B1(men_men_n141_), .Y(men_men_n468_));
  AOI210     u452(.A0(men_men_n468_), .A1(men_men_n460_), .B0(men_men_n246_), .Y(men_men_n469_));
  NA2        u453(.A(x9), .B(x5), .Y(men_men_n470_));
  NO4        u454(.A(men_men_n109_), .B(men_men_n470_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n471_));
  NO4        u455(.A(men_men_n471_), .B(men_men_n469_), .C(men_men_n457_), .D(men_men_n453_), .Y(men_men_n472_));
  NA3        u456(.A(men_men_n472_), .B(men_men_n451_), .C(men_men_n410_), .Y(men_men_n473_));
  AOI210     u457(.A0(men_men_n396_), .A1(men_men_n25_), .B0(men_men_n473_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule