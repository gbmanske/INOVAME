// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n118_, new_new_n119_,
    new_new_n121_, new_new_n122_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n271_, new_new_n272_, new_new_n273_,
    new_new_n274_, new_new_n275_, new_new_n276_, new_new_n277_,
    new_new_n278_, new_new_n279_, new_new_n280_, new_new_n281_,
    new_new_n282_, new_new_n283_, new_new_n284_, new_new_n285_,
    new_new_n286_, new_new_n287_, new_new_n288_, new_new_n289_,
    new_new_n290_, new_new_n291_, new_new_n292_, new_new_n293_,
    new_new_n294_, new_new_n295_, new_new_n296_, new_new_n297_,
    new_new_n298_, new_new_n299_, new_new_n300_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n314_, new_new_n315_, new_new_n316_, new_new_n317_,
    new_new_n318_, new_new_n319_, new_new_n320_, new_new_n321_,
    new_new_n322_, new_new_n323_, new_new_n324_, new_new_n325_,
    new_new_n326_, new_new_n327_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n336_, new_new_n337_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n352_, new_new_n353_,
    new_new_n355_, new_new_n356_, new_new_n357_, new_new_n358_,
    new_new_n359_, new_new_n360_, new_new_n361_, new_new_n362_,
    new_new_n363_, new_new_n364_, new_new_n365_, new_new_n366_,
    new_new_n367_, new_new_n368_, new_new_n369_, new_new_n370_,
    new_new_n371_, new_new_n372_, new_new_n373_, new_new_n374_,
    new_new_n375_, new_new_n376_, new_new_n377_, new_new_n378_,
    new_new_n379_, new_new_n381_, new_new_n382_, new_new_n383_,
    new_new_n384_, new_new_n385_, new_new_n386_, new_new_n387_,
    new_new_n388_, new_new_n389_, new_new_n390_, new_new_n391_,
    new_new_n392_, new_new_n393_, new_new_n394_, new_new_n395_,
    new_new_n396_, new_new_n397_, new_new_n398_, new_new_n399_,
    new_new_n400_, new_new_n401_, new_new_n402_, new_new_n403_,
    new_new_n404_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n479_,
    new_new_n480_, new_new_n481_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(ori1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_5_), .A1(new_new_n46_), .B0(new_new_n45_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n50_), .B(new_new_n44_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  INV        g034(.A(new_new_n56_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA2        g039(.A(i_1_), .B(i_10_), .Y(new_new_n62_));
  NO2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NAi21      g041(.An(new_new_n63_), .B(new_new_n58_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n49_), .B(i_2_), .Y(new_new_n65_));
  AOI210     g043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n68_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n66_), .A1(new_new_n65_), .B0(new_new_n73_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n74_), .A1(new_new_n64_), .B0(i_0_), .Y(new_new_n75_));
  NA2        g053(.A(i_12_), .B(i_5_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_9_), .Y(new_new_n77_));
  NO2        g055(.A(i_3_), .B(i_7_), .Y(new_new_n78_));
  NO2        g056(.A(new_new_n77_), .B(new_new_n60_), .Y(new_new_n79_));
  INV        g057(.A(i_6_), .Y(new_new_n80_));
  NO2        g058(.A(i_2_), .B(i_7_), .Y(new_new_n81_));
  INV        g059(.A(new_new_n81_), .Y(new_new_n82_));
  OAI210     g060(.A0(new_new_n79_), .A1(i_8_), .B0(new_new_n82_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_10_), .Y(new_new_n84_));
  NA2        g062(.A(i_6_), .B(i_9_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n84_), .B0(new_new_n60_), .Y(new_new_n86_));
  NA2        g064(.A(i_2_), .B(i_6_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n88_));
  NO2        g066(.A(new_new_n88_), .B(new_new_n86_), .Y(new_new_n89_));
  AOI210     g067(.A0(new_new_n89_), .A1(new_new_n83_), .B0(new_new_n76_), .Y(new_new_n90_));
  AN3        g068(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n91_));
  NAi21      g069(.An(i_6_), .B(i_11_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n45_), .B(new_new_n93_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n80_), .Y(new_new_n96_));
  NA2        g074(.A(i_12_), .B(i_3_), .Y(new_new_n97_));
  INV        g075(.A(new_new_n97_), .Y(new_new_n98_));
  NA3        g076(.A(new_new_n98_), .B(new_new_n96_), .C(new_new_n94_), .Y(new_new_n99_));
  NAi21      g077(.An(i_7_), .B(i_11_), .Y(new_new_n100_));
  AN2        g078(.A(i_2_), .B(i_10_), .Y(new_new_n101_));
  BUFFER     g079(.A(new_new_n76_), .Y(new_new_n102_));
  NO2        g080(.A(new_new_n60_), .B(new_new_n26_), .Y(new_new_n103_));
  NA2        g081(.A(i_11_), .B(i_12_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n104_), .B(new_new_n99_), .Y(new_new_n105_));
  NA2        g083(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n106_));
  NA2        g084(.A(i_7_), .B(new_new_n25_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n107_), .B(new_new_n106_), .Y(new_new_n108_));
  NO2        g086(.A(new_new_n108_), .B(new_new_n45_), .Y(new_new_n109_));
  NA2        g087(.A(new_new_n85_), .B(new_new_n84_), .Y(new_new_n110_));
  NAi21      g088(.An(i_3_), .B(i_8_), .Y(new_new_n111_));
  NO2        g089(.A(i_1_), .B(new_new_n80_), .Y(new_new_n112_));
  NO2        g090(.A(i_6_), .B(i_5_), .Y(new_new_n113_));
  AO210      g091(.A0(i_5_), .A1(new_new_n46_), .B0(new_new_n112_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n114_), .B(new_new_n100_), .Y(new_new_n115_));
  NO3        g093(.A(new_new_n115_), .B(new_new_n105_), .C(new_new_n90_), .Y(new_new_n116_));
  NA3        g094(.A(new_new_n116_), .B(new_new_n75_), .C(new_new_n54_), .Y(ori2));
  NO2        g095(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n479_), .B(new_new_n118_), .Y(new_new_n119_));
  NA4        g097(.A(new_new_n119_), .B(new_new_n73_), .C(new_new_n65_), .D(new_new_n30_), .Y(ori0));
  NA2        g098(.A(i_7_), .B(i_6_), .Y(new_new_n121_));
  NO2        g099(.A(i_12_), .B(i_13_), .Y(new_new_n122_));
  NAi21      g100(.An(i_5_), .B(i_11_), .Y(new_new_n123_));
  NO2        g101(.A(i_0_), .B(i_1_), .Y(new_new_n124_));
  AN2        g102(.A(new_new_n122_), .B(new_new_n77_), .Y(new_new_n125_));
  NA2        g103(.A(i_1_), .B(i_5_), .Y(new_new_n126_));
  OR2        g104(.A(i_0_), .B(i_1_), .Y(new_new_n127_));
  NOi21      g105(.An(i_4_), .B(i_10_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n40_), .Y(new_new_n129_));
  NOi21      g107(.An(i_4_), .B(i_9_), .Y(new_new_n130_));
  NOi21      g108(.An(i_11_), .B(i_13_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(new_new_n130_), .Y(new_new_n132_));
  NO2        g110(.A(new_new_n69_), .B(new_new_n60_), .Y(new_new_n133_));
  NO2        g111(.A(new_new_n69_), .B(i_5_), .Y(new_new_n134_));
  NO2        g112(.A(i_2_), .B(i_1_), .Y(new_new_n135_));
  NAi21      g113(.An(i_4_), .B(i_12_), .Y(new_new_n136_));
  INV        g114(.A(i_8_), .Y(new_new_n137_));
  NO2        g115(.A(i_3_), .B(i_8_), .Y(new_new_n138_));
  NO3        g116(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n139_));
  NO2        g117(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n140_));
  NO2        g118(.A(i_13_), .B(i_9_), .Y(new_new_n141_));
  NO2        g119(.A(new_new_n43_), .B(i_5_), .Y(new_new_n142_));
  NA2        g120(.A(i_0_), .B(i_5_), .Y(new_new_n143_));
  NAi31      g121(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n144_));
  INV        g122(.A(i_13_), .Y(new_new_n145_));
  NO2        g123(.A(i_12_), .B(new_new_n145_), .Y(new_new_n146_));
  INV        g124(.A(i_12_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n43_), .B(new_new_n147_), .Y(new_new_n148_));
  NO3        g126(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n149_));
  NA2        g127(.A(i_2_), .B(i_1_), .Y(new_new_n150_));
  NO3        g128(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n151_));
  NAi21      g129(.An(i_4_), .B(i_3_), .Y(new_new_n152_));
  NOi41      g130(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n153_));
  NO2        g131(.A(i_11_), .B(new_new_n145_), .Y(new_new_n154_));
  NOi21      g132(.An(i_1_), .B(i_6_), .Y(new_new_n155_));
  INV        g133(.A(i_7_), .Y(new_new_n156_));
  NA2        g134(.A(new_new_n147_), .B(i_9_), .Y(new_new_n157_));
  OR4        g135(.A(new_new_n157_), .B(new_new_n156_), .C(new_new_n155_), .D(new_new_n134_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n69_), .B(i_5_), .Y(new_new_n159_));
  NA2        g137(.A(i_3_), .B(i_9_), .Y(new_new_n160_));
  NAi21      g138(.An(i_7_), .B(i_10_), .Y(new_new_n161_));
  NO2        g139(.A(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NA3        g140(.A(new_new_n162_), .B(new_new_n159_), .C(new_new_n61_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n163_), .B(new_new_n158_), .Y(new_new_n164_));
  INV        g142(.A(new_new_n121_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n147_), .B(i_13_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n166_), .B(new_new_n71_), .Y(new_new_n167_));
  AOI220     g145(.A0(new_new_n167_), .A1(new_new_n165_), .B0(new_new_n164_), .B1(new_new_n154_), .Y(new_new_n168_));
  NA2        g146(.A(i_12_), .B(i_6_), .Y(new_new_n169_));
  OR2        g147(.A(i_13_), .B(i_9_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n152_), .B(i_2_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n154_), .B(i_9_), .Y(new_new_n172_));
  NO3        g150(.A(i_12_), .B(new_new_n145_), .C(new_new_n37_), .Y(new_new_n173_));
  AN2        g151(.A(i_3_), .B(i_10_), .Y(new_new_n174_));
  NO2        g152(.A(i_5_), .B(new_new_n37_), .Y(new_new_n175_));
  NO2        g153(.A(new_new_n45_), .B(new_new_n26_), .Y(new_new_n176_));
  NO3        g154(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n177_));
  NO2        g155(.A(i_2_), .B(i_3_), .Y(new_new_n178_));
  NO2        g156(.A(i_12_), .B(i_10_), .Y(new_new_n179_));
  NOi21      g157(.An(i_5_), .B(i_0_), .Y(new_new_n180_));
  NOi21      g158(.An(new_new_n126_), .B(new_new_n96_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n181_), .B(new_new_n107_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(i_3_), .Y(new_new_n183_));
  NO2        g161(.A(new_new_n137_), .B(i_9_), .Y(new_new_n184_));
  NA2        g162(.A(new_new_n184_), .B(new_new_n140_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(new_new_n45_), .Y(new_new_n186_));
  INV        g164(.A(new_new_n186_), .Y(new_new_n187_));
  AOI210     g165(.A0(new_new_n187_), .A1(new_new_n183_), .B0(new_new_n129_), .Y(new_new_n188_));
  INV        g166(.A(new_new_n188_), .Y(new_new_n189_));
  NOi32      g167(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n190_));
  INV        g168(.A(new_new_n190_), .Y(new_new_n191_));
  NOi32      g169(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n192_));
  NO2        g170(.A(i_1_), .B(new_new_n93_), .Y(new_new_n193_));
  NAi21      g171(.An(i_3_), .B(i_4_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n194_), .B(i_9_), .Y(new_new_n195_));
  AN2        g173(.A(i_6_), .B(i_7_), .Y(new_new_n196_));
  OAI210     g174(.A0(new_new_n196_), .A1(new_new_n193_), .B0(new_new_n195_), .Y(new_new_n197_));
  NA2        g175(.A(i_2_), .B(i_7_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n194_), .B(i_10_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n197_), .B(new_new_n134_), .Y(new_new_n200_));
  AOI210     g178(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n201_));
  OAI210     g179(.A0(new_new_n201_), .A1(new_new_n135_), .B0(new_new_n199_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n202_), .B(i_5_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n203_), .B(new_new_n200_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n204_), .B(new_new_n191_), .Y(new_new_n205_));
  AN2        g183(.A(i_12_), .B(i_5_), .Y(new_new_n206_));
  NO2        g184(.A(i_11_), .B(i_6_), .Y(new_new_n207_));
  NO2        g185(.A(i_5_), .B(i_10_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n209_));
  NO3        g187(.A(i_1_), .B(i_12_), .C(new_new_n80_), .Y(new_new_n210_));
  NO2        g188(.A(i_0_), .B(i_11_), .Y(new_new_n211_));
  BUFFER     g189(.A(i_6_), .Y(new_new_n212_));
  NAi21      g190(.An(i_9_), .B(i_4_), .Y(new_new_n213_));
  OR2        g191(.A(i_13_), .B(i_10_), .Y(new_new_n214_));
  NO3        g192(.A(new_new_n214_), .B(new_new_n104_), .C(new_new_n213_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n173_), .B(new_new_n216_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n217_), .B(new_new_n181_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n137_), .B(i_10_), .Y(new_new_n219_));
  NA3        g197(.A(new_new_n159_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  INV        g199(.A(new_new_n221_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n222_), .B(new_new_n172_), .Y(new_new_n223_));
  NO3        g201(.A(new_new_n223_), .B(new_new_n218_), .C(new_new_n205_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n69_), .B(i_13_), .Y(new_new_n225_));
  NO2        g203(.A(i_10_), .B(i_9_), .Y(new_new_n226_));
  NO3        g204(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n169_), .B(new_new_n92_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  NA2        g207(.A(i_8_), .B(i_9_), .Y(new_new_n230_));
  NO2        g208(.A(i_7_), .B(i_2_), .Y(new_new_n231_));
  OR2        g209(.A(new_new_n231_), .B(new_new_n230_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n173_), .B(new_new_n140_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n154_), .B(new_new_n175_), .Y(new_new_n235_));
  NO3        g213(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n236_));
  INV        g214(.A(new_new_n236_), .Y(new_new_n237_));
  NA3        g215(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n238_));
  NA4        g216(.A(new_new_n123_), .B(new_new_n103_), .C(new_new_n76_), .D(new_new_n23_), .Y(new_new_n239_));
  OAI220     g217(.A0(new_new_n239_), .A1(new_new_n238_), .B0(new_new_n237_), .B1(new_new_n235_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n240_), .B(new_new_n234_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n91_), .B(i_13_), .Y(new_new_n242_));
  NO2        g220(.A(i_11_), .B(i_1_), .Y(new_new_n243_));
  NA3        g221(.A(new_new_n153_), .B(new_new_n131_), .C(new_new_n113_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n45_), .B(new_new_n43_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n127_), .B(i_3_), .Y(new_new_n246_));
  NAi31      g224(.An(new_new_n245_), .B(new_new_n246_), .C(new_new_n146_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n247_), .B(new_new_n244_), .Y(new_new_n248_));
  INV        g226(.A(new_new_n248_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n227_), .B(new_new_n206_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n236_), .B(new_new_n208_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n27_), .B(i_10_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n177_), .B(new_new_n149_), .Y(new_new_n253_));
  OAI220     g231(.A0(new_new_n253_), .A1(new_new_n220_), .B0(new_new_n252_), .B1(new_new_n242_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n254_), .Y(new_new_n255_));
  NA3        g233(.A(new_new_n255_), .B(new_new_n249_), .C(new_new_n241_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n206_), .B(new_new_n145_), .Y(new_new_n257_));
  NA2        g235(.A(new_new_n196_), .B(new_new_n192_), .Y(new_new_n258_));
  OR2        g236(.A(new_new_n257_), .B(new_new_n258_), .Y(new_new_n259_));
  AOI210     g237(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n215_), .Y(new_new_n260_));
  NA2        g238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  NA3        g239(.A(new_new_n143_), .B(new_new_n67_), .C(new_new_n43_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n173_), .B(new_new_n78_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n262_), .B(new_new_n263_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n214_), .B(i_1_), .Y(new_new_n265_));
  NOi31      g243(.An(new_new_n265_), .B(new_new_n228_), .C(new_new_n69_), .Y(new_new_n266_));
  NOi21      g244(.An(i_10_), .B(i_6_), .Y(new_new_n267_));
  OR2        g245(.A(i_2_), .B(i_5_), .Y(new_new_n268_));
  NO3        g246(.A(new_new_n264_), .B(new_new_n261_), .C(new_new_n256_), .Y(new_new_n269_));
  NA4        g247(.A(new_new_n269_), .B(new_new_n224_), .C(new_new_n189_), .D(new_new_n168_), .Y(ori7));
  NO2        g248(.A(new_new_n87_), .B(new_new_n52_), .Y(new_new_n271_));
  NA2        g249(.A(i_11_), .B(new_new_n137_), .Y(new_new_n272_));
  NA3        g250(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n147_), .B(i_4_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n274_), .B(i_8_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n97_), .B(new_new_n273_), .Y(new_new_n276_));
  NA2        g254(.A(i_2_), .B(new_new_n80_), .Y(new_new_n277_));
  OAI210     g255(.A0(new_new_n81_), .A1(new_new_n138_), .B0(new_new_n139_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n276_), .B(new_new_n271_), .Y(new_new_n279_));
  AOI210     g257(.A0(new_new_n111_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n280_));
  AOI210     g258(.A0(new_new_n280_), .A1(new_new_n147_), .B0(new_new_n128_), .Y(new_new_n281_));
  OR2        g259(.A(i_6_), .B(i_10_), .Y(new_new_n282_));
  OR3        g260(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n283_));
  OR2        g261(.A(new_new_n281_), .B(new_new_n170_), .Y(new_new_n284_));
  AOI210     g262(.A0(new_new_n284_), .A1(new_new_n279_), .B0(new_new_n60_), .Y(new_new_n285_));
  NOi21      g263(.An(i_11_), .B(i_7_), .Y(new_new_n286_));
  AO210      g264(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(new_new_n286_), .Y(new_new_n288_));
  NA2        g266(.A(new_new_n288_), .B(new_new_n141_), .Y(new_new_n289_));
  NA3        g267(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n289_), .B(new_new_n60_), .Y(new_new_n291_));
  NA2        g269(.A(new_new_n146_), .B(new_new_n60_), .Y(new_new_n292_));
  NO2        g270(.A(i_1_), .B(i_12_), .Y(new_new_n293_));
  INV        g271(.A(new_new_n292_), .Y(new_new_n294_));
  OAI210     g272(.A0(new_new_n294_), .A1(new_new_n291_), .B0(i_6_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n290_), .B(new_new_n100_), .Y(new_new_n296_));
  NA2        g274(.A(new_new_n296_), .B(i_6_), .Y(new_new_n297_));
  NO2        g275(.A(i_6_), .B(i_11_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n297_), .B(new_new_n229_), .Y(new_new_n299_));
  NO3        g277(.A(new_new_n282_), .B(i_7_), .C(new_new_n23_), .Y(new_new_n300_));
  AOI210     g278(.A0(i_1_), .A1(new_new_n162_), .B0(new_new_n300_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(new_new_n43_), .Y(new_new_n302_));
  INV        g280(.A(i_2_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n118_), .B(i_9_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n304_), .B(new_new_n303_), .Y(new_new_n305_));
  AOI210     g283(.A0(new_new_n243_), .A1(new_new_n216_), .B0(new_new_n151_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(new_new_n277_), .Y(new_new_n307_));
  OR2        g285(.A(new_new_n307_), .B(new_new_n305_), .Y(new_new_n308_));
  NO3        g286(.A(new_new_n308_), .B(new_new_n302_), .C(new_new_n299_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n147_), .B(new_new_n93_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n310_), .B(new_new_n286_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n311_), .B(i_1_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n312_), .B(new_new_n283_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n213_), .B(new_new_n80_), .Y(new_new_n314_));
  NA2        g292(.A(new_new_n313_), .B(new_new_n45_), .Y(new_new_n315_));
  NO2        g293(.A(i_7_), .B(new_new_n43_), .Y(new_new_n316_));
  NO3        g294(.A(new_new_n316_), .B(new_new_n176_), .C(new_new_n148_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n318_));
  NO2        g296(.A(new_new_n318_), .B(i_6_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n80_), .B(i_9_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(new_new_n60_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n321_), .B(new_new_n293_), .Y(new_new_n322_));
  NO4        g300(.A(new_new_n322_), .B(new_new_n319_), .C(new_new_n317_), .D(i_4_), .Y(new_new_n323_));
  INV        g301(.A(new_new_n323_), .Y(new_new_n324_));
  NA4        g302(.A(new_new_n324_), .B(new_new_n315_), .C(new_new_n309_), .D(new_new_n295_), .Y(new_new_n325_));
  AOI210     g303(.A0(new_new_n169_), .A1(new_new_n92_), .B0(i_1_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n194_), .B(i_2_), .Y(new_new_n327_));
  NA2        g305(.A(new_new_n327_), .B(new_new_n326_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n328_), .B(i_13_), .Y(new_new_n329_));
  OR2        g307(.A(i_11_), .B(i_7_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n52_), .B(i_12_), .Y(new_new_n331_));
  INV        g309(.A(new_new_n331_), .Y(new_new_n332_));
  NA2        g310(.A(i_7_), .B(new_new_n314_), .Y(new_new_n333_));
  OAI220     g311(.A0(new_new_n333_), .A1(new_new_n41_), .B0(new_new_n332_), .B1(new_new_n87_), .Y(new_new_n334_));
  INV        g312(.A(new_new_n334_), .Y(new_new_n335_));
  NA2        g313(.A(new_new_n110_), .B(i_13_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n336_), .B(new_new_n326_), .Y(new_new_n337_));
  INV        g315(.A(i_7_), .Y(new_new_n338_));
  AOI220     g316(.A0(new_new_n207_), .A1(new_new_n481_), .B0(new_new_n86_), .B1(new_new_n94_), .Y(new_new_n339_));
  NO2        g317(.A(new_new_n339_), .B(new_new_n275_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n340_), .B(new_new_n337_), .Y(new_new_n341_));
  OR2        g319(.A(i_11_), .B(i_6_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n274_), .B(i_7_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n343_), .B(new_new_n342_), .Y(new_new_n344_));
  NA2        g322(.A(new_new_n298_), .B(i_13_), .Y(new_new_n345_));
  INV        g323(.A(new_new_n345_), .Y(new_new_n346_));
  OAI210     g324(.A0(new_new_n346_), .A1(new_new_n344_), .B0(new_new_n60_), .Y(new_new_n347_));
  NO2        g325(.A(i_2_), .B(i_12_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n193_), .B(new_new_n348_), .Y(new_new_n349_));
  NA2        g327(.A(new_new_n195_), .B(new_new_n193_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n350_), .B(new_new_n349_), .Y(new_new_n351_));
  NA3        g329(.A(new_new_n351_), .B(new_new_n44_), .C(new_new_n145_), .Y(new_new_n352_));
  NA4        g330(.A(new_new_n352_), .B(new_new_n347_), .C(new_new_n341_), .D(new_new_n335_), .Y(new_new_n353_));
  OR4        g331(.A(new_new_n353_), .B(new_new_n329_), .C(new_new_n325_), .D(new_new_n285_), .Y(ori5));
  NA2        g332(.A(new_new_n311_), .B(new_new_n171_), .Y(new_new_n355_));
  NA3        g333(.A(new_new_n24_), .B(new_new_n348_), .C(new_new_n100_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n356_), .B(new_new_n355_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n107_), .B(new_new_n23_), .Y(new_new_n358_));
  INV        g336(.A(new_new_n226_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n358_), .B(new_new_n357_), .Y(new_new_n360_));
  INV        g338(.A(new_new_n153_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(i_13_), .Y(new_new_n362_));
  INV        g340(.A(new_new_n362_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n136_), .B(new_new_n108_), .Y(new_new_n364_));
  OAI210     g342(.A0(new_new_n364_), .A1(new_new_n358_), .B0(i_2_), .Y(new_new_n365_));
  INV        g343(.A(new_new_n132_), .Y(new_new_n366_));
  NO3        g344(.A(new_new_n287_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n366_), .B(new_new_n367_), .Y(new_new_n368_));
  AOI210     g346(.A0(new_new_n368_), .A1(new_new_n365_), .B0(new_new_n137_), .Y(new_new_n369_));
  OA210      g347(.A0(new_new_n288_), .A1(new_new_n109_), .B0(i_13_), .Y(new_new_n370_));
  INV        g348(.A(new_new_n125_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n371_), .B(new_new_n198_), .Y(new_new_n372_));
  NA3        g350(.A(i_2_), .B(new_new_n174_), .C(new_new_n107_), .Y(new_new_n373_));
  INV        g351(.A(new_new_n373_), .Y(new_new_n374_));
  NO4        g352(.A(new_new_n374_), .B(new_new_n372_), .C(new_new_n370_), .D(new_new_n369_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n59_), .B(i_12_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(new_new_n109_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n377_), .B(new_new_n272_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n378_), .B(new_new_n36_), .Y(new_new_n379_));
  NA4        g357(.A(new_new_n379_), .B(new_new_n375_), .C(new_new_n363_), .D(new_new_n360_), .Y(ori6));
  NO2        g358(.A(new_new_n144_), .B(new_new_n245_), .Y(new_new_n381_));
  INV        g359(.A(new_new_n180_), .Y(new_new_n382_));
  OR2        g360(.A(new_new_n382_), .B(i_12_), .Y(new_new_n383_));
  INV        g361(.A(new_new_n179_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n71_), .B(new_new_n112_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n155_), .B(i_9_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n387_), .B(new_new_n376_), .Y(new_new_n388_));
  AOI210     g366(.A0(new_new_n388_), .A1(new_new_n258_), .B0(new_new_n134_), .Y(new_new_n389_));
  NAi32      g367(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n342_), .B(new_new_n390_), .Y(new_new_n391_));
  OR3        g369(.A(new_new_n391_), .B(new_new_n389_), .C(new_new_n386_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n330_), .B(i_2_), .Y(new_new_n393_));
  BUFFER     g371(.A(new_new_n288_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n394_), .B(new_new_n124_), .Y(new_new_n395_));
  AO210      g373(.A0(new_new_n251_), .A1(new_new_n359_), .B0(new_new_n36_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n396_), .B(new_new_n395_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n381_), .B(new_new_n338_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n398_), .B(new_new_n278_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n282_), .B(new_new_n94_), .Y(new_new_n400_));
  OAI210     g378(.A0(new_new_n400_), .A1(new_new_n102_), .B0(new_new_n211_), .Y(new_new_n401_));
  NA3        g379(.A(new_new_n480_), .B(new_new_n179_), .C(i_7_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n402_), .B(new_new_n401_), .Y(new_new_n403_));
  NO4        g381(.A(new_new_n403_), .B(new_new_n399_), .C(new_new_n397_), .D(new_new_n392_), .Y(new_new_n404_));
  NA3        g382(.A(new_new_n404_), .B(new_new_n383_), .C(new_new_n204_), .Y(ori3));
  NA2        g383(.A(i_12_), .B(i_10_), .Y(new_new_n406_));
  NO2        g384(.A(i_11_), .B(new_new_n147_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n278_), .B(new_new_n197_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n408_), .B(new_new_n40_), .Y(new_new_n409_));
  NOi21      g387(.An(new_new_n91_), .B(new_new_n25_), .Y(new_new_n410_));
  AN2        g388(.A(new_new_n228_), .B(new_new_n53_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(new_new_n410_), .Y(new_new_n412_));
  AOI210     g390(.A0(new_new_n412_), .A1(new_new_n409_), .B0(new_new_n47_), .Y(new_new_n413_));
  NO3        g391(.A(new_new_n206_), .B(new_new_n38_), .C(i_0_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n134_), .B(new_new_n267_), .Y(new_new_n415_));
  NOi21      g393(.An(new_new_n415_), .B(new_new_n414_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n416_), .B(new_new_n60_), .Y(new_new_n417_));
  NOi21      g395(.An(i_5_), .B(i_9_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n418_), .B(new_new_n225_), .Y(new_new_n419_));
  BUFFER     g397(.A(new_new_n169_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n420_), .B(new_new_n243_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n421_), .B(new_new_n419_), .Y(new_new_n422_));
  NO3        g400(.A(new_new_n422_), .B(new_new_n417_), .C(new_new_n413_), .Y(new_new_n423_));
  NO4        g401(.A(new_new_n268_), .B(i_12_), .C(new_new_n214_), .D(new_new_n212_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n424_), .B(i_11_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n157_), .B(new_new_n126_), .Y(new_new_n426_));
  NA2        g404(.A(i_0_), .B(i_10_), .Y(new_new_n427_));
  AN2        g405(.A(new_new_n426_), .B(i_6_), .Y(new_new_n428_));
  INV        g406(.A(new_new_n428_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n425_), .Y(new_new_n430_));
  NA2        g408(.A(i_11_), .B(i_9_), .Y(new_new_n431_));
  NO3        g409(.A(i_12_), .B(new_new_n431_), .C(new_new_n277_), .Y(new_new_n432_));
  AN2        g410(.A(new_new_n432_), .B(i_5_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n209_), .B(new_new_n133_), .Y(new_new_n434_));
  INV        g412(.A(new_new_n434_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n431_), .B(new_new_n69_), .Y(new_new_n436_));
  INV        g414(.A(new_new_n210_), .Y(new_new_n437_));
  NO2        g415(.A(new_new_n437_), .B(new_new_n419_), .Y(new_new_n438_));
  NO3        g416(.A(new_new_n438_), .B(new_new_n435_), .C(new_new_n433_), .Y(new_new_n439_));
  INV        g417(.A(new_new_n439_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n406_), .B(new_new_n178_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n441_), .B(new_new_n436_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n259_), .B(new_new_n442_), .Y(new_new_n443_));
  NO3        g421(.A(new_new_n443_), .B(new_new_n440_), .C(new_new_n430_), .Y(new_new_n444_));
  NO3        g422(.A(new_new_n427_), .B(new_new_n418_), .C(new_new_n136_), .Y(new_new_n445_));
  AOI220     g423(.A0(new_new_n445_), .A1(i_11_), .B0(new_new_n266_), .B1(new_new_n71_), .Y(new_new_n446_));
  NO3        g424(.A(new_new_n142_), .B(new_new_n206_), .C(i_0_), .Y(new_new_n447_));
  OAI210     g425(.A0(new_new_n447_), .A1(new_new_n72_), .B0(i_13_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n448_), .B(new_new_n446_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n250_), .B(new_new_n244_), .Y(new_new_n450_));
  INV        g428(.A(new_new_n450_), .Y(new_new_n451_));
  NA3        g429(.A(new_new_n208_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n452_));
  INV        g430(.A(new_new_n452_), .Y(new_new_n453_));
  NO3        g431(.A(new_new_n431_), .B(new_new_n143_), .C(new_new_n136_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(new_new_n451_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n80_), .B(i_5_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n407_), .B(new_new_n101_), .Y(new_new_n458_));
  INV        g436(.A(new_new_n458_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n459_), .B(new_new_n457_), .Y(new_new_n460_));
  NAi21      g438(.An(new_new_n151_), .B(new_new_n152_), .Y(new_new_n461_));
  NO4        g439(.A(new_new_n150_), .B(new_new_n142_), .C(i_0_), .D(i_12_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n462_), .B(new_new_n461_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n463_), .B(new_new_n460_), .Y(new_new_n464_));
  NO3        g442(.A(new_new_n464_), .B(new_new_n456_), .C(new_new_n449_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n393_), .B(new_new_n37_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n466_), .B(new_new_n281_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n467_), .B(new_new_n141_), .Y(new_new_n468_));
  NA2        g446(.A(i_2_), .B(i_10_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n66_), .B(new_new_n469_), .Y(new_new_n470_));
  AOI210     g448(.A0(new_new_n470_), .A1(new_new_n47_), .B0(new_new_n424_), .Y(new_new_n471_));
  AOI210     g449(.A0(new_new_n471_), .A1(new_new_n468_), .B0(new_new_n69_), .Y(new_new_n472_));
  INV        g450(.A(new_new_n203_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n473_), .B(i_13_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n472_), .Y(new_new_n475_));
  NA4        g453(.A(new_new_n475_), .B(new_new_n465_), .C(new_new_n444_), .D(new_new_n423_), .Y(ori4));
  INV        g454(.A(i_6_), .Y(new_new_n479_));
  INV        g455(.A(new_new_n268_), .Y(new_new_n480_));
  INV        g456(.A(i_1_), .Y(new_new_n481_));
endmodule


