//Benchmark atmr_misex3_1774_0.0625

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1586_, men_men_n1587_, men_men_n1588_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o000(.A(f), .B(e), .Y(ori_ori_n29_));
  NOi32      o001(.An(m), .Bn(l), .C(n), .Y(ori_ori_n30_));
  NOi32      o002(.An(i), .Bn(g), .C(h), .Y(ori_ori_n31_));
  NA2        o003(.A(ori_ori_n31_), .B(ori_ori_n30_), .Y(ori_ori_n32_));
  AN2        o004(.A(m), .B(l), .Y(ori_ori_n33_));
  NOi32      o005(.An(j), .Bn(g), .C(k), .Y(ori_ori_n34_));
  NA2        o006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  INV        o007(.A(h), .Y(ori_ori_n36_));
  NAi21      o008(.An(j), .B(l), .Y(ori_ori_n37_));
  INV        o009(.A(i), .Y(ori_ori_n38_));
  AN2        o010(.A(h), .B(g), .Y(ori_ori_n39_));
  NAi21      o011(.An(n), .B(m), .Y(ori_ori_n40_));
  NOi32      o012(.An(k), .Bn(h), .C(l), .Y(ori_ori_n41_));
  NOi32      o013(.An(k), .Bn(h), .C(g), .Y(ori_ori_n42_));
  INV        o014(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o015(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o016(.A(c), .Y(ori_ori_n45_));
  NA2        o017(.A(e), .B(b), .Y(ori_ori_n46_));
  NO2        o018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  INV        o019(.A(d), .Y(ori_ori_n48_));
  NAi21      o020(.An(i), .B(h), .Y(ori_ori_n49_));
  INV        o021(.A(f), .Y(ori_ori_n50_));
  NAi32      o022(.An(n), .Bn(k), .C(m), .Y(ori_ori_n51_));
  NAi21      o023(.An(e), .B(h), .Y(ori_ori_n52_));
  INV        o024(.A(m), .Y(ori_ori_n53_));
  NOi21      o025(.An(k), .B(l), .Y(ori_ori_n54_));
  NA2        o026(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  AN4        o027(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n56_));
  NOi21      o028(.An(h), .B(f), .Y(ori_ori_n57_));
  NA2        o029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  NAi32      o030(.An(m), .Bn(k), .C(j), .Y(ori_ori_n59_));
  NOi32      o031(.An(h), .Bn(g), .C(f), .Y(ori_ori_n60_));
  OR2        o032(.A(ori_ori_n58_), .B(ori_ori_n55_), .Y(ori_ori_n61_));
  INV        o033(.A(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o034(.A(n), .Y(ori_ori_n63_));
  NOi32      o035(.An(e), .Bn(b), .C(d), .Y(ori_ori_n64_));
  INV        o036(.A(j), .Y(ori_ori_n65_));
  AN3        o037(.A(m), .B(k), .C(i), .Y(ori_ori_n66_));
  NA3        o038(.A(ori_ori_n66_), .B(ori_ori_n65_), .C(g), .Y(ori_ori_n67_));
  NAi32      o039(.An(g), .Bn(f), .C(h), .Y(ori_ori_n68_));
  NA2        o040(.A(m), .B(l), .Y(ori_ori_n69_));
  AN2        o041(.A(j), .B(g), .Y(ori_ori_n70_));
  NOi32      o042(.An(m), .Bn(l), .C(i), .Y(ori_ori_n71_));
  NOi21      o043(.An(g), .B(i), .Y(ori_ori_n72_));
  NOi32      o044(.An(m), .Bn(j), .C(k), .Y(ori_ori_n73_));
  AOI220     o045(.A0(ori_ori_n73_), .A1(ori_ori_n72_), .B0(ori_ori_n71_), .B1(ori_ori_n70_), .Y(ori_ori_n74_));
  NAi41      o046(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n75_));
  AN2        o047(.A(e), .B(b), .Y(ori_ori_n76_));
  NOi31      o048(.An(c), .B(h), .C(f), .Y(ori_ori_n77_));
  NA2        o049(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n78_));
  NO2        o050(.A(ori_ori_n78_), .B(ori_ori_n75_), .Y(ori_ori_n79_));
  NOi21      o051(.An(g), .B(f), .Y(ori_ori_n80_));
  NOi21      o052(.An(i), .B(h), .Y(ori_ori_n81_));
  INV        o053(.A(a), .Y(ori_ori_n82_));
  NA2        o054(.A(ori_ori_n76_), .B(ori_ori_n82_), .Y(ori_ori_n83_));
  INV        o055(.A(l), .Y(ori_ori_n84_));
  NOi21      o056(.An(m), .B(n), .Y(ori_ori_n85_));
  AN2        o057(.A(k), .B(h), .Y(ori_ori_n86_));
  INV        o058(.A(b), .Y(ori_ori_n87_));
  AN2        o059(.A(k), .B(i), .Y(ori_ori_n88_));
  NOi31      o060(.An(k), .B(m), .C(j), .Y(ori_ori_n89_));
  NA3        o061(.A(ori_ori_n89_), .B(ori_ori_n57_), .C(ori_ori_n56_), .Y(ori_ori_n90_));
  NOi31      o062(.An(k), .B(m), .C(i), .Y(ori_ori_n91_));
  INV        o063(.A(ori_ori_n90_), .Y(ori_ori_n92_));
  NOi32      o064(.An(f), .Bn(b), .C(e), .Y(ori_ori_n93_));
  NAi21      o065(.An(g), .B(h), .Y(ori_ori_n94_));
  NAi21      o066(.An(m), .B(n), .Y(ori_ori_n95_));
  NAi21      o067(.An(j), .B(k), .Y(ori_ori_n96_));
  NO3        o068(.A(ori_ori_n96_), .B(ori_ori_n95_), .C(ori_ori_n94_), .Y(ori_ori_n97_));
  NAi31      o069(.An(j), .B(k), .C(h), .Y(ori_ori_n98_));
  NA2        o070(.A(ori_ori_n97_), .B(ori_ori_n93_), .Y(ori_ori_n99_));
  NO2        o071(.A(k), .B(j), .Y(ori_ori_n100_));
  NO2        o072(.A(ori_ori_n100_), .B(ori_ori_n95_), .Y(ori_ori_n101_));
  AN2        o073(.A(k), .B(j), .Y(ori_ori_n102_));
  NAi21      o074(.An(c), .B(b), .Y(ori_ori_n103_));
  NA2        o075(.A(f), .B(d), .Y(ori_ori_n104_));
  NO4        o076(.A(ori_ori_n104_), .B(ori_ori_n103_), .C(ori_ori_n102_), .D(ori_ori_n94_), .Y(ori_ori_n105_));
  NAi31      o077(.An(f), .B(e), .C(b), .Y(ori_ori_n106_));
  NA2        o078(.A(ori_ori_n105_), .B(ori_ori_n101_), .Y(ori_ori_n107_));
  NA2        o079(.A(d), .B(b), .Y(ori_ori_n108_));
  NAi21      o080(.An(e), .B(f), .Y(ori_ori_n109_));
  NAi21      o081(.An(e), .B(g), .Y(ori_ori_n110_));
  NAi21      o082(.An(c), .B(d), .Y(ori_ori_n111_));
  NAi31      o083(.An(l), .B(k), .C(h), .Y(ori_ori_n112_));
  NO2        o084(.A(ori_ori_n95_), .B(ori_ori_n112_), .Y(ori_ori_n113_));
  NAi31      o085(.An(ori_ori_n92_), .B(ori_ori_n107_), .C(ori_ori_n99_), .Y(ori_ori_n114_));
  NAi31      o086(.An(e), .B(f), .C(b), .Y(ori_ori_n115_));
  BUFFER     o087(.A(g), .Y(ori_ori_n116_));
  NO2        o088(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NOi21      o089(.An(h), .B(i), .Y(ori_ori_n118_));
  NOi21      o090(.An(k), .B(m), .Y(ori_ori_n119_));
  NA3        o091(.A(ori_ori_n119_), .B(ori_ori_n118_), .C(n), .Y(ori_ori_n120_));
  NOi21      o092(.An(ori_ori_n117_), .B(ori_ori_n120_), .Y(ori_ori_n121_));
  NOi21      o093(.An(h), .B(g), .Y(ori_ori_n122_));
  NOi32      o094(.An(n), .Bn(k), .C(m), .Y(ori_ori_n123_));
  INV        o095(.A(l), .Y(ori_ori_n124_));
  NAi31      o096(.An(d), .B(f), .C(c), .Y(ori_ori_n125_));
  NAi31      o097(.An(e), .B(f), .C(c), .Y(ori_ori_n126_));
  NA2        o098(.A(ori_ori_n126_), .B(ori_ori_n125_), .Y(ori_ori_n127_));
  NA2        o099(.A(j), .B(h), .Y(ori_ori_n128_));
  OR3        o100(.A(n), .B(m), .C(k), .Y(ori_ori_n129_));
  NO2        o101(.A(ori_ori_n129_), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  NAi32      o102(.An(m), .Bn(k), .C(n), .Y(ori_ori_n131_));
  NO2        o103(.A(ori_ori_n131_), .B(ori_ori_n128_), .Y(ori_ori_n132_));
  AOI220     o104(.A0(ori_ori_n132_), .A1(ori_ori_n117_), .B0(ori_ori_n130_), .B1(ori_ori_n127_), .Y(ori_ori_n133_));
  NO2        o105(.A(n), .B(m), .Y(ori_ori_n134_));
  NA2        o106(.A(ori_ori_n134_), .B(ori_ori_n41_), .Y(ori_ori_n135_));
  NAi21      o107(.An(f), .B(e), .Y(ori_ori_n136_));
  NA2        o108(.A(d), .B(c), .Y(ori_ori_n137_));
  NO2        o109(.A(ori_ori_n137_), .B(ori_ori_n136_), .Y(ori_ori_n138_));
  NOi21      o110(.An(ori_ori_n138_), .B(ori_ori_n135_), .Y(ori_ori_n139_));
  NAi31      o111(.An(m), .B(n), .C(b), .Y(ori_ori_n140_));
  NA2        o112(.A(k), .B(i), .Y(ori_ori_n141_));
  NAi21      o113(.An(h), .B(f), .Y(ori_ori_n142_));
  NO2        o114(.A(ori_ori_n142_), .B(ori_ori_n141_), .Y(ori_ori_n143_));
  NO2        o115(.A(ori_ori_n140_), .B(ori_ori_n111_), .Y(ori_ori_n144_));
  NA2        o116(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n145_));
  NOi32      o117(.An(f), .Bn(c), .C(d), .Y(ori_ori_n146_));
  NOi32      o118(.An(f), .Bn(c), .C(e), .Y(ori_ori_n147_));
  NO2        o119(.A(ori_ori_n147_), .B(ori_ori_n146_), .Y(ori_ori_n148_));
  NO3        o120(.A(n), .B(m), .C(j), .Y(ori_ori_n149_));
  NA2        o121(.A(ori_ori_n149_), .B(ori_ori_n86_), .Y(ori_ori_n150_));
  AO210      o122(.A0(ori_ori_n150_), .A1(ori_ori_n135_), .B0(ori_ori_n148_), .Y(ori_ori_n151_));
  NAi41      o123(.An(ori_ori_n139_), .B(ori_ori_n151_), .C(ori_ori_n145_), .D(ori_ori_n133_), .Y(ori_ori_n152_));
  OR3        o124(.A(ori_ori_n152_), .B(ori_ori_n121_), .C(ori_ori_n114_), .Y(ori_ori_n153_));
  NO3        o125(.A(ori_ori_n153_), .B(ori_ori_n79_), .C(ori_ori_n62_), .Y(ori_ori_n154_));
  NA3        o126(.A(m), .B(ori_ori_n84_), .C(j), .Y(ori_ori_n155_));
  NAi31      o127(.An(n), .B(h), .C(g), .Y(ori_ori_n156_));
  NO2        o128(.A(ori_ori_n156_), .B(ori_ori_n155_), .Y(ori_ori_n157_));
  NOi21      o129(.An(k), .B(j), .Y(ori_ori_n158_));
  NA4        o130(.A(ori_ori_n158_), .B(ori_ori_n85_), .C(i), .D(g), .Y(ori_ori_n159_));
  NAi41      o131(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n160_));
  INV        o132(.A(f), .Y(ori_ori_n161_));
  INV        o133(.A(g), .Y(ori_ori_n162_));
  NOi31      o134(.An(i), .B(j), .C(h), .Y(ori_ori_n163_));
  NOi21      o135(.An(l), .B(m), .Y(ori_ori_n164_));
  NA2        o136(.A(ori_ori_n164_), .B(ori_ori_n163_), .Y(ori_ori_n165_));
  NOi21      o137(.An(n), .B(m), .Y(ori_ori_n166_));
  OR2        o138(.A(ori_ori_n59_), .B(ori_ori_n58_), .Y(ori_ori_n167_));
  NAi21      o139(.An(j), .B(h), .Y(ori_ori_n168_));
  XN2        o140(.A(i), .B(h), .Y(ori_ori_n169_));
  NA2        o141(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  NOi31      o142(.An(k), .B(n), .C(m), .Y(ori_ori_n171_));
  NOi31      o143(.An(ori_ori_n171_), .B(ori_ori_n137_), .C(ori_ori_n136_), .Y(ori_ori_n172_));
  NA2        o144(.A(ori_ori_n172_), .B(ori_ori_n170_), .Y(ori_ori_n173_));
  NAi31      o145(.An(f), .B(e), .C(c), .Y(ori_ori_n174_));
  NO4        o146(.A(ori_ori_n174_), .B(ori_ori_n129_), .C(ori_ori_n128_), .D(ori_ori_n48_), .Y(ori_ori_n175_));
  NA3        o147(.A(e), .B(c), .C(b), .Y(ori_ori_n176_));
  NAi32      o148(.An(m), .Bn(i), .C(k), .Y(ori_ori_n177_));
  INV        o149(.A(k), .Y(ori_ori_n178_));
  INV        o150(.A(ori_ori_n175_), .Y(ori_ori_n179_));
  NAi21      o151(.An(n), .B(a), .Y(ori_ori_n180_));
  NO2        o152(.A(ori_ori_n180_), .B(ori_ori_n108_), .Y(ori_ori_n181_));
  NAi41      o153(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n182_));
  NO2        o154(.A(ori_ori_n182_), .B(e), .Y(ori_ori_n183_));
  NA2        o155(.A(ori_ori_n183_), .B(ori_ori_n181_), .Y(ori_ori_n184_));
  AN4        o156(.A(ori_ori_n184_), .B(ori_ori_n179_), .C(ori_ori_n173_), .D(ori_ori_n167_), .Y(ori_ori_n185_));
  OR2        o157(.A(h), .B(g), .Y(ori_ori_n186_));
  NO2        o158(.A(ori_ori_n186_), .B(ori_ori_n75_), .Y(ori_ori_n187_));
  NA2        o159(.A(ori_ori_n187_), .B(ori_ori_n93_), .Y(ori_ori_n188_));
  NA2        o160(.A(ori_ori_n119_), .B(ori_ori_n81_), .Y(ori_ori_n189_));
  NO2        o161(.A(n), .B(a), .Y(ori_ori_n190_));
  NAi31      o162(.An(ori_ori_n182_), .B(ori_ori_n190_), .C(ori_ori_n76_), .Y(ori_ori_n191_));
  NAi21      o163(.An(h), .B(i), .Y(ori_ori_n192_));
  NA2        o164(.A(ori_ori_n134_), .B(k), .Y(ori_ori_n193_));
  NO2        o165(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NA2        o166(.A(ori_ori_n194_), .B(ori_ori_n146_), .Y(ori_ori_n195_));
  NA3        o167(.A(ori_ori_n195_), .B(ori_ori_n191_), .C(ori_ori_n188_), .Y(ori_ori_n196_));
  NOi21      o168(.An(g), .B(e), .Y(ori_ori_n197_));
  NOi21      o169(.An(ori_ori_n185_), .B(ori_ori_n196_), .Y(ori_ori_n198_));
  INV        o170(.A(ori_ori_n157_), .Y(ori_ori_n199_));
  NO2        o171(.A(ori_ori_n199_), .B(ori_ori_n83_), .Y(ori_ori_n200_));
  NA3        o172(.A(ori_ori_n48_), .B(c), .C(b), .Y(ori_ori_n201_));
  NAi21      o173(.An(h), .B(g), .Y(ori_ori_n202_));
  NAi31      o174(.An(g), .B(k), .C(h), .Y(ori_ori_n203_));
  NA3        o175(.A(ori_ori_n119_), .B(ori_ori_n118_), .C(ori_ori_n63_), .Y(ori_ori_n204_));
  NO2        o176(.A(ori_ori_n204_), .B(ori_ori_n148_), .Y(ori_ori_n205_));
  NA3        o177(.A(e), .B(c), .C(b), .Y(ori_ori_n206_));
  NAi21      o178(.An(l), .B(k), .Y(ori_ori_n207_));
  NO2        o179(.A(ori_ori_n207_), .B(ori_ori_n40_), .Y(ori_ori_n208_));
  NAi32      o180(.An(j), .Bn(h), .C(i), .Y(ori_ori_n209_));
  NAi21      o181(.An(m), .B(l), .Y(ori_ori_n210_));
  NO3        o182(.A(ori_ori_n210_), .B(ori_ori_n209_), .C(ori_ori_n63_), .Y(ori_ori_n211_));
  NA2        o183(.A(h), .B(g), .Y(ori_ori_n212_));
  NO2        o184(.A(ori_ori_n106_), .B(d), .Y(ori_ori_n213_));
  NA2        o185(.A(ori_ori_n213_), .B(ori_ori_n44_), .Y(ori_ori_n214_));
  NO2        o186(.A(ori_ori_n78_), .B(ori_ori_n75_), .Y(ori_ori_n215_));
  NAi32      o187(.An(n), .Bn(m), .C(l), .Y(ori_ori_n216_));
  NO2        o188(.A(ori_ori_n216_), .B(ori_ori_n209_), .Y(ori_ori_n217_));
  NA2        o189(.A(ori_ori_n217_), .B(ori_ori_n138_), .Y(ori_ori_n218_));
  NA2        o190(.A(ori_ori_n218_), .B(ori_ori_n214_), .Y(ori_ori_n219_));
  NO3        o191(.A(ori_ori_n219_), .B(ori_ori_n205_), .C(ori_ori_n200_), .Y(ori_ori_n220_));
  NA2        o192(.A(ori_ori_n194_), .B(ori_ori_n147_), .Y(ori_ori_n221_));
  NAi21      o193(.An(m), .B(k), .Y(ori_ori_n222_));
  NO2        o194(.A(ori_ori_n169_), .B(ori_ori_n222_), .Y(ori_ori_n223_));
  NAi41      o195(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n224_));
  NO2        o196(.A(ori_ori_n224_), .B(ori_ori_n110_), .Y(ori_ori_n225_));
  NA2        o197(.A(ori_ori_n225_), .B(ori_ori_n223_), .Y(ori_ori_n226_));
  NA2        o198(.A(e), .B(c), .Y(ori_ori_n227_));
  NO3        o199(.A(ori_ori_n227_), .B(n), .C(d), .Y(ori_ori_n228_));
  NOi21      o200(.An(f), .B(h), .Y(ori_ori_n229_));
  NA2        o201(.A(ori_ori_n229_), .B(ori_ori_n88_), .Y(ori_ori_n230_));
  NO2        o202(.A(ori_ori_n230_), .B(ori_ori_n162_), .Y(ori_ori_n231_));
  NAi31      o203(.An(d), .B(e), .C(b), .Y(ori_ori_n232_));
  NO2        o204(.A(ori_ori_n95_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NA2        o205(.A(ori_ori_n233_), .B(ori_ori_n231_), .Y(ori_ori_n234_));
  NA3        o206(.A(ori_ori_n234_), .B(ori_ori_n226_), .C(ori_ori_n221_), .Y(ori_ori_n235_));
  NO4        o207(.A(ori_ori_n224_), .B(ori_ori_n59_), .C(ori_ori_n52_), .D(ori_ori_n162_), .Y(ori_ori_n236_));
  NA2        o208(.A(ori_ori_n190_), .B(ori_ori_n76_), .Y(ori_ori_n237_));
  NOi31      o209(.An(l), .B(n), .C(m), .Y(ori_ori_n238_));
  NA2        o210(.A(ori_ori_n238_), .B(ori_ori_n163_), .Y(ori_ori_n239_));
  NO2        o211(.A(ori_ori_n239_), .B(ori_ori_n148_), .Y(ori_ori_n240_));
  OR2        o212(.A(ori_ori_n240_), .B(ori_ori_n236_), .Y(ori_ori_n241_));
  NAi32      o213(.An(m), .Bn(j), .C(k), .Y(ori_ori_n242_));
  NAi41      o214(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n243_));
  NA2        o215(.A(ori_ori_n160_), .B(ori_ori_n243_), .Y(ori_ori_n244_));
  NOi31      o216(.An(j), .B(m), .C(k), .Y(ori_ori_n245_));
  NO2        o217(.A(ori_ori_n89_), .B(ori_ori_n245_), .Y(ori_ori_n246_));
  AN3        o218(.A(h), .B(g), .C(f), .Y(ori_ori_n247_));
  NAi31      o219(.An(ori_ori_n246_), .B(ori_ori_n247_), .C(ori_ori_n244_), .Y(ori_ori_n248_));
  NOi32      o220(.An(m), .Bn(j), .C(l), .Y(ori_ori_n249_));
  NO2        o221(.A(ori_ori_n210_), .B(ori_ori_n209_), .Y(ori_ori_n250_));
  INV        o222(.A(ori_ori_n248_), .Y(ori_ori_n251_));
  NA3        o223(.A(h), .B(g), .C(f), .Y(ori_ori_n252_));
  NO2        o224(.A(ori_ori_n252_), .B(ori_ori_n55_), .Y(ori_ori_n253_));
  NA2        o225(.A(ori_ori_n243_), .B(ori_ori_n160_), .Y(ori_ori_n254_));
  NA2        o226(.A(ori_ori_n122_), .B(e), .Y(ori_ori_n255_));
  NA2        o227(.A(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n256_));
  NOi32      o228(.An(j), .Bn(g), .C(i), .Y(ori_ori_n257_));
  NA3        o229(.A(ori_ori_n257_), .B(ori_ori_n207_), .C(ori_ori_n85_), .Y(ori_ori_n258_));
  OR2        o230(.A(ori_ori_n83_), .B(ori_ori_n258_), .Y(ori_ori_n259_));
  NOi32      o231(.An(e), .Bn(b), .C(a), .Y(ori_ori_n260_));
  AN2        o232(.A(l), .B(j), .Y(ori_ori_n261_));
  NO2        o233(.A(ori_ori_n222_), .B(ori_ori_n261_), .Y(ori_ori_n262_));
  NO3        o234(.A(ori_ori_n224_), .B(ori_ori_n52_), .C(ori_ori_n162_), .Y(ori_ori_n263_));
  NA2        o235(.A(ori_ori_n159_), .B(ori_ori_n32_), .Y(ori_ori_n264_));
  AOI220     o236(.A0(ori_ori_n264_), .A1(ori_ori_n260_), .B0(ori_ori_n263_), .B1(ori_ori_n262_), .Y(ori_ori_n265_));
  NA2        o237(.A(ori_ori_n42_), .B(ori_ori_n85_), .Y(ori_ori_n266_));
  NA3        o238(.A(ori_ori_n265_), .B(ori_ori_n259_), .C(ori_ori_n256_), .Y(ori_ori_n267_));
  NO4        o239(.A(ori_ori_n267_), .B(ori_ori_n251_), .C(ori_ori_n241_), .D(ori_ori_n235_), .Y(ori_ori_n268_));
  NA4        o240(.A(ori_ori_n268_), .B(ori_ori_n220_), .C(ori_ori_n198_), .D(ori_ori_n154_), .Y(ori10));
  NA3        o241(.A(m), .B(k), .C(i), .Y(ori_ori_n270_));
  NOi21      o242(.An(e), .B(f), .Y(ori_ori_n271_));
  NO3        o243(.A(ori_ori_n111_), .B(n), .C(ori_ori_n82_), .Y(ori_ori_n272_));
  NAi31      o244(.An(b), .B(f), .C(c), .Y(ori_ori_n273_));
  INV        o245(.A(ori_ori_n273_), .Y(ori_ori_n274_));
  NOi32      o246(.An(k), .Bn(h), .C(j), .Y(ori_ori_n275_));
  NA2        o247(.A(ori_ori_n275_), .B(ori_ori_n166_), .Y(ori_ori_n276_));
  NA2        o248(.A(ori_ori_n120_), .B(ori_ori_n276_), .Y(ori_ori_n277_));
  NA2        o249(.A(ori_ori_n277_), .B(ori_ori_n274_), .Y(ori_ori_n278_));
  AN2        o250(.A(j), .B(h), .Y(ori_ori_n279_));
  NO3        o251(.A(n), .B(m), .C(k), .Y(ori_ori_n280_));
  NA2        o252(.A(ori_ori_n280_), .B(ori_ori_n279_), .Y(ori_ori_n281_));
  NO3        o253(.A(ori_ori_n281_), .B(ori_ori_n111_), .C(ori_ori_n161_), .Y(ori_ori_n282_));
  OR2        o254(.A(m), .B(k), .Y(ori_ori_n283_));
  NO2        o255(.A(ori_ori_n128_), .B(ori_ori_n283_), .Y(ori_ori_n284_));
  NA4        o256(.A(n), .B(f), .C(c), .D(ori_ori_n87_), .Y(ori_ori_n285_));
  NOi21      o257(.An(ori_ori_n284_), .B(ori_ori_n285_), .Y(ori_ori_n286_));
  NOi32      o258(.An(d), .Bn(a), .C(c), .Y(ori_ori_n287_));
  NA2        o259(.A(ori_ori_n287_), .B(ori_ori_n136_), .Y(ori_ori_n288_));
  NO2        o260(.A(ori_ori_n286_), .B(ori_ori_n282_), .Y(ori_ori_n289_));
  NO2        o261(.A(ori_ori_n285_), .B(ori_ori_n210_), .Y(ori_ori_n290_));
  NOi32      o262(.An(f), .Bn(d), .C(c), .Y(ori_ori_n291_));
  AOI220     o263(.A0(ori_ori_n291_), .A1(ori_ori_n217_), .B0(ori_ori_n290_), .B1(ori_ori_n163_), .Y(ori_ori_n292_));
  NA3        o264(.A(ori_ori_n292_), .B(ori_ori_n289_), .C(ori_ori_n278_), .Y(ori_ori_n293_));
  NO2        o265(.A(ori_ori_n48_), .B(ori_ori_n87_), .Y(ori_ori_n294_));
  NA2        o266(.A(ori_ori_n190_), .B(ori_ori_n294_), .Y(ori_ori_n295_));
  INV        o267(.A(e), .Y(ori_ori_n296_));
  NA2        o268(.A(ori_ori_n39_), .B(e), .Y(ori_ori_n297_));
  NO2        o269(.A(ori_ori_n297_), .B(ori_ori_n155_), .Y(ori_ori_n298_));
  NO2        o270(.A(ori_ori_n67_), .B(ori_ori_n296_), .Y(ori_ori_n299_));
  NO2        o271(.A(ori_ori_n74_), .B(ori_ori_n296_), .Y(ori_ori_n300_));
  NO3        o272(.A(ori_ori_n300_), .B(ori_ori_n299_), .C(ori_ori_n298_), .Y(ori_ori_n301_));
  NOi21      o273(.An(g), .B(h), .Y(ori_ori_n302_));
  AN3        o274(.A(m), .B(l), .C(i), .Y(ori_ori_n303_));
  NA3        o275(.A(ori_ori_n303_), .B(ori_ori_n302_), .C(e), .Y(ori_ori_n304_));
  AN3        o276(.A(h), .B(g), .C(e), .Y(ori_ori_n305_));
  AOI210     o277(.A0(ori_ori_n304_), .A1(ori_ori_n301_), .B0(ori_ori_n295_), .Y(ori_ori_n306_));
  NO2        o278(.A(ori_ori_n306_), .B(ori_ori_n293_), .Y(ori_ori_n307_));
  NOi21      o279(.An(d), .B(c), .Y(ori_ori_n308_));
  OR2        o280(.A(n), .B(m), .Y(ori_ori_n309_));
  NO2        o281(.A(ori_ori_n309_), .B(ori_ori_n112_), .Y(ori_ori_n310_));
  NO2        o282(.A(ori_ori_n137_), .B(ori_ori_n109_), .Y(ori_ori_n311_));
  OAI210     o283(.A0(ori_ori_n310_), .A1(ori_ori_n130_), .B0(ori_ori_n311_), .Y(ori_ori_n312_));
  INV        o284(.A(ori_ori_n266_), .Y(ori_ori_n313_));
  NA3        o285(.A(ori_ori_n313_), .B(ori_ori_n260_), .C(d), .Y(ori_ori_n314_));
  NAi21      o286(.An(k), .B(j), .Y(ori_ori_n315_));
  NAi21      o287(.An(e), .B(d), .Y(ori_ori_n316_));
  INV        o288(.A(ori_ori_n316_), .Y(ori_ori_n317_));
  NO2        o289(.A(ori_ori_n193_), .B(ori_ori_n161_), .Y(ori_ori_n318_));
  NA3        o290(.A(ori_ori_n318_), .B(ori_ori_n317_), .C(ori_ori_n170_), .Y(ori_ori_n319_));
  NA3        o291(.A(ori_ori_n319_), .B(ori_ori_n314_), .C(ori_ori_n312_), .Y(ori_ori_n320_));
  NO2        o292(.A(ori_ori_n239_), .B(ori_ori_n161_), .Y(ori_ori_n321_));
  NA2        o293(.A(ori_ori_n321_), .B(ori_ori_n317_), .Y(ori_ori_n322_));
  NOi31      o294(.An(n), .B(m), .C(k), .Y(ori_ori_n323_));
  AOI220     o295(.A0(ori_ori_n323_), .A1(ori_ori_n279_), .B0(ori_ori_n166_), .B1(ori_ori_n41_), .Y(ori_ori_n324_));
  NAi31      o296(.An(g), .B(f), .C(c), .Y(ori_ori_n325_));
  OR3        o297(.A(ori_ori_n325_), .B(ori_ori_n324_), .C(e), .Y(ori_ori_n326_));
  NA3        o298(.A(ori_ori_n326_), .B(ori_ori_n322_), .C(ori_ori_n218_), .Y(ori_ori_n327_));
  NO2        o299(.A(ori_ori_n327_), .B(ori_ori_n320_), .Y(ori_ori_n328_));
  INV        o300(.A(ori_ori_n203_), .Y(ori_ori_n329_));
  AN2        o301(.A(e), .B(d), .Y(ori_ori_n330_));
  NO2        o302(.A(ori_ori_n50_), .B(e), .Y(ori_ori_n331_));
  NO4        o303(.A(ori_ori_n142_), .B(ori_ori_n75_), .C(ori_ori_n45_), .D(b), .Y(ori_ori_n332_));
  NA2        o304(.A(ori_ori_n274_), .B(ori_ori_n113_), .Y(ori_ori_n333_));
  OR2        o305(.A(k), .B(j), .Y(ori_ori_n334_));
  NA2        o306(.A(l), .B(k), .Y(ori_ori_n335_));
  NA3        o307(.A(ori_ori_n335_), .B(ori_ori_n334_), .C(ori_ori_n166_), .Y(ori_ori_n336_));
  AOI210     o308(.A0(ori_ori_n177_), .A1(ori_ori_n242_), .B0(ori_ori_n63_), .Y(ori_ori_n337_));
  NOi21      o309(.An(ori_ori_n336_), .B(ori_ori_n337_), .Y(ori_ori_n338_));
  INV        o310(.A(ori_ori_n90_), .Y(ori_ori_n339_));
  NA2        o311(.A(ori_ori_n90_), .B(ori_ori_n333_), .Y(ori_ori_n340_));
  NO2        o312(.A(ori_ori_n340_), .B(ori_ori_n332_), .Y(ori_ori_n341_));
  INV        o313(.A(e), .Y(ori_ori_n342_));
  NO2        o314(.A(ori_ori_n142_), .B(ori_ori_n45_), .Y(ori_ori_n343_));
  INV        o315(.A(ori_ori_n75_), .Y(ori_ori_n344_));
  NA3        o316(.A(ori_ori_n344_), .B(ori_ori_n343_), .C(ori_ori_n342_), .Y(ori_ori_n345_));
  NO2        o317(.A(ori_ori_n288_), .B(ori_ori_n266_), .Y(ori_ori_n346_));
  NO3        o318(.A(ori_ori_n346_), .B(ori_ori_n139_), .C(ori_ori_n215_), .Y(ori_ori_n347_));
  NA3        o319(.A(ori_ori_n347_), .B(ori_ori_n345_), .C(ori_ori_n185_), .Y(ori_ori_n348_));
  OAI210     o320(.A0(ori_ori_n91_), .A1(ori_ori_n89_), .B0(n), .Y(ori_ori_n349_));
  NO2        o321(.A(ori_ori_n349_), .B(ori_ori_n94_), .Y(ori_ori_n350_));
  AN2        o322(.A(ori_ori_n350_), .B(ori_ori_n147_), .Y(ori_ori_n351_));
  XO2        o323(.A(i), .B(h), .Y(ori_ori_n352_));
  NA3        o324(.A(ori_ori_n352_), .B(ori_ori_n119_), .C(n), .Y(ori_ori_n353_));
  NAi41      o325(.An(ori_ori_n211_), .B(ori_ori_n353_), .C(ori_ori_n324_), .D(ori_ori_n276_), .Y(ori_ori_n354_));
  NOi32      o326(.An(ori_ori_n354_), .Bn(ori_ori_n331_), .C(ori_ori_n201_), .Y(ori_ori_n355_));
  NAi31      o327(.An(c), .B(f), .C(d), .Y(ori_ori_n356_));
  AOI210     o328(.A0(ori_ori_n204_), .A1(ori_ori_n150_), .B0(ori_ori_n356_), .Y(ori_ori_n357_));
  NOi21      o329(.An(ori_ori_n61_), .B(ori_ori_n357_), .Y(ori_ori_n358_));
  NA2        o330(.A(ori_ori_n171_), .B(ori_ori_n81_), .Y(ori_ori_n359_));
  AOI210     o331(.A0(ori_ori_n359_), .A1(ori_ori_n135_), .B0(ori_ori_n356_), .Y(ori_ori_n360_));
  INV        o332(.A(ori_ori_n360_), .Y(ori_ori_n361_));
  NA2        o333(.A(ori_ori_n361_), .B(ori_ori_n358_), .Y(ori_ori_n362_));
  NO4        o334(.A(ori_ori_n362_), .B(ori_ori_n355_), .C(ori_ori_n351_), .D(ori_ori_n348_), .Y(ori_ori_n363_));
  NA4        o335(.A(ori_ori_n363_), .B(ori_ori_n341_), .C(ori_ori_n328_), .D(ori_ori_n307_), .Y(ori11));
  NA2        o336(.A(j), .B(g), .Y(ori_ori_n365_));
  NAi31      o337(.An(i), .B(m), .C(l), .Y(ori_ori_n366_));
  NA3        o338(.A(m), .B(k), .C(j), .Y(ori_ori_n367_));
  NOi32      o339(.An(e), .Bn(b), .C(f), .Y(ori_ori_n368_));
  NA2        o340(.A(ori_ori_n39_), .B(j), .Y(ori_ori_n369_));
  NAi31      o341(.An(d), .B(e), .C(a), .Y(ori_ori_n370_));
  NA2        o342(.A(j), .B(i), .Y(ori_ori_n371_));
  NAi31      o343(.An(n), .B(m), .C(k), .Y(ori_ori_n372_));
  NO3        o344(.A(ori_ori_n372_), .B(ori_ori_n371_), .C(ori_ori_n84_), .Y(ori_ori_n373_));
  NO2        o345(.A(ori_ori_n203_), .B(ori_ori_n40_), .Y(ori_ori_n374_));
  NA2        o346(.A(ori_ori_n102_), .B(ori_ori_n31_), .Y(ori_ori_n375_));
  OAI220     o347(.A0(ori_ori_n375_), .A1(m), .B0(ori_ori_n369_), .B1(ori_ori_n177_), .Y(ori_ori_n376_));
  NOi41      o348(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n377_));
  NAi32      o349(.An(e), .Bn(b), .C(c), .Y(ori_ori_n378_));
  OR2        o350(.A(ori_ori_n378_), .B(ori_ori_n63_), .Y(ori_ori_n379_));
  AN2        o351(.A(ori_ori_n243_), .B(ori_ori_n224_), .Y(ori_ori_n380_));
  NA2        o352(.A(ori_ori_n380_), .B(ori_ori_n379_), .Y(ori_ori_n381_));
  OA210      o353(.A0(ori_ori_n381_), .A1(ori_ori_n377_), .B0(ori_ori_n376_), .Y(ori_ori_n382_));
  NO2        o354(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n383_));
  NA2        o355(.A(ori_ori_n383_), .B(f), .Y(ori_ori_n384_));
  NO3        o356(.A(ori_ori_n131_), .B(ori_ori_n128_), .C(g), .Y(ori_ori_n385_));
  NA2        o357(.A(ori_ori_n385_), .B(ori_ori_n47_), .Y(ori_ori_n386_));
  INV        o358(.A(ori_ori_n386_), .Y(ori_ori_n387_));
  AN3        o359(.A(j), .B(h), .C(g), .Y(ori_ori_n388_));
  NO2        o360(.A(ori_ori_n108_), .B(c), .Y(ori_ori_n389_));
  NA3        o361(.A(ori_ori_n389_), .B(ori_ori_n388_), .C(ori_ori_n323_), .Y(ori_ori_n390_));
  NA3        o362(.A(f), .B(d), .C(b), .Y(ori_ori_n391_));
  NO4        o363(.A(ori_ori_n391_), .B(ori_ori_n131_), .C(ori_ori_n128_), .D(g), .Y(ori_ori_n392_));
  NAi21      o364(.An(ori_ori_n392_), .B(ori_ori_n390_), .Y(ori_ori_n393_));
  NO3        o365(.A(ori_ori_n393_), .B(ori_ori_n387_), .C(ori_ori_n382_), .Y(ori_ori_n394_));
  INV        o366(.A(k), .Y(ori_ori_n395_));
  NAi41      o367(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n396_));
  OAI210     o368(.A0(ori_ori_n370_), .A1(n), .B0(ori_ori_n396_), .Y(ori_ori_n397_));
  NAi31      o369(.An(h), .B(g), .C(f), .Y(ori_ori_n398_));
  NAi31      o370(.An(f), .B(h), .C(g), .Y(ori_ori_n399_));
  NOi32      o371(.An(d), .Bn(a), .C(e), .Y(ori_ori_n400_));
  NOi32      o372(.An(e), .Bn(a), .C(d), .Y(ori_ori_n401_));
  INV        o373(.A(ori_ori_n401_), .Y(ori_ori_n402_));
  NO3        o374(.A(ori_ori_n222_), .B(ori_ori_n49_), .C(n), .Y(ori_ori_n403_));
  NA3        o375(.A(ori_ori_n356_), .B(ori_ori_n126_), .C(ori_ori_n125_), .Y(ori_ori_n404_));
  NA2        o376(.A(ori_ori_n325_), .B(ori_ori_n174_), .Y(ori_ori_n405_));
  OR2        o377(.A(ori_ori_n405_), .B(ori_ori_n404_), .Y(ori_ori_n406_));
  NA2        o378(.A(ori_ori_n406_), .B(ori_ori_n403_), .Y(ori_ori_n407_));
  NO2        o379(.A(ori_ori_n407_), .B(ori_ori_n65_), .Y(ori_ori_n408_));
  NA3        o380(.A(ori_ori_n377_), .B(ori_ori_n245_), .C(ori_ori_n39_), .Y(ori_ori_n409_));
  NOi32      o381(.An(e), .Bn(c), .C(f), .Y(ori_ori_n410_));
  NOi21      o382(.An(f), .B(g), .Y(ori_ori_n411_));
  NO2        o383(.A(ori_ori_n411_), .B(ori_ori_n160_), .Y(ori_ori_n412_));
  AOI220     o384(.A0(ori_ori_n412_), .A1(ori_ori_n284_), .B0(ori_ori_n410_), .B1(ori_ori_n130_), .Y(ori_ori_n413_));
  NA3        o385(.A(ori_ori_n413_), .B(ori_ori_n409_), .C(ori_ori_n133_), .Y(ori_ori_n414_));
  NA2        o386(.A(ori_ori_n81_), .B(ori_ori_n33_), .Y(ori_ori_n415_));
  NO2        o387(.A(k), .B(ori_ori_n162_), .Y(ori_ori_n416_));
  INV        o388(.A(ori_ori_n260_), .Y(ori_ori_n417_));
  NO2        o389(.A(ori_ori_n417_), .B(n), .Y(ori_ori_n418_));
  NAi31      o390(.An(ori_ori_n415_), .B(ori_ori_n418_), .C(ori_ori_n416_), .Y(ori_ori_n419_));
  NO2        o391(.A(ori_ori_n369_), .B(ori_ori_n131_), .Y(ori_ori_n420_));
  NA3        o392(.A(ori_ori_n378_), .B(ori_ori_n201_), .C(ori_ori_n106_), .Y(ori_ori_n421_));
  NA2        o393(.A(ori_ori_n352_), .B(ori_ori_n119_), .Y(ori_ori_n422_));
  NO3        o394(.A(ori_ori_n285_), .B(ori_ori_n422_), .C(ori_ori_n65_), .Y(ori_ori_n423_));
  AOI210     o395(.A0(ori_ori_n421_), .A1(ori_ori_n420_), .B0(ori_ori_n423_), .Y(ori_ori_n424_));
  AN3        o396(.A(f), .B(d), .C(b), .Y(ori_ori_n425_));
  OAI210     o397(.A0(ori_ori_n425_), .A1(ori_ori_n93_), .B0(n), .Y(ori_ori_n426_));
  NA3        o398(.A(ori_ori_n352_), .B(ori_ori_n119_), .C(ori_ori_n162_), .Y(ori_ori_n427_));
  AOI210     o399(.A0(ori_ori_n426_), .A1(ori_ori_n176_), .B0(ori_ori_n427_), .Y(ori_ori_n428_));
  NAi31      o400(.An(m), .B(n), .C(k), .Y(ori_ori_n429_));
  INV        o401(.A(ori_ori_n191_), .Y(ori_ori_n430_));
  OAI210     o402(.A0(ori_ori_n430_), .A1(ori_ori_n428_), .B0(j), .Y(ori_ori_n431_));
  NA3        o403(.A(ori_ori_n431_), .B(ori_ori_n424_), .C(ori_ori_n419_), .Y(ori_ori_n432_));
  NO3        o404(.A(ori_ori_n432_), .B(ori_ori_n414_), .C(ori_ori_n408_), .Y(ori_ori_n433_));
  NA2        o405(.A(ori_ori_n272_), .B(ori_ori_n122_), .Y(ori_ori_n434_));
  NAi31      o406(.An(g), .B(h), .C(f), .Y(ori_ori_n435_));
  OA210      o407(.A0(ori_ori_n370_), .A1(n), .B0(ori_ori_n396_), .Y(ori_ori_n436_));
  NO2        o408(.A(ori_ori_n436_), .B(ori_ori_n68_), .Y(ori_ori_n437_));
  INV        o409(.A(ori_ori_n437_), .Y(ori_ori_n438_));
  AOI210     o410(.A0(ori_ori_n438_), .A1(ori_ori_n434_), .B0(ori_ori_n367_), .Y(ori_ori_n439_));
  NO3        o411(.A(g), .B(ori_ori_n161_), .C(ori_ori_n45_), .Y(ori_ori_n440_));
  NO2        o412(.A(ori_ori_n359_), .B(ori_ori_n65_), .Y(ori_ori_n441_));
  OAI210     o413(.A0(ori_ori_n441_), .A1(ori_ori_n284_), .B0(ori_ori_n440_), .Y(ori_ori_n442_));
  AN2        o414(.A(h), .B(f), .Y(ori_ori_n443_));
  NA2        o415(.A(ori_ori_n443_), .B(ori_ori_n34_), .Y(ori_ori_n444_));
  NA2        o416(.A(ori_ori_n73_), .B(ori_ori_n39_), .Y(ori_ori_n445_));
  NO2        o417(.A(ori_ori_n445_), .B(ori_ori_n237_), .Y(ori_ori_n446_));
  INV        o418(.A(ori_ori_n446_), .Y(ori_ori_n447_));
  NA2        o419(.A(ori_ori_n447_), .B(ori_ori_n442_), .Y(ori_ori_n448_));
  NO2        o420(.A(ori_ori_n411_), .B(ori_ori_n49_), .Y(ori_ori_n449_));
  NO2        o421(.A(ori_ori_n449_), .B(ori_ori_n31_), .Y(ori_ori_n450_));
  NA2        o422(.A(ori_ori_n233_), .B(ori_ori_n102_), .Y(ori_ori_n451_));
  NA2        o423(.A(ori_ori_n95_), .B(ori_ori_n40_), .Y(ori_ori_n452_));
  NA2        o424(.A(ori_ori_n260_), .B(ori_ori_n85_), .Y(ori_ori_n453_));
  OA220      o425(.A0(ori_ori_n453_), .A1(ori_ori_n375_), .B0(ori_ori_n258_), .B1(ori_ori_n83_), .Y(ori_ori_n454_));
  OAI210     o426(.A0(ori_ori_n451_), .A1(ori_ori_n450_), .B0(ori_ori_n454_), .Y(ori_ori_n455_));
  NO3        o427(.A(ori_ori_n291_), .B(ori_ori_n147_), .C(ori_ori_n146_), .Y(ori_ori_n456_));
  NA2        o428(.A(ori_ori_n456_), .B(ori_ori_n174_), .Y(ori_ori_n457_));
  NA3        o429(.A(ori_ori_n457_), .B(ori_ori_n194_), .C(j), .Y(ori_ori_n458_));
  NO3        o430(.A(ori_ori_n325_), .B(ori_ori_n128_), .C(i), .Y(ori_ori_n459_));
  NA2        o431(.A(ori_ori_n458_), .B(ori_ori_n289_), .Y(ori_ori_n460_));
  NO4        o432(.A(ori_ori_n460_), .B(ori_ori_n455_), .C(ori_ori_n448_), .D(ori_ori_n439_), .Y(ori_ori_n461_));
  NA3        o433(.A(ori_ori_n461_), .B(ori_ori_n433_), .C(ori_ori_n394_), .Y(ori08));
  NO2        o434(.A(k), .B(h), .Y(ori_ori_n463_));
  AO210      o435(.A0(ori_ori_n192_), .A1(ori_ori_n315_), .B0(ori_ori_n463_), .Y(ori_ori_n464_));
  NO2        o436(.A(ori_ori_n464_), .B(ori_ori_n210_), .Y(ori_ori_n465_));
  NA2        o437(.A(ori_ori_n410_), .B(ori_ori_n63_), .Y(ori_ori_n466_));
  NA2        o438(.A(ori_ori_n466_), .B(ori_ori_n325_), .Y(ori_ori_n467_));
  NA2        o439(.A(ori_ori_n467_), .B(ori_ori_n465_), .Y(ori_ori_n468_));
  NA2        o440(.A(ori_ori_n63_), .B(ori_ori_n82_), .Y(ori_ori_n469_));
  NO2        o441(.A(ori_ori_n469_), .B(ori_ori_n46_), .Y(ori_ori_n470_));
  NO4        o442(.A(ori_ori_n270_), .B(ori_ori_n84_), .C(j), .D(ori_ori_n162_), .Y(ori_ori_n471_));
  NA2        o443(.A(ori_ori_n391_), .B(ori_ori_n176_), .Y(ori_ori_n472_));
  NA2        o444(.A(ori_ori_n471_), .B(ori_ori_n470_), .Y(ori_ori_n473_));
  AOI210     o445(.A0(ori_ori_n391_), .A1(ori_ori_n115_), .B0(ori_ori_n63_), .Y(ori_ori_n474_));
  NA4        o446(.A(ori_ori_n164_), .B(ori_ori_n102_), .C(ori_ori_n38_), .D(h), .Y(ori_ori_n475_));
  AN2        o447(.A(l), .B(k), .Y(ori_ori_n476_));
  NA4        o448(.A(ori_ori_n476_), .B(ori_ori_n81_), .C(ori_ori_n53_), .D(ori_ori_n162_), .Y(ori_ori_n477_));
  OAI210     o449(.A0(ori_ori_n475_), .A1(g), .B0(ori_ori_n477_), .Y(ori_ori_n478_));
  NA2        o450(.A(ori_ori_n478_), .B(ori_ori_n474_), .Y(ori_ori_n479_));
  NA3        o451(.A(ori_ori_n479_), .B(ori_ori_n473_), .C(ori_ori_n468_), .Y(ori_ori_n480_));
  NO4        o452(.A(ori_ori_n128_), .B(ori_ori_n283_), .C(ori_ori_n84_), .D(g), .Y(ori_ori_n481_));
  NA2        o453(.A(ori_ori_n481_), .B(ori_ori_n472_), .Y(ori_ori_n482_));
  NA2        o454(.A(ori_ori_n412_), .B(ori_ori_n250_), .Y(ori_ori_n483_));
  NA2        o455(.A(ori_ori_n483_), .B(ori_ori_n482_), .Y(ori_ori_n484_));
  NO3        o456(.A(ori_ori_n222_), .B(ori_ori_n94_), .C(ori_ori_n37_), .Y(ori_ori_n485_));
  NAi21      o457(.An(ori_ori_n485_), .B(ori_ori_n477_), .Y(ori_ori_n486_));
  NA2        o458(.A(ori_ori_n464_), .B(ori_ori_n98_), .Y(ori_ori_n487_));
  AOI220     o459(.A0(ori_ori_n487_), .A1(ori_ori_n290_), .B0(ori_ori_n486_), .B1(ori_ori_n56_), .Y(ori_ori_n488_));
  INV        o460(.A(ori_ori_n488_), .Y(ori_ori_n489_));
  NA3        o461(.A(ori_ori_n457_), .B(ori_ori_n238_), .C(ori_ori_n275_), .Y(ori_ori_n490_));
  NA3        o462(.A(m), .B(l), .C(k), .Y(ori_ori_n491_));
  INV        o463(.A(ori_ori_n490_), .Y(ori_ori_n492_));
  NO4        o464(.A(ori_ori_n492_), .B(ori_ori_n489_), .C(ori_ori_n484_), .D(ori_ori_n480_), .Y(ori_ori_n493_));
  NA2        o465(.A(ori_ori_n412_), .B(ori_ori_n284_), .Y(ori_ori_n494_));
  INV        o466(.A(ori_ori_n346_), .Y(ori_ori_n495_));
  NA3        o467(.A(ori_ori_n495_), .B(ori_ori_n494_), .C(ori_ori_n191_), .Y(ori_ori_n496_));
  NA2        o468(.A(ori_ori_n476_), .B(ori_ori_n53_), .Y(ori_ori_n497_));
  NO4        o469(.A(ori_ori_n456_), .B(ori_ori_n128_), .C(n), .D(i), .Y(ori_ori_n498_));
  NOi21      o470(.An(h), .B(j), .Y(ori_ori_n499_));
  NO2        o471(.A(ori_ori_n498_), .B(ori_ori_n459_), .Y(ori_ori_n500_));
  NO2        o472(.A(ori_ori_n500_), .B(ori_ori_n497_), .Y(ori_ori_n501_));
  AOI210     o473(.A0(ori_ori_n496_), .A1(l), .B0(ori_ori_n501_), .Y(ori_ori_n502_));
  NO2        o474(.A(j), .B(i), .Y(ori_ori_n503_));
  NA2        o475(.A(ori_ori_n503_), .B(ori_ori_n30_), .Y(ori_ori_n504_));
  INV        o476(.A(j), .Y(ori_ori_n505_));
  NO3        o477(.A(ori_ori_n210_), .B(ori_ori_n505_), .C(ori_ori_n36_), .Y(ori_ori_n506_));
  AOI210     o478(.A0(ori_ori_n368_), .A1(n), .B0(ori_ori_n377_), .Y(ori_ori_n507_));
  NA2        o479(.A(ori_ori_n507_), .B(ori_ori_n380_), .Y(ori_ori_n508_));
  AN3        o480(.A(ori_ori_n508_), .B(ori_ori_n506_), .C(ori_ori_n72_), .Y(ori_ori_n509_));
  NA2        o481(.A(ori_ori_n405_), .B(ori_ori_n217_), .Y(ori_ori_n510_));
  INV        o482(.A(ori_ori_n510_), .Y(ori_ori_n511_));
  NO2        o483(.A(ori_ori_n210_), .B(ori_ori_n98_), .Y(ori_ori_n512_));
  AOI220     o484(.A0(ori_ori_n512_), .A1(ori_ori_n412_), .B0(ori_ori_n485_), .B1(ori_ori_n474_), .Y(ori_ori_n513_));
  NO2        o485(.A(ori_ori_n491_), .B(ori_ori_n68_), .Y(ori_ori_n514_));
  NA2        o486(.A(ori_ori_n514_), .B(ori_ori_n397_), .Y(ori_ori_n515_));
  NA2        o487(.A(ori_ori_n515_), .B(ori_ori_n513_), .Y(ori_ori_n516_));
  OR3        o488(.A(ori_ori_n516_), .B(ori_ori_n511_), .C(ori_ori_n509_), .Y(ori_ori_n517_));
  NA3        o489(.A(ori_ori_n507_), .B(ori_ori_n380_), .C(ori_ori_n379_), .Y(ori_ori_n518_));
  NA4        o490(.A(ori_ori_n518_), .B(ori_ori_n164_), .C(ori_ori_n315_), .D(ori_ori_n31_), .Y(ori_ori_n519_));
  OAI220     o491(.A0(ori_ori_n475_), .A1(ori_ori_n466_), .B0(ori_ori_n237_), .B1(ori_ori_n35_), .Y(ori_ori_n520_));
  INV        o492(.A(ori_ori_n520_), .Y(ori_ori_n521_));
  NA2        o493(.A(ori_ori_n521_), .B(ori_ori_n519_), .Y(ori_ori_n522_));
  NO3        o494(.A(ori_ori_n240_), .B(ori_ori_n522_), .C(ori_ori_n517_), .Y(ori_ori_n523_));
  NO3        o495(.A(ori_ori_n246_), .B(ori_ori_n212_), .C(ori_ori_n84_), .Y(ori_ori_n524_));
  NA2        o496(.A(ori_ori_n524_), .B(ori_ori_n508_), .Y(ori_ori_n525_));
  NO3        o497(.A(ori_ori_n365_), .B(ori_ori_n69_), .C(h), .Y(ori_ori_n526_));
  NA2        o498(.A(ori_ori_n526_), .B(ori_ori_n470_), .Y(ori_ori_n527_));
  NA3        o499(.A(ori_ori_n527_), .B(ori_ori_n525_), .C(ori_ori_n292_), .Y(ori_ori_n528_));
  INV        o500(.A(ori_ori_n400_), .Y(ori_ori_n529_));
  NO2        o501(.A(ori_ori_n378_), .B(ori_ori_n63_), .Y(ori_ori_n530_));
  NA2        o502(.A(ori_ori_n524_), .B(ori_ori_n530_), .Y(ori_ori_n531_));
  OAI210     o503(.A0(ori_ori_n475_), .A1(ori_ori_n285_), .B0(ori_ori_n531_), .Y(ori_ori_n532_));
  NO2        o504(.A(ori_ori_n456_), .B(n), .Y(ori_ori_n533_));
  BUFFER     o505(.A(ori_ori_n512_), .Y(ori_ori_n534_));
  AOI220     o506(.A0(ori_ori_n534_), .A1(ori_ori_n440_), .B0(ori_ori_n533_), .B1(ori_ori_n465_), .Y(ori_ori_n535_));
  INV        o507(.A(ori_ori_n535_), .Y(ori_ori_n536_));
  NO3        o508(.A(ori_ori_n536_), .B(ori_ori_n532_), .C(ori_ori_n528_), .Y(ori_ori_n537_));
  NA4        o509(.A(ori_ori_n537_), .B(ori_ori_n523_), .C(ori_ori_n502_), .D(ori_ori_n493_), .Y(ori09));
  NA2        o510(.A(ori_ori_n310_), .B(e), .Y(ori_ori_n539_));
  NO2        o511(.A(ori_ori_n539_), .B(ori_ori_n356_), .Y(ori_ori_n540_));
  INV        o512(.A(ori_ori_n540_), .Y(ori_ori_n541_));
  NA3        o513(.A(m), .B(l), .C(i), .Y(ori_ori_n542_));
  NO2        o514(.A(ori_ori_n398_), .B(ori_ori_n542_), .Y(ori_ori_n543_));
  INV        o515(.A(ori_ori_n384_), .Y(ori_ori_n544_));
  INV        o516(.A(ori_ori_n243_), .Y(ori_ori_n545_));
  NO2        o517(.A(ori_ori_n91_), .B(ori_ori_n89_), .Y(ori_ori_n546_));
  NOi31      o518(.An(k), .B(m), .C(l), .Y(ori_ori_n547_));
  NO2        o519(.A(ori_ori_n245_), .B(ori_ori_n547_), .Y(ori_ori_n548_));
  AOI210     o520(.A0(ori_ori_n548_), .A1(ori_ori_n546_), .B0(ori_ori_n399_), .Y(ori_ori_n549_));
  INV        o521(.A(ori_ori_n237_), .Y(ori_ori_n550_));
  NA2        o522(.A(ori_ori_n247_), .B(ori_ori_n249_), .Y(ori_ori_n551_));
  INV        o523(.A(ori_ori_n551_), .Y(ori_ori_n552_));
  AOI220     o524(.A0(ori_ori_n552_), .A1(ori_ori_n550_), .B0(ori_ori_n549_), .B1(ori_ori_n545_), .Y(ori_ori_n553_));
  NA2        o525(.A(ori_ori_n124_), .B(ori_ori_n86_), .Y(ori_ori_n554_));
  NA3        o526(.A(ori_ori_n554_), .B(ori_ori_n464_), .C(ori_ori_n98_), .Y(ori_ori_n555_));
  NA3        o527(.A(ori_ori_n555_), .B(ori_ori_n144_), .C(ori_ori_n29_), .Y(ori_ori_n556_));
  NA4        o528(.A(ori_ori_n556_), .B(ori_ori_n553_), .C(ori_ori_n413_), .D(ori_ori_n61_), .Y(ori_ori_n557_));
  NO4        o529(.A(ori_ori_n411_), .B(ori_ori_n95_), .C(ori_ori_n232_), .D(ori_ori_n112_), .Y(ori_ori_n558_));
  NO2        o530(.A(ori_ori_n429_), .B(ori_ori_n232_), .Y(ori_ori_n559_));
  INV        o531(.A(ori_ori_n558_), .Y(ori_ori_n560_));
  NA3        o532(.A(ori_ori_n119_), .B(ori_ori_n81_), .C(ori_ori_n80_), .Y(ori_ori_n561_));
  NO2        o533(.A(ori_ori_n243_), .B(ori_ori_n561_), .Y(ori_ori_n562_));
  NOi31      o534(.An(ori_ori_n167_), .B(ori_ori_n562_), .C(ori_ori_n215_), .Y(ori_ori_n563_));
  NA2        o535(.A(c), .B(ori_ori_n87_), .Y(ori_ori_n564_));
  NO2        o536(.A(ori_ori_n564_), .B(ori_ori_n296_), .Y(ori_ori_n565_));
  NA3        o537(.A(ori_ori_n565_), .B(ori_ori_n354_), .C(f), .Y(ori_ori_n566_));
  OR2        o538(.A(ori_ori_n435_), .B(ori_ori_n372_), .Y(ori_ori_n567_));
  INV        o539(.A(ori_ori_n567_), .Y(ori_ori_n568_));
  NA2        o540(.A(ori_ori_n529_), .B(ori_ori_n83_), .Y(ori_ori_n569_));
  NA2        o541(.A(ori_ori_n569_), .B(ori_ori_n568_), .Y(ori_ori_n570_));
  NA4        o542(.A(ori_ori_n570_), .B(ori_ori_n566_), .C(ori_ori_n563_), .D(ori_ori_n560_), .Y(ori_ori_n571_));
  NO3        o543(.A(ori_ori_n571_), .B(ori_ori_n339_), .C(ori_ori_n557_), .Y(ori_ori_n572_));
  NO2        o544(.A(ori_ori_n98_), .B(ori_ori_n95_), .Y(ori_ori_n573_));
  NO2        o545(.A(ori_ori_n174_), .B(ori_ori_n168_), .Y(ori_ori_n574_));
  AOI220     o546(.A0(ori_ori_n574_), .A1(ori_ori_n171_), .B0(ori_ori_n213_), .B1(ori_ori_n573_), .Y(ori_ori_n575_));
  INV        o547(.A(ori_ori_n575_), .Y(ori_ori_n576_));
  NA2        o548(.A(e), .B(d), .Y(ori_ori_n577_));
  OAI220     o549(.A0(ori_ori_n577_), .A1(c), .B0(ori_ori_n227_), .B1(d), .Y(ori_ori_n578_));
  NA3        o550(.A(ori_ori_n578_), .B(ori_ori_n318_), .C(ori_ori_n352_), .Y(ori_ori_n579_));
  AOI210     o551(.A0(ori_ori_n359_), .A1(ori_ori_n135_), .B0(ori_ori_n174_), .Y(ori_ori_n580_));
  INV        o552(.A(ori_ori_n580_), .Y(ori_ori_n581_));
  NA3        o553(.A(ori_ori_n123_), .B(ori_ori_n64_), .C(ori_ori_n31_), .Y(ori_ori_n582_));
  NA3        o554(.A(ori_ori_n582_), .B(ori_ori_n581_), .C(ori_ori_n579_), .Y(ori_ori_n583_));
  NO2        o555(.A(ori_ori_n583_), .B(ori_ori_n576_), .Y(ori_ori_n584_));
  OR2        o556(.A(ori_ori_n466_), .B(ori_ori_n165_), .Y(ori_ori_n585_));
  OAI220     o557(.A0(ori_ori_n411_), .A1(ori_ori_n49_), .B0(ori_ori_n212_), .B1(j), .Y(ori_ori_n586_));
  AOI220     o558(.A0(ori_ori_n586_), .A1(ori_ori_n559_), .B0(ori_ori_n403_), .B1(ori_ori_n410_), .Y(ori_ori_n587_));
  OAI210     o559(.A0(ori_ori_n539_), .A1(ori_ori_n125_), .B0(ori_ori_n587_), .Y(ori_ori_n588_));
  AN2        o560(.A(ori_ori_n550_), .B(ori_ori_n543_), .Y(ori_ori_n589_));
  NO2        o561(.A(ori_ori_n589_), .B(ori_ori_n588_), .Y(ori_ori_n590_));
  AO220      o562(.A0(ori_ori_n318_), .A1(ori_ori_n499_), .B0(ori_ori_n130_), .B1(f), .Y(ori_ori_n591_));
  OAI210     o563(.A0(ori_ori_n591_), .A1(ori_ori_n321_), .B0(ori_ori_n578_), .Y(ori_ori_n592_));
  NA2        o564(.A(ori_ori_n544_), .B(ori_ori_n470_), .Y(ori_ori_n593_));
  AN4        o565(.A(ori_ori_n593_), .B(ori_ori_n592_), .C(ori_ori_n590_), .D(ori_ori_n585_), .Y(ori_ori_n594_));
  NA4        o566(.A(ori_ori_n594_), .B(ori_ori_n584_), .C(ori_ori_n572_), .D(ori_ori_n541_), .Y(ori12));
  NO2        o567(.A(ori_ori_n316_), .B(c), .Y(ori_ori_n596_));
  NO4        o568(.A(ori_ori_n309_), .B(ori_ori_n192_), .C(ori_ori_n395_), .D(ori_ori_n162_), .Y(ori_ori_n597_));
  NA2        o569(.A(ori_ori_n597_), .B(ori_ori_n596_), .Y(ori_ori_n598_));
  NO2        o570(.A(ori_ori_n316_), .B(ori_ori_n87_), .Y(ori_ori_n599_));
  NO2        o571(.A(ori_ori_n546_), .B(ori_ori_n252_), .Y(ori_ori_n600_));
  NA2        o572(.A(ori_ori_n600_), .B(ori_ori_n599_), .Y(ori_ori_n601_));
  NA2        o573(.A(ori_ori_n601_), .B(ori_ori_n598_), .Y(ori_ori_n602_));
  AOI210     o574(.A0(ori_ori_n177_), .A1(ori_ori_n242_), .B0(ori_ori_n156_), .Y(ori_ori_n603_));
  OR2        o575(.A(ori_ori_n603_), .B(ori_ori_n597_), .Y(ori_ori_n604_));
  AOI210     o576(.A0(ori_ori_n239_), .A1(ori_ori_n281_), .B0(ori_ori_n162_), .Y(ori_ori_n605_));
  OAI210     o577(.A0(ori_ori_n605_), .A1(ori_ori_n604_), .B0(ori_ori_n291_), .Y(ori_ori_n606_));
  NO2        o578(.A(ori_ori_n111_), .B(ori_ori_n180_), .Y(ori_ori_n607_));
  NA3        o579(.A(ori_ori_n607_), .B(ori_ori_n183_), .C(i), .Y(ori_ori_n608_));
  NA2        o580(.A(ori_ori_n608_), .B(ori_ori_n606_), .Y(ori_ori_n609_));
  NA2        o581(.A(ori_ori_n228_), .B(ori_ori_n253_), .Y(ori_ori_n610_));
  NO3        o582(.A(ori_ori_n95_), .B(ori_ori_n112_), .C(ori_ori_n162_), .Y(ori_ori_n611_));
  NA2        o583(.A(ori_ori_n611_), .B(ori_ori_n368_), .Y(ori_ori_n612_));
  NA4        o584(.A(ori_ori_n310_), .B(ori_ori_n308_), .C(ori_ori_n136_), .D(g), .Y(ori_ori_n613_));
  NA3        o585(.A(ori_ori_n613_), .B(ori_ori_n612_), .C(ori_ori_n610_), .Y(ori_ori_n614_));
  NO3        o586(.A(ori_ori_n614_), .B(ori_ori_n609_), .C(ori_ori_n602_), .Y(ori_ori_n615_));
  NA2        o587(.A(ori_ori_n378_), .B(ori_ori_n106_), .Y(ori_ori_n616_));
  NOi21      o588(.An(ori_ori_n31_), .B(ori_ori_n429_), .Y(ori_ori_n617_));
  NA2        o589(.A(ori_ori_n617_), .B(ori_ori_n616_), .Y(ori_ori_n618_));
  OAI210     o590(.A0(ori_ori_n191_), .A1(ori_ori_n38_), .B0(ori_ori_n618_), .Y(ori_ori_n619_));
  INV        o591(.A(ori_ori_n226_), .Y(ori_ori_n620_));
  NO2        o592(.A(ori_ori_n349_), .B(ori_ori_n212_), .Y(ori_ori_n621_));
  INV        o593(.A(ori_ori_n621_), .Y(ori_ori_n622_));
  NO2        o594(.A(ori_ori_n622_), .B(ori_ori_n106_), .Y(ori_ori_n623_));
  INV        o595(.A(ori_ori_n265_), .Y(ori_ori_n624_));
  NO4        o596(.A(ori_ori_n624_), .B(ori_ori_n623_), .C(ori_ori_n620_), .D(ori_ori_n619_), .Y(ori_ori_n625_));
  NA2        o597(.A(ori_ori_n250_), .B(g), .Y(ori_ori_n626_));
  NA2        o598(.A(ori_ori_n122_), .B(i), .Y(ori_ori_n627_));
  NA2        o599(.A(ori_ori_n39_), .B(i), .Y(ori_ori_n628_));
  NO2        o600(.A(ori_ori_n628_), .B(ori_ori_n155_), .Y(ori_ori_n629_));
  INV        o601(.A(ori_ori_n629_), .Y(ori_ori_n630_));
  NA2        o602(.A(ori_ori_n378_), .B(ori_ori_n273_), .Y(ori_ori_n631_));
  AOI210     o603(.A0(ori_ori_n631_), .A1(n), .B0(ori_ori_n377_), .Y(ori_ori_n632_));
  OAI220     o604(.A0(ori_ori_n632_), .A1(ori_ori_n626_), .B0(ori_ori_n630_), .B1(ori_ori_n237_), .Y(ori_ori_n633_));
  NA3        o605(.A(ori_ori_n229_), .B(ori_ori_n88_), .C(g), .Y(ori_ori_n634_));
  AOI210     o606(.A0(ori_ori_n444_), .A1(ori_ori_n634_), .B0(m), .Y(ori_ori_n635_));
  OAI210     o607(.A0(ori_ori_n635_), .A1(ori_ori_n600_), .B0(ori_ori_n228_), .Y(ori_ori_n636_));
  INV        o608(.A(ori_ori_n636_), .Y(ori_ori_n637_));
  NA2        o609(.A(ori_ori_n437_), .B(ori_ori_n66_), .Y(ori_ori_n638_));
  NO2        o610(.A(ori_ori_n324_), .B(ori_ori_n162_), .Y(ori_ori_n639_));
  NA2        o611(.A(ori_ori_n639_), .B(ori_ori_n274_), .Y(ori_ori_n640_));
  NA2        o612(.A(ori_ori_n640_), .B(ori_ori_n638_), .Y(ori_ori_n641_));
  NA2        o613(.A(ori_ori_n635_), .B(ori_ori_n599_), .Y(ori_ori_n642_));
  NA2        o614(.A(ori_ori_n420_), .B(ori_ori_n368_), .Y(ori_ori_n643_));
  NA2        o615(.A(ori_ori_n643_), .B(ori_ori_n642_), .Y(ori_ori_n644_));
  NO4        o616(.A(ori_ori_n644_), .B(ori_ori_n641_), .C(ori_ori_n637_), .D(ori_ori_n633_), .Y(ori_ori_n645_));
  NAi31      o617(.An(ori_ori_n103_), .B(ori_ori_n305_), .C(n), .Y(ori_ori_n646_));
  NO3        o618(.A(ori_ori_n89_), .B(ori_ori_n245_), .C(ori_ori_n547_), .Y(ori_ori_n647_));
  NO2        o619(.A(ori_ori_n647_), .B(ori_ori_n646_), .Y(ori_ori_n648_));
  NO3        o620(.A(ori_ori_n202_), .B(ori_ori_n103_), .C(ori_ori_n296_), .Y(ori_ori_n649_));
  AOI210     o621(.A0(ori_ori_n649_), .A1(ori_ori_n344_), .B0(ori_ori_n648_), .Y(ori_ori_n650_));
  INV        o622(.A(ori_ori_n650_), .Y(ori_ori_n651_));
  NA2        o623(.A(ori_ori_n174_), .B(ori_ori_n126_), .Y(ori_ori_n652_));
  NO3        o624(.A(ori_ori_n217_), .B(ori_ori_n310_), .C(ori_ori_n130_), .Y(ori_ori_n653_));
  NOi31      o625(.An(ori_ori_n652_), .B(ori_ori_n653_), .C(ori_ori_n162_), .Y(ori_ori_n654_));
  NAi21      o626(.An(ori_ori_n378_), .B(ori_ori_n639_), .Y(ori_ori_n655_));
  NA2        o627(.A(ori_ori_n332_), .B(g), .Y(ori_ori_n656_));
  NA2        o628(.A(ori_ori_n656_), .B(ori_ori_n655_), .Y(ori_ori_n657_));
  NA2        o629(.A(ori_ori_n603_), .B(ori_ori_n596_), .Y(ori_ori_n658_));
  NA2        o630(.A(ori_ori_n658_), .B(ori_ori_n409_), .Y(ori_ori_n659_));
  OAI210     o631(.A0(ori_ori_n603_), .A1(ori_ori_n597_), .B0(ori_ori_n652_), .Y(ori_ori_n660_));
  NA3        o632(.A(ori_ori_n631_), .B(ori_ori_n337_), .C(ori_ori_n39_), .Y(ori_ori_n661_));
  INV        o633(.A(ori_ori_n236_), .Y(ori_ori_n662_));
  NA3        o634(.A(ori_ori_n662_), .B(ori_ori_n661_), .C(ori_ori_n660_), .Y(ori_ori_n663_));
  OR2        o635(.A(ori_ori_n663_), .B(ori_ori_n659_), .Y(ori_ori_n664_));
  NO4        o636(.A(ori_ori_n664_), .B(ori_ori_n657_), .C(ori_ori_n654_), .D(ori_ori_n651_), .Y(ori_ori_n665_));
  NA4        o637(.A(ori_ori_n665_), .B(ori_ori_n645_), .C(ori_ori_n625_), .D(ori_ori_n615_), .Y(ori13));
  AN2        o638(.A(c), .B(b), .Y(ori_ori_n667_));
  NAi32      o639(.An(d), .Bn(c), .C(e), .Y(ori_ori_n668_));
  AN2        o640(.A(d), .B(c), .Y(ori_ori_n669_));
  NA2        o641(.A(ori_ori_n669_), .B(ori_ori_n87_), .Y(ori_ori_n670_));
  NAi32      o642(.An(f), .Bn(e), .C(c), .Y(ori_ori_n671_));
  NO3        o643(.A(m), .B(i), .C(h), .Y(ori_ori_n672_));
  NA3        o644(.A(k), .B(j), .C(i), .Y(ori_ori_n673_));
  NO2        o645(.A(f), .B(c), .Y(ori_ori_n674_));
  NOi21      o646(.An(ori_ori_n674_), .B(ori_ori_n309_), .Y(ori_ori_n675_));
  AN3        o647(.A(g), .B(f), .C(c), .Y(ori_ori_n676_));
  NA3        o648(.A(l), .B(k), .C(j), .Y(ori_ori_n677_));
  NA2        o649(.A(i), .B(h), .Y(ori_ori_n678_));
  NO3        o650(.A(ori_ori_n678_), .B(ori_ori_n677_), .C(ori_ori_n95_), .Y(ori_ori_n679_));
  NO3        o651(.A(ori_ori_n104_), .B(ori_ori_n206_), .C(ori_ori_n162_), .Y(ori_ori_n680_));
  NOi31      o652(.An(m), .B(n), .C(f), .Y(ori_ori_n681_));
  NA2        o653(.A(ori_ori_n681_), .B(ori_ori_n42_), .Y(ori_ori_n682_));
  AN2        o654(.A(e), .B(c), .Y(ori_ori_n683_));
  NA2        o655(.A(ori_ori_n683_), .B(a), .Y(ori_ori_n684_));
  NO2        o656(.A(ori_ori_n684_), .B(ori_ori_n682_), .Y(ori_ori_n685_));
  NO2        o657(.A(ori_ori_n206_), .B(a), .Y(ori_ori_n686_));
  INV        o658(.A(ori_ori_n685_), .Y(ori_ori_n687_));
  NA2        o659(.A(c), .B(b), .Y(ori_ori_n688_));
  NO2        o660(.A(ori_ori_n469_), .B(ori_ori_n688_), .Y(ori_ori_n689_));
  INV        o661(.A(ori_ori_n301_), .Y(ori_ori_n690_));
  NA2        o662(.A(ori_ori_n690_), .B(ori_ori_n689_), .Y(ori_ori_n691_));
  NAi21      o663(.An(ori_ori_n304_), .B(ori_ori_n689_), .Y(ori_ori_n692_));
  NA2        o664(.A(ori_ori_n374_), .B(ori_ori_n686_), .Y(ori_ori_n693_));
  NA2        o665(.A(ori_ori_n693_), .B(ori_ori_n692_), .Y(ori_ori_n694_));
  INV        o666(.A(ori_ori_n694_), .Y(ori_ori_n695_));
  NA3        o667(.A(ori_ori_n695_), .B(ori_ori_n691_), .C(ori_ori_n687_), .Y(ori00));
  NA2        o668(.A(ori_ori_n354_), .B(f), .Y(ori_ori_n697_));
  OAI210     o669(.A0(ori_ori_n647_), .A1(ori_ori_n36_), .B0(ori_ori_n422_), .Y(ori_ori_n698_));
  NA3        o670(.A(ori_ori_n698_), .B(ori_ori_n197_), .C(n), .Y(ori_ori_n699_));
  AOI210     o671(.A0(ori_ori_n699_), .A1(ori_ori_n697_), .B0(ori_ori_n670_), .Y(ori_ori_n700_));
  INV        o672(.A(ori_ori_n700_), .Y(ori_ori_n701_));
  NA3        o673(.A(ori_ori_n123_), .B(ori_ori_n39_), .C(ori_ori_n38_), .Y(ori_ori_n702_));
  NA3        o674(.A(d), .B(ori_ori_n45_), .C(b), .Y(ori_ori_n703_));
  NO2        o675(.A(ori_ori_n703_), .B(ori_ori_n702_), .Y(ori_ori_n704_));
  NO4        o676(.A(ori_ori_n338_), .B(ori_ori_n255_), .C(ori_ori_n688_), .D(ori_ori_n48_), .Y(ori_ori_n705_));
  NA3        o677(.A(ori_ori_n275_), .B(ori_ori_n166_), .C(g), .Y(ori_ori_n706_));
  OR2        o678(.A(ori_ori_n706_), .B(ori_ori_n703_), .Y(ori_ori_n707_));
  NO2        o679(.A(h), .B(g), .Y(ori_ori_n708_));
  NA4        o680(.A(ori_ori_n344_), .B(ori_ori_n330_), .C(ori_ori_n708_), .D(ori_ori_n667_), .Y(ori_ori_n709_));
  NA2        o681(.A(ori_ori_n611_), .B(ori_ori_n389_), .Y(ori_ori_n710_));
  NA3        o682(.A(ori_ori_n710_), .B(ori_ori_n709_), .C(ori_ori_n707_), .Y(ori_ori_n711_));
  NO2        o683(.A(ori_ori_n711_), .B(ori_ori_n705_), .Y(ori_ori_n712_));
  INV        o684(.A(ori_ori_n392_), .Y(ori_ori_n713_));
  AN3        o685(.A(ori_ori_n713_), .B(ori_ori_n712_), .C(ori_ori_n390_), .Y(ori_ori_n714_));
  NA3        o686(.A(ori_ori_n681_), .B(ori_ori_n401_), .C(ori_ori_n329_), .Y(ori_ori_n715_));
  NA2        o687(.A(ori_ori_n715_), .B(ori_ori_n184_), .Y(ori_ori_n716_));
  NA4        o688(.A(ori_ori_n425_), .B(ori_ori_n158_), .C(ori_ori_n166_), .D(ori_ori_n122_), .Y(ori_ori_n717_));
  INV        o689(.A(ori_ori_n717_), .Y(ori_ori_n718_));
  NA2        o690(.A(n), .B(e), .Y(ori_ori_n719_));
  NO2        o691(.A(ori_ori_n719_), .B(ori_ori_n108_), .Y(ori_ori_n720_));
  NA2        o692(.A(ori_ori_n720_), .B(ori_ori_n549_), .Y(ori_ori_n721_));
  AOI220     o693(.A0(ori_ori_n617_), .A1(ori_ori_n389_), .B0(ori_ori_n425_), .B1(ori_ori_n187_), .Y(ori_ori_n722_));
  NO2        o694(.A(i), .B(h), .Y(ori_ori_n723_));
  NA2        o695(.A(ori_ori_n722_), .B(ori_ori_n721_), .Y(ori_ori_n724_));
  NO3        o696(.A(ori_ori_n724_), .B(ori_ori_n718_), .C(ori_ori_n716_), .Y(ori_ori_n725_));
  NA3        o697(.A(ori_ori_n725_), .B(ori_ori_n714_), .C(ori_ori_n701_), .Y(ori01));
  INV        o698(.A(ori_ori_n205_), .Y(ori_ori_n727_));
  NA2        o699(.A(ori_ori_n286_), .B(i), .Y(ori_ori_n728_));
  NA3        o700(.A(ori_ori_n728_), .B(ori_ori_n727_), .C(ori_ori_n658_), .Y(ori_ori_n729_));
  NA2        o701(.A(ori_ori_n378_), .B(ori_ori_n201_), .Y(ori_ori_n730_));
  NA2        o702(.A(ori_ori_n621_), .B(ori_ori_n730_), .Y(ori_ori_n731_));
  NA2        o703(.A(ori_ori_n731_), .B(ori_ori_n587_), .Y(ori_ori_n732_));
  NAi31      o704(.An(ori_ori_n121_), .B(ori_ori_n717_), .C(ori_ori_n575_), .Y(ori_ori_n733_));
  NO2        o705(.A(ori_ori_n446_), .B(ori_ori_n357_), .Y(ori_ori_n734_));
  OR2        o706(.A(ori_ori_n150_), .B(ori_ori_n148_), .Y(ori_ori_n735_));
  NA3        o707(.A(ori_ori_n735_), .B(ori_ori_n734_), .C(ori_ori_n99_), .Y(ori_ori_n736_));
  NO4        o708(.A(ori_ori_n736_), .B(ori_ori_n733_), .C(ori_ori_n732_), .D(ori_ori_n729_), .Y(ori_ori_n737_));
  INV        o709(.A(ori_ori_n706_), .Y(ori_ori_n738_));
  NA2        o710(.A(ori_ori_n738_), .B(ori_ori_n368_), .Y(ori_ori_n739_));
  AN3        o711(.A(m), .B(l), .C(k), .Y(ori_ori_n740_));
  OAI210     o712(.A0(ori_ori_n257_), .A1(ori_ori_n31_), .B0(ori_ori_n740_), .Y(ori_ori_n741_));
  OR2        o713(.A(ori_ori_n741_), .B(ori_ori_n237_), .Y(ori_ori_n742_));
  NA2        o714(.A(ori_ori_n742_), .B(ori_ori_n739_), .Y(ori_ori_n743_));
  NA2        o715(.A(ori_ori_n204_), .B(ori_ori_n150_), .Y(ori_ori_n744_));
  NA2        o716(.A(ori_ori_n744_), .B(ori_ori_n440_), .Y(ori_ori_n745_));
  INV        o717(.A(ori_ori_n745_), .Y(ori_ori_n746_));
  NO2        o718(.A(ori_ori_n746_), .B(ori_ori_n743_), .Y(ori_ori_n747_));
  NA2        o719(.A(ori_ori_n350_), .B(ori_ori_n47_), .Y(ori_ori_n748_));
  NO2        o720(.A(ori_ori_n159_), .B(ori_ori_n83_), .Y(ori_ori_n749_));
  NO2        o721(.A(ori_ori_n749_), .B(ori_ori_n704_), .Y(ori_ori_n750_));
  NA2        o722(.A(ori_ori_n750_), .B(ori_ori_n748_), .Y(ori_ori_n751_));
  NO2        o723(.A(ori_ori_n627_), .B(ori_ori_n176_), .Y(ori_ori_n752_));
  NO2        o724(.A(ori_ori_n628_), .B(ori_ori_n380_), .Y(ori_ori_n753_));
  OAI210     o725(.A0(ori_ori_n753_), .A1(ori_ori_n752_), .B0(ori_ori_n245_), .Y(ori_ori_n754_));
  NO3        o726(.A(ori_ori_n59_), .B(ori_ori_n212_), .C(ori_ori_n38_), .Y(ori_ori_n755_));
  NA2        o727(.A(ori_ori_n755_), .B(ori_ori_n377_), .Y(ori_ori_n756_));
  INV        o728(.A(ori_ori_n756_), .Y(ori_ori_n757_));
  OR2        o729(.A(ori_ori_n706_), .B(ori_ori_n703_), .Y(ori_ori_n758_));
  NA2        o730(.A(ori_ori_n755_), .B(ori_ori_n530_), .Y(ori_ori_n759_));
  NA3        o731(.A(ori_ori_n759_), .B(ori_ori_n758_), .C(ori_ori_n278_), .Y(ori_ori_n760_));
  NOi41      o732(.An(ori_ori_n754_), .B(ori_ori_n760_), .C(ori_ori_n757_), .D(ori_ori_n751_), .Y(ori_ori_n761_));
  NO2        o733(.A(ori_ori_n94_), .B(ori_ori_n38_), .Y(ori_ori_n762_));
  NO2        o734(.A(ori_ori_n38_), .B(ori_ori_n36_), .Y(ori_ori_n763_));
  AO220      o735(.A0(ori_ori_n763_), .A1(ori_ori_n412_), .B0(ori_ori_n762_), .B1(ori_ori_n474_), .Y(ori_ori_n764_));
  NA2        o736(.A(ori_ori_n764_), .B(ori_ori_n245_), .Y(ori_ori_n765_));
  NO3        o737(.A(ori_ori_n678_), .B(ori_ori_n131_), .C(ori_ori_n65_), .Y(ori_ori_n766_));
  INV        o738(.A(ori_ori_n765_), .Y(ori_ori_n767_));
  NO2        o739(.A(ori_ori_n405_), .B(ori_ori_n404_), .Y(ori_ori_n768_));
  NO4        o740(.A(ori_ori_n678_), .B(ori_ori_n768_), .C(ori_ori_n129_), .D(ori_ori_n65_), .Y(ori_ori_n769_));
  NO2        o741(.A(ori_ori_n769_), .B(ori_ori_n767_), .Y(ori_ori_n770_));
  NA4        o742(.A(ori_ori_n770_), .B(ori_ori_n761_), .C(ori_ori_n747_), .D(ori_ori_n737_), .Y(ori06));
  NO2        o743(.A(ori_ori_n168_), .B(ori_ori_n75_), .Y(ori_ori_n772_));
  OAI210     o744(.A0(ori_ori_n772_), .A1(ori_ori_n766_), .B0(ori_ori_n274_), .Y(ori_ori_n773_));
  NA2        o745(.A(ori_ori_n773_), .B(ori_ori_n754_), .Y(ori_ori_n774_));
  NO3        o746(.A(ori_ori_n774_), .B(ori_ori_n757_), .C(ori_ori_n196_), .Y(ori_ori_n775_));
  NO2        o747(.A(ori_ori_n212_), .B(ori_ori_n38_), .Y(ori_ori_n776_));
  AOI210     o748(.A0(ori_ori_n776_), .A1(ori_ori_n377_), .B0(ori_ori_n752_), .Y(ori_ori_n777_));
  AOI210     o749(.A0(ori_ori_n776_), .A1(ori_ori_n381_), .B0(ori_ori_n764_), .Y(ori_ori_n778_));
  AOI210     o750(.A0(ori_ori_n778_), .A1(ori_ori_n777_), .B0(ori_ori_n242_), .Y(ori_ori_n779_));
  OAI210     o751(.A0(ori_ori_n67_), .A1(ori_ori_n36_), .B0(ori_ori_n445_), .Y(ori_ori_n780_));
  NA2        o752(.A(ori_ori_n780_), .B(ori_ori_n418_), .Y(ori_ori_n781_));
  NO2        o753(.A(ori_ori_n359_), .B(ori_ori_n126_), .Y(ori_ori_n782_));
  NO2        o754(.A(ori_ori_n402_), .B(ori_ori_n682_), .Y(ori_ori_n783_));
  OAI210     o755(.A0(ori_ori_n325_), .A1(ori_ori_n189_), .B0(ori_ori_n582_), .Y(ori_ori_n784_));
  NO3        o756(.A(ori_ori_n784_), .B(ori_ori_n783_), .C(ori_ori_n782_), .Y(ori_ori_n785_));
  NA2        o757(.A(ori_ori_n785_), .B(ori_ori_n781_), .Y(ori_ori_n786_));
  AN2        o758(.A(ori_ori_n617_), .B(ori_ori_n421_), .Y(ori_ori_n787_));
  NO3        o759(.A(ori_ori_n787_), .B(ori_ori_n786_), .C(ori_ori_n779_), .Y(ori_ori_n788_));
  NO3        o760(.A(ori_ori_n186_), .B(ori_ori_n75_), .C(ori_ori_n206_), .Y(ori_ori_n789_));
  OAI220     o761(.A0(ori_ori_n466_), .A1(ori_ori_n189_), .B0(ori_ori_n356_), .B1(ori_ori_n359_), .Y(ori_ori_n790_));
  NO3        o762(.A(ori_ori_n790_), .B(ori_ori_n789_), .C(ori_ori_n685_), .Y(ori_ori_n791_));
  NA2        o763(.A(ori_ori_n791_), .B(ori_ori_n722_), .Y(ori_ori_n792_));
  AN2        o764(.A(ori_ori_n597_), .B(ori_ori_n596_), .Y(ori_ori_n793_));
  NO3        o765(.A(ori_ori_n793_), .B(ori_ori_n346_), .C(ori_ori_n332_), .Y(ori_ori_n794_));
  NA2        o766(.A(ori_ori_n794_), .B(ori_ori_n759_), .Y(ori_ori_n795_));
  NAi21      o767(.An(j), .B(i), .Y(ori_ori_n796_));
  NO4        o768(.A(ori_ori_n768_), .B(ori_ori_n796_), .C(ori_ori_n309_), .D(ori_ori_n178_), .Y(ori_ori_n797_));
  NO3        o769(.A(ori_ori_n797_), .B(ori_ori_n795_), .C(ori_ori_n792_), .Y(ori_ori_n798_));
  NA4        o770(.A(ori_ori_n798_), .B(ori_ori_n788_), .C(ori_ori_n775_), .D(ori_ori_n770_), .Y(ori07));
  NAi32      o771(.An(m), .Bn(b), .C(n), .Y(ori_ori_n800_));
  NO3        o772(.A(ori_ori_n800_), .B(g), .C(f), .Y(ori_ori_n801_));
  NAi21      o773(.An(f), .B(c), .Y(ori_ori_n802_));
  NOi31      o774(.An(n), .B(m), .C(b), .Y(ori_ori_n803_));
  NO3        o775(.A(ori_ori_n95_), .B(ori_ori_n315_), .C(h), .Y(ori_ori_n804_));
  NO3        o776(.A(n), .B(m), .C(h), .Y(ori_ori_n805_));
  NO2        o777(.A(ori_ori_n671_), .B(ori_ori_n309_), .Y(ori_ori_n806_));
  INV        o778(.A(ori_ori_n806_), .Y(ori_ori_n807_));
  NO2        o779(.A(ori_ori_n673_), .B(ori_ori_n216_), .Y(ori_ori_n808_));
  NA2        o780(.A(ori_ori_n373_), .B(ori_ori_n60_), .Y(ori_ori_n809_));
  NA2        o781(.A(ori_ori_n723_), .B(ori_ori_n208_), .Y(ori_ori_n810_));
  NA3        o782(.A(ori_ori_n810_), .B(ori_ori_n809_), .C(ori_ori_n807_), .Y(ori_ori_n811_));
  NO2        o783(.A(ori_ori_n811_), .B(ori_ori_n801_), .Y(ori_ori_n812_));
  NO3        o784(.A(e), .B(d), .C(c), .Y(ori_ori_n813_));
  NO2        o785(.A(ori_ori_n95_), .B(ori_ori_n162_), .Y(ori_ori_n814_));
  NA2        o786(.A(ori_ori_n814_), .B(ori_ori_n813_), .Y(ori_ori_n815_));
  INV        o787(.A(ori_ori_n815_), .Y(ori_ori_n816_));
  NA3        o788(.A(ori_ori_n463_), .B(ori_ori_n452_), .C(ori_ori_n84_), .Y(ori_ori_n817_));
  NO2        o789(.A(ori_ori_n817_), .B(ori_ori_n38_), .Y(ori_ori_n818_));
  NO2        o790(.A(l), .B(k), .Y(ori_ori_n819_));
  NO3        o791(.A(ori_ori_n309_), .B(d), .C(c), .Y(ori_ori_n820_));
  NO2        o792(.A(ori_ori_n818_), .B(ori_ori_n816_), .Y(ori_ori_n821_));
  NO2        o793(.A(g), .B(c), .Y(ori_ori_n822_));
  NO2        o794(.A(ori_ori_n316_), .B(a), .Y(ori_ori_n823_));
  NA2        o795(.A(ori_ori_n823_), .B(ori_ori_n85_), .Y(ori_ori_n824_));
  NO2        o796(.A(ori_ori_n504_), .B(ori_ori_n142_), .Y(ori_ori_n825_));
  NOi31      o797(.An(m), .B(n), .C(b), .Y(ori_ori_n826_));
  NOi31      o798(.An(f), .B(d), .C(c), .Y(ori_ori_n827_));
  NA2        o799(.A(ori_ori_n827_), .B(ori_ori_n826_), .Y(ori_ori_n828_));
  INV        o800(.A(ori_ori_n828_), .Y(ori_ori_n829_));
  NO2        o801(.A(ori_ori_n829_), .B(ori_ori_n825_), .Y(ori_ori_n830_));
  NA2        o802(.A(ori_ori_n676_), .B(ori_ori_n330_), .Y(ori_ori_n831_));
  NO2        o803(.A(ori_ori_n831_), .B(ori_ori_n309_), .Y(ori_ori_n832_));
  NO3        o804(.A(ori_ori_n37_), .B(i), .C(h), .Y(ori_ori_n833_));
  NO2        o805(.A(ori_ori_n672_), .B(ori_ori_n832_), .Y(ori_ori_n834_));
  AN3        o806(.A(ori_ori_n834_), .B(ori_ori_n830_), .C(ori_ori_n824_), .Y(ori_ori_n835_));
  NA2        o807(.A(ori_ori_n803_), .B(ori_ori_n271_), .Y(ori_ori_n836_));
  INV        o808(.A(ori_ori_n836_), .Y(ori_ori_n837_));
  INV        o809(.A(ori_ori_n679_), .Y(ori_ori_n838_));
  NAi21      o810(.An(ori_ori_n837_), .B(ori_ori_n838_), .Y(ori_ori_n839_));
  NO4        o811(.A(ori_ori_n95_), .B(g), .C(f), .D(e), .Y(ori_ori_n840_));
  NA2        o812(.A(ori_ori_n805_), .B(ori_ori_n819_), .Y(ori_ori_n841_));
  INV        o813(.A(ori_ori_n841_), .Y(ori_ori_n842_));
  OR3        o814(.A(ori_ori_n372_), .B(ori_ori_n371_), .C(ori_ori_n84_), .Y(ori_ori_n843_));
  NA2        o815(.A(ori_ori_n681_), .B(ori_ori_n296_), .Y(ori_ori_n844_));
  NO2        o816(.A(ori_ori_n844_), .B(ori_ori_n308_), .Y(ori_ori_n845_));
  OR2        o817(.A(ori_ori_n845_), .B(ori_ori_n842_), .Y(ori_ori_n846_));
  NO2        o818(.A(ori_ori_n846_), .B(ori_ori_n839_), .Y(ori_ori_n847_));
  NA4        o819(.A(ori_ori_n847_), .B(ori_ori_n835_), .C(ori_ori_n821_), .D(ori_ori_n812_), .Y(ori_ori_n848_));
  NO2        o820(.A(ori_ori_n688_), .B(ori_ori_n82_), .Y(ori_ori_n849_));
  NO2        o821(.A(ori_ori_n283_), .B(j), .Y(ori_ori_n850_));
  NA2        o822(.A(ori_ori_n833_), .B(ori_ori_n681_), .Y(ori_ori_n851_));
  NA2        o823(.A(ori_ori_n675_), .B(ori_ori_n110_), .Y(ori_ori_n852_));
  NA2        o824(.A(ori_ori_n852_), .B(ori_ori_n851_), .Y(ori_ori_n853_));
  NA2        o825(.A(ori_ori_n850_), .B(ori_ori_n118_), .Y(ori_ori_n854_));
  INV        o826(.A(ori_ori_n854_), .Y(ori_ori_n855_));
  NO2        o827(.A(ori_ori_n855_), .B(ori_ori_n853_), .Y(ori_ori_n856_));
  INV        o828(.A(ori_ori_n40_), .Y(ori_ori_n857_));
  NA2        o829(.A(ori_ori_n857_), .B(ori_ori_n708_), .Y(ori_ori_n858_));
  INV        o830(.A(ori_ori_n858_), .Y(ori_ori_n859_));
  NO2        o831(.A(ori_ori_n168_), .B(ori_ori_n131_), .Y(ori_ori_n860_));
  NO2        o832(.A(ori_ori_n843_), .B(ori_ori_n252_), .Y(ori_ori_n861_));
  NO3        o833(.A(ori_ori_n861_), .B(ori_ori_n860_), .C(ori_ori_n859_), .Y(ori_ori_n862_));
  NA2        o834(.A(ori_ori_n849_), .B(f), .Y(ori_ori_n863_));
  NO2        o835(.A(ori_ori_n902_), .B(ori_ori_n863_), .Y(ori_ori_n864_));
  NO2        o836(.A(ori_ori_n796_), .B(ori_ori_n129_), .Y(ori_ori_n865_));
  NOi21      o837(.An(d), .B(f), .Y(ori_ori_n866_));
  NA2        o838(.A(h), .B(ori_ori_n865_), .Y(ori_ori_n867_));
  INV        o839(.A(ori_ori_n867_), .Y(ori_ori_n868_));
  NO2        o840(.A(ori_ori_n868_), .B(ori_ori_n864_), .Y(ori_ori_n869_));
  NA3        o841(.A(ori_ori_n869_), .B(ori_ori_n862_), .C(ori_ori_n856_), .Y(ori_ori_n870_));
  NA2        o842(.A(h), .B(ori_ori_n808_), .Y(ori_ori_n871_));
  OAI210     o843(.A0(ori_ori_n840_), .A1(ori_ori_n803_), .B0(ori_ori_n564_), .Y(ori_ori_n872_));
  NO2        o844(.A(ori_ori_n668_), .B(ori_ori_n95_), .Y(ori_ori_n873_));
  NA2        o845(.A(ori_ori_n873_), .B(ori_ori_n411_), .Y(ori_ori_n874_));
  NA3        o846(.A(ori_ori_n874_), .B(ori_ori_n872_), .C(ori_ori_n871_), .Y(ori_ori_n875_));
  NA2        o847(.A(ori_ori_n822_), .B(ori_ori_n866_), .Y(ori_ori_n876_));
  NO2        o848(.A(ori_ori_n876_), .B(m), .Y(ori_ori_n877_));
  NA2        o849(.A(ori_ori_n680_), .B(ori_ori_n166_), .Y(ori_ori_n878_));
  NO2        o850(.A(ori_ori_n111_), .B(ori_ori_n136_), .Y(ori_ori_n879_));
  OAI210     o851(.A0(ori_ori_n879_), .A1(ori_ori_n82_), .B0(ori_ori_n826_), .Y(ori_ori_n880_));
  NA2        o852(.A(ori_ori_n880_), .B(ori_ori_n878_), .Y(ori_ori_n881_));
  NO3        o853(.A(ori_ori_n881_), .B(ori_ori_n877_), .C(ori_ori_n875_), .Y(ori_ori_n882_));
  NO2        o854(.A(ori_ori_n802_), .B(e), .Y(ori_ori_n883_));
  NA2        o855(.A(ori_ori_n883_), .B(ori_ori_n294_), .Y(ori_ori_n884_));
  NO2        o856(.A(ori_ori_n95_), .B(ori_ori_n884_), .Y(ori_ori_n885_));
  INV        o857(.A(ori_ori_n885_), .Y(ori_ori_n886_));
  INV        o858(.A(ori_ori_n820_), .Y(ori_ori_n887_));
  OAI210     o859(.A0(g), .A1(ori_ori_n51_), .B0(ori_ori_n887_), .Y(ori_ori_n888_));
  OR2        o860(.A(h), .B(ori_ori_n371_), .Y(ori_ori_n889_));
  NO2        o861(.A(ori_ori_n889_), .B(ori_ori_n129_), .Y(ori_ori_n890_));
  NO2        o862(.A(ori_ori_n40_), .B(l), .Y(ori_ori_n891_));
  INV        o863(.A(ori_ori_n334_), .Y(ori_ori_n892_));
  NA2        o864(.A(ori_ori_n892_), .B(ori_ori_n891_), .Y(ori_ori_n893_));
  INV        o865(.A(ori_ori_n893_), .Y(ori_ori_n894_));
  NO3        o866(.A(ori_ori_n894_), .B(ori_ori_n890_), .C(ori_ori_n888_), .Y(ori_ori_n895_));
  NA3        o867(.A(ori_ori_n895_), .B(ori_ori_n886_), .C(ori_ori_n882_), .Y(ori_ori_n896_));
  NA3        o868(.A(ori_ori_n904_), .B(ori_ori_n100_), .C(ori_ori_n39_), .Y(ori_ori_n897_));
  NA2        o869(.A(ori_ori_n903_), .B(ori_ori_n897_), .Y(ori_ori_n898_));
  OR4        o870(.A(ori_ori_n898_), .B(ori_ori_n896_), .C(ori_ori_n870_), .D(ori_ori_n848_), .Y(ori04));
  INV        o871(.A(ori_ori_n85_), .Y(ori_ori_n902_));
  INV        o872(.A(ori_ori_n804_), .Y(ori_ori_n903_));
  INV        o873(.A(n), .Y(ori_ori_n904_));
  ZERO       o874(.Y(ori02));
  ZERO       o875(.Y(ori03));
  ZERO       o876(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  NO2        m0026(.A(mai_mai_n54_), .B(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(g), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi41      m0043(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n72_));
  NA2        m0044(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n73_));
  INV        m0045(.A(m), .Y(mai_mai_n74_));
  NOi21      m0046(.An(k), .B(l), .Y(mai_mai_n75_));
  NA2        m0047(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  AN4        m0048(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n77_));
  NAi32      m0049(.An(m), .Bn(k), .C(j), .Y(mai_mai_n78_));
  NOi32      m0050(.An(h), .Bn(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n73_), .B(mai_mai_n64_), .Y(mai_mai_n80_));
  INV        m0052(.A(n), .Y(mai_mai_n81_));
  NOi32      m0053(.An(e), .Bn(b), .C(d), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n83_));
  INV        m0055(.A(j), .Y(mai_mai_n84_));
  AN3        m0056(.A(m), .B(k), .C(i), .Y(mai_mai_n85_));
  NA3        m0057(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .Y(mai_mai_n86_));
  NO2        m0058(.A(mai_mai_n86_), .B(f), .Y(mai_mai_n87_));
  NAi32      m0059(.An(g), .Bn(f), .C(h), .Y(mai_mai_n88_));
  NAi31      m0060(.An(j), .B(m), .C(l), .Y(mai_mai_n89_));
  NO2        m0061(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n90_));
  NA2        m0062(.A(m), .B(l), .Y(mai_mai_n91_));
  NAi31      m0063(.An(k), .B(j), .C(g), .Y(mai_mai_n92_));
  NO3        m0064(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(f), .Y(mai_mai_n93_));
  AN2        m0065(.A(j), .B(g), .Y(mai_mai_n94_));
  NOi32      m0066(.An(m), .Bn(l), .C(i), .Y(mai_mai_n95_));
  NOi21      m0067(.An(g), .B(i), .Y(mai_mai_n96_));
  NOi32      m0068(.An(m), .Bn(j), .C(k), .Y(mai_mai_n97_));
  AOI220     m0069(.A0(mai_mai_n97_), .A1(mai_mai_n96_), .B0(mai_mai_n95_), .B1(mai_mai_n94_), .Y(mai_mai_n98_));
  NO2        m0070(.A(mai_mai_n98_), .B(f), .Y(mai_mai_n99_));
  NO4        m0071(.A(mai_mai_n99_), .B(mai_mai_n93_), .C(mai_mai_n90_), .D(mai_mai_n87_), .Y(mai_mai_n100_));
  NAi41      m0072(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n101_));
  AN2        m0073(.A(e), .B(b), .Y(mai_mai_n102_));
  NOi31      m0074(.An(c), .B(h), .C(f), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NOi21      m0076(.An(i), .B(h), .Y(mai_mai_n105_));
  NA3        m0077(.A(mai_mai_n105_), .B(g), .C(mai_mai_n36_), .Y(mai_mai_n106_));
  INV        m0078(.A(a), .Y(mai_mai_n107_));
  NA2        m0079(.A(mai_mai_n102_), .B(mai_mai_n107_), .Y(mai_mai_n108_));
  INV        m0080(.A(l), .Y(mai_mai_n109_));
  NOi21      m0081(.An(m), .B(n), .Y(mai_mai_n110_));
  AN2        m0082(.A(k), .B(h), .Y(mai_mai_n111_));
  NO2        m0083(.A(mai_mai_n106_), .B(mai_mai_n83_), .Y(mai_mai_n112_));
  INV        m0084(.A(b), .Y(mai_mai_n113_));
  NA2        m0085(.A(l), .B(j), .Y(mai_mai_n114_));
  AN2        m0086(.A(k), .B(i), .Y(mai_mai_n115_));
  NA2        m0087(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NA2        m0088(.A(g), .B(e), .Y(mai_mai_n117_));
  NOi32      m0089(.An(c), .Bn(a), .C(d), .Y(mai_mai_n118_));
  NA2        m0090(.A(mai_mai_n118_), .B(mai_mai_n110_), .Y(mai_mai_n119_));
  NO4        m0091(.A(mai_mai_n119_), .B(mai_mai_n117_), .C(mai_mai_n116_), .D(mai_mai_n113_), .Y(mai_mai_n120_));
  NO2        m0092(.A(mai_mai_n120_), .B(mai_mai_n112_), .Y(mai_mai_n121_));
  OAI210     m0093(.A0(mai_mai_n100_), .A1(mai_mai_n83_), .B0(mai_mai_n121_), .Y(mai_mai_n122_));
  NOi31      m0094(.An(k), .B(m), .C(j), .Y(mai_mai_n123_));
  NOi31      m0095(.An(k), .B(m), .C(i), .Y(mai_mai_n124_));
  NA3        m0096(.A(mai_mai_n124_), .B(mai_mai_n79_), .C(mai_mai_n77_), .Y(mai_mai_n125_));
  INV        m0097(.A(mai_mai_n125_), .Y(mai_mai_n126_));
  NOi32      m0098(.An(f), .Bn(b), .C(e), .Y(mai_mai_n127_));
  NAi21      m0099(.An(g), .B(h), .Y(mai_mai_n128_));
  NAi21      m0100(.An(m), .B(n), .Y(mai_mai_n129_));
  NAi21      m0101(.An(j), .B(k), .Y(mai_mai_n130_));
  NAi41      m0102(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n131_));
  NAi31      m0103(.An(j), .B(k), .C(h), .Y(mai_mai_n132_));
  NO3        m0104(.A(mai_mai_n132_), .B(mai_mai_n131_), .C(mai_mai_n129_), .Y(mai_mai_n133_));
  INV        m0105(.A(mai_mai_n133_), .Y(mai_mai_n134_));
  NO2        m0106(.A(k), .B(j), .Y(mai_mai_n135_));
  AN2        m0107(.A(k), .B(j), .Y(mai_mai_n136_));
  NAi21      m0108(.An(c), .B(b), .Y(mai_mai_n137_));
  NA2        m0109(.A(f), .B(d), .Y(mai_mai_n138_));
  NA2        m0110(.A(h), .B(c), .Y(mai_mai_n139_));
  NAi31      m0111(.An(f), .B(e), .C(b), .Y(mai_mai_n140_));
  NA2        m0112(.A(d), .B(b), .Y(mai_mai_n141_));
  NAi21      m0113(.An(e), .B(f), .Y(mai_mai_n142_));
  NO2        m0114(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  NA2        m0115(.A(b), .B(a), .Y(mai_mai_n144_));
  NAi21      m0116(.An(c), .B(d), .Y(mai_mai_n145_));
  NAi31      m0117(.An(l), .B(k), .C(h), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n129_), .B(mai_mai_n146_), .Y(mai_mai_n147_));
  NA2        m0119(.A(mai_mai_n147_), .B(mai_mai_n143_), .Y(mai_mai_n148_));
  NAi31      m0120(.An(mai_mai_n126_), .B(mai_mai_n148_), .C(mai_mai_n134_), .Y(mai_mai_n149_));
  NAi31      m0121(.An(e), .B(f), .C(b), .Y(mai_mai_n150_));
  NOi21      m0122(.An(g), .B(d), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  NOi21      m0124(.An(h), .B(i), .Y(mai_mai_n153_));
  NOi21      m0125(.An(k), .B(m), .Y(mai_mai_n154_));
  NA3        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .C(n), .Y(mai_mai_n155_));
  NOi21      m0127(.An(mai_mai_n152_), .B(mai_mai_n155_), .Y(mai_mai_n156_));
  NOi21      m0128(.An(h), .B(g), .Y(mai_mai_n157_));
  NO2        m0129(.A(mai_mai_n138_), .B(mai_mai_n137_), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NAi31      m0131(.An(l), .B(j), .C(h), .Y(mai_mai_n160_));
  NO2        m0132(.A(mai_mai_n160_), .B(mai_mai_n49_), .Y(mai_mai_n161_));
  NA2        m0133(.A(mai_mai_n161_), .B(mai_mai_n67_), .Y(mai_mai_n162_));
  NOi32      m0134(.An(n), .Bn(k), .C(m), .Y(mai_mai_n163_));
  NA2        m0135(.A(l), .B(i), .Y(mai_mai_n164_));
  INV        m0136(.A(mai_mai_n163_), .Y(mai_mai_n165_));
  OAI210     m0137(.A0(mai_mai_n165_), .A1(mai_mai_n159_), .B0(mai_mai_n162_), .Y(mai_mai_n166_));
  NAi31      m0138(.An(d), .B(f), .C(c), .Y(mai_mai_n167_));
  NAi31      m0139(.An(e), .B(f), .C(c), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  NA2        m0141(.A(j), .B(h), .Y(mai_mai_n170_));
  OR3        m0142(.A(n), .B(m), .C(k), .Y(mai_mai_n171_));
  NO2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NAi32      m0144(.An(m), .Bn(k), .C(n), .Y(mai_mai_n173_));
  NO2        m0145(.A(mai_mai_n173_), .B(mai_mai_n170_), .Y(mai_mai_n174_));
  AOI220     m0146(.A0(mai_mai_n174_), .A1(mai_mai_n152_), .B0(mai_mai_n172_), .B1(mai_mai_n169_), .Y(mai_mai_n175_));
  NO2        m0147(.A(n), .B(m), .Y(mai_mai_n176_));
  NA2        m0148(.A(mai_mai_n176_), .B(mai_mai_n50_), .Y(mai_mai_n177_));
  NAi21      m0149(.An(f), .B(e), .Y(mai_mai_n178_));
  NA2        m0150(.A(d), .B(c), .Y(mai_mai_n179_));
  NAi21      m0151(.An(d), .B(c), .Y(mai_mai_n180_));
  NAi31      m0152(.An(m), .B(n), .C(b), .Y(mai_mai_n181_));
  NA2        m0153(.A(k), .B(i), .Y(mai_mai_n182_));
  NAi21      m0154(.An(h), .B(f), .Y(mai_mai_n183_));
  NO2        m0155(.A(mai_mai_n181_), .B(mai_mai_n145_), .Y(mai_mai_n184_));
  NOi32      m0156(.An(f), .Bn(c), .C(d), .Y(mai_mai_n185_));
  NOi32      m0157(.An(f), .Bn(c), .C(e), .Y(mai_mai_n186_));
  NO2        m0158(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NO3        m0159(.A(n), .B(m), .C(j), .Y(mai_mai_n188_));
  NA2        m0160(.A(mai_mai_n188_), .B(mai_mai_n111_), .Y(mai_mai_n189_));
  AO210      m0161(.A0(mai_mai_n189_), .A1(mai_mai_n177_), .B0(mai_mai_n187_), .Y(mai_mai_n190_));
  NA2        m0162(.A(mai_mai_n190_), .B(mai_mai_n175_), .Y(mai_mai_n191_));
  OR4        m0163(.A(mai_mai_n191_), .B(mai_mai_n166_), .C(mai_mai_n156_), .D(mai_mai_n149_), .Y(mai_mai_n192_));
  NO4        m0164(.A(mai_mai_n192_), .B(mai_mai_n122_), .C(mai_mai_n80_), .D(mai_mai_n55_), .Y(mai_mai_n193_));
  NA3        m0165(.A(m), .B(mai_mai_n109_), .C(j), .Y(mai_mai_n194_));
  NAi31      m0166(.An(n), .B(h), .C(g), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NOi32      m0168(.An(m), .Bn(k), .C(l), .Y(mai_mai_n197_));
  NA3        m0169(.A(mai_mai_n197_), .B(mai_mai_n84_), .C(g), .Y(mai_mai_n198_));
  NO2        m0170(.A(mai_mai_n198_), .B(n), .Y(mai_mai_n199_));
  NA4        m0171(.A(k), .B(mai_mai_n110_), .C(i), .D(g), .Y(mai_mai_n200_));
  AN2        m0172(.A(i), .B(g), .Y(mai_mai_n201_));
  INV        m0173(.A(mai_mai_n200_), .Y(mai_mai_n202_));
  NO3        m0174(.A(mai_mai_n202_), .B(mai_mai_n199_), .C(mai_mai_n196_), .Y(mai_mai_n203_));
  NAi41      m0175(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n204_));
  INV        m0176(.A(mai_mai_n204_), .Y(mai_mai_n205_));
  INV        m0177(.A(f), .Y(mai_mai_n206_));
  INV        m0178(.A(g), .Y(mai_mai_n207_));
  NOi31      m0179(.An(i), .B(j), .C(h), .Y(mai_mai_n208_));
  NOi21      m0180(.An(l), .B(m), .Y(mai_mai_n209_));
  NA2        m0181(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  NO3        m0182(.A(mai_mai_n210_), .B(mai_mai_n207_), .C(mai_mai_n206_), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n205_), .Y(mai_mai_n212_));
  OAI210     m0184(.A0(mai_mai_n203_), .A1(mai_mai_n32_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  NOi21      m0185(.An(n), .B(m), .Y(mai_mai_n214_));
  NOi32      m0186(.An(l), .Bn(i), .C(j), .Y(mai_mai_n215_));
  NA2        m0187(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n216_));
  OR2        m0188(.A(mai_mai_n216_), .B(mai_mai_n104_), .Y(mai_mai_n217_));
  NAi21      m0189(.An(j), .B(h), .Y(mai_mai_n218_));
  XN2        m0190(.A(i), .B(h), .Y(mai_mai_n219_));
  NA2        m0191(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  NOi31      m0192(.An(k), .B(n), .C(m), .Y(mai_mai_n221_));
  NOi31      m0193(.An(mai_mai_n221_), .B(mai_mai_n179_), .C(mai_mai_n178_), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n220_), .Y(mai_mai_n223_));
  NAi31      m0195(.An(f), .B(e), .C(c), .Y(mai_mai_n224_));
  NO4        m0196(.A(mai_mai_n224_), .B(mai_mai_n171_), .C(mai_mai_n170_), .D(mai_mai_n59_), .Y(mai_mai_n225_));
  NA4        m0197(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n226_));
  NAi32      m0198(.An(m), .Bn(i), .C(k), .Y(mai_mai_n227_));
  NO3        m0199(.A(mai_mai_n227_), .B(mai_mai_n88_), .C(mai_mai_n226_), .Y(mai_mai_n228_));
  INV        m0200(.A(k), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n228_), .B(mai_mai_n225_), .Y(mai_mai_n230_));
  NAi21      m0202(.An(n), .B(a), .Y(mai_mai_n231_));
  NO2        m0203(.A(mai_mai_n231_), .B(mai_mai_n141_), .Y(mai_mai_n232_));
  NAi41      m0204(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n233_));
  NO2        m0205(.A(mai_mai_n233_), .B(e), .Y(mai_mai_n234_));
  NO3        m0206(.A(mai_mai_n142_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n235_));
  OAI210     m0207(.A0(mai_mai_n235_), .A1(mai_mai_n234_), .B0(mai_mai_n232_), .Y(mai_mai_n236_));
  AN4        m0208(.A(mai_mai_n236_), .B(mai_mai_n230_), .C(mai_mai_n223_), .D(mai_mai_n217_), .Y(mai_mai_n237_));
  OR2        m0209(.A(h), .B(g), .Y(mai_mai_n238_));
  NAi41      m0210(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(mai_mai_n206_), .Y(mai_mai_n240_));
  NA2        m0212(.A(mai_mai_n154_), .B(mai_mai_n105_), .Y(mai_mai_n241_));
  NAi21      m0213(.An(mai_mai_n241_), .B(mai_mai_n240_), .Y(mai_mai_n242_));
  NO2        m0214(.A(n), .B(a), .Y(mai_mai_n243_));
  NAi31      m0215(.An(mai_mai_n233_), .B(mai_mai_n243_), .C(mai_mai_n102_), .Y(mai_mai_n244_));
  AN2        m0216(.A(mai_mai_n244_), .B(mai_mai_n242_), .Y(mai_mai_n245_));
  NAi21      m0217(.An(h), .B(i), .Y(mai_mai_n246_));
  NA2        m0218(.A(mai_mai_n176_), .B(k), .Y(mai_mai_n247_));
  NO2        m0219(.A(mai_mai_n247_), .B(mai_mai_n246_), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n248_), .B(mai_mai_n185_), .Y(mai_mai_n249_));
  NA2        m0221(.A(mai_mai_n249_), .B(mai_mai_n245_), .Y(mai_mai_n250_));
  NOi21      m0222(.An(g), .B(e), .Y(mai_mai_n251_));
  NO2        m0223(.A(mai_mai_n72_), .B(mai_mai_n74_), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n252_), .B(mai_mai_n251_), .Y(mai_mai_n253_));
  NOi32      m0225(.An(l), .Bn(j), .C(i), .Y(mai_mai_n254_));
  AOI210     m0226(.A0(mai_mai_n75_), .A1(mai_mai_n84_), .B0(mai_mai_n254_), .Y(mai_mai_n255_));
  NO2        m0227(.A(mai_mai_n246_), .B(mai_mai_n44_), .Y(mai_mai_n256_));
  NAi21      m0228(.An(f), .B(g), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n65_), .Y(mai_mai_n258_));
  NO2        m0230(.A(mai_mai_n69_), .B(mai_mai_n114_), .Y(mai_mai_n259_));
  AOI220     m0231(.A0(mai_mai_n259_), .A1(mai_mai_n258_), .B0(mai_mai_n256_), .B1(mai_mai_n67_), .Y(mai_mai_n260_));
  OAI210     m0232(.A0(mai_mai_n255_), .A1(mai_mai_n253_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  NO3        m0233(.A(mai_mai_n130_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n262_));
  NOi41      m0234(.An(mai_mai_n237_), .B(mai_mai_n261_), .C(mai_mai_n250_), .D(mai_mai_n213_), .Y(mai_mai_n263_));
  NO4        m0235(.A(mai_mai_n196_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n264_), .B(mai_mai_n108_), .Y(mai_mai_n265_));
  NA3        m0237(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n266_));
  NAi21      m0238(.An(h), .B(g), .Y(mai_mai_n267_));
  OR4        m0239(.A(mai_mai_n267_), .B(mai_mai_n266_), .C(mai_mai_n216_), .D(e), .Y(mai_mai_n268_));
  NO2        m0240(.A(mai_mai_n241_), .B(mai_mai_n257_), .Y(mai_mai_n269_));
  NA2        m0241(.A(mai_mai_n269_), .B(mai_mai_n77_), .Y(mai_mai_n270_));
  NAi31      m0242(.An(g), .B(k), .C(h), .Y(mai_mai_n271_));
  NO3        m0243(.A(mai_mai_n129_), .B(mai_mai_n271_), .C(l), .Y(mai_mai_n272_));
  NAi31      m0244(.An(e), .B(d), .C(a), .Y(mai_mai_n273_));
  NA2        m0245(.A(mai_mai_n272_), .B(mai_mai_n127_), .Y(mai_mai_n274_));
  NA3        m0246(.A(mai_mai_n274_), .B(mai_mai_n270_), .C(mai_mai_n268_), .Y(mai_mai_n275_));
  NA3        m0247(.A(mai_mai_n154_), .B(mai_mai_n153_), .C(mai_mai_n81_), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n276_), .B(mai_mai_n187_), .Y(mai_mai_n277_));
  INV        m0249(.A(mai_mai_n277_), .Y(mai_mai_n278_));
  NA3        m0250(.A(e), .B(c), .C(b), .Y(mai_mai_n279_));
  NO2        m0251(.A(mai_mai_n60_), .B(mai_mai_n279_), .Y(mai_mai_n280_));
  NAi32      m0252(.An(k), .Bn(i), .C(j), .Y(mai_mai_n281_));
  NAi31      m0253(.An(h), .B(l), .C(i), .Y(mai_mai_n282_));
  NA3        m0254(.A(mai_mai_n282_), .B(mai_mai_n281_), .C(mai_mai_n160_), .Y(mai_mai_n283_));
  NOi21      m0255(.An(mai_mai_n283_), .B(mai_mai_n49_), .Y(mai_mai_n284_));
  OAI210     m0256(.A0(mai_mai_n258_), .A1(mai_mai_n280_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  NAi21      m0257(.An(l), .B(k), .Y(mai_mai_n286_));
  NO2        m0258(.A(mai_mai_n286_), .B(mai_mai_n49_), .Y(mai_mai_n287_));
  NOi21      m0259(.An(l), .B(j), .Y(mai_mai_n288_));
  NA2        m0260(.A(mai_mai_n157_), .B(mai_mai_n288_), .Y(mai_mai_n289_));
  NA3        m0261(.A(mai_mai_n115_), .B(mai_mai_n114_), .C(g), .Y(mai_mai_n290_));
  OR3        m0262(.A(mai_mai_n72_), .B(mai_mai_n74_), .C(e), .Y(mai_mai_n291_));
  AOI210     m0263(.A0(mai_mai_n290_), .A1(mai_mai_n289_), .B0(mai_mai_n291_), .Y(mai_mai_n292_));
  INV        m0264(.A(mai_mai_n292_), .Y(mai_mai_n293_));
  NAi32      m0265(.An(j), .Bn(h), .C(i), .Y(mai_mai_n294_));
  NAi21      m0266(.An(m), .B(l), .Y(mai_mai_n295_));
  NO3        m0267(.A(mai_mai_n295_), .B(mai_mai_n294_), .C(mai_mai_n81_), .Y(mai_mai_n296_));
  NA2        m0268(.A(h), .B(g), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n163_), .B(mai_mai_n45_), .Y(mai_mai_n298_));
  NO2        m0270(.A(mai_mai_n298_), .B(mai_mai_n297_), .Y(mai_mai_n299_));
  OAI210     m0271(.A0(mai_mai_n299_), .A1(mai_mai_n296_), .B0(mai_mai_n158_), .Y(mai_mai_n300_));
  NA4        m0272(.A(mai_mai_n300_), .B(mai_mai_n293_), .C(mai_mai_n285_), .D(mai_mai_n278_), .Y(mai_mai_n301_));
  NO2        m0273(.A(mai_mai_n140_), .B(d), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n303_));
  NAi32      m0275(.An(n), .Bn(m), .C(l), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n119_), .B(mai_mai_n113_), .Y(mai_mai_n305_));
  NAi31      m0277(.An(k), .B(l), .C(j), .Y(mai_mai_n306_));
  OAI210     m0278(.A0(mai_mai_n286_), .A1(j), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  NOi21      m0279(.An(mai_mai_n307_), .B(mai_mai_n117_), .Y(mai_mai_n308_));
  NA2        m0280(.A(mai_mai_n308_), .B(mai_mai_n305_), .Y(mai_mai_n309_));
  INV        m0281(.A(mai_mai_n309_), .Y(mai_mai_n310_));
  NO4        m0282(.A(mai_mai_n310_), .B(mai_mai_n301_), .C(mai_mai_n275_), .D(mai_mai_n265_), .Y(mai_mai_n311_));
  NA2        m0283(.A(mai_mai_n248_), .B(mai_mai_n186_), .Y(mai_mai_n312_));
  NAi21      m0284(.An(m), .B(k), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n219_), .B(mai_mai_n313_), .Y(mai_mai_n314_));
  NAi31      m0286(.An(i), .B(l), .C(h), .Y(mai_mai_n315_));
  NO4        m0287(.A(mai_mai_n315_), .B(e), .C(mai_mai_n72_), .D(mai_mai_n74_), .Y(mai_mai_n316_));
  NA2        m0288(.A(e), .B(c), .Y(mai_mai_n317_));
  NO3        m0289(.A(mai_mai_n317_), .B(n), .C(d), .Y(mai_mai_n318_));
  NOi21      m0290(.An(f), .B(h), .Y(mai_mai_n319_));
  NA2        m0291(.A(mai_mai_n319_), .B(mai_mai_n115_), .Y(mai_mai_n320_));
  NO2        m0292(.A(mai_mai_n320_), .B(mai_mai_n207_), .Y(mai_mai_n321_));
  NAi31      m0293(.An(d), .B(e), .C(b), .Y(mai_mai_n322_));
  NO2        m0294(.A(mai_mai_n129_), .B(mai_mai_n322_), .Y(mai_mai_n323_));
  NA2        m0295(.A(mai_mai_n323_), .B(mai_mai_n321_), .Y(mai_mai_n324_));
  NAi31      m0296(.An(mai_mai_n316_), .B(mai_mai_n324_), .C(mai_mai_n312_), .Y(mai_mai_n325_));
  NA2        m0297(.A(mai_mai_n243_), .B(mai_mai_n102_), .Y(mai_mai_n326_));
  OR2        m0298(.A(mai_mai_n326_), .B(mai_mai_n198_), .Y(mai_mai_n327_));
  NOi31      m0299(.An(l), .B(n), .C(m), .Y(mai_mai_n328_));
  INV        m0300(.A(mai_mai_n327_), .Y(mai_mai_n329_));
  NAi32      m0301(.An(m), .Bn(j), .C(k), .Y(mai_mai_n330_));
  NAi41      m0302(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n331_));
  AN3        m0303(.A(h), .B(g), .C(f), .Y(mai_mai_n332_));
  NOi32      m0304(.An(m), .Bn(j), .C(l), .Y(mai_mai_n333_));
  NO2        m0305(.A(mai_mai_n333_), .B(mai_mai_n95_), .Y(mai_mai_n334_));
  NAi32      m0306(.An(mai_mai_n334_), .Bn(mai_mai_n195_), .C(mai_mai_n302_), .Y(mai_mai_n335_));
  NO2        m0307(.A(mai_mai_n295_), .B(mai_mai_n294_), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n210_), .B(g), .Y(mai_mai_n337_));
  NO2        m0309(.A(mai_mai_n150_), .B(mai_mai_n81_), .Y(mai_mai_n338_));
  AOI220     m0310(.A0(mai_mai_n338_), .A1(mai_mai_n337_), .B0(mai_mai_n240_), .B1(mai_mai_n336_), .Y(mai_mai_n339_));
  INV        m0311(.A(mai_mai_n227_), .Y(mai_mai_n340_));
  NA3        m0312(.A(mai_mai_n340_), .B(mai_mai_n332_), .C(mai_mai_n205_), .Y(mai_mai_n341_));
  NA3        m0313(.A(mai_mai_n341_), .B(mai_mai_n339_), .C(mai_mai_n335_), .Y(mai_mai_n342_));
  NA3        m0314(.A(h), .B(g), .C(f), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n343_), .B(mai_mai_n76_), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n157_), .B(e), .Y(mai_mai_n345_));
  NO2        m0317(.A(mai_mai_n345_), .B(mai_mai_n41_), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n346_), .B(mai_mai_n305_), .Y(mai_mai_n347_));
  NOi32      m0319(.An(j), .Bn(g), .C(i), .Y(mai_mai_n348_));
  NA3        m0320(.A(mai_mai_n348_), .B(mai_mai_n286_), .C(mai_mai_n110_), .Y(mai_mai_n349_));
  AO210      m0321(.A0(mai_mai_n108_), .A1(mai_mai_n32_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NOi32      m0322(.An(e), .Bn(b), .C(a), .Y(mai_mai_n351_));
  AN2        m0323(.A(l), .B(j), .Y(mai_mai_n352_));
  NA2        m0324(.A(mai_mai_n200_), .B(mai_mai_n35_), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n353_), .B(mai_mai_n351_), .Y(mai_mai_n354_));
  NO2        m0326(.A(mai_mai_n322_), .B(n), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n201_), .B(k), .Y(mai_mai_n356_));
  NA3        m0328(.A(m), .B(mai_mai_n109_), .C(mai_mai_n206_), .Y(mai_mai_n357_));
  NA4        m0329(.A(mai_mai_n197_), .B(mai_mai_n84_), .C(g), .D(mai_mai_n206_), .Y(mai_mai_n358_));
  OAI210     m0330(.A0(mai_mai_n357_), .A1(mai_mai_n356_), .B0(mai_mai_n358_), .Y(mai_mai_n359_));
  NAi41      m0331(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n360_));
  NA2        m0332(.A(mai_mai_n51_), .B(mai_mai_n110_), .Y(mai_mai_n361_));
  NO2        m0333(.A(mai_mai_n361_), .B(mai_mai_n360_), .Y(mai_mai_n362_));
  AOI220     m0334(.A0(mai_mai_n362_), .A1(b), .B0(mai_mai_n359_), .B1(mai_mai_n355_), .Y(mai_mai_n363_));
  NA4        m0335(.A(mai_mai_n363_), .B(mai_mai_n354_), .C(mai_mai_n350_), .D(mai_mai_n347_), .Y(mai_mai_n364_));
  NO4        m0336(.A(mai_mai_n364_), .B(mai_mai_n342_), .C(mai_mai_n329_), .D(mai_mai_n325_), .Y(mai_mai_n365_));
  NA4        m0337(.A(mai_mai_n365_), .B(mai_mai_n311_), .C(mai_mai_n263_), .D(mai_mai_n193_), .Y(mai10));
  NA3        m0338(.A(m), .B(k), .C(i), .Y(mai_mai_n367_));
  NO3        m0339(.A(mai_mai_n367_), .B(j), .C(mai_mai_n207_), .Y(mai_mai_n368_));
  NOi21      m0340(.An(e), .B(f), .Y(mai_mai_n369_));
  NO4        m0341(.A(mai_mai_n145_), .B(mai_mai_n369_), .C(n), .D(mai_mai_n107_), .Y(mai_mai_n370_));
  NAi31      m0342(.An(b), .B(f), .C(c), .Y(mai_mai_n371_));
  INV        m0343(.A(mai_mai_n371_), .Y(mai_mai_n372_));
  NOi32      m0344(.An(k), .Bn(h), .C(j), .Y(mai_mai_n373_));
  NA2        m0345(.A(mai_mai_n373_), .B(mai_mai_n214_), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n155_), .B(mai_mai_n374_), .Y(mai_mai_n375_));
  AOI220     m0347(.A0(mai_mai_n375_), .A1(mai_mai_n372_), .B0(mai_mai_n370_), .B1(mai_mai_n368_), .Y(mai_mai_n376_));
  AN2        m0348(.A(j), .B(h), .Y(mai_mai_n377_));
  NO3        m0349(.A(n), .B(m), .C(k), .Y(mai_mai_n378_));
  NA2        m0350(.A(mai_mai_n378_), .B(mai_mai_n377_), .Y(mai_mai_n379_));
  NO3        m0351(.A(mai_mai_n379_), .B(mai_mai_n145_), .C(mai_mai_n206_), .Y(mai_mai_n380_));
  OR2        m0352(.A(m), .B(k), .Y(mai_mai_n381_));
  NO2        m0353(.A(mai_mai_n170_), .B(mai_mai_n381_), .Y(mai_mai_n382_));
  NA4        m0354(.A(n), .B(f), .C(c), .D(mai_mai_n113_), .Y(mai_mai_n383_));
  NOi21      m0355(.An(mai_mai_n382_), .B(mai_mai_n383_), .Y(mai_mai_n384_));
  NOi32      m0356(.An(d), .Bn(a), .C(c), .Y(mai_mai_n385_));
  NA2        m0357(.A(mai_mai_n385_), .B(mai_mai_n178_), .Y(mai_mai_n386_));
  NAi21      m0358(.An(i), .B(g), .Y(mai_mai_n387_));
  NAi31      m0359(.An(k), .B(m), .C(j), .Y(mai_mai_n388_));
  NO3        m0360(.A(mai_mai_n388_), .B(mai_mai_n387_), .C(n), .Y(mai_mai_n389_));
  NOi21      m0361(.An(mai_mai_n389_), .B(mai_mai_n386_), .Y(mai_mai_n390_));
  NO3        m0362(.A(mai_mai_n390_), .B(mai_mai_n384_), .C(mai_mai_n380_), .Y(mai_mai_n391_));
  NO2        m0363(.A(mai_mai_n383_), .B(mai_mai_n295_), .Y(mai_mai_n392_));
  NOi32      m0364(.An(f), .Bn(d), .C(c), .Y(mai_mai_n393_));
  NA2        m0365(.A(mai_mai_n392_), .B(mai_mai_n208_), .Y(mai_mai_n394_));
  NA3        m0366(.A(mai_mai_n394_), .B(mai_mai_n391_), .C(mai_mai_n376_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n59_), .B(mai_mai_n113_), .Y(mai_mai_n396_));
  NA2        m0368(.A(mai_mai_n243_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  INV        m0369(.A(e), .Y(mai_mai_n398_));
  NA2        m0370(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n399_));
  OAI220     m0371(.A0(mai_mai_n399_), .A1(mai_mai_n194_), .B0(mai_mai_n198_), .B1(mai_mai_n398_), .Y(mai_mai_n400_));
  AN2        m0372(.A(g), .B(e), .Y(mai_mai_n401_));
  NA3        m0373(.A(mai_mai_n401_), .B(mai_mai_n197_), .C(i), .Y(mai_mai_n402_));
  INV        m0374(.A(mai_mai_n402_), .Y(mai_mai_n403_));
  NO2        m0375(.A(mai_mai_n403_), .B(mai_mai_n400_), .Y(mai_mai_n404_));
  NOi32      m0376(.An(h), .Bn(e), .C(g), .Y(mai_mai_n405_));
  NA3        m0377(.A(mai_mai_n405_), .B(mai_mai_n288_), .C(m), .Y(mai_mai_n406_));
  NOi21      m0378(.An(g), .B(h), .Y(mai_mai_n407_));
  AN3        m0379(.A(m), .B(l), .C(i), .Y(mai_mai_n408_));
  AN3        m0380(.A(h), .B(g), .C(e), .Y(mai_mai_n409_));
  NA2        m0381(.A(mai_mai_n409_), .B(mai_mai_n95_), .Y(mai_mai_n410_));
  AN2        m0382(.A(mai_mai_n410_), .B(mai_mai_n406_), .Y(mai_mai_n411_));
  AOI210     m0383(.A0(mai_mai_n411_), .A1(mai_mai_n404_), .B0(mai_mai_n397_), .Y(mai_mai_n412_));
  NA3        m0384(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n413_), .B(mai_mai_n397_), .Y(mai_mai_n414_));
  NA3        m0386(.A(mai_mai_n385_), .B(mai_mai_n178_), .C(mai_mai_n81_), .Y(mai_mai_n415_));
  NAi31      m0387(.An(b), .B(c), .C(a), .Y(mai_mai_n416_));
  NO2        m0388(.A(mai_mai_n416_), .B(n), .Y(mai_mai_n417_));
  OAI210     m0389(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n418_));
  NO2        m0390(.A(mai_mai_n418_), .B(mai_mai_n142_), .Y(mai_mai_n419_));
  NA2        m0391(.A(mai_mai_n419_), .B(mai_mai_n417_), .Y(mai_mai_n420_));
  INV        m0392(.A(mai_mai_n420_), .Y(mai_mai_n421_));
  NO4        m0393(.A(mai_mai_n421_), .B(mai_mai_n414_), .C(mai_mai_n412_), .D(mai_mai_n395_), .Y(mai_mai_n422_));
  NA2        m0394(.A(i), .B(g), .Y(mai_mai_n423_));
  NO3        m0395(.A(mai_mai_n273_), .B(mai_mai_n423_), .C(c), .Y(mai_mai_n424_));
  NOi21      m0396(.An(a), .B(n), .Y(mai_mai_n425_));
  NOi21      m0397(.An(d), .B(c), .Y(mai_mai_n426_));
  NA2        m0398(.A(mai_mai_n426_), .B(mai_mai_n425_), .Y(mai_mai_n427_));
  NA3        m0399(.A(i), .B(g), .C(f), .Y(mai_mai_n428_));
  OR2        m0400(.A(mai_mai_n428_), .B(mai_mai_n71_), .Y(mai_mai_n429_));
  NA3        m0401(.A(mai_mai_n408_), .B(mai_mai_n407_), .C(mai_mai_n178_), .Y(mai_mai_n430_));
  AOI210     m0402(.A0(mai_mai_n430_), .A1(mai_mai_n429_), .B0(mai_mai_n427_), .Y(mai_mai_n431_));
  AOI210     m0403(.A0(mai_mai_n424_), .A1(mai_mai_n287_), .B0(mai_mai_n431_), .Y(mai_mai_n432_));
  OR2        m0404(.A(n), .B(m), .Y(mai_mai_n433_));
  NO2        m0405(.A(mai_mai_n433_), .B(mai_mai_n146_), .Y(mai_mai_n434_));
  NO2        m0406(.A(mai_mai_n179_), .B(mai_mai_n142_), .Y(mai_mai_n435_));
  OAI210     m0407(.A0(mai_mai_n434_), .A1(mai_mai_n172_), .B0(mai_mai_n435_), .Y(mai_mai_n436_));
  INV        m0408(.A(mai_mai_n361_), .Y(mai_mai_n437_));
  NA3        m0409(.A(mai_mai_n437_), .B(mai_mai_n351_), .C(d), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n416_), .B(mai_mai_n49_), .Y(mai_mai_n439_));
  NO3        m0411(.A(mai_mai_n66_), .B(mai_mai_n109_), .C(e), .Y(mai_mai_n440_));
  NAi21      m0412(.An(k), .B(j), .Y(mai_mai_n441_));
  NA3        m0413(.A(i), .B(mai_mai_n440_), .C(mai_mai_n439_), .Y(mai_mai_n442_));
  NAi21      m0414(.An(e), .B(d), .Y(mai_mai_n443_));
  INV        m0415(.A(mai_mai_n443_), .Y(mai_mai_n444_));
  NO2        m0416(.A(mai_mai_n247_), .B(mai_mai_n206_), .Y(mai_mai_n445_));
  NA3        m0417(.A(mai_mai_n445_), .B(mai_mai_n444_), .C(mai_mai_n220_), .Y(mai_mai_n446_));
  NA4        m0418(.A(mai_mai_n446_), .B(mai_mai_n442_), .C(mai_mai_n438_), .D(mai_mai_n436_), .Y(mai_mai_n447_));
  NOi31      m0419(.An(n), .B(m), .C(k), .Y(mai_mai_n448_));
  AOI220     m0420(.A0(mai_mai_n448_), .A1(mai_mai_n377_), .B0(mai_mai_n214_), .B1(mai_mai_n50_), .Y(mai_mai_n449_));
  NAi31      m0421(.An(g), .B(f), .C(c), .Y(mai_mai_n450_));
  NOi31      m0422(.An(mai_mai_n432_), .B(mai_mai_n447_), .C(mai_mai_n261_), .Y(mai_mai_n451_));
  NOi32      m0423(.An(c), .Bn(a), .C(b), .Y(mai_mai_n452_));
  NA2        m0424(.A(mai_mai_n452_), .B(mai_mai_n110_), .Y(mai_mai_n453_));
  INV        m0425(.A(mai_mai_n271_), .Y(mai_mai_n454_));
  AN2        m0426(.A(e), .B(d), .Y(mai_mai_n455_));
  NA2        m0427(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n456_));
  INV        m0428(.A(mai_mai_n142_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n128_), .B(mai_mai_n41_), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n459_));
  NOi31      m0431(.An(j), .B(k), .C(i), .Y(mai_mai_n460_));
  NOi21      m0432(.An(mai_mai_n160_), .B(mai_mai_n460_), .Y(mai_mai_n461_));
  NA4        m0433(.A(mai_mai_n315_), .B(mai_mai_n461_), .C(mai_mai_n255_), .D(mai_mai_n116_), .Y(mai_mai_n462_));
  AOI220     m0434(.A0(mai_mai_n462_), .A1(mai_mai_n459_), .B0(mai_mai_n458_), .B1(mai_mai_n457_), .Y(mai_mai_n463_));
  AOI210     m0435(.A0(mai_mai_n463_), .A1(mai_mai_n456_), .B0(mai_mai_n453_), .Y(mai_mai_n464_));
  NO2        m0436(.A(mai_mai_n202_), .B(mai_mai_n199_), .Y(mai_mai_n465_));
  NOi21      m0437(.An(a), .B(b), .Y(mai_mai_n466_));
  NA3        m0438(.A(e), .B(d), .C(c), .Y(mai_mai_n467_));
  NAi21      m0439(.An(mai_mai_n467_), .B(mai_mai_n466_), .Y(mai_mai_n468_));
  NO2        m0440(.A(mai_mai_n415_), .B(mai_mai_n198_), .Y(mai_mai_n469_));
  NOi21      m0441(.An(mai_mai_n468_), .B(mai_mai_n469_), .Y(mai_mai_n470_));
  AOI210     m0442(.A0(mai_mai_n264_), .A1(mai_mai_n465_), .B0(mai_mai_n470_), .Y(mai_mai_n471_));
  NO4        m0443(.A(mai_mai_n183_), .B(mai_mai_n101_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n472_));
  NA2        m0444(.A(mai_mai_n372_), .B(mai_mai_n147_), .Y(mai_mai_n473_));
  OR2        m0445(.A(k), .B(j), .Y(mai_mai_n474_));
  NA2        m0446(.A(l), .B(k), .Y(mai_mai_n475_));
  NA3        m0447(.A(mai_mai_n475_), .B(mai_mai_n474_), .C(mai_mai_n214_), .Y(mai_mai_n476_));
  AOI210     m0448(.A0(mai_mai_n227_), .A1(mai_mai_n330_), .B0(mai_mai_n81_), .Y(mai_mai_n477_));
  NOi21      m0449(.An(mai_mai_n476_), .B(mai_mai_n477_), .Y(mai_mai_n478_));
  OR3        m0450(.A(mai_mai_n478_), .B(mai_mai_n139_), .C(mai_mai_n131_), .Y(mai_mai_n479_));
  INV        m0451(.A(mai_mai_n125_), .Y(mai_mai_n480_));
  NA2        m0452(.A(mai_mai_n385_), .B(mai_mai_n110_), .Y(mai_mai_n481_));
  NO4        m0453(.A(mai_mai_n481_), .B(mai_mai_n92_), .C(mai_mai_n109_), .D(e), .Y(mai_mai_n482_));
  NO3        m0454(.A(mai_mai_n415_), .B(mai_mai_n89_), .C(mai_mai_n128_), .Y(mai_mai_n483_));
  NO4        m0455(.A(mai_mai_n483_), .B(mai_mai_n482_), .C(mai_mai_n480_), .D(mai_mai_n316_), .Y(mai_mai_n484_));
  NA3        m0456(.A(mai_mai_n484_), .B(mai_mai_n479_), .C(mai_mai_n473_), .Y(mai_mai_n485_));
  NO4        m0457(.A(mai_mai_n485_), .B(mai_mai_n472_), .C(mai_mai_n471_), .D(mai_mai_n464_), .Y(mai_mai_n486_));
  NA2        m0458(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n487_));
  NOi21      m0459(.An(d), .B(e), .Y(mai_mai_n488_));
  NO2        m0460(.A(mai_mai_n183_), .B(mai_mai_n56_), .Y(mai_mai_n489_));
  NAi31      m0461(.An(j), .B(l), .C(i), .Y(mai_mai_n490_));
  OAI210     m0462(.A0(mai_mai_n490_), .A1(mai_mai_n129_), .B0(mai_mai_n101_), .Y(mai_mai_n491_));
  NA3        m0463(.A(mai_mai_n491_), .B(mai_mai_n489_), .C(mai_mai_n488_), .Y(mai_mai_n492_));
  NO3        m0464(.A(mai_mai_n386_), .B(mai_mai_n334_), .C(mai_mai_n195_), .Y(mai_mai_n493_));
  NO2        m0465(.A(mai_mai_n386_), .B(mai_mai_n361_), .Y(mai_mai_n494_));
  NO3        m0466(.A(mai_mai_n494_), .B(mai_mai_n493_), .C(mai_mai_n303_), .Y(mai_mai_n495_));
  NA4        m0467(.A(mai_mai_n495_), .B(mai_mai_n492_), .C(mai_mai_n487_), .D(mai_mai_n237_), .Y(mai_mai_n496_));
  OAI210     m0468(.A0(mai_mai_n124_), .A1(mai_mai_n123_), .B0(n), .Y(mai_mai_n497_));
  NO2        m0469(.A(mai_mai_n497_), .B(mai_mai_n128_), .Y(mai_mai_n498_));
  XO2        m0470(.A(i), .B(h), .Y(mai_mai_n499_));
  NA3        m0471(.A(mai_mai_n499_), .B(mai_mai_n154_), .C(n), .Y(mai_mai_n500_));
  NAi41      m0472(.An(mai_mai_n296_), .B(mai_mai_n500_), .C(mai_mai_n449_), .D(mai_mai_n374_), .Y(mai_mai_n501_));
  NAi31      m0473(.An(c), .B(f), .C(d), .Y(mai_mai_n502_));
  AOI210     m0474(.A0(mai_mai_n276_), .A1(mai_mai_n189_), .B0(mai_mai_n502_), .Y(mai_mai_n503_));
  INV        m0475(.A(mai_mai_n503_), .Y(mai_mai_n504_));
  NA3        m0476(.A(mai_mai_n370_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n505_));
  NA2        m0477(.A(mai_mai_n221_), .B(mai_mai_n105_), .Y(mai_mai_n506_));
  AOI210     m0478(.A0(mai_mai_n506_), .A1(mai_mai_n177_), .B0(mai_mai_n502_), .Y(mai_mai_n507_));
  AOI210     m0479(.A0(mai_mai_n349_), .A1(mai_mai_n35_), .B0(mai_mai_n468_), .Y(mai_mai_n508_));
  NOi31      m0480(.An(mai_mai_n505_), .B(mai_mai_n508_), .C(mai_mai_n507_), .Y(mai_mai_n509_));
  AO220      m0481(.A0(mai_mai_n284_), .A1(mai_mai_n258_), .B0(mai_mai_n161_), .B1(mai_mai_n67_), .Y(mai_mai_n510_));
  NA3        m0482(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n511_), .B(mai_mai_n427_), .Y(mai_mai_n512_));
  NO2        m0484(.A(mai_mai_n512_), .B(mai_mai_n292_), .Y(mai_mai_n513_));
  NAi41      m0485(.An(mai_mai_n510_), .B(mai_mai_n513_), .C(mai_mai_n509_), .D(mai_mai_n504_), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n514_), .B(mai_mai_n496_), .Y(mai_mai_n515_));
  NA4        m0487(.A(mai_mai_n515_), .B(mai_mai_n486_), .C(mai_mai_n451_), .D(mai_mai_n422_), .Y(mai11));
  NO2        m0488(.A(mai_mai_n72_), .B(f), .Y(mai_mai_n517_));
  NA2        m0489(.A(j), .B(g), .Y(mai_mai_n518_));
  NAi31      m0490(.An(i), .B(m), .C(l), .Y(mai_mai_n519_));
  NA3        m0491(.A(m), .B(k), .C(j), .Y(mai_mai_n520_));
  OAI220     m0492(.A0(mai_mai_n520_), .A1(mai_mai_n128_), .B0(mai_mai_n519_), .B1(mai_mai_n518_), .Y(mai_mai_n521_));
  NA2        m0493(.A(mai_mai_n521_), .B(mai_mai_n517_), .Y(mai_mai_n522_));
  NOi32      m0494(.An(e), .Bn(b), .C(f), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n254_), .B(mai_mai_n110_), .Y(mai_mai_n524_));
  NA2        m0496(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n525_));
  NO2        m0497(.A(mai_mai_n525_), .B(mai_mai_n298_), .Y(mai_mai_n526_));
  NAi31      m0498(.An(d), .B(e), .C(a), .Y(mai_mai_n527_));
  NO2        m0499(.A(mai_mai_n527_), .B(n), .Y(mai_mai_n528_));
  AOI220     m0500(.A0(mai_mai_n528_), .A1(mai_mai_n99_), .B0(mai_mai_n526_), .B1(mai_mai_n523_), .Y(mai_mai_n529_));
  NAi41      m0501(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n530_));
  AN2        m0502(.A(mai_mai_n530_), .B(mai_mai_n360_), .Y(mai_mai_n531_));
  AOI210     m0503(.A0(mai_mai_n531_), .A1(mai_mai_n386_), .B0(mai_mai_n267_), .Y(mai_mai_n532_));
  NA2        m0504(.A(j), .B(i), .Y(mai_mai_n533_));
  NAi31      m0505(.An(n), .B(m), .C(k), .Y(mai_mai_n534_));
  NO3        m0506(.A(mai_mai_n534_), .B(mai_mai_n533_), .C(mai_mai_n109_), .Y(mai_mai_n535_));
  NO4        m0507(.A(n), .B(d), .C(mai_mai_n113_), .D(a), .Y(mai_mai_n536_));
  OR2        m0508(.A(n), .B(c), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n537_), .B(mai_mai_n144_), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n538_), .B(mai_mai_n536_), .Y(mai_mai_n539_));
  NOi32      m0511(.An(g), .Bn(f), .C(i), .Y(mai_mai_n540_));
  AOI220     m0512(.A0(mai_mai_n540_), .A1(mai_mai_n97_), .B0(mai_mai_n521_), .B1(f), .Y(mai_mai_n541_));
  NO2        m0513(.A(mai_mai_n271_), .B(mai_mai_n49_), .Y(mai_mai_n542_));
  NO2        m0514(.A(mai_mai_n541_), .B(mai_mai_n539_), .Y(mai_mai_n543_));
  AOI210     m0515(.A0(mai_mai_n535_), .A1(mai_mai_n532_), .B0(mai_mai_n543_), .Y(mai_mai_n544_));
  NA2        m0516(.A(mai_mai_n136_), .B(mai_mai_n34_), .Y(mai_mai_n545_));
  NAi32      m0517(.An(e), .Bn(b), .C(c), .Y(mai_mai_n546_));
  OR2        m0518(.A(mai_mai_n546_), .B(mai_mai_n81_), .Y(mai_mai_n547_));
  OAI220     m0519(.A0(mai_mai_n388_), .A1(mai_mai_n387_), .B0(mai_mai_n519_), .B1(mai_mai_n518_), .Y(mai_mai_n548_));
  NAi31      m0520(.An(d), .B(c), .C(a), .Y(mai_mai_n549_));
  NO2        m0521(.A(mai_mai_n549_), .B(n), .Y(mai_mai_n550_));
  NA3        m0522(.A(mai_mai_n550_), .B(mai_mai_n548_), .C(e), .Y(mai_mai_n551_));
  NO3        m0523(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n207_), .Y(mai_mai_n552_));
  NO2        m0524(.A(mai_mai_n224_), .B(mai_mai_n107_), .Y(mai_mai_n553_));
  OAI210     m0525(.A0(mai_mai_n552_), .A1(mai_mai_n389_), .B0(mai_mai_n553_), .Y(mai_mai_n554_));
  NA2        m0526(.A(mai_mai_n554_), .B(mai_mai_n551_), .Y(mai_mai_n555_));
  NO2        m0527(.A(mai_mai_n273_), .B(n), .Y(mai_mai_n556_));
  NO2        m0528(.A(mai_mai_n417_), .B(mai_mai_n556_), .Y(mai_mai_n557_));
  NA2        m0529(.A(mai_mai_n548_), .B(f), .Y(mai_mai_n558_));
  NAi32      m0530(.An(d), .Bn(a), .C(b), .Y(mai_mai_n559_));
  NO2        m0531(.A(mai_mai_n559_), .B(mai_mai_n49_), .Y(mai_mai_n560_));
  NA2        m0532(.A(h), .B(f), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n561_), .B(mai_mai_n92_), .Y(mai_mai_n562_));
  NA2        m0534(.A(mai_mai_n562_), .B(mai_mai_n560_), .Y(mai_mai_n563_));
  OAI210     m0535(.A0(mai_mai_n558_), .A1(mai_mai_n557_), .B0(mai_mai_n563_), .Y(mai_mai_n564_));
  AN3        m0536(.A(j), .B(h), .C(g), .Y(mai_mai_n565_));
  NA3        m0537(.A(f), .B(d), .C(b), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n564_), .B(mai_mai_n555_), .Y(mai_mai_n567_));
  AN4        m0539(.A(mai_mai_n567_), .B(mai_mai_n544_), .C(mai_mai_n529_), .D(mai_mai_n522_), .Y(mai_mai_n568_));
  INV        m0540(.A(k), .Y(mai_mai_n569_));
  NA3        m0541(.A(l), .B(mai_mai_n569_), .C(i), .Y(mai_mai_n570_));
  INV        m0542(.A(mai_mai_n570_), .Y(mai_mai_n571_));
  NA4        m0543(.A(mai_mai_n385_), .B(mai_mai_n407_), .C(mai_mai_n178_), .D(mai_mai_n110_), .Y(mai_mai_n572_));
  NAi32      m0544(.An(h), .Bn(f), .C(g), .Y(mai_mai_n573_));
  NAi41      m0545(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n574_));
  OAI210     m0546(.A0(mai_mai_n527_), .A1(n), .B0(mai_mai_n574_), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n575_), .B(m), .Y(mai_mai_n576_));
  NAi31      m0548(.An(h), .B(g), .C(f), .Y(mai_mai_n577_));
  OR3        m0549(.A(mai_mai_n577_), .B(mai_mai_n273_), .C(mai_mai_n49_), .Y(mai_mai_n578_));
  NA4        m0550(.A(mai_mai_n407_), .B(mai_mai_n118_), .C(mai_mai_n110_), .D(e), .Y(mai_mai_n579_));
  AN2        m0551(.A(mai_mai_n579_), .B(mai_mai_n578_), .Y(mai_mai_n580_));
  OA210      m0552(.A0(mai_mai_n576_), .A1(mai_mai_n573_), .B0(mai_mai_n580_), .Y(mai_mai_n581_));
  NO3        m0553(.A(mai_mai_n573_), .B(mai_mai_n72_), .C(mai_mai_n74_), .Y(mai_mai_n582_));
  NO4        m0554(.A(mai_mai_n577_), .B(mai_mai_n537_), .C(mai_mai_n144_), .D(mai_mai_n74_), .Y(mai_mai_n583_));
  OR2        m0555(.A(mai_mai_n583_), .B(mai_mai_n582_), .Y(mai_mai_n584_));
  NAi31      m0556(.An(mai_mai_n584_), .B(mai_mai_n581_), .C(mai_mai_n572_), .Y(mai_mai_n585_));
  NAi31      m0557(.An(f), .B(h), .C(g), .Y(mai_mai_n586_));
  NO4        m0558(.A(mai_mai_n306_), .B(mai_mai_n586_), .C(mai_mai_n72_), .D(mai_mai_n74_), .Y(mai_mai_n587_));
  NOi32      m0559(.An(b), .Bn(a), .C(c), .Y(mai_mai_n588_));
  NOi41      m0560(.An(mai_mai_n588_), .B(mai_mai_n343_), .C(mai_mai_n69_), .D(mai_mai_n114_), .Y(mai_mai_n589_));
  OR2        m0561(.A(mai_mai_n589_), .B(mai_mai_n587_), .Y(mai_mai_n590_));
  NOi32      m0562(.An(d), .Bn(a), .C(e), .Y(mai_mai_n591_));
  NA2        m0563(.A(mai_mai_n591_), .B(mai_mai_n110_), .Y(mai_mai_n592_));
  NO2        m0564(.A(n), .B(c), .Y(mai_mai_n593_));
  NA3        m0565(.A(mai_mai_n593_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n594_));
  NAi32      m0566(.An(n), .Bn(f), .C(m), .Y(mai_mai_n595_));
  NA3        m0567(.A(mai_mai_n595_), .B(mai_mai_n594_), .C(mai_mai_n592_), .Y(mai_mai_n596_));
  NOi32      m0568(.An(e), .Bn(a), .C(d), .Y(mai_mai_n597_));
  AOI210     m0569(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n597_), .Y(mai_mai_n598_));
  AOI210     m0570(.A0(mai_mai_n598_), .A1(mai_mai_n206_), .B0(mai_mai_n545_), .Y(mai_mai_n599_));
  AOI210     m0571(.A0(mai_mai_n599_), .A1(mai_mai_n596_), .B0(mai_mai_n590_), .Y(mai_mai_n600_));
  OAI210     m0572(.A0(mai_mai_n242_), .A1(mai_mai_n84_), .B0(mai_mai_n600_), .Y(mai_mai_n601_));
  AOI210     m0573(.A0(mai_mai_n585_), .A1(mai_mai_n571_), .B0(mai_mai_n601_), .Y(mai_mai_n602_));
  NO3        m0574(.A(mai_mai_n313_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n603_));
  NA3        m0575(.A(mai_mai_n502_), .B(mai_mai_n168_), .C(mai_mai_n167_), .Y(mai_mai_n604_));
  NA2        m0576(.A(mai_mai_n450_), .B(mai_mai_n224_), .Y(mai_mai_n605_));
  OR2        m0577(.A(mai_mai_n605_), .B(mai_mai_n604_), .Y(mai_mai_n606_));
  NA2        m0578(.A(mai_mai_n75_), .B(mai_mai_n110_), .Y(mai_mai_n607_));
  NO2        m0579(.A(mai_mai_n607_), .B(mai_mai_n45_), .Y(mai_mai_n608_));
  AOI220     m0580(.A0(mai_mai_n608_), .A1(mai_mai_n532_), .B0(mai_mai_n606_), .B1(mai_mai_n603_), .Y(mai_mai_n609_));
  NO2        m0581(.A(mai_mai_n609_), .B(mai_mai_n84_), .Y(mai_mai_n610_));
  NOi32      m0582(.An(e), .Bn(c), .C(f), .Y(mai_mai_n611_));
  NOi21      m0583(.An(f), .B(g), .Y(mai_mai_n612_));
  NO2        m0584(.A(mai_mai_n612_), .B(mai_mai_n204_), .Y(mai_mai_n613_));
  NA2        m0585(.A(mai_mai_n611_), .B(mai_mai_n172_), .Y(mai_mai_n614_));
  NA2        m0586(.A(mai_mai_n614_), .B(mai_mai_n175_), .Y(mai_mai_n615_));
  AOI210     m0587(.A0(mai_mai_n531_), .A1(mai_mai_n386_), .B0(mai_mai_n297_), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n616_), .B(mai_mai_n259_), .Y(mai_mai_n617_));
  NOi21      m0589(.An(j), .B(l), .Y(mai_mai_n618_));
  NAi21      m0590(.An(k), .B(h), .Y(mai_mai_n619_));
  NO2        m0591(.A(mai_mai_n619_), .B(mai_mai_n257_), .Y(mai_mai_n620_));
  NA2        m0592(.A(mai_mai_n620_), .B(mai_mai_n618_), .Y(mai_mai_n621_));
  OR2        m0593(.A(mai_mai_n621_), .B(mai_mai_n576_), .Y(mai_mai_n622_));
  NOi31      m0594(.An(m), .B(n), .C(k), .Y(mai_mai_n623_));
  NA2        m0595(.A(mai_mai_n618_), .B(mai_mai_n623_), .Y(mai_mai_n624_));
  AOI210     m0596(.A0(mai_mai_n386_), .A1(mai_mai_n360_), .B0(mai_mai_n297_), .Y(mai_mai_n625_));
  NAi21      m0597(.An(mai_mai_n624_), .B(mai_mai_n625_), .Y(mai_mai_n626_));
  NO2        m0598(.A(mai_mai_n273_), .B(mai_mai_n49_), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n306_), .B(mai_mai_n586_), .Y(mai_mai_n628_));
  NO2        m0600(.A(mai_mai_n527_), .B(mai_mai_n49_), .Y(mai_mai_n629_));
  AOI220     m0601(.A0(mai_mai_n629_), .A1(mai_mai_n628_), .B0(mai_mai_n627_), .B1(mai_mai_n562_), .Y(mai_mai_n630_));
  NA4        m0602(.A(mai_mai_n630_), .B(mai_mai_n626_), .C(mai_mai_n622_), .D(mai_mai_n617_), .Y(mai_mai_n631_));
  NA2        m0603(.A(mai_mai_n105_), .B(mai_mai_n36_), .Y(mai_mai_n632_));
  NO2        m0604(.A(mai_mai_n523_), .B(mai_mai_n351_), .Y(mai_mai_n633_));
  NO2        m0605(.A(mai_mai_n633_), .B(n), .Y(mai_mai_n634_));
  NA2        m0606(.A(mai_mai_n546_), .B(mai_mai_n140_), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n499_), .B(mai_mai_n154_), .Y(mai_mai_n636_));
  NO3        m0608(.A(mai_mai_n383_), .B(mai_mai_n636_), .C(mai_mai_n84_), .Y(mai_mai_n637_));
  INV        m0609(.A(mai_mai_n637_), .Y(mai_mai_n638_));
  AN3        m0610(.A(f), .B(d), .C(b), .Y(mai_mai_n639_));
  NA3        m0611(.A(mai_mai_n499_), .B(mai_mai_n154_), .C(mai_mai_n207_), .Y(mai_mai_n640_));
  NO2        m0612(.A(mai_mai_n226_), .B(mai_mai_n640_), .Y(mai_mai_n641_));
  NAi31      m0613(.An(m), .B(n), .C(k), .Y(mai_mai_n642_));
  OR2        m0614(.A(mai_mai_n131_), .B(mai_mai_n61_), .Y(mai_mai_n643_));
  OAI210     m0615(.A0(mai_mai_n643_), .A1(mai_mai_n642_), .B0(mai_mai_n244_), .Y(mai_mai_n644_));
  OAI210     m0616(.A0(mai_mai_n644_), .A1(mai_mai_n641_), .B0(j), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n645_), .B(mai_mai_n638_), .Y(mai_mai_n646_));
  NO4        m0618(.A(mai_mai_n646_), .B(mai_mai_n631_), .C(mai_mai_n615_), .D(mai_mai_n610_), .Y(mai_mai_n647_));
  NAi31      m0619(.An(g), .B(h), .C(f), .Y(mai_mai_n648_));
  OR3        m0620(.A(mai_mai_n648_), .B(mai_mai_n273_), .C(n), .Y(mai_mai_n649_));
  OA210      m0621(.A0(mai_mai_n527_), .A1(n), .B0(mai_mai_n574_), .Y(mai_mai_n650_));
  NA3        m0622(.A(mai_mai_n405_), .B(mai_mai_n118_), .C(mai_mai_n81_), .Y(mai_mai_n651_));
  OAI210     m0623(.A0(mai_mai_n650_), .A1(mai_mai_n88_), .B0(mai_mai_n651_), .Y(mai_mai_n652_));
  NOi21      m0624(.An(mai_mai_n649_), .B(mai_mai_n652_), .Y(mai_mai_n653_));
  NO2        m0625(.A(mai_mai_n653_), .B(mai_mai_n520_), .Y(mai_mai_n654_));
  NO3        m0626(.A(g), .B(mai_mai_n206_), .C(mai_mai_n56_), .Y(mai_mai_n655_));
  NO2        m0627(.A(mai_mai_n506_), .B(mai_mai_n84_), .Y(mai_mai_n656_));
  OAI210     m0628(.A0(mai_mai_n656_), .A1(mai_mai_n382_), .B0(mai_mai_n655_), .Y(mai_mai_n657_));
  OR2        m0629(.A(mai_mai_n72_), .B(mai_mai_n74_), .Y(mai_mai_n658_));
  NA2        m0630(.A(mai_mai_n588_), .B(mai_mai_n332_), .Y(mai_mai_n659_));
  OA220      m0631(.A0(mai_mai_n624_), .A1(mai_mai_n659_), .B0(mai_mai_n621_), .B1(mai_mai_n658_), .Y(mai_mai_n660_));
  NA3        m0632(.A(mai_mai_n517_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n661_));
  AN2        m0633(.A(h), .B(f), .Y(mai_mai_n662_));
  NA2        m0634(.A(mai_mai_n662_), .B(mai_mai_n37_), .Y(mai_mai_n663_));
  NO2        m0635(.A(mai_mai_n663_), .B(mai_mai_n453_), .Y(mai_mai_n664_));
  AOI210     m0636(.A0(mai_mai_n559_), .A1(mai_mai_n416_), .B0(mai_mai_n49_), .Y(mai_mai_n665_));
  OAI220     m0637(.A0(mai_mai_n577_), .A1(mai_mai_n570_), .B0(mai_mai_n320_), .B1(mai_mai_n518_), .Y(mai_mai_n666_));
  AOI210     m0638(.A0(mai_mai_n666_), .A1(mai_mai_n665_), .B0(mai_mai_n664_), .Y(mai_mai_n667_));
  NA4        m0639(.A(mai_mai_n667_), .B(mai_mai_n661_), .C(mai_mai_n660_), .D(mai_mai_n657_), .Y(mai_mai_n668_));
  NO2        m0640(.A(mai_mai_n246_), .B(f), .Y(mai_mai_n669_));
  INV        m0641(.A(mai_mai_n61_), .Y(mai_mai_n670_));
  NO3        m0642(.A(mai_mai_n670_), .B(mai_mai_n669_), .C(mai_mai_n34_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n323_), .B(mai_mai_n136_), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n129_), .B(mai_mai_n49_), .Y(mai_mai_n673_));
  NA2        m0645(.A(mai_mai_n673_), .B(mai_mai_n523_), .Y(mai_mai_n674_));
  OA220      m0646(.A0(mai_mai_n674_), .A1(mai_mai_n545_), .B0(mai_mai_n349_), .B1(mai_mai_n108_), .Y(mai_mai_n675_));
  OAI210     m0647(.A0(mai_mai_n672_), .A1(mai_mai_n671_), .B0(mai_mai_n675_), .Y(mai_mai_n676_));
  NO3        m0648(.A(mai_mai_n393_), .B(mai_mai_n186_), .C(mai_mai_n185_), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n677_), .B(mai_mai_n224_), .Y(mai_mai_n678_));
  NA3        m0650(.A(mai_mai_n678_), .B(mai_mai_n248_), .C(j), .Y(mai_mai_n679_));
  NA2        m0651(.A(mai_mai_n452_), .B(mai_mai_n81_), .Y(mai_mai_n680_));
  NO4        m0652(.A(mai_mai_n520_), .B(mai_mai_n680_), .C(mai_mai_n128_), .D(mai_mai_n206_), .Y(mai_mai_n681_));
  INV        m0653(.A(mai_mai_n681_), .Y(mai_mai_n682_));
  NA4        m0654(.A(mai_mai_n682_), .B(mai_mai_n679_), .C(mai_mai_n505_), .D(mai_mai_n391_), .Y(mai_mai_n683_));
  NO4        m0655(.A(mai_mai_n683_), .B(mai_mai_n676_), .C(mai_mai_n668_), .D(mai_mai_n654_), .Y(mai_mai_n684_));
  NA4        m0656(.A(mai_mai_n684_), .B(mai_mai_n647_), .C(mai_mai_n602_), .D(mai_mai_n568_), .Y(mai08));
  NO2        m0657(.A(k), .B(h), .Y(mai_mai_n686_));
  AO210      m0658(.A0(mai_mai_n246_), .A1(mai_mai_n441_), .B0(mai_mai_n686_), .Y(mai_mai_n687_));
  NO2        m0659(.A(mai_mai_n687_), .B(mai_mai_n295_), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n611_), .B(mai_mai_n81_), .Y(mai_mai_n689_));
  NA2        m0661(.A(mai_mai_n689_), .B(mai_mai_n450_), .Y(mai_mai_n690_));
  AOI210     m0662(.A0(mai_mai_n690_), .A1(mai_mai_n688_), .B0(mai_mai_n483_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n81_), .B(mai_mai_n107_), .Y(mai_mai_n692_));
  NO2        m0664(.A(mai_mai_n692_), .B(mai_mai_n57_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n566_), .B(mai_mai_n226_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n337_), .Y(mai_mai_n695_));
  NA4        m0667(.A(mai_mai_n209_), .B(mai_mai_n136_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n696_));
  AN2        m0668(.A(l), .B(k), .Y(mai_mai_n697_));
  NA3        m0669(.A(mai_mai_n695_), .B(mai_mai_n691_), .C(mai_mai_n339_), .Y(mai_mai_n698_));
  AN2        m0670(.A(mai_mai_n528_), .B(mai_mai_n93_), .Y(mai_mai_n699_));
  NO4        m0671(.A(mai_mai_n170_), .B(mai_mai_n381_), .C(mai_mai_n109_), .D(g), .Y(mai_mai_n700_));
  INV        m0672(.A(mai_mai_n512_), .Y(mai_mai_n701_));
  NO2        m0673(.A(mai_mai_n38_), .B(mai_mai_n206_), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n702_), .B(mai_mai_n556_), .Y(mai_mai_n703_));
  NAi31      m0675(.An(mai_mai_n699_), .B(mai_mai_n703_), .C(mai_mai_n701_), .Y(mai_mai_n704_));
  NO2        m0676(.A(mai_mai_n531_), .B(mai_mai_n35_), .Y(mai_mai_n705_));
  OAI210     m0677(.A0(mai_mai_n546_), .A1(mai_mai_n47_), .B0(mai_mai_n643_), .Y(mai_mai_n706_));
  NO2        m0678(.A(mai_mai_n475_), .B(mai_mai_n129_), .Y(mai_mai_n707_));
  AOI210     m0679(.A0(mai_mai_n707_), .A1(mai_mai_n706_), .B0(mai_mai_n705_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n687_), .B(mai_mai_n132_), .Y(mai_mai_n709_));
  NA2        m0681(.A(mai_mai_n709_), .B(mai_mai_n392_), .Y(mai_mai_n710_));
  NA2        m0682(.A(mai_mai_n708_), .B(mai_mai_n710_), .Y(mai_mai_n711_));
  NA2        m0683(.A(mai_mai_n351_), .B(mai_mai_n43_), .Y(mai_mai_n712_));
  NA3        m0684(.A(mai_mai_n678_), .B(mai_mai_n328_), .C(mai_mai_n373_), .Y(mai_mai_n713_));
  NA2        m0685(.A(mai_mai_n697_), .B(mai_mai_n214_), .Y(mai_mai_n714_));
  NO2        m0686(.A(mai_mai_n714_), .B(mai_mai_n322_), .Y(mai_mai_n715_));
  AOI210     m0687(.A0(mai_mai_n715_), .A1(mai_mai_n669_), .B0(mai_mai_n482_), .Y(mai_mai_n716_));
  NA3        m0688(.A(m), .B(l), .C(k), .Y(mai_mai_n717_));
  AOI210     m0689(.A0(mai_mai_n651_), .A1(mai_mai_n649_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  NO2        m0690(.A(mai_mai_n530_), .B(mai_mai_n267_), .Y(mai_mai_n719_));
  NOi21      m0691(.An(mai_mai_n719_), .B(mai_mai_n524_), .Y(mai_mai_n720_));
  NA4        m0692(.A(mai_mai_n110_), .B(l), .C(k), .D(mai_mai_n84_), .Y(mai_mai_n721_));
  NA3        m0693(.A(mai_mai_n118_), .B(mai_mai_n401_), .C(i), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n722_), .B(mai_mai_n721_), .Y(mai_mai_n723_));
  NO3        m0695(.A(mai_mai_n723_), .B(mai_mai_n720_), .C(mai_mai_n718_), .Y(mai_mai_n724_));
  NA4        m0696(.A(mai_mai_n724_), .B(mai_mai_n716_), .C(mai_mai_n713_), .D(mai_mai_n712_), .Y(mai_mai_n725_));
  NO4        m0697(.A(mai_mai_n725_), .B(mai_mai_n711_), .C(mai_mai_n704_), .D(mai_mai_n698_), .Y(mai_mai_n726_));
  NOi31      m0698(.An(g), .B(h), .C(f), .Y(mai_mai_n727_));
  NA2        m0699(.A(mai_mai_n629_), .B(mai_mai_n727_), .Y(mai_mai_n728_));
  OR2        m0700(.A(mai_mai_n728_), .B(mai_mai_n533_), .Y(mai_mai_n729_));
  NO3        m0701(.A(mai_mai_n386_), .B(mai_mai_n518_), .C(h), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n730_), .B(mai_mai_n110_), .Y(mai_mai_n731_));
  NA3        m0703(.A(mai_mai_n731_), .B(mai_mai_n729_), .C(mai_mai_n245_), .Y(mai_mai_n732_));
  NA2        m0704(.A(mai_mai_n697_), .B(mai_mai_n74_), .Y(mai_mai_n733_));
  NO3        m0705(.A(mai_mai_n677_), .B(mai_mai_n170_), .C(i), .Y(mai_mai_n734_));
  NOi21      m0706(.An(h), .B(j), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n735_), .B(f), .Y(mai_mai_n736_));
  NO2        m0708(.A(mai_mai_n736_), .B(mai_mai_n239_), .Y(mai_mai_n737_));
  NO2        m0709(.A(mai_mai_n737_), .B(mai_mai_n734_), .Y(mai_mai_n738_));
  OAI220     m0710(.A0(mai_mai_n738_), .A1(mai_mai_n733_), .B0(mai_mai_n580_), .B1(mai_mai_n62_), .Y(mai_mai_n739_));
  AOI210     m0711(.A0(mai_mai_n732_), .A1(l), .B0(mai_mai_n739_), .Y(mai_mai_n740_));
  NO2        m0712(.A(j), .B(i), .Y(mai_mai_n741_));
  NA3        m0713(.A(mai_mai_n741_), .B(mai_mai_n79_), .C(l), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n741_), .B(mai_mai_n33_), .Y(mai_mai_n743_));
  NA2        m0715(.A(mai_mai_n409_), .B(mai_mai_n118_), .Y(mai_mai_n744_));
  OA220      m0716(.A0(mai_mai_n744_), .A1(mai_mai_n743_), .B0(mai_mai_n742_), .B1(mai_mai_n576_), .Y(mai_mai_n745_));
  NO3        m0717(.A(mai_mai_n145_), .B(mai_mai_n49_), .C(mai_mai_n107_), .Y(mai_mai_n746_));
  NO3        m0718(.A(mai_mai_n537_), .B(mai_mai_n144_), .C(mai_mai_n74_), .Y(mai_mai_n747_));
  NO2        m0719(.A(mai_mai_n475_), .B(mai_mai_n428_), .Y(mai_mai_n748_));
  OAI210     m0720(.A0(mai_mai_n747_), .A1(mai_mai_n746_), .B0(mai_mai_n748_), .Y(mai_mai_n749_));
  OAI210     m0721(.A0(mai_mai_n728_), .A1(mai_mai_n62_), .B0(mai_mai_n749_), .Y(mai_mai_n750_));
  NA2        m0722(.A(k), .B(j), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n523_), .B(n), .Y(mai_mai_n752_));
  NO3        m0724(.A(mai_mai_n170_), .B(mai_mai_n381_), .C(mai_mai_n109_), .Y(mai_mai_n753_));
  NA2        m0725(.A(mai_mai_n753_), .B(mai_mai_n240_), .Y(mai_mai_n754_));
  NAi31      m0726(.An(mai_mai_n598_), .B(mai_mai_n90_), .C(mai_mai_n81_), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n755_), .B(mai_mai_n754_), .Y(mai_mai_n756_));
  NO2        m0728(.A(mai_mai_n295_), .B(mai_mai_n132_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n717_), .B(mai_mai_n88_), .Y(mai_mai_n758_));
  NO2        m0730(.A(mai_mai_n577_), .B(mai_mai_n114_), .Y(mai_mai_n759_));
  OAI210     m0731(.A0(mai_mai_n759_), .A1(mai_mai_n748_), .B0(mai_mai_n665_), .Y(mai_mai_n760_));
  INV        m0732(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  OR3        m0733(.A(mai_mai_n761_), .B(mai_mai_n756_), .C(mai_mai_n750_), .Y(mai_mai_n762_));
  NA3        m0734(.A(mai_mai_n752_), .B(mai_mai_n331_), .C(mai_mai_n547_), .Y(mai_mai_n763_));
  NA4        m0735(.A(mai_mai_n763_), .B(mai_mai_n209_), .C(mai_mai_n441_), .D(mai_mai_n34_), .Y(mai_mai_n764_));
  NO4        m0736(.A(mai_mai_n475_), .B(mai_mai_n423_), .C(j), .D(f), .Y(mai_mai_n765_));
  OAI220     m0737(.A0(mai_mai_n696_), .A1(mai_mai_n689_), .B0(mai_mai_n326_), .B1(mai_mai_n38_), .Y(mai_mai_n766_));
  AOI210     m0738(.A0(mai_mai_n765_), .A1(mai_mai_n252_), .B0(mai_mai_n766_), .Y(mai_mai_n767_));
  NA3        m0739(.A(mai_mai_n540_), .B(mai_mai_n288_), .C(h), .Y(mai_mai_n768_));
  NOi21      m0740(.An(mai_mai_n665_), .B(mai_mai_n768_), .Y(mai_mai_n769_));
  NO2        m0741(.A(mai_mai_n89_), .B(mai_mai_n47_), .Y(mai_mai_n770_));
  OAI220     m0742(.A0(mai_mai_n768_), .A1(mai_mai_n594_), .B0(mai_mai_n742_), .B1(mai_mai_n658_), .Y(mai_mai_n771_));
  AOI210     m0743(.A0(mai_mai_n770_), .A1(mai_mai_n634_), .B0(mai_mai_n771_), .Y(mai_mai_n772_));
  NAi41      m0744(.An(mai_mai_n769_), .B(mai_mai_n772_), .C(mai_mai_n767_), .D(mai_mai_n764_), .Y(mai_mai_n773_));
  OR2        m0745(.A(mai_mai_n758_), .B(mai_mai_n93_), .Y(mai_mai_n774_));
  AOI220     m0746(.A0(mai_mai_n774_), .A1(mai_mai_n232_), .B0(mai_mai_n748_), .B1(mai_mai_n627_), .Y(mai_mai_n775_));
  NO2        m0747(.A(mai_mai_n650_), .B(mai_mai_n74_), .Y(mai_mai_n776_));
  NA2        m0748(.A(mai_mai_n765_), .B(mai_mai_n776_), .Y(mai_mai_n777_));
  OAI210     m0749(.A0(mai_mai_n717_), .A1(mai_mai_n648_), .B0(mai_mai_n511_), .Y(mai_mai_n778_));
  NA3        m0750(.A(mai_mai_n243_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n779_));
  AOI220     m0751(.A0(mai_mai_n593_), .A1(mai_mai_n29_), .B0(mai_mai_n452_), .B1(mai_mai_n81_), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n780_), .B(mai_mai_n779_), .Y(mai_mai_n781_));
  NO2        m0753(.A(mai_mai_n768_), .B(mai_mai_n481_), .Y(mai_mai_n782_));
  AOI210     m0754(.A0(mai_mai_n781_), .A1(mai_mai_n778_), .B0(mai_mai_n782_), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n783_), .B(mai_mai_n777_), .C(mai_mai_n775_), .Y(mai_mai_n784_));
  NOi41      m0756(.An(mai_mai_n745_), .B(mai_mai_n784_), .C(mai_mai_n773_), .D(mai_mai_n762_), .Y(mai_mai_n785_));
  OR2        m0757(.A(mai_mai_n696_), .B(mai_mai_n226_), .Y(mai_mai_n786_));
  NA2        m0758(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n787_));
  NO3        m0759(.A(mai_mai_n787_), .B(mai_mai_n743_), .C(mai_mai_n273_), .Y(mai_mai_n788_));
  INV        m0760(.A(mai_mai_n788_), .Y(mai_mai_n789_));
  NA3        m0761(.A(mai_mai_n789_), .B(mai_mai_n786_), .C(mai_mai_n394_), .Y(mai_mai_n790_));
  OR2        m0762(.A(mai_mai_n648_), .B(mai_mai_n89_), .Y(mai_mai_n791_));
  NOi31      m0763(.An(b), .B(d), .C(a), .Y(mai_mai_n792_));
  NO2        m0764(.A(mai_mai_n792_), .B(mai_mai_n591_), .Y(mai_mai_n793_));
  NO2        m0765(.A(mai_mai_n793_), .B(n), .Y(mai_mai_n794_));
  NOi21      m0766(.An(mai_mai_n780_), .B(mai_mai_n794_), .Y(mai_mai_n795_));
  OAI220     m0767(.A0(mai_mai_n795_), .A1(mai_mai_n791_), .B0(mai_mai_n768_), .B1(mai_mai_n592_), .Y(mai_mai_n796_));
  NO2        m0768(.A(mai_mai_n322_), .B(mai_mai_n114_), .Y(mai_mai_n797_));
  NOi21      m0769(.An(mai_mai_n797_), .B(mai_mai_n155_), .Y(mai_mai_n798_));
  NO2        m0770(.A(mai_mai_n677_), .B(n), .Y(mai_mai_n799_));
  AOI220     m0771(.A0(mai_mai_n757_), .A1(mai_mai_n655_), .B0(mai_mai_n799_), .B1(mai_mai_n688_), .Y(mai_mai_n800_));
  NO2        m0772(.A(mai_mai_n317_), .B(mai_mai_n231_), .Y(mai_mai_n801_));
  OAI210     m0773(.A0(mai_mai_n93_), .A1(mai_mai_n90_), .B0(mai_mai_n801_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n118_), .B(mai_mai_n81_), .Y(mai_mai_n803_));
  AOI210     m0775(.A0(mai_mai_n413_), .A1(mai_mai_n406_), .B0(mai_mai_n803_), .Y(mai_mai_n804_));
  NAi21      m0776(.An(mai_mai_n804_), .B(mai_mai_n802_), .Y(mai_mai_n805_));
  NA2        m0777(.A(mai_mai_n715_), .B(mai_mai_n34_), .Y(mai_mai_n806_));
  NAi21      m0778(.An(mai_mai_n721_), .B(mai_mai_n424_), .Y(mai_mai_n807_));
  NO2        m0779(.A(mai_mai_n267_), .B(i), .Y(mai_mai_n808_));
  NA2        m0780(.A(mai_mai_n700_), .B(mai_mai_n338_), .Y(mai_mai_n809_));
  OAI210     m0781(.A0(mai_mai_n583_), .A1(mai_mai_n582_), .B0(mai_mai_n352_), .Y(mai_mai_n810_));
  AN3        m0782(.A(mai_mai_n810_), .B(mai_mai_n809_), .C(mai_mai_n807_), .Y(mai_mai_n811_));
  NAi41      m0783(.An(mai_mai_n805_), .B(mai_mai_n811_), .C(mai_mai_n806_), .D(mai_mai_n800_), .Y(mai_mai_n812_));
  NO4        m0784(.A(mai_mai_n812_), .B(mai_mai_n798_), .C(mai_mai_n796_), .D(mai_mai_n790_), .Y(mai_mai_n813_));
  NA4        m0785(.A(mai_mai_n813_), .B(mai_mai_n785_), .C(mai_mai_n740_), .D(mai_mai_n726_), .Y(mai09));
  INV        m0786(.A(mai_mai_n119_), .Y(mai_mai_n815_));
  NA2        m0787(.A(f), .B(e), .Y(mai_mai_n816_));
  NO2        m0788(.A(mai_mai_n219_), .B(mai_mai_n109_), .Y(mai_mai_n817_));
  NA2        m0789(.A(mai_mai_n817_), .B(g), .Y(mai_mai_n818_));
  NA4        m0790(.A(mai_mai_n306_), .B(mai_mai_n461_), .C(mai_mai_n255_), .D(mai_mai_n116_), .Y(mai_mai_n819_));
  AOI210     m0791(.A0(mai_mai_n819_), .A1(g), .B0(mai_mai_n458_), .Y(mai_mai_n820_));
  AOI210     m0792(.A0(mai_mai_n820_), .A1(mai_mai_n818_), .B0(mai_mai_n816_), .Y(mai_mai_n821_));
  NA2        m0793(.A(mai_mai_n821_), .B(mai_mai_n815_), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n198_), .B(mai_mai_n206_), .Y(mai_mai_n823_));
  NA3        m0795(.A(m), .B(l), .C(i), .Y(mai_mai_n824_));
  OAI220     m0796(.A0(mai_mai_n577_), .A1(mai_mai_n824_), .B0(mai_mai_n343_), .B1(mai_mai_n519_), .Y(mai_mai_n825_));
  NA4        m0797(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .D(f), .Y(mai_mai_n826_));
  NAi31      m0798(.An(mai_mai_n825_), .B(mai_mai_n826_), .C(mai_mai_n429_), .Y(mai_mai_n827_));
  OR2        m0799(.A(mai_mai_n827_), .B(mai_mai_n823_), .Y(mai_mai_n828_));
  NA3        m0800(.A(mai_mai_n791_), .B(mai_mai_n558_), .C(mai_mai_n511_), .Y(mai_mai_n829_));
  OA210      m0801(.A0(mai_mai_n829_), .A1(mai_mai_n828_), .B0(mai_mai_n794_), .Y(mai_mai_n830_));
  INV        m0802(.A(mai_mai_n331_), .Y(mai_mai_n831_));
  NO2        m0803(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n832_));
  NO2        m0804(.A(mai_mai_n832_), .B(mai_mai_n586_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n779_), .B(mai_mai_n326_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n332_), .B(mai_mai_n333_), .Y(mai_mai_n835_));
  OAI210     m0807(.A0(mai_mai_n198_), .A1(mai_mai_n206_), .B0(mai_mai_n835_), .Y(mai_mai_n836_));
  AOI220     m0808(.A0(mai_mai_n836_), .A1(mai_mai_n834_), .B0(mai_mai_n833_), .B1(mai_mai_n831_), .Y(mai_mai_n837_));
  NA3        m0809(.A(mai_mai_n111_), .B(mai_mai_n184_), .C(mai_mai_n31_), .Y(mai_mai_n838_));
  NA3        m0810(.A(mai_mai_n838_), .B(mai_mai_n837_), .C(mai_mai_n614_), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n573_), .B(mai_mai_n490_), .Y(mai_mai_n840_));
  NA2        m0812(.A(mai_mai_n840_), .B(mai_mai_n184_), .Y(mai_mai_n841_));
  NOi21      m0813(.An(f), .B(d), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n842_), .B(m), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n843_), .B(mai_mai_n52_), .Y(mai_mai_n844_));
  NOi32      m0816(.An(g), .Bn(f), .C(d), .Y(mai_mai_n845_));
  NA4        m0817(.A(mai_mai_n845_), .B(mai_mai_n593_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n846_));
  NOi21      m0818(.An(mai_mai_n307_), .B(mai_mai_n846_), .Y(mai_mai_n847_));
  AOI210     m0819(.A0(mai_mai_n844_), .A1(mai_mai_n538_), .B0(mai_mai_n847_), .Y(mai_mai_n848_));
  NA3        m0820(.A(mai_mai_n306_), .B(mai_mai_n255_), .C(mai_mai_n116_), .Y(mai_mai_n849_));
  AN2        m0821(.A(f), .B(d), .Y(mai_mai_n850_));
  NA3        m0822(.A(mai_mai_n466_), .B(mai_mai_n850_), .C(mai_mai_n81_), .Y(mai_mai_n851_));
  NO3        m0823(.A(mai_mai_n851_), .B(mai_mai_n74_), .C(mai_mai_n207_), .Y(mai_mai_n852_));
  NO2        m0824(.A(mai_mai_n281_), .B(mai_mai_n56_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n849_), .B(mai_mai_n852_), .Y(mai_mai_n854_));
  NAi41      m0826(.An(mai_mai_n480_), .B(mai_mai_n854_), .C(mai_mai_n848_), .D(mai_mai_n841_), .Y(mai_mai_n855_));
  NO2        m0827(.A(mai_mai_n642_), .B(mai_mai_n322_), .Y(mai_mai_n856_));
  AN2        m0828(.A(mai_mai_n856_), .B(mai_mai_n669_), .Y(mai_mai_n857_));
  NO2        m0829(.A(mai_mai_n857_), .B(mai_mai_n228_), .Y(mai_mai_n858_));
  NA2        m0830(.A(mai_mai_n591_), .B(mai_mai_n81_), .Y(mai_mai_n859_));
  NO2        m0831(.A(mai_mai_n835_), .B(mai_mai_n859_), .Y(mai_mai_n860_));
  NO2        m0832(.A(mai_mai_n851_), .B(mai_mai_n418_), .Y(mai_mai_n861_));
  NOi41      m0833(.An(mai_mai_n217_), .B(mai_mai_n861_), .C(mai_mai_n860_), .D(mai_mai_n303_), .Y(mai_mai_n862_));
  NA2        m0834(.A(c), .B(mai_mai_n113_), .Y(mai_mai_n863_));
  NO2        m0835(.A(mai_mai_n863_), .B(mai_mai_n398_), .Y(mai_mai_n864_));
  NA3        m0836(.A(mai_mai_n864_), .B(mai_mai_n501_), .C(f), .Y(mai_mai_n865_));
  OR2        m0837(.A(mai_mai_n648_), .B(mai_mai_n534_), .Y(mai_mai_n866_));
  INV        m0838(.A(mai_mai_n866_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n793_), .B(mai_mai_n108_), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n868_), .B(mai_mai_n867_), .Y(mai_mai_n869_));
  NA4        m0841(.A(mai_mai_n869_), .B(mai_mai_n865_), .C(mai_mai_n862_), .D(mai_mai_n858_), .Y(mai_mai_n870_));
  NO4        m0842(.A(mai_mai_n870_), .B(mai_mai_n855_), .C(mai_mai_n839_), .D(mai_mai_n830_), .Y(mai_mai_n871_));
  OR2        m0843(.A(mai_mai_n851_), .B(mai_mai_n74_), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n109_), .B(j), .Y(mai_mai_n873_));
  NA2        m0845(.A(mai_mai_n817_), .B(g), .Y(mai_mai_n874_));
  AOI210     m0846(.A0(mai_mai_n874_), .A1(mai_mai_n289_), .B0(mai_mai_n872_), .Y(mai_mai_n875_));
  NO2        m0847(.A(mai_mai_n326_), .B(mai_mai_n826_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n224_), .B(mai_mai_n218_), .Y(mai_mai_n877_));
  NA2        m0849(.A(mai_mai_n877_), .B(mai_mai_n221_), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n418_), .B(mai_mai_n816_), .Y(mai_mai_n879_));
  NA2        m0851(.A(mai_mai_n879_), .B(mai_mai_n550_), .Y(mai_mai_n880_));
  NA2        m0852(.A(mai_mai_n880_), .B(mai_mai_n878_), .Y(mai_mai_n881_));
  NA2        m0853(.A(e), .B(d), .Y(mai_mai_n882_));
  OAI220     m0854(.A0(mai_mai_n882_), .A1(c), .B0(mai_mai_n317_), .B1(d), .Y(mai_mai_n883_));
  NA3        m0855(.A(mai_mai_n883_), .B(mai_mai_n445_), .C(mai_mai_n499_), .Y(mai_mai_n884_));
  AOI210     m0856(.A0(mai_mai_n506_), .A1(mai_mai_n177_), .B0(mai_mai_n224_), .Y(mai_mai_n885_));
  AOI210     m0857(.A0(mai_mai_n613_), .A1(mai_mai_n336_), .B0(mai_mai_n885_), .Y(mai_mai_n886_));
  NA2        m0858(.A(mai_mai_n281_), .B(mai_mai_n160_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n852_), .B(mai_mai_n887_), .Y(mai_mai_n888_));
  NA3        m0860(.A(mai_mai_n163_), .B(mai_mai_n82_), .C(mai_mai_n34_), .Y(mai_mai_n889_));
  NA4        m0861(.A(mai_mai_n889_), .B(mai_mai_n888_), .C(mai_mai_n886_), .D(mai_mai_n884_), .Y(mai_mai_n890_));
  NO4        m0862(.A(mai_mai_n890_), .B(mai_mai_n881_), .C(mai_mai_n876_), .D(mai_mai_n875_), .Y(mai_mai_n891_));
  NA2        m0863(.A(mai_mai_n831_), .B(mai_mai_n31_), .Y(mai_mai_n892_));
  OR2        m0864(.A(mai_mai_n892_), .B(mai_mai_n210_), .Y(mai_mai_n893_));
  NO2        m0865(.A(mai_mai_n612_), .B(mai_mai_n61_), .Y(mai_mai_n894_));
  AOI220     m0866(.A0(mai_mai_n894_), .A1(mai_mai_n856_), .B0(mai_mai_n603_), .B1(mai_mai_n611_), .Y(mai_mai_n895_));
  INV        m0867(.A(mai_mai_n895_), .Y(mai_mai_n896_));
  OAI210     m0868(.A0(mai_mai_n817_), .A1(mai_mai_n887_), .B0(mai_mai_n845_), .Y(mai_mai_n897_));
  NO2        m0869(.A(mai_mai_n897_), .B(mai_mai_n594_), .Y(mai_mai_n898_));
  AOI210     m0870(.A0(mai_mai_n115_), .A1(mai_mai_n114_), .B0(mai_mai_n254_), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n899_), .B(mai_mai_n846_), .Y(mai_mai_n900_));
  AO210      m0872(.A0(mai_mai_n834_), .A1(mai_mai_n825_), .B0(mai_mai_n900_), .Y(mai_mai_n901_));
  NOi31      m0873(.An(mai_mai_n538_), .B(mai_mai_n843_), .C(mai_mai_n289_), .Y(mai_mai_n902_));
  NO4        m0874(.A(mai_mai_n902_), .B(mai_mai_n901_), .C(mai_mai_n898_), .D(mai_mai_n896_), .Y(mai_mai_n903_));
  AO220      m0875(.A0(mai_mai_n445_), .A1(mai_mai_n735_), .B0(mai_mai_n172_), .B1(f), .Y(mai_mai_n904_));
  NA2        m0876(.A(mai_mai_n904_), .B(mai_mai_n883_), .Y(mai_mai_n905_));
  NO2        m0877(.A(mai_mai_n428_), .B(mai_mai_n71_), .Y(mai_mai_n906_));
  OAI210     m0878(.A0(mai_mai_n829_), .A1(mai_mai_n906_), .B0(mai_mai_n693_), .Y(mai_mai_n907_));
  AN4        m0879(.A(mai_mai_n907_), .B(mai_mai_n905_), .C(mai_mai_n903_), .D(mai_mai_n893_), .Y(mai_mai_n908_));
  NA4        m0880(.A(mai_mai_n908_), .B(mai_mai_n891_), .C(mai_mai_n871_), .D(mai_mai_n822_), .Y(mai12));
  NO4        m0881(.A(mai_mai_n433_), .B(mai_mai_n246_), .C(mai_mai_n569_), .D(mai_mai_n207_), .Y(mai_mai_n910_));
  NA2        m0882(.A(mai_mai_n538_), .B(mai_mai_n906_), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n443_), .B(mai_mai_n113_), .Y(mai_mai_n912_));
  NO2        m0884(.A(mai_mai_n832_), .B(mai_mai_n343_), .Y(mai_mai_n913_));
  NO2        m0885(.A(mai_mai_n648_), .B(mai_mai_n367_), .Y(mai_mai_n914_));
  AOI220     m0886(.A0(mai_mai_n914_), .A1(mai_mai_n536_), .B0(mai_mai_n913_), .B1(mai_mai_n912_), .Y(mai_mai_n915_));
  NA3        m0887(.A(mai_mai_n915_), .B(mai_mai_n911_), .C(mai_mai_n432_), .Y(mai_mai_n916_));
  AOI210     m0888(.A0(mai_mai_n227_), .A1(mai_mai_n330_), .B0(mai_mai_n195_), .Y(mai_mai_n917_));
  OR2        m0889(.A(mai_mai_n917_), .B(mai_mai_n910_), .Y(mai_mai_n918_));
  NO2        m0890(.A(mai_mai_n379_), .B(mai_mai_n207_), .Y(mai_mai_n919_));
  OAI210     m0891(.A0(mai_mai_n919_), .A1(mai_mai_n918_), .B0(mai_mai_n393_), .Y(mai_mai_n920_));
  NO2        m0892(.A(mai_mai_n632_), .B(mai_mai_n257_), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n577_), .B(mai_mai_n824_), .Y(mai_mai_n922_));
  AOI220     m0894(.A0(mai_mai_n922_), .A1(mai_mai_n556_), .B0(mai_mai_n801_), .B1(mai_mai_n921_), .Y(mai_mai_n923_));
  NO2        m0895(.A(mai_mai_n145_), .B(mai_mai_n231_), .Y(mai_mai_n924_));
  NA2        m0896(.A(mai_mai_n923_), .B(mai_mai_n920_), .Y(mai_mai_n925_));
  OR2        m0897(.A(mai_mai_n318_), .B(mai_mai_n912_), .Y(mai_mai_n926_));
  NA2        m0898(.A(mai_mai_n926_), .B(mai_mai_n344_), .Y(mai_mai_n927_));
  INV        m0899(.A(mai_mai_n927_), .Y(mai_mai_n928_));
  NO3        m0900(.A(mai_mai_n653_), .B(mai_mai_n89_), .C(mai_mai_n45_), .Y(mai_mai_n929_));
  NO4        m0901(.A(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n925_), .D(mai_mai_n916_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n357_), .B(mai_mai_n356_), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n574_), .B(mai_mai_n72_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n546_), .B(mai_mai_n140_), .Y(mai_mai_n933_));
  NOi21      m0905(.An(mai_mai_n34_), .B(mai_mai_n642_), .Y(mai_mai_n934_));
  AOI220     m0906(.A0(mai_mai_n934_), .A1(mai_mai_n933_), .B0(mai_mai_n932_), .B1(mai_mai_n931_), .Y(mai_mai_n935_));
  OAI210     m0907(.A0(mai_mai_n244_), .A1(mai_mai_n45_), .B0(mai_mai_n935_), .Y(mai_mai_n936_));
  NA2        m0908(.A(mai_mai_n424_), .B(mai_mai_n259_), .Y(mai_mai_n937_));
  NO3        m0909(.A(mai_mai_n803_), .B(mai_mai_n86_), .C(mai_mai_n398_), .Y(mai_mai_n938_));
  NAi21      m0910(.An(mai_mai_n938_), .B(mai_mai_n937_), .Y(mai_mai_n939_));
  NO2        m0911(.A(mai_mai_n497_), .B(mai_mai_n297_), .Y(mai_mai_n940_));
  INV        m0912(.A(mai_mai_n940_), .Y(mai_mai_n941_));
  NO2        m0913(.A(mai_mai_n941_), .B(mai_mai_n140_), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n623_), .B(mai_mai_n352_), .Y(mai_mai_n943_));
  OAI210     m0915(.A0(mai_mai_n722_), .A1(mai_mai_n943_), .B0(mai_mai_n354_), .Y(mai_mai_n944_));
  NO4        m0916(.A(mai_mai_n944_), .B(mai_mai_n942_), .C(mai_mai_n939_), .D(mai_mai_n936_), .Y(mai_mai_n945_));
  NA2        m0917(.A(mai_mai_n336_), .B(g), .Y(mai_mai_n946_));
  NA2        m0918(.A(mai_mai_n157_), .B(i), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n947_), .B(mai_mai_n89_), .Y(mai_mai_n948_));
  AOI210     m0920(.A0(mai_mai_n408_), .A1(mai_mai_n37_), .B0(mai_mai_n948_), .Y(mai_mai_n949_));
  NO2        m0921(.A(mai_mai_n140_), .B(mai_mai_n81_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n546_), .B(mai_mai_n371_), .Y(mai_mai_n951_));
  AOI210     m0923(.A0(mai_mai_n951_), .A1(n), .B0(mai_mai_n950_), .Y(mai_mai_n952_));
  OAI220     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n946_), .B0(mai_mai_n949_), .B1(mai_mai_n326_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n648_), .B(mai_mai_n490_), .Y(mai_mai_n954_));
  NA3        m0926(.A(mai_mai_n332_), .B(mai_mai_n618_), .C(i), .Y(mai_mai_n955_));
  OAI210     m0927(.A0(mai_mai_n428_), .A1(mai_mai_n306_), .B0(mai_mai_n955_), .Y(mai_mai_n956_));
  OAI220     m0928(.A0(mai_mai_n956_), .A1(mai_mai_n954_), .B0(mai_mai_n665_), .B1(mai_mai_n747_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n597_), .B(mai_mai_n110_), .Y(mai_mai_n958_));
  OR3        m0930(.A(mai_mai_n306_), .B(mai_mai_n423_), .C(f), .Y(mai_mai_n959_));
  NA3        m0931(.A(mai_mai_n618_), .B(mai_mai_n79_), .C(i), .Y(mai_mai_n960_));
  OA220      m0932(.A0(mai_mai_n960_), .A1(mai_mai_n958_), .B0(mai_mai_n959_), .B1(mai_mai_n576_), .Y(mai_mai_n961_));
  NA3        m0933(.A(mai_mai_n319_), .B(mai_mai_n115_), .C(g), .Y(mai_mai_n962_));
  AOI210     m0934(.A0(mai_mai_n663_), .A1(mai_mai_n962_), .B0(m), .Y(mai_mai_n963_));
  OAI210     m0935(.A0(mai_mai_n963_), .A1(mai_mai_n913_), .B0(mai_mai_n318_), .Y(mai_mai_n964_));
  NA2        m0936(.A(mai_mai_n680_), .B(mai_mai_n859_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n826_), .B(mai_mai_n429_), .Y(mai_mai_n966_));
  NA2        m0938(.A(mai_mai_n215_), .B(h), .Y(mai_mai_n967_));
  NA3        m0939(.A(mai_mai_n967_), .B(mai_mai_n960_), .C(mai_mai_n959_), .Y(mai_mai_n968_));
  AOI220     m0940(.A0(mai_mai_n968_), .A1(mai_mai_n252_), .B0(mai_mai_n966_), .B1(mai_mai_n965_), .Y(mai_mai_n969_));
  NA4        m0941(.A(mai_mai_n969_), .B(mai_mai_n964_), .C(mai_mai_n961_), .D(mai_mai_n957_), .Y(mai_mai_n970_));
  NO2        m0942(.A(mai_mai_n367_), .B(mai_mai_n88_), .Y(mai_mai_n971_));
  OAI210     m0943(.A0(mai_mai_n971_), .A1(mai_mai_n921_), .B0(mai_mai_n232_), .Y(mai_mai_n972_));
  NA2        m0944(.A(mai_mai_n652_), .B(mai_mai_n85_), .Y(mai_mai_n973_));
  NO2        m0945(.A(mai_mai_n449_), .B(mai_mai_n207_), .Y(mai_mai_n974_));
  AOI220     m0946(.A0(mai_mai_n974_), .A1(mai_mai_n372_), .B0(mai_mai_n926_), .B1(mai_mai_n211_), .Y(mai_mai_n975_));
  AOI220     m0947(.A0(mai_mai_n914_), .A1(mai_mai_n924_), .B0(mai_mai_n575_), .B1(mai_mai_n87_), .Y(mai_mai_n976_));
  NA4        m0948(.A(mai_mai_n976_), .B(mai_mai_n975_), .C(mai_mai_n973_), .D(mai_mai_n972_), .Y(mai_mai_n977_));
  OAI210     m0949(.A0(mai_mai_n966_), .A1(mai_mai_n922_), .B0(mai_mai_n536_), .Y(mai_mai_n978_));
  NO2        m0950(.A(mai_mai_n402_), .B(mai_mai_n803_), .Y(mai_mai_n979_));
  OAI210     m0951(.A0(mai_mai_n357_), .A1(mai_mai_n356_), .B0(mai_mai_n106_), .Y(mai_mai_n980_));
  AOI210     m0952(.A0(mai_mai_n980_), .A1(mai_mai_n528_), .B0(mai_mai_n979_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n963_), .B(mai_mai_n912_), .Y(mai_mai_n982_));
  NO3        m0954(.A(mai_mai_n873_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n983_), .B(mai_mai_n616_), .Y(mai_mai_n984_));
  NA4        m0956(.A(mai_mai_n984_), .B(mai_mai_n982_), .C(mai_mai_n981_), .D(mai_mai_n978_), .Y(mai_mai_n985_));
  NO4        m0957(.A(mai_mai_n985_), .B(mai_mai_n977_), .C(mai_mai_n970_), .D(mai_mai_n953_), .Y(mai_mai_n986_));
  NAi31      m0958(.An(mai_mai_n137_), .B(mai_mai_n409_), .C(n), .Y(mai_mai_n987_));
  NO3        m0959(.A(mai_mai_n267_), .B(mai_mai_n137_), .C(mai_mai_n398_), .Y(mai_mai_n988_));
  NA2        m0960(.A(mai_mai_n988_), .B(mai_mai_n491_), .Y(mai_mai_n989_));
  NA2        m0961(.A(mai_mai_n483_), .B(i), .Y(mai_mai_n990_));
  NA2        m0962(.A(mai_mai_n990_), .B(mai_mai_n989_), .Y(mai_mai_n991_));
  NA2        m0963(.A(mai_mai_n224_), .B(mai_mai_n168_), .Y(mai_mai_n992_));
  NO2        m0964(.A(mai_mai_n434_), .B(mai_mai_n172_), .Y(mai_mai_n993_));
  NOi31      m0965(.An(mai_mai_n992_), .B(mai_mai_n993_), .C(mai_mai_n207_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n427_), .B(mai_mai_n859_), .Y(mai_mai_n995_));
  NO3        m0967(.A(mai_mai_n428_), .B(mai_mai_n306_), .C(mai_mai_n74_), .Y(mai_mai_n996_));
  AOI220     m0968(.A0(mai_mai_n996_), .A1(mai_mai_n995_), .B0(mai_mai_n472_), .B1(g), .Y(mai_mai_n997_));
  INV        m0969(.A(mai_mai_n997_), .Y(mai_mai_n998_));
  OAI220     m0970(.A0(mai_mai_n987_), .A1(mai_mai_n227_), .B0(mai_mai_n955_), .B1(mai_mai_n592_), .Y(mai_mai_n999_));
  NO2        m0971(.A(mai_mai_n649_), .B(mai_mai_n367_), .Y(mai_mai_n1000_));
  NO3        m0972(.A(mai_mai_n537_), .B(mai_mai_n144_), .C(mai_mai_n206_), .Y(mai_mai_n1001_));
  OAI210     m0973(.A0(mai_mai_n1001_), .A1(mai_mai_n517_), .B0(mai_mai_n368_), .Y(mai_mai_n1002_));
  OAI220     m0974(.A0(mai_mai_n914_), .A1(mai_mai_n922_), .B0(mai_mai_n538_), .B1(mai_mai_n417_), .Y(mai_mai_n1003_));
  NA2        m0975(.A(mai_mai_n1003_), .B(mai_mai_n1002_), .Y(mai_mai_n1004_));
  OAI210     m0976(.A0(mai_mai_n917_), .A1(mai_mai_n910_), .B0(mai_mai_n992_), .Y(mai_mai_n1005_));
  NA3        m0977(.A(mai_mai_n951_), .B(mai_mai_n477_), .C(mai_mai_n46_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n370_), .B(mai_mai_n368_), .Y(mai_mai_n1007_));
  NA4        m0979(.A(mai_mai_n1007_), .B(mai_mai_n1006_), .C(mai_mai_n1005_), .D(mai_mai_n268_), .Y(mai_mai_n1008_));
  OR4        m0980(.A(mai_mai_n1008_), .B(mai_mai_n1004_), .C(mai_mai_n1000_), .D(mai_mai_n999_), .Y(mai_mai_n1009_));
  NO4        m0981(.A(mai_mai_n1009_), .B(mai_mai_n998_), .C(mai_mai_n994_), .D(mai_mai_n991_), .Y(mai_mai_n1010_));
  NA4        m0982(.A(mai_mai_n1010_), .B(mai_mai_n986_), .C(mai_mai_n945_), .D(mai_mai_n930_), .Y(mai13));
  AN2        m0983(.A(c), .B(b), .Y(mai_mai_n1012_));
  NA3        m0984(.A(mai_mai_n243_), .B(mai_mai_n1012_), .C(m), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n488_), .B(f), .Y(mai_mai_n1014_));
  NO3        m0986(.A(mai_mai_n1014_), .B(mai_mai_n1013_), .C(mai_mai_n570_), .Y(mai_mai_n1015_));
  NAi32      m0987(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1016_));
  NA2        m0988(.A(mai_mai_n136_), .B(mai_mai_n45_), .Y(mai_mai_n1017_));
  NO4        m0989(.A(mai_mai_n1017_), .B(mai_mai_n1016_), .C(mai_mai_n577_), .D(mai_mai_n304_), .Y(mai_mai_n1018_));
  NA2        m0990(.A(mai_mai_n401_), .B(mai_mai_n206_), .Y(mai_mai_n1019_));
  AN2        m0991(.A(d), .B(c), .Y(mai_mai_n1020_));
  NA2        m0992(.A(mai_mai_n1020_), .B(mai_mai_n113_), .Y(mai_mai_n1021_));
  NO4        m0993(.A(mai_mai_n1021_), .B(mai_mai_n1019_), .C(mai_mai_n173_), .D(mai_mai_n164_), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n488_), .B(c), .Y(mai_mai_n1023_));
  NO4        m0995(.A(mai_mai_n1017_), .B(mai_mai_n573_), .C(mai_mai_n1023_), .D(mai_mai_n304_), .Y(mai_mai_n1024_));
  OR2        m0996(.A(mai_mai_n1022_), .B(mai_mai_n1024_), .Y(mai_mai_n1025_));
  OR3        m0997(.A(mai_mai_n1025_), .B(mai_mai_n1018_), .C(mai_mai_n1015_), .Y(mai_mai_n1026_));
  NAi32      m0998(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n1027_), .B(mai_mai_n141_), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n1028_), .B(g), .Y(mai_mai_n1029_));
  OR3        m1001(.A(mai_mai_n218_), .B(mai_mai_n173_), .C(mai_mai_n164_), .Y(mai_mai_n1030_));
  NO2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1029_), .Y(mai_mai_n1031_));
  NO2        m1003(.A(mai_mai_n1023_), .B(mai_mai_n304_), .Y(mai_mai_n1032_));
  NO2        m1004(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n620_), .B(mai_mai_n1033_), .Y(mai_mai_n1034_));
  NOi21      m1006(.An(mai_mai_n1032_), .B(mai_mai_n1034_), .Y(mai_mai_n1035_));
  NO2        m1007(.A(mai_mai_n751_), .B(mai_mai_n109_), .Y(mai_mai_n1036_));
  NOi41      m1008(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1037_));
  NA2        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1036_), .Y(mai_mai_n1038_));
  NO2        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1029_), .Y(mai_mai_n1039_));
  OR3        m1011(.A(e), .B(d), .C(c), .Y(mai_mai_n1040_));
  NA3        m1012(.A(k), .B(j), .C(i), .Y(mai_mai_n1041_));
  NO3        m1013(.A(mai_mai_n1041_), .B(mai_mai_n304_), .C(mai_mai_n88_), .Y(mai_mai_n1042_));
  NOi21      m1014(.An(mai_mai_n1042_), .B(mai_mai_n1040_), .Y(mai_mai_n1043_));
  OR4        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1039_), .C(mai_mai_n1035_), .D(mai_mai_n1031_), .Y(mai_mai_n1044_));
  NA3        m1016(.A(mai_mai_n455_), .B(mai_mai_n328_), .C(mai_mai_n56_), .Y(mai_mai_n1045_));
  NO2        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1034_), .Y(mai_mai_n1046_));
  NO3        m1018(.A(mai_mai_n1045_), .B(mai_mai_n573_), .C(mai_mai_n441_), .Y(mai_mai_n1047_));
  NO2        m1019(.A(f), .B(c), .Y(mai_mai_n1048_));
  NOi21      m1020(.An(mai_mai_n1048_), .B(mai_mai_n433_), .Y(mai_mai_n1049_));
  NA2        m1021(.A(mai_mai_n1049_), .B(mai_mai_n59_), .Y(mai_mai_n1050_));
  OR2        m1022(.A(k), .B(i), .Y(mai_mai_n1051_));
  NO3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n238_), .C(l), .Y(mai_mai_n1052_));
  NOi31      m1024(.An(mai_mai_n1052_), .B(mai_mai_n1050_), .C(j), .Y(mai_mai_n1053_));
  OR3        m1025(.A(mai_mai_n1053_), .B(mai_mai_n1047_), .C(mai_mai_n1046_), .Y(mai_mai_n1054_));
  OR3        m1026(.A(mai_mai_n1054_), .B(mai_mai_n1044_), .C(mai_mai_n1026_), .Y(mai02));
  OR2        m1027(.A(l), .B(k), .Y(mai_mai_n1056_));
  OR3        m1028(.A(h), .B(g), .C(f), .Y(mai_mai_n1057_));
  OR3        m1029(.A(n), .B(m), .C(i), .Y(mai_mai_n1058_));
  NO4        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1057_), .C(mai_mai_n1056_), .D(mai_mai_n1040_), .Y(mai_mai_n1059_));
  NOi31      m1031(.An(e), .B(d), .C(c), .Y(mai_mai_n1060_));
  AOI210     m1032(.A0(mai_mai_n1042_), .A1(mai_mai_n1060_), .B0(mai_mai_n1018_), .Y(mai_mai_n1061_));
  AN3        m1033(.A(g), .B(f), .C(c), .Y(mai_mai_n1062_));
  NA2        m1034(.A(mai_mai_n1062_), .B(mai_mai_n455_), .Y(mai_mai_n1063_));
  OR2        m1035(.A(mai_mai_n1041_), .B(mai_mai_n304_), .Y(mai_mai_n1064_));
  OR2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n1063_), .Y(mai_mai_n1065_));
  NO3        m1037(.A(mai_mai_n1045_), .B(mai_mai_n1017_), .C(mai_mai_n573_), .Y(mai_mai_n1066_));
  NO2        m1038(.A(mai_mai_n1066_), .B(mai_mai_n1031_), .Y(mai_mai_n1067_));
  NA3        m1039(.A(l), .B(k), .C(j), .Y(mai_mai_n1068_));
  NA2        m1040(.A(i), .B(h), .Y(mai_mai_n1069_));
  NO3        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1068_), .C(mai_mai_n129_), .Y(mai_mai_n1070_));
  NO3        m1042(.A(mai_mai_n138_), .B(mai_mai_n279_), .C(mai_mai_n207_), .Y(mai_mai_n1071_));
  AOI210     m1043(.A0(mai_mai_n1071_), .A1(mai_mai_n1070_), .B0(mai_mai_n1035_), .Y(mai_mai_n1072_));
  NA3        m1044(.A(c), .B(b), .C(a), .Y(mai_mai_n1073_));
  NO3        m1045(.A(mai_mai_n1073_), .B(mai_mai_n882_), .C(mai_mai_n206_), .Y(mai_mai_n1074_));
  NO3        m1046(.A(mai_mai_n297_), .B(mai_mai_n49_), .C(mai_mai_n109_), .Y(mai_mai_n1075_));
  AOI210     m1047(.A0(mai_mai_n1075_), .A1(mai_mai_n1074_), .B0(mai_mai_n1046_), .Y(mai_mai_n1076_));
  AN4        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1072_), .C(mai_mai_n1067_), .D(mai_mai_n1065_), .Y(mai_mai_n1077_));
  NO2        m1049(.A(mai_mai_n1021_), .B(mai_mai_n1019_), .Y(mai_mai_n1078_));
  NA2        m1050(.A(mai_mai_n1038_), .B(mai_mai_n1030_), .Y(mai_mai_n1079_));
  AOI210     m1051(.A0(mai_mai_n1079_), .A1(mai_mai_n1078_), .B0(mai_mai_n1015_), .Y(mai_mai_n1080_));
  NAi41      m1052(.An(mai_mai_n1059_), .B(mai_mai_n1080_), .C(mai_mai_n1077_), .D(mai_mai_n1061_), .Y(mai03));
  NO2        m1053(.A(mai_mai_n519_), .B(mai_mai_n586_), .Y(mai_mai_n1082_));
  NA4        m1054(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .D(mai_mai_n206_), .Y(mai_mai_n1083_));
  NA4        m1055(.A(mai_mai_n565_), .B(m), .C(mai_mai_n109_), .D(mai_mai_n206_), .Y(mai_mai_n1084_));
  NA3        m1056(.A(mai_mai_n1084_), .B(mai_mai_n358_), .C(mai_mai_n1083_), .Y(mai_mai_n1085_));
  NO3        m1057(.A(mai_mai_n1085_), .B(mai_mai_n1082_), .C(mai_mai_n980_), .Y(mai_mai_n1086_));
  NOi41      m1058(.An(mai_mai_n791_), .B(mai_mai_n836_), .C(mai_mai_n827_), .D(mai_mai_n702_), .Y(mai_mai_n1087_));
  OAI220     m1059(.A0(mai_mai_n1087_), .A1(mai_mai_n680_), .B0(mai_mai_n1086_), .B1(mai_mai_n574_), .Y(mai_mai_n1088_));
  NA4        m1060(.A(i), .B(mai_mai_n1060_), .C(mai_mai_n332_), .D(mai_mai_n328_), .Y(mai_mai_n1089_));
  OAI210     m1061(.A0(mai_mai_n803_), .A1(mai_mai_n410_), .B0(mai_mai_n1089_), .Y(mai_mai_n1090_));
  NOi31      m1062(.An(m), .B(n), .C(f), .Y(mai_mai_n1091_));
  NA2        m1063(.A(mai_mai_n1091_), .B(mai_mai_n51_), .Y(mai_mai_n1092_));
  NO2        m1064(.A(mai_mai_n866_), .B(mai_mai_n416_), .Y(mai_mai_n1093_));
  NA2        m1065(.A(mai_mai_n499_), .B(l), .Y(mai_mai_n1094_));
  NOi31      m1066(.An(mai_mai_n845_), .B(mai_mai_n1013_), .C(mai_mai_n1094_), .Y(mai_mai_n1095_));
  NO4        m1067(.A(mai_mai_n1095_), .B(mai_mai_n1093_), .C(mai_mai_n1090_), .D(mai_mai_n979_), .Y(mai_mai_n1096_));
  NO2        m1068(.A(mai_mai_n279_), .B(a), .Y(mai_mai_n1097_));
  INV        m1069(.A(mai_mai_n1018_), .Y(mai_mai_n1098_));
  NO2        m1070(.A(mai_mai_n1069_), .B(mai_mai_n475_), .Y(mai_mai_n1099_));
  NO2        m1071(.A(mai_mai_n84_), .B(g), .Y(mai_mai_n1100_));
  AOI210     m1072(.A0(mai_mai_n1100_), .A1(mai_mai_n1099_), .B0(mai_mai_n1052_), .Y(mai_mai_n1101_));
  OR2        m1073(.A(mai_mai_n1101_), .B(mai_mai_n1050_), .Y(mai_mai_n1102_));
  NA3        m1074(.A(mai_mai_n1102_), .B(mai_mai_n1098_), .C(mai_mai_n1096_), .Y(mai_mai_n1103_));
  NO4        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1088_), .C(mai_mai_n805_), .D(mai_mai_n555_), .Y(mai_mai_n1104_));
  NA2        m1076(.A(c), .B(b), .Y(mai_mai_n1105_));
  NO2        m1077(.A(mai_mai_n692_), .B(mai_mai_n1105_), .Y(mai_mai_n1106_));
  OAI210     m1078(.A0(mai_mai_n843_), .A1(mai_mai_n820_), .B0(mai_mai_n404_), .Y(mai_mai_n1107_));
  OAI210     m1079(.A0(mai_mai_n1107_), .A1(mai_mai_n844_), .B0(mai_mai_n1106_), .Y(mai_mai_n1108_));
  NAi21      m1080(.An(mai_mai_n411_), .B(mai_mai_n1106_), .Y(mai_mai_n1109_));
  NA3        m1081(.A(mai_mai_n417_), .B(mai_mai_n548_), .C(f), .Y(mai_mai_n1110_));
  OAI210     m1082(.A0(mai_mai_n542_), .A1(mai_mai_n39_), .B0(mai_mai_n1097_), .Y(mai_mai_n1111_));
  NA3        m1083(.A(mai_mai_n1111_), .B(mai_mai_n1110_), .C(mai_mai_n1109_), .Y(mai_mai_n1112_));
  NA2        m1084(.A(mai_mai_n255_), .B(mai_mai_n116_), .Y(mai_mai_n1113_));
  OAI210     m1085(.A0(mai_mai_n1113_), .A1(mai_mai_n283_), .B0(g), .Y(mai_mai_n1114_));
  NAi21      m1086(.An(f), .B(d), .Y(mai_mai_n1115_));
  NO2        m1087(.A(mai_mai_n1115_), .B(mai_mai_n1073_), .Y(mai_mai_n1116_));
  INV        m1088(.A(mai_mai_n1116_), .Y(mai_mai_n1117_));
  AOI210     m1089(.A0(mai_mai_n1114_), .A1(mai_mai_n289_), .B0(mai_mai_n1117_), .Y(mai_mai_n1118_));
  AOI210     m1090(.A0(mai_mai_n1118_), .A1(mai_mai_n110_), .B0(mai_mai_n1112_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n458_), .B(mai_mai_n457_), .Y(mai_mai_n1120_));
  NO2        m1092(.A(mai_mai_n179_), .B(mai_mai_n231_), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n1121_), .B(m), .Y(mai_mai_n1122_));
  NA3        m1094(.A(mai_mai_n899_), .B(mai_mai_n1094_), .C(mai_mai_n461_), .Y(mai_mai_n1123_));
  OAI210     m1095(.A0(mai_mai_n1123_), .A1(mai_mai_n307_), .B0(mai_mai_n459_), .Y(mai_mai_n1124_));
  AOI210     m1096(.A0(mai_mai_n1124_), .A1(mai_mai_n1120_), .B0(mai_mai_n1122_), .Y(mai_mai_n1125_));
  NA2        m1097(.A(mai_mai_n550_), .B(mai_mai_n400_), .Y(mai_mai_n1126_));
  NA2        m1098(.A(mai_mai_n153_), .B(mai_mai_n33_), .Y(mai_mai_n1127_));
  AOI210     m1099(.A0(mai_mai_n943_), .A1(mai_mai_n1127_), .B0(mai_mai_n207_), .Y(mai_mai_n1128_));
  OAI210     m1100(.A0(mai_mai_n1128_), .A1(mai_mai_n437_), .B0(mai_mai_n1116_), .Y(mai_mai_n1129_));
  NO2        m1101(.A(mai_mai_n361_), .B(mai_mai_n360_), .Y(mai_mai_n1130_));
  AOI210     m1102(.A0(mai_mai_n1121_), .A1(mai_mai_n419_), .B0(mai_mai_n938_), .Y(mai_mai_n1131_));
  NAi41      m1103(.An(mai_mai_n1130_), .B(mai_mai_n1131_), .C(mai_mai_n1129_), .D(mai_mai_n1126_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1125_), .Y(mai_mai_n1133_));
  NA4        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1119_), .C(mai_mai_n1108_), .D(mai_mai_n1104_), .Y(mai00));
  AOI210     m1106(.A0(mai_mai_n296_), .A1(mai_mai_n207_), .B0(mai_mai_n272_), .Y(mai_mai_n1135_));
  NO2        m1107(.A(mai_mai_n1135_), .B(mai_mai_n566_), .Y(mai_mai_n1136_));
  AOI210     m1108(.A0(mai_mai_n879_), .A1(mai_mai_n924_), .B0(mai_mai_n1090_), .Y(mai_mai_n1137_));
  NO3        m1109(.A(mai_mai_n1066_), .B(mai_mai_n938_), .C(mai_mai_n699_), .Y(mai_mai_n1138_));
  NA3        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1137_), .C(mai_mai_n981_), .Y(mai_mai_n1139_));
  NA2        m1111(.A(mai_mai_n501_), .B(f), .Y(mai_mai_n1140_));
  NO2        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1021_), .Y(mai_mai_n1141_));
  NO4        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1139_), .C(mai_mai_n1136_), .D(mai_mai_n1044_), .Y(mai_mai_n1142_));
  NA3        m1114(.A(mai_mai_n163_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1143_));
  NA3        m1115(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1144_));
  NOi31      m1116(.An(n), .B(m), .C(i), .Y(mai_mai_n1145_));
  NA3        m1117(.A(mai_mai_n1145_), .B(mai_mai_n639_), .C(mai_mai_n51_), .Y(mai_mai_n1146_));
  OAI210     m1118(.A0(mai_mai_n1144_), .A1(mai_mai_n1143_), .B0(mai_mai_n1146_), .Y(mai_mai_n1147_));
  NO3        m1119(.A(mai_mai_n1147_), .B(mai_mai_n1130_), .C(mai_mai_n902_), .Y(mai_mai_n1148_));
  NO4        m1120(.A(mai_mai_n478_), .B(mai_mai_n345_), .C(mai_mai_n1105_), .D(mai_mai_n59_), .Y(mai_mai_n1149_));
  OR2        m1121(.A(mai_mai_n374_), .B(mai_mai_n131_), .Y(mai_mai_n1150_));
  NO2        m1122(.A(h), .B(g), .Y(mai_mai_n1151_));
  NA4        m1123(.A(mai_mai_n491_), .B(mai_mai_n455_), .C(mai_mai_n1151_), .D(mai_mai_n1012_), .Y(mai_mai_n1152_));
  OAI220     m1124(.A0(mai_mai_n519_), .A1(mai_mai_n586_), .B0(mai_mai_n89_), .B1(mai_mai_n88_), .Y(mai_mai_n1153_));
  NA2        m1125(.A(mai_mai_n1153_), .B(mai_mai_n528_), .Y(mai_mai_n1154_));
  AOI220     m1126(.A0(mai_mai_n314_), .A1(mai_mai_n240_), .B0(mai_mai_n174_), .B1(mai_mai_n143_), .Y(mai_mai_n1155_));
  NA4        m1127(.A(mai_mai_n1155_), .B(mai_mai_n1154_), .C(mai_mai_n1152_), .D(mai_mai_n1150_), .Y(mai_mai_n1156_));
  NO3        m1128(.A(mai_mai_n1156_), .B(mai_mai_n1149_), .C(mai_mai_n261_), .Y(mai_mai_n1157_));
  INV        m1129(.A(mai_mai_n316_), .Y(mai_mai_n1158_));
  NA2        m1130(.A(mai_mai_n240_), .B(mai_mai_n336_), .Y(mai_mai_n1159_));
  NA3        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1158_), .C(mai_mai_n148_), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n233_), .B(mai_mai_n178_), .Y(mai_mai_n1161_));
  NA2        m1133(.A(mai_mai_n1161_), .B(mai_mai_n417_), .Y(mai_mai_n1162_));
  NA3        m1134(.A(mai_mai_n176_), .B(mai_mai_n109_), .C(g), .Y(mai_mai_n1163_));
  NA2        m1135(.A(mai_mai_n455_), .B(f), .Y(mai_mai_n1164_));
  NOi31      m1136(.An(mai_mai_n853_), .B(mai_mai_n1164_), .C(mai_mai_n1163_), .Y(mai_mai_n1165_));
  NAi31      m1137(.An(mai_mai_n181_), .B(mai_mai_n840_), .C(mai_mai_n455_), .Y(mai_mai_n1166_));
  NAi31      m1138(.An(mai_mai_n1165_), .B(mai_mai_n1166_), .C(mai_mai_n1162_), .Y(mai_mai_n1167_));
  NO2        m1139(.A(mai_mai_n271_), .B(mai_mai_n74_), .Y(mai_mai_n1168_));
  NO3        m1140(.A(mai_mai_n416_), .B(mai_mai_n816_), .C(n), .Y(mai_mai_n1169_));
  AOI210     m1141(.A0(mai_mai_n1169_), .A1(mai_mai_n1168_), .B0(mai_mai_n1059_), .Y(mai_mai_n1170_));
  NAi31      m1142(.An(mai_mai_n1024_), .B(mai_mai_n1170_), .C(mai_mai_n73_), .Y(mai_mai_n1171_));
  NO4        m1143(.A(mai_mai_n1171_), .B(mai_mai_n1167_), .C(mai_mai_n1160_), .D(mai_mai_n510_), .Y(mai_mai_n1172_));
  AN3        m1144(.A(mai_mai_n1172_), .B(mai_mai_n1157_), .C(mai_mai_n1148_), .Y(mai_mai_n1173_));
  NA2        m1145(.A(mai_mai_n528_), .B(mai_mai_n99_), .Y(mai_mai_n1174_));
  NA3        m1146(.A(mai_mai_n551_), .B(mai_mai_n1174_), .C(mai_mai_n236_), .Y(mai_mai_n1175_));
  NA2        m1147(.A(mai_mai_n1085_), .B(mai_mai_n528_), .Y(mai_mai_n1176_));
  NA2        m1148(.A(mai_mai_n1176_), .B(mai_mai_n293_), .Y(mai_mai_n1177_));
  OAI210     m1149(.A0(mai_mai_n453_), .A1(mai_mai_n117_), .B0(mai_mai_n846_), .Y(mai_mai_n1178_));
  AOI220     m1150(.A0(mai_mai_n1178_), .A1(mai_mai_n1123_), .B0(mai_mai_n550_), .B1(mai_mai_n400_), .Y(mai_mai_n1179_));
  OR3        m1151(.A(mai_mai_n1021_), .B(mai_mai_n267_), .C(mai_mai_n216_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n210_), .B(mai_mai_n207_), .Y(mai_mai_n1181_));
  NA2        m1153(.A(n), .B(e), .Y(mai_mai_n1182_));
  NO2        m1154(.A(mai_mai_n1182_), .B(mai_mai_n141_), .Y(mai_mai_n1183_));
  AOI220     m1155(.A0(mai_mai_n1183_), .A1(mai_mai_n269_), .B0(mai_mai_n831_), .B1(mai_mai_n1181_), .Y(mai_mai_n1184_));
  OAI210     m1156(.A0(mai_mai_n346_), .A1(mai_mai_n308_), .B0(mai_mai_n439_), .Y(mai_mai_n1185_));
  NA4        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1184_), .C(mai_mai_n1180_), .D(mai_mai_n1179_), .Y(mai_mai_n1186_));
  AOI210     m1158(.A0(mai_mai_n1183_), .A1(mai_mai_n833_), .B0(mai_mai_n804_), .Y(mai_mai_n1187_));
  NO2        m1159(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n1021_), .B(mai_mai_n1019_), .C(mai_mai_n714_), .Y(mai_mai_n1189_));
  INV        m1161(.A(mai_mai_n129_), .Y(mai_mai_n1190_));
  AN2        m1162(.A(mai_mai_n1190_), .B(mai_mai_n1071_), .Y(mai_mai_n1191_));
  OAI210     m1163(.A0(mai_mai_n1191_), .A1(mai_mai_n1189_), .B0(mai_mai_n1188_), .Y(mai_mai_n1192_));
  NA3        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1187_), .C(mai_mai_n848_), .Y(mai_mai_n1193_));
  NO4        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1186_), .C(mai_mai_n1177_), .D(mai_mai_n1175_), .Y(mai_mai_n1194_));
  NA2        m1166(.A(mai_mai_n821_), .B(mai_mai_n746_), .Y(mai_mai_n1195_));
  NA4        m1167(.A(mai_mai_n1195_), .B(mai_mai_n1194_), .C(mai_mai_n1173_), .D(mai_mai_n1142_), .Y(mai01));
  NO4        m1168(.A(mai_mai_n788_), .B(mai_mai_n782_), .C(mai_mai_n469_), .D(mai_mai_n277_), .Y(mai_mai_n1197_));
  NA2        m1169(.A(mai_mai_n384_), .B(i), .Y(mai_mai_n1198_));
  NA3        m1170(.A(mai_mai_n1198_), .B(mai_mai_n1197_), .C(mai_mai_n1002_), .Y(mai_mai_n1199_));
  NA2        m1171(.A(mai_mai_n575_), .B(mai_mai_n87_), .Y(mai_mai_n1200_));
  NA3        m1172(.A(mai_mai_n1200_), .B(mai_mai_n895_), .C(mai_mai_n327_), .Y(mai_mai_n1201_));
  NA2        m1173(.A(mai_mai_n697_), .B(mai_mai_n94_), .Y(mai_mai_n1202_));
  NO2        m1174(.A(mai_mai_n1202_), .B(mai_mai_n1470_), .Y(mai_mai_n1203_));
  NO2        m1175(.A(mai_mai_n768_), .B(mai_mai_n592_), .Y(mai_mai_n1204_));
  AOI210     m1176(.A0(mai_mai_n1203_), .A1(mai_mai_n627_), .B0(mai_mai_n1204_), .Y(mai_mai_n1205_));
  INV        m1177(.A(mai_mai_n115_), .Y(mai_mai_n1206_));
  OA220      m1178(.A0(mai_mai_n1206_), .A1(mai_mai_n572_), .B0(mai_mai_n650_), .B1(mai_mai_n358_), .Y(mai_mai_n1207_));
  NAi41      m1179(.An(mai_mai_n156_), .B(mai_mai_n1207_), .C(mai_mai_n1205_), .D(mai_mai_n878_), .Y(mai_mai_n1208_));
  NO3        m1180(.A(mai_mai_n769_), .B(mai_mai_n664_), .C(mai_mai_n503_), .Y(mai_mai_n1209_));
  NA4        m1181(.A(mai_mai_n697_), .B(mai_mai_n94_), .C(mai_mai_n45_), .D(mai_mai_n206_), .Y(mai_mai_n1210_));
  OA220      m1182(.A0(mai_mai_n1210_), .A1(mai_mai_n658_), .B0(mai_mai_n189_), .B1(mai_mai_n187_), .Y(mai_mai_n1211_));
  NA3        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1209_), .C(mai_mai_n134_), .Y(mai_mai_n1212_));
  NO4        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1208_), .C(mai_mai_n1201_), .D(mai_mai_n1199_), .Y(mai_mai_n1213_));
  NA2        m1185(.A(mai_mai_n299_), .B(mai_mai_n523_), .Y(mai_mai_n1214_));
  NA2        m1186(.A(mai_mai_n531_), .B(mai_mai_n386_), .Y(mai_mai_n1215_));
  NOi21      m1187(.An(mai_mai_n552_), .B(mai_mai_n569_), .Y(mai_mai_n1216_));
  NA2        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1215_), .Y(mai_mai_n1217_));
  AOI210     m1189(.A0(mai_mai_n198_), .A1(mai_mai_n86_), .B0(mai_mai_n206_), .Y(mai_mai_n1218_));
  OAI210     m1190(.A0(mai_mai_n794_), .A1(mai_mai_n417_), .B0(mai_mai_n1218_), .Y(mai_mai_n1219_));
  NA2        m1191(.A(mai_mai_n197_), .B(mai_mai_n34_), .Y(mai_mai_n1220_));
  OR2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n326_), .Y(mai_mai_n1221_));
  NA4        m1193(.A(mai_mai_n1221_), .B(mai_mai_n1219_), .C(mai_mai_n1217_), .D(mai_mai_n1214_), .Y(mai_mai_n1222_));
  AOI210     m1194(.A0(mai_mai_n584_), .A1(mai_mai_n115_), .B0(mai_mai_n590_), .Y(mai_mai_n1223_));
  OAI210     m1195(.A0(mai_mai_n1206_), .A1(mai_mai_n581_), .B0(mai_mai_n1223_), .Y(mai_mai_n1224_));
  NA2        m1196(.A(mai_mai_n276_), .B(mai_mai_n189_), .Y(mai_mai_n1225_));
  NA2        m1197(.A(mai_mai_n1225_), .B(mai_mai_n655_), .Y(mai_mai_n1226_));
  NO3        m1198(.A(mai_mai_n803_), .B(mai_mai_n198_), .C(mai_mai_n398_), .Y(mai_mai_n1227_));
  NO2        m1199(.A(mai_mai_n1227_), .B(mai_mai_n938_), .Y(mai_mai_n1228_));
  OAI210     m1200(.A0(mai_mai_n1203_), .A1(mai_mai_n321_), .B0(mai_mai_n665_), .Y(mai_mai_n1229_));
  NA4        m1201(.A(mai_mai_n1229_), .B(mai_mai_n1228_), .C(mai_mai_n1226_), .D(mai_mai_n772_), .Y(mai_mai_n1230_));
  NO3        m1202(.A(mai_mai_n1230_), .B(mai_mai_n1224_), .C(mai_mai_n1222_), .Y(mai_mai_n1231_));
  NA3        m1203(.A(mai_mai_n593_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1232_));
  NO2        m1204(.A(mai_mai_n1232_), .B(mai_mai_n198_), .Y(mai_mai_n1233_));
  AOI210     m1205(.A0(mai_mai_n498_), .A1(mai_mai_n58_), .B0(mai_mai_n1233_), .Y(mai_mai_n1234_));
  OR3        m1206(.A(mai_mai_n1202_), .B(mai_mai_n594_), .C(mai_mai_n1470_), .Y(mai_mai_n1235_));
  NO2        m1207(.A(mai_mai_n1210_), .B(mai_mai_n958_), .Y(mai_mai_n1236_));
  NO2        m1208(.A(mai_mai_n1236_), .B(mai_mai_n1147_), .Y(mai_mai_n1237_));
  NA4        m1209(.A(mai_mai_n1237_), .B(mai_mai_n1235_), .C(mai_mai_n1234_), .D(mai_mai_n745_), .Y(mai_mai_n1238_));
  NO2        m1210(.A(mai_mai_n947_), .B(mai_mai_n226_), .Y(mai_mai_n1239_));
  NA2        m1211(.A(mai_mai_n562_), .B(mai_mai_n560_), .Y(mai_mai_n1240_));
  NO3        m1212(.A(mai_mai_n78_), .B(mai_mai_n297_), .C(mai_mai_n45_), .Y(mai_mai_n1241_));
  NA2        m1213(.A(mai_mai_n1240_), .B(mai_mai_n660_), .Y(mai_mai_n1242_));
  NO2        m1214(.A(mai_mai_n358_), .B(mai_mai_n72_), .Y(mai_mai_n1243_));
  INV        m1215(.A(mai_mai_n1243_), .Y(mai_mai_n1244_));
  NA2        m1216(.A(mai_mai_n1244_), .B(mai_mai_n376_), .Y(mai_mai_n1245_));
  NO3        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1242_), .C(mai_mai_n1238_), .Y(mai_mai_n1246_));
  INV        m1218(.A(mai_mai_n131_), .Y(mai_mai_n1247_));
  NO3        m1219(.A(mai_mai_n1069_), .B(mai_mai_n173_), .C(mai_mai_n84_), .Y(mai_mai_n1248_));
  AOI220     m1220(.A0(mai_mai_n1248_), .A1(mai_mai_n1247_), .B0(mai_mai_n1241_), .B1(mai_mai_n950_), .Y(mai_mai_n1249_));
  INV        m1221(.A(mai_mai_n1249_), .Y(mai_mai_n1250_));
  NO2        m1222(.A(mai_mai_n605_), .B(mai_mai_n604_), .Y(mai_mai_n1251_));
  NO4        m1223(.A(mai_mai_n1069_), .B(mai_mai_n1251_), .C(mai_mai_n171_), .D(mai_mai_n84_), .Y(mai_mai_n1252_));
  NO3        m1224(.A(mai_mai_n1252_), .B(mai_mai_n1250_), .C(mai_mai_n631_), .Y(mai_mai_n1253_));
  NA4        m1225(.A(mai_mai_n1253_), .B(mai_mai_n1246_), .C(mai_mai_n1231_), .D(mai_mai_n1213_), .Y(mai06));
  NO2        m1226(.A(mai_mai_n399_), .B(mai_mai_n549_), .Y(mai_mai_n1255_));
  INV        m1227(.A(mai_mai_n721_), .Y(mai_mai_n1256_));
  OAI210     m1228(.A0(mai_mai_n1256_), .A1(mai_mai_n262_), .B0(mai_mai_n1255_), .Y(mai_mai_n1257_));
  NO2        m1229(.A(mai_mai_n218_), .B(mai_mai_n101_), .Y(mai_mai_n1258_));
  OAI210     m1230(.A0(mai_mai_n1258_), .A1(mai_mai_n1248_), .B0(mai_mai_n372_), .Y(mai_mai_n1259_));
  NO3        m1231(.A(mai_mai_n588_), .B(mai_mai_n792_), .C(mai_mai_n591_), .Y(mai_mai_n1260_));
  OR2        m1232(.A(mai_mai_n1260_), .B(mai_mai_n866_), .Y(mai_mai_n1261_));
  NA3        m1233(.A(mai_mai_n1261_), .B(mai_mai_n1259_), .C(mai_mai_n1257_), .Y(mai_mai_n1262_));
  NO3        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1242_), .C(mai_mai_n250_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n297_), .B(mai_mai_n45_), .Y(mai_mai_n1264_));
  AOI210     m1236(.A0(mai_mai_n1264_), .A1(mai_mai_n950_), .B0(mai_mai_n1239_), .Y(mai_mai_n1265_));
  NO2        m1237(.A(mai_mai_n1265_), .B(mai_mai_n330_), .Y(mai_mai_n1266_));
  NO2        m1238(.A(mai_mai_n506_), .B(mai_mai_n168_), .Y(mai_mai_n1267_));
  NOi21      m1239(.An(mai_mai_n133_), .B(mai_mai_n45_), .Y(mai_mai_n1268_));
  NO2        m1240(.A(mai_mai_n598_), .B(mai_mai_n1092_), .Y(mai_mai_n1269_));
  OAI210     m1241(.A0(mai_mai_n450_), .A1(mai_mai_n241_), .B0(mai_mai_n889_), .Y(mai_mai_n1270_));
  NO4        m1242(.A(mai_mai_n1270_), .B(mai_mai_n1269_), .C(mai_mai_n1268_), .D(mai_mai_n1267_), .Y(mai_mai_n1271_));
  OR2        m1243(.A(mai_mai_n589_), .B(mai_mai_n587_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n357_), .B(mai_mai_n132_), .Y(mai_mai_n1273_));
  AOI210     m1245(.A0(mai_mai_n1273_), .A1(mai_mai_n575_), .B0(mai_mai_n1272_), .Y(mai_mai_n1274_));
  NA2        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1271_), .Y(mai_mai_n1275_));
  NO2        m1247(.A(mai_mai_n736_), .B(mai_mai_n356_), .Y(mai_mai_n1276_));
  NO3        m1248(.A(mai_mai_n665_), .B(mai_mai_n747_), .C(mai_mai_n627_), .Y(mai_mai_n1277_));
  NOi21      m1249(.An(mai_mai_n1276_), .B(mai_mai_n1277_), .Y(mai_mai_n1278_));
  AN2        m1250(.A(mai_mai_n934_), .B(mai_mai_n635_), .Y(mai_mai_n1279_));
  NO4        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1278_), .C(mai_mai_n1275_), .D(mai_mai_n1266_), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n787_), .B(mai_mai_n273_), .Y(mai_mai_n1281_));
  OAI220     m1253(.A0(mai_mai_n721_), .A1(mai_mai_n47_), .B0(mai_mai_n218_), .B1(mai_mai_n607_), .Y(mai_mai_n1282_));
  OAI210     m1254(.A0(mai_mai_n273_), .A1(c), .B0(mai_mai_n633_), .Y(mai_mai_n1283_));
  AOI220     m1255(.A0(mai_mai_n1283_), .A1(mai_mai_n1282_), .B0(mai_mai_n1281_), .B1(mai_mai_n262_), .Y(mai_mai_n1284_));
  OAI220     m1256(.A0(mai_mai_n689_), .A1(mai_mai_n241_), .B0(mai_mai_n502_), .B1(mai_mai_n506_), .Y(mai_mai_n1285_));
  OAI210     m1257(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1286_));
  NO3        m1258(.A(mai_mai_n1286_), .B(mai_mai_n586_), .C(j), .Y(mai_mai_n1287_));
  NOi21      m1259(.An(mai_mai_n1287_), .B(mai_mai_n658_), .Y(mai_mai_n1288_));
  NO3        m1260(.A(mai_mai_n1288_), .B(mai_mai_n1285_), .C(mai_mai_n1093_), .Y(mai_mai_n1289_));
  NA4        m1261(.A(mai_mai_n780_), .B(mai_mai_n779_), .C(mai_mai_n427_), .D(mai_mai_n859_), .Y(mai_mai_n1290_));
  NAi31      m1262(.An(mai_mai_n736_), .B(mai_mai_n1290_), .C(mai_mai_n197_), .Y(mai_mai_n1291_));
  NA3        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1289_), .C(mai_mai_n1284_), .Y(mai_mai_n1292_));
  NOi31      m1264(.An(mai_mai_n1260_), .B(mai_mai_n452_), .C(mai_mai_n385_), .Y(mai_mai_n1293_));
  OR3        m1265(.A(mai_mai_n1293_), .B(mai_mai_n768_), .C(mai_mai_n534_), .Y(mai_mai_n1294_));
  OR3        m1266(.A(mai_mai_n360_), .B(mai_mai_n218_), .C(mai_mai_n607_), .Y(mai_mai_n1295_));
  AOI210     m1267(.A0(mai_mai_n562_), .A1(mai_mai_n439_), .B0(mai_mai_n362_), .Y(mai_mai_n1296_));
  NA2        m1268(.A(mai_mai_n1287_), .B(mai_mai_n776_), .Y(mai_mai_n1297_));
  NA4        m1269(.A(mai_mai_n1297_), .B(mai_mai_n1296_), .C(mai_mai_n1295_), .D(mai_mai_n1294_), .Y(mai_mai_n1298_));
  AOI220     m1270(.A0(mai_mai_n1276_), .A1(mai_mai_n746_), .B0(mai_mai_n1273_), .B1(mai_mai_n232_), .Y(mai_mai_n1299_));
  NO3        m1271(.A(mai_mai_n857_), .B(mai_mai_n494_), .C(mai_mai_n472_), .Y(mai_mai_n1300_));
  NA2        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1299_), .Y(mai_mai_n1301_));
  NAi21      m1273(.An(j), .B(i), .Y(mai_mai_n1302_));
  NO4        m1274(.A(mai_mai_n1251_), .B(mai_mai_n1302_), .C(mai_mai_n433_), .D(mai_mai_n229_), .Y(mai_mai_n1303_));
  NO4        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1301_), .C(mai_mai_n1298_), .D(mai_mai_n1292_), .Y(mai_mai_n1304_));
  NA4        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1280_), .C(mai_mai_n1263_), .D(mai_mai_n1253_), .Y(mai07));
  NOi21      m1277(.An(j), .B(k), .Y(mai_mai_n1306_));
  NA4        m1278(.A(mai_mai_n176_), .B(mai_mai_n105_), .C(mai_mai_n1306_), .D(f), .Y(mai_mai_n1307_));
  NAi32      m1279(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1308_));
  NO3        m1280(.A(mai_mai_n1308_), .B(g), .C(f), .Y(mai_mai_n1309_));
  OAI210     m1281(.A0(mai_mai_n315_), .A1(mai_mai_n474_), .B0(mai_mai_n1309_), .Y(mai_mai_n1310_));
  NAi21      m1282(.An(f), .B(c), .Y(mai_mai_n1311_));
  OR2        m1283(.A(e), .B(d), .Y(mai_mai_n1312_));
  OAI220     m1284(.A0(mai_mai_n1312_), .A1(mai_mai_n1311_), .B0(mai_mai_n619_), .B1(mai_mai_n317_), .Y(mai_mai_n1313_));
  NA3        m1285(.A(mai_mai_n1313_), .B(mai_mai_n1033_), .C(mai_mai_n176_), .Y(mai_mai_n1314_));
  NOi31      m1286(.An(n), .B(m), .C(b), .Y(mai_mai_n1315_));
  NO3        m1287(.A(mai_mai_n129_), .B(mai_mai_n441_), .C(h), .Y(mai_mai_n1316_));
  NA3        m1288(.A(mai_mai_n1314_), .B(mai_mai_n1310_), .C(mai_mai_n1307_), .Y(mai_mai_n1317_));
  NOi41      m1289(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1318_));
  NO2        m1290(.A(k), .B(i), .Y(mai_mai_n1319_));
  NA3        m1291(.A(mai_mai_n1319_), .B(mai_mai_n877_), .C(mai_mai_n176_), .Y(mai_mai_n1320_));
  NA2        m1292(.A(mai_mai_n84_), .B(mai_mai_n45_), .Y(mai_mai_n1321_));
  NO2        m1293(.A(mai_mai_n1027_), .B(mai_mai_n433_), .Y(mai_mai_n1322_));
  NA3        m1294(.A(mai_mai_n1322_), .B(mai_mai_n1321_), .C(mai_mai_n207_), .Y(mai_mai_n1323_));
  NO2        m1295(.A(mai_mai_n1041_), .B(mai_mai_n304_), .Y(mai_mai_n1324_));
  NA2        m1296(.A(mai_mai_n535_), .B(mai_mai_n79_), .Y(mai_mai_n1325_));
  NA2        m1297(.A(mai_mai_n1188_), .B(mai_mai_n287_), .Y(mai_mai_n1326_));
  NA4        m1298(.A(mai_mai_n1326_), .B(mai_mai_n1325_), .C(mai_mai_n1323_), .D(mai_mai_n1320_), .Y(mai_mai_n1327_));
  NO2        m1299(.A(mai_mai_n1327_), .B(mai_mai_n1317_), .Y(mai_mai_n1328_));
  NO3        m1300(.A(e), .B(d), .C(c), .Y(mai_mai_n1329_));
  NA2        m1301(.A(mai_mai_n1468_), .B(mai_mai_n1329_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n1330_), .B(mai_mai_n207_), .Y(mai_mai_n1331_));
  NA3        m1303(.A(mai_mai_n686_), .B(mai_mai_n673_), .C(mai_mai_n109_), .Y(mai_mai_n1332_));
  NO2        m1304(.A(mai_mai_n1332_), .B(mai_mai_n45_), .Y(mai_mai_n1333_));
  NO2        m1305(.A(l), .B(k), .Y(mai_mai_n1334_));
  NOi41      m1306(.An(mai_mai_n540_), .B(mai_mai_n1334_), .C(mai_mai_n467_), .D(mai_mai_n433_), .Y(mai_mai_n1335_));
  NO3        m1307(.A(mai_mai_n433_), .B(d), .C(c), .Y(mai_mai_n1336_));
  NO3        m1308(.A(mai_mai_n1335_), .B(mai_mai_n1333_), .C(mai_mai_n1331_), .Y(mai_mai_n1337_));
  NO2        m1309(.A(mai_mai_n142_), .B(h), .Y(mai_mai_n1338_));
  NO2        m1310(.A(g), .B(c), .Y(mai_mai_n1339_));
  NA3        m1311(.A(mai_mai_n1339_), .B(mai_mai_n138_), .C(mai_mai_n182_), .Y(mai_mai_n1340_));
  NO2        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1467_), .Y(mai_mai_n1341_));
  NA2        m1313(.A(mai_mai_n1341_), .B(mai_mai_n176_), .Y(mai_mai_n1342_));
  NO2        m1314(.A(mai_mai_n443_), .B(a), .Y(mai_mai_n1343_));
  NA3        m1315(.A(mai_mai_n1343_), .B(k), .C(mai_mai_n110_), .Y(mai_mai_n1344_));
  NO2        m1316(.A(i), .B(h), .Y(mai_mai_n1345_));
  NA2        m1317(.A(mai_mai_n1115_), .B(h), .Y(mai_mai_n1346_));
  NA2        m1318(.A(mai_mai_n135_), .B(mai_mai_n214_), .Y(mai_mai_n1347_));
  NO2        m1319(.A(mai_mai_n1347_), .B(mai_mai_n1346_), .Y(mai_mai_n1348_));
  NO2        m1320(.A(mai_mai_n743_), .B(mai_mai_n183_), .Y(mai_mai_n1349_));
  NOi31      m1321(.An(m), .B(n), .C(b), .Y(mai_mai_n1350_));
  NOi31      m1322(.An(f), .B(d), .C(c), .Y(mai_mai_n1351_));
  NA2        m1323(.A(mai_mai_n1351_), .B(mai_mai_n1350_), .Y(mai_mai_n1352_));
  INV        m1324(.A(mai_mai_n1352_), .Y(mai_mai_n1353_));
  NO3        m1325(.A(mai_mai_n1353_), .B(mai_mai_n1349_), .C(mai_mai_n1348_), .Y(mai_mai_n1354_));
  NA2        m1326(.A(mai_mai_n1062_), .B(mai_mai_n455_), .Y(mai_mai_n1355_));
  NO4        m1327(.A(mai_mai_n1355_), .B(mai_mai_n1036_), .C(mai_mai_n433_), .D(mai_mai_n45_), .Y(mai_mai_n1356_));
  OAI210     m1328(.A0(mai_mai_n179_), .A1(mai_mai_n518_), .B0(mai_mai_n1037_), .Y(mai_mai_n1357_));
  NO3        m1329(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1358_));
  INV        m1330(.A(mai_mai_n1357_), .Y(mai_mai_n1359_));
  NO2        m1331(.A(mai_mai_n1359_), .B(mai_mai_n1356_), .Y(mai_mai_n1360_));
  AN4        m1332(.A(mai_mai_n1360_), .B(mai_mai_n1354_), .C(mai_mai_n1344_), .D(mai_mai_n1342_), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n1315_), .B(mai_mai_n369_), .Y(mai_mai_n1362_));
  NA2        m1334(.A(mai_mai_n1336_), .B(mai_mai_n208_), .Y(mai_mai_n1363_));
  NA2        m1335(.A(mai_mai_n1070_), .B(mai_mai_n1355_), .Y(mai_mai_n1364_));
  NA2        m1336(.A(mai_mai_n1364_), .B(mai_mai_n1363_), .Y(mai_mai_n1365_));
  NO4        m1337(.A(mai_mai_n129_), .B(g), .C(f), .D(e), .Y(mai_mai_n1366_));
  NA3        m1338(.A(mai_mai_n1319_), .B(mai_mai_n288_), .C(h), .Y(mai_mai_n1367_));
  OR2        m1339(.A(e), .B(a), .Y(mai_mai_n1368_));
  NO2        m1340(.A(mai_mai_n1312_), .B(mai_mai_n1311_), .Y(mai_mai_n1369_));
  AOI210     m1341(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1369_), .Y(mai_mai_n1370_));
  NO2        m1342(.A(mai_mai_n1370_), .B(mai_mai_n1058_), .Y(mai_mai_n1371_));
  NA2        m1343(.A(mai_mai_n1318_), .B(mai_mai_n1334_), .Y(mai_mai_n1372_));
  INV        m1344(.A(mai_mai_n1372_), .Y(mai_mai_n1373_));
  NA2        m1345(.A(mai_mai_n1091_), .B(mai_mai_n398_), .Y(mai_mai_n1374_));
  NO2        m1346(.A(mai_mai_n1374_), .B(mai_mai_n426_), .Y(mai_mai_n1375_));
  AO210      m1347(.A0(mai_mai_n1375_), .A1(mai_mai_n113_), .B0(mai_mai_n1373_), .Y(mai_mai_n1376_));
  NO3        m1348(.A(mai_mai_n1376_), .B(mai_mai_n1371_), .C(mai_mai_n1365_), .Y(mai_mai_n1377_));
  NA4        m1349(.A(mai_mai_n1377_), .B(mai_mai_n1361_), .C(mai_mai_n1337_), .D(mai_mai_n1328_), .Y(mai_mai_n1378_));
  NO2        m1350(.A(mai_mai_n381_), .B(j), .Y(mai_mai_n1379_));
  NA3        m1351(.A(mai_mai_n1358_), .B(mai_mai_n1312_), .C(mai_mai_n1091_), .Y(mai_mai_n1380_));
  NAi31      m1352(.An(mai_mai_n1345_), .B(mai_mai_n1049_), .C(mai_mai_n164_), .Y(mai_mai_n1381_));
  NA2        m1353(.A(mai_mai_n1381_), .B(mai_mai_n1380_), .Y(mai_mai_n1382_));
  NA3        m1354(.A(g), .B(mai_mai_n1379_), .C(mai_mai_n153_), .Y(mai_mai_n1383_));
  INV        m1355(.A(mai_mai_n1383_), .Y(mai_mai_n1384_));
  NO3        m1356(.A(mai_mai_n736_), .B(mai_mai_n171_), .C(mai_mai_n401_), .Y(mai_mai_n1385_));
  NO3        m1357(.A(mai_mai_n1385_), .B(mai_mai_n1384_), .C(mai_mai_n1382_), .Y(mai_mai_n1386_));
  OR2        m1358(.A(n), .B(i), .Y(mai_mai_n1387_));
  OAI210     m1359(.A0(mai_mai_n1387_), .A1(mai_mai_n1048_), .B0(mai_mai_n49_), .Y(mai_mai_n1388_));
  AOI220     m1360(.A0(mai_mai_n1388_), .A1(mai_mai_n1151_), .B0(mai_mai_n808_), .B1(mai_mai_n188_), .Y(mai_mai_n1389_));
  INV        m1361(.A(mai_mai_n1389_), .Y(mai_mai_n1390_));
  NO2        m1362(.A(mai_mai_n129_), .B(l), .Y(mai_mai_n1391_));
  NO2        m1363(.A(mai_mai_n218_), .B(k), .Y(mai_mai_n1392_));
  OAI210     m1364(.A0(mai_mai_n1392_), .A1(mai_mai_n1345_), .B0(mai_mai_n1391_), .Y(mai_mai_n1393_));
  NO2        m1365(.A(mai_mai_n1393_), .B(mai_mai_n31_), .Y(mai_mai_n1394_));
  NO2        m1366(.A(mai_mai_n1394_), .B(mai_mai_n1390_), .Y(mai_mai_n1395_));
  NO3        m1367(.A(mai_mai_n1073_), .B(mai_mai_n1312_), .C(mai_mai_n49_), .Y(mai_mai_n1396_));
  NO2        m1368(.A(mai_mai_n1058_), .B(h), .Y(mai_mai_n1397_));
  NA3        m1369(.A(mai_mai_n1397_), .B(d), .C(mai_mai_n1019_), .Y(mai_mai_n1398_));
  NO2        m1370(.A(mai_mai_n1398_), .B(c), .Y(mai_mai_n1399_));
  NA2        m1371(.A(mai_mai_n176_), .B(mai_mai_n109_), .Y(mai_mai_n1400_));
  NOi21      m1372(.An(d), .B(f), .Y(mai_mai_n1401_));
  NO2        m1373(.A(mai_mai_n1312_), .B(f), .Y(mai_mai_n1402_));
  INV        m1374(.A(mai_mai_n1399_), .Y(mai_mai_n1403_));
  NA3        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1395_), .C(mai_mai_n1386_), .Y(mai_mai_n1404_));
  NO3        m1376(.A(mai_mai_n1062_), .B(mai_mai_n1048_), .C(mai_mai_n40_), .Y(mai_mai_n1405_));
  OAI220     m1377(.A0(mai_mai_n455_), .A1(mai_mai_n297_), .B0(mai_mai_n128_), .B1(mai_mai_n59_), .Y(mai_mai_n1406_));
  OAI210     m1378(.A0(mai_mai_n1406_), .A1(mai_mai_n1405_), .B0(mai_mai_n1324_), .Y(mai_mai_n1407_));
  OAI210     m1379(.A0(mai_mai_n1366_), .A1(mai_mai_n1315_), .B0(mai_mai_n863_), .Y(mai_mai_n1408_));
  NO2        m1380(.A(mai_mai_n1016_), .B(mai_mai_n129_), .Y(mai_mai_n1409_));
  NA2        m1381(.A(mai_mai_n1409_), .B(mai_mai_n612_), .Y(mai_mai_n1410_));
  NA3        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1408_), .C(mai_mai_n1407_), .Y(mai_mai_n1411_));
  NA2        m1383(.A(mai_mai_n1339_), .B(mai_mai_n1401_), .Y(mai_mai_n1412_));
  NO2        m1384(.A(mai_mai_n1412_), .B(m), .Y(mai_mai_n1413_));
  NO2        m1385(.A(mai_mai_n145_), .B(mai_mai_n178_), .Y(mai_mai_n1414_));
  OAI210     m1386(.A0(mai_mai_n1414_), .A1(mai_mai_n107_), .B0(mai_mai_n1350_), .Y(mai_mai_n1415_));
  INV        m1387(.A(mai_mai_n1415_), .Y(mai_mai_n1416_));
  NO3        m1388(.A(mai_mai_n1416_), .B(mai_mai_n1413_), .C(mai_mai_n1411_), .Y(mai_mai_n1417_));
  NO2        m1389(.A(mai_mai_n1311_), .B(e), .Y(mai_mai_n1418_));
  NA2        m1390(.A(mai_mai_n1418_), .B(mai_mai_n396_), .Y(mai_mai_n1419_));
  OAI210     m1391(.A0(mai_mai_n1402_), .A1(mai_mai_n1100_), .B0(mai_mai_n623_), .Y(mai_mai_n1420_));
  OR3        m1392(.A(mai_mai_n1392_), .B(mai_mai_n1188_), .C(mai_mai_n129_), .Y(mai_mai_n1421_));
  OAI220     m1393(.A0(mai_mai_n1421_), .A1(mai_mai_n1419_), .B0(mai_mai_n1420_), .B1(mai_mai_n435_), .Y(mai_mai_n1422_));
  INV        m1394(.A(mai_mai_n1422_), .Y(mai_mai_n1423_));
  NO2        m1395(.A(mai_mai_n178_), .B(c), .Y(mai_mai_n1424_));
  OAI210     m1396(.A0(mai_mai_n1424_), .A1(mai_mai_n1418_), .B0(mai_mai_n176_), .Y(mai_mai_n1425_));
  AOI220     m1397(.A0(mai_mai_n1425_), .A1(mai_mai_n1050_), .B0(mai_mai_n525_), .B1(mai_mai_n356_), .Y(mai_mai_n1426_));
  NA2        m1398(.A(mai_mai_n533_), .B(g), .Y(mai_mai_n1427_));
  AOI210     m1399(.A0(mai_mai_n1427_), .A1(mai_mai_n1336_), .B0(mai_mai_n1396_), .Y(mai_mai_n1428_));
  NO2        m1400(.A(mai_mai_n1368_), .B(f), .Y(mai_mai_n1429_));
  NO2        m1401(.A(mai_mai_n1428_), .B(mai_mai_n206_), .Y(mai_mai_n1430_));
  NA2        m1402(.A(mai_mai_n1429_), .B(mai_mai_n1321_), .Y(mai_mai_n1431_));
  OAI220     m1403(.A0(mai_mai_n1431_), .A1(mai_mai_n49_), .B0(mai_mai_n1469_), .B1(mai_mai_n171_), .Y(mai_mai_n1432_));
  NA4        m1404(.A(mai_mai_n1071_), .B(mai_mai_n1068_), .C(mai_mai_n214_), .D(mai_mai_n68_), .Y(mai_mai_n1433_));
  NA2        m1405(.A(mai_mai_n1316_), .B(mai_mai_n179_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1435_));
  OAI210     m1407(.A0(mai_mai_n1368_), .A1(mai_mai_n842_), .B0(mai_mai_n474_), .Y(mai_mai_n1436_));
  OAI210     m1408(.A0(mai_mai_n1436_), .A1(mai_mai_n1074_), .B0(mai_mai_n1435_), .Y(mai_mai_n1437_));
  NO2        m1409(.A(m), .B(i), .Y(mai_mai_n1438_));
  BUFFER     m1410(.A(mai_mai_n1438_), .Y(mai_mai_n1439_));
  NA2        m1411(.A(mai_mai_n1439_), .B(mai_mai_n1338_), .Y(mai_mai_n1440_));
  NA4        m1412(.A(mai_mai_n1440_), .B(mai_mai_n1437_), .C(mai_mai_n1434_), .D(mai_mai_n1433_), .Y(mai_mai_n1441_));
  NO4        m1413(.A(mai_mai_n1441_), .B(mai_mai_n1432_), .C(mai_mai_n1430_), .D(mai_mai_n1426_), .Y(mai_mai_n1442_));
  NA3        m1414(.A(mai_mai_n1442_), .B(mai_mai_n1423_), .C(mai_mai_n1417_), .Y(mai_mai_n1443_));
  OAI210     m1415(.A0(mai_mai_n569_), .A1(g), .B0(mai_mai_n180_), .Y(mai_mai_n1444_));
  NA2        m1416(.A(mai_mai_n1444_), .B(mai_mai_n1397_), .Y(mai_mai_n1445_));
  AOI210     m1417(.A0(mai_mai_n151_), .A1(mai_mai_n56_), .B0(mai_mai_n1418_), .Y(mai_mai_n1446_));
  NO2        m1418(.A(mai_mai_n1446_), .B(mai_mai_n1400_), .Y(mai_mai_n1447_));
  NOi21      m1419(.An(mai_mai_n1316_), .B(e), .Y(mai_mai_n1448_));
  NO2        m1420(.A(mai_mai_n1448_), .B(mai_mai_n1447_), .Y(mai_mai_n1449_));
  NA2        m1421(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1450_));
  NO2        m1422(.A(mai_mai_n1319_), .B(mai_mai_n115_), .Y(mai_mai_n1451_));
  OAI220     m1423(.A0(mai_mai_n1451_), .A1(mai_mai_n1362_), .B0(mai_mai_n1374_), .B1(mai_mai_n1450_), .Y(mai_mai_n1452_));
  INV        m1424(.A(mai_mai_n1452_), .Y(mai_mai_n1453_));
  NA3        m1425(.A(mai_mai_n1453_), .B(mai_mai_n1449_), .C(mai_mai_n1445_), .Y(mai_mai_n1454_));
  OR4        m1426(.A(mai_mai_n1454_), .B(mai_mai_n1443_), .C(mai_mai_n1404_), .D(mai_mai_n1378_), .Y(mai04));
  NOi31      m1427(.An(mai_mai_n1366_), .B(mai_mai_n1367_), .C(mai_mai_n1021_), .Y(mai_mai_n1456_));
  NA2        m1428(.A(mai_mai_n1402_), .B(mai_mai_n808_), .Y(mai_mai_n1457_));
  NO3        m1429(.A(mai_mai_n1457_), .B(mai_mai_n1013_), .C(mai_mai_n475_), .Y(mai_mai_n1458_));
  OR3        m1430(.A(mai_mai_n1458_), .B(mai_mai_n1456_), .C(mai_mai_n1039_), .Y(mai_mai_n1459_));
  NO2        m1431(.A(mai_mai_n1321_), .B(mai_mai_n88_), .Y(mai_mai_n1460_));
  AOI210     m1432(.A0(mai_mai_n1460_), .A1(mai_mai_n1032_), .B0(mai_mai_n1165_), .Y(mai_mai_n1461_));
  NA2        m1433(.A(mai_mai_n1461_), .B(mai_mai_n1192_), .Y(mai_mai_n1462_));
  NO4        m1434(.A(mai_mai_n1462_), .B(mai_mai_n1459_), .C(mai_mai_n1047_), .D(mai_mai_n1026_), .Y(mai_mai_n1463_));
  NA4        m1435(.A(mai_mai_n1463_), .B(mai_mai_n1102_), .C(mai_mai_n1089_), .D(mai_mai_n1077_), .Y(mai05));
  INV        m1436(.A(l), .Y(mai_mai_n1467_));
  INV        m1437(.A(m), .Y(mai_mai_n1468_));
  INV        m1438(.A(mai_mai_n103_), .Y(mai_mai_n1469_));
  INV        m1439(.A(f), .Y(mai_mai_n1470_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  NAi41      u0034(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n63_));
  NA2        u0035(.A(g), .B(f), .Y(men_men_n64_));
  NO2        u0036(.A(men_men_n64_), .B(men_men_n63_), .Y(men_men_n65_));
  NAi21      u0037(.An(i), .B(j), .Y(men_men_n66_));
  NAi32      u0038(.An(n), .Bn(k), .C(m), .Y(men_men_n67_));
  NO2        u0039(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n68_));
  NAi31      u0040(.An(l), .B(m), .C(k), .Y(men_men_n69_));
  NAi21      u0041(.An(e), .B(h), .Y(men_men_n70_));
  NAi41      u0042(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n71_));
  NA2        u0043(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n72_));
  INV        u0044(.A(m), .Y(men_men_n73_));
  NOi21      u0045(.An(k), .B(l), .Y(men_men_n74_));
  NA2        u0046(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n75_));
  AN4        u0047(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n76_));
  NOi31      u0048(.An(h), .B(g), .C(f), .Y(men_men_n77_));
  NA2        u0049(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NAi32      u0050(.An(m), .Bn(k), .C(j), .Y(men_men_n79_));
  NOi32      u0051(.An(h), .Bn(g), .C(f), .Y(men_men_n80_));
  NA2        u0052(.A(men_men_n80_), .B(men_men_n76_), .Y(men_men_n81_));
  OA220      u0053(.A0(men_men_n81_), .A1(men_men_n79_), .B0(men_men_n78_), .B1(men_men_n75_), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n72_), .Y(men_men_n83_));
  INV        u0055(.A(n), .Y(men_men_n84_));
  NOi32      u0056(.An(e), .Bn(b), .C(d), .Y(men_men_n85_));
  NA2        u0057(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n86_));
  INV        u0058(.A(j), .Y(men_men_n87_));
  AN3        u0059(.A(m), .B(k), .C(i), .Y(men_men_n88_));
  NA3        u0060(.A(men_men_n88_), .B(men_men_n87_), .C(g), .Y(men_men_n89_));
  NO2        u0061(.A(men_men_n89_), .B(f), .Y(men_men_n90_));
  NAi32      u0062(.An(g), .Bn(f), .C(h), .Y(men_men_n91_));
  NAi31      u0063(.An(j), .B(m), .C(l), .Y(men_men_n92_));
  NO2        u0064(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  NA2        u0065(.A(m), .B(l), .Y(men_men_n94_));
  NAi31      u0066(.An(k), .B(j), .C(g), .Y(men_men_n95_));
  NO3        u0067(.A(men_men_n95_), .B(men_men_n94_), .C(f), .Y(men_men_n96_));
  AN2        u0068(.A(j), .B(g), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(l), .C(i), .Y(men_men_n98_));
  NOi21      u0070(.An(g), .B(i), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(j), .C(k), .Y(men_men_n100_));
  AOI220     u0072(.A0(men_men_n100_), .A1(men_men_n99_), .B0(men_men_n98_), .B1(men_men_n97_), .Y(men_men_n101_));
  NO2        u0073(.A(men_men_n101_), .B(f), .Y(men_men_n102_));
  NO4        u0074(.A(men_men_n102_), .B(men_men_n96_), .C(men_men_n93_), .D(men_men_n90_), .Y(men_men_n103_));
  NAi41      u0075(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n104_));
  AN2        u0076(.A(e), .B(b), .Y(men_men_n105_));
  NOi31      u0077(.An(c), .B(h), .C(f), .Y(men_men_n106_));
  NA2        u0078(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NO3        u0079(.A(men_men_n107_), .B(men_men_n104_), .C(g), .Y(men_men_n108_));
  NOi21      u0080(.An(g), .B(f), .Y(men_men_n109_));
  NOi21      u0081(.An(i), .B(h), .Y(men_men_n110_));
  NA3        u0082(.A(men_men_n110_), .B(men_men_n109_), .C(men_men_n36_), .Y(men_men_n111_));
  INV        u0083(.A(a), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n105_), .B(men_men_n112_), .Y(men_men_n113_));
  INV        u0085(.A(l), .Y(men_men_n114_));
  NOi21      u0086(.An(m), .B(n), .Y(men_men_n115_));
  AN2        u0087(.A(k), .B(h), .Y(men_men_n116_));
  NO2        u0088(.A(men_men_n111_), .B(men_men_n86_), .Y(men_men_n117_));
  INV        u0089(.A(b), .Y(men_men_n118_));
  NA2        u0090(.A(l), .B(j), .Y(men_men_n119_));
  AN2        u0091(.A(k), .B(i), .Y(men_men_n120_));
  NA2        u0092(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NA2        u0093(.A(g), .B(e), .Y(men_men_n122_));
  NOi32      u0094(.An(c), .Bn(a), .C(d), .Y(men_men_n123_));
  NA2        u0095(.A(men_men_n123_), .B(men_men_n115_), .Y(men_men_n124_));
  NO2        u0096(.A(men_men_n117_), .B(men_men_n108_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n103_), .A1(men_men_n86_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n77_), .C(men_men_n76_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(i), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n80_), .C(men_men_n76_), .Y(men_men_n130_));
  NA2        u0102(.A(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NOi32      u0103(.An(f), .Bn(b), .C(e), .Y(men_men_n132_));
  NAi21      u0104(.An(g), .B(h), .Y(men_men_n133_));
  NAi21      u0105(.An(m), .B(n), .Y(men_men_n134_));
  NAi21      u0106(.An(j), .B(k), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n136_));
  NAi41      u0108(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n137_));
  NAi31      u0109(.An(j), .B(k), .C(h), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n139_));
  AOI210     u0111(.A0(men_men_n136_), .A1(men_men_n132_), .B0(men_men_n139_), .Y(men_men_n140_));
  NO2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n141_), .B(men_men_n134_), .Y(men_men_n142_));
  AN2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  NAi21      u0115(.An(c), .B(b), .Y(men_men_n144_));
  NA2        u0116(.A(f), .B(d), .Y(men_men_n145_));
  NO4        u0117(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .D(men_men_n133_), .Y(men_men_n146_));
  NA2        u0118(.A(h), .B(c), .Y(men_men_n147_));
  NAi31      u0119(.An(f), .B(e), .C(b), .Y(men_men_n148_));
  NA2        u0120(.A(men_men_n146_), .B(men_men_n142_), .Y(men_men_n149_));
  NA2        u0121(.A(d), .B(b), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(f), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NA2        u0124(.A(b), .B(a), .Y(men_men_n153_));
  NAi21      u0125(.An(e), .B(g), .Y(men_men_n154_));
  NAi21      u0126(.An(c), .B(d), .Y(men_men_n155_));
  NAi31      u0127(.An(l), .B(k), .C(h), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n134_), .B(men_men_n156_), .Y(men_men_n157_));
  NA2        u0129(.A(men_men_n157_), .B(men_men_n152_), .Y(men_men_n158_));
  NAi41      u0130(.An(men_men_n131_), .B(men_men_n158_), .C(men_men_n149_), .D(men_men_n140_), .Y(men_men_n159_));
  NAi31      u0131(.An(e), .B(f), .C(b), .Y(men_men_n160_));
  NOi21      u0132(.An(g), .B(d), .Y(men_men_n161_));
  NO2        u0133(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NOi21      u0134(.An(h), .B(i), .Y(men_men_n163_));
  NOi21      u0135(.An(k), .B(m), .Y(men_men_n164_));
  NA3        u0136(.A(men_men_n164_), .B(men_men_n163_), .C(n), .Y(men_men_n165_));
  NOi21      u0137(.An(men_men_n162_), .B(men_men_n165_), .Y(men_men_n166_));
  NOi21      u0138(.An(h), .B(g), .Y(men_men_n167_));
  NO2        u0139(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n168_));
  NA2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NAi31      u0141(.An(l), .B(j), .C(h), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n170_), .B(men_men_n49_), .Y(men_men_n171_));
  NA2        u0143(.A(men_men_n171_), .B(men_men_n65_), .Y(men_men_n172_));
  NOi32      u0144(.An(n), .Bn(k), .C(m), .Y(men_men_n173_));
  NA2        u0145(.A(l), .B(i), .Y(men_men_n174_));
  NA2        u0146(.A(men_men_n174_), .B(men_men_n173_), .Y(men_men_n175_));
  OAI210     u0147(.A0(men_men_n175_), .A1(men_men_n169_), .B0(men_men_n172_), .Y(men_men_n176_));
  NAi31      u0148(.An(d), .B(f), .C(c), .Y(men_men_n177_));
  NAi31      u0149(.An(e), .B(f), .C(c), .Y(men_men_n178_));
  NA2        u0150(.A(men_men_n178_), .B(men_men_n177_), .Y(men_men_n179_));
  NA2        u0151(.A(j), .B(h), .Y(men_men_n180_));
  OR3        u0152(.A(n), .B(m), .C(k), .Y(men_men_n181_));
  NO2        u0153(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  NAi32      u0154(.An(m), .Bn(k), .C(n), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n180_), .Y(men_men_n184_));
  AOI220     u0156(.A0(men_men_n184_), .A1(men_men_n162_), .B0(men_men_n182_), .B1(men_men_n179_), .Y(men_men_n185_));
  NO2        u0157(.A(n), .B(m), .Y(men_men_n186_));
  NA2        u0158(.A(men_men_n186_), .B(men_men_n50_), .Y(men_men_n187_));
  NAi21      u0159(.An(f), .B(e), .Y(men_men_n188_));
  NA2        u0160(.A(d), .B(c), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NOi21      u0162(.An(men_men_n190_), .B(men_men_n187_), .Y(men_men_n191_));
  NAi21      u0163(.An(d), .B(c), .Y(men_men_n192_));
  NAi31      u0164(.An(m), .B(n), .C(b), .Y(men_men_n193_));
  NA2        u0165(.A(k), .B(i), .Y(men_men_n194_));
  NAi21      u0166(.An(h), .B(f), .Y(men_men_n195_));
  NO2        u0167(.A(men_men_n195_), .B(men_men_n194_), .Y(men_men_n196_));
  NO2        u0168(.A(men_men_n193_), .B(men_men_n155_), .Y(men_men_n197_));
  NA2        u0169(.A(men_men_n197_), .B(men_men_n196_), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(d), .Y(men_men_n199_));
  NOi32      u0171(.An(f), .Bn(c), .C(e), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n200_), .B(men_men_n199_), .Y(men_men_n201_));
  NO3        u0173(.A(n), .B(m), .C(j), .Y(men_men_n202_));
  NA2        u0174(.A(men_men_n202_), .B(men_men_n116_), .Y(men_men_n203_));
  AO210      u0175(.A0(men_men_n203_), .A1(men_men_n187_), .B0(men_men_n201_), .Y(men_men_n204_));
  NAi41      u0176(.An(men_men_n191_), .B(men_men_n204_), .C(men_men_n198_), .D(men_men_n185_), .Y(men_men_n205_));
  OR4        u0177(.A(men_men_n205_), .B(men_men_n176_), .C(men_men_n166_), .D(men_men_n159_), .Y(men_men_n206_));
  NO4        u0178(.A(men_men_n206_), .B(men_men_n126_), .C(men_men_n83_), .D(men_men_n55_), .Y(men_men_n207_));
  NA3        u0179(.A(m), .B(men_men_n114_), .C(j), .Y(men_men_n208_));
  NAi31      u0180(.An(n), .B(h), .C(g), .Y(men_men_n209_));
  NO2        u0181(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  NOi32      u0182(.An(m), .Bn(k), .C(l), .Y(men_men_n211_));
  NA3        u0183(.A(men_men_n211_), .B(men_men_n87_), .C(g), .Y(men_men_n212_));
  NO2        u0184(.A(men_men_n212_), .B(n), .Y(men_men_n213_));
  NOi21      u0185(.An(k), .B(j), .Y(men_men_n214_));
  NA4        u0186(.A(men_men_n214_), .B(men_men_n115_), .C(i), .D(g), .Y(men_men_n215_));
  AN2        u0187(.A(i), .B(g), .Y(men_men_n216_));
  NA3        u0188(.A(men_men_n74_), .B(men_men_n216_), .C(men_men_n115_), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n215_), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n213_), .C(men_men_n210_), .Y(men_men_n219_));
  NAi41      u0191(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n220_));
  INV        u0192(.A(men_men_n220_), .Y(men_men_n221_));
  INV        u0193(.A(f), .Y(men_men_n222_));
  INV        u0194(.A(g), .Y(men_men_n223_));
  NOi31      u0195(.An(i), .B(j), .C(h), .Y(men_men_n224_));
  NOi21      u0196(.An(l), .B(m), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NO3        u0198(.A(men_men_n226_), .B(men_men_n223_), .C(men_men_n222_), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n221_), .Y(men_men_n228_));
  OAI210     u0200(.A0(men_men_n219_), .A1(men_men_n32_), .B0(men_men_n228_), .Y(men_men_n229_));
  NOi21      u0201(.An(n), .B(m), .Y(men_men_n230_));
  NOi32      u0202(.An(l), .Bn(i), .C(j), .Y(men_men_n231_));
  NA2        u0203(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  OA220      u0204(.A0(men_men_n232_), .A1(men_men_n107_), .B0(men_men_n79_), .B1(men_men_n78_), .Y(men_men_n233_));
  NAi21      u0205(.An(j), .B(h), .Y(men_men_n234_));
  XN2        u0206(.A(i), .B(h), .Y(men_men_n235_));
  NA2        u0207(.A(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  NOi31      u0208(.An(k), .B(n), .C(m), .Y(men_men_n237_));
  NOi31      u0209(.An(men_men_n237_), .B(men_men_n189_), .C(men_men_n188_), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n238_), .B(men_men_n236_), .Y(men_men_n239_));
  NAi31      u0211(.An(f), .B(e), .C(c), .Y(men_men_n240_));
  NO4        u0212(.A(men_men_n240_), .B(men_men_n181_), .C(men_men_n180_), .D(men_men_n59_), .Y(men_men_n241_));
  NA4        u0213(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n242_));
  NAi32      u0214(.An(m), .Bn(i), .C(k), .Y(men_men_n243_));
  NO3        u0215(.A(men_men_n243_), .B(men_men_n91_), .C(men_men_n242_), .Y(men_men_n244_));
  INV        u0216(.A(k), .Y(men_men_n245_));
  NO2        u0217(.A(men_men_n244_), .B(men_men_n241_), .Y(men_men_n246_));
  NAi21      u0218(.An(n), .B(a), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n247_), .B(men_men_n150_), .Y(men_men_n248_));
  NAi41      u0220(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(e), .Y(men_men_n250_));
  NO3        u0222(.A(men_men_n151_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n251_));
  OAI210     u0223(.A0(men_men_n251_), .A1(men_men_n250_), .B0(men_men_n248_), .Y(men_men_n252_));
  AN4        u0224(.A(men_men_n252_), .B(men_men_n246_), .C(men_men_n239_), .D(men_men_n233_), .Y(men_men_n253_));
  OR2        u0225(.A(h), .B(g), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n254_), .B(men_men_n104_), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n255_), .B(men_men_n132_), .Y(men_men_n256_));
  NAi41      u0228(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n257_), .B(men_men_n222_), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n164_), .B(men_men_n110_), .Y(men_men_n259_));
  NAi21      u0231(.An(men_men_n259_), .B(men_men_n258_), .Y(men_men_n260_));
  NO2        u0232(.A(n), .B(a), .Y(men_men_n261_));
  NAi31      u0233(.An(men_men_n249_), .B(men_men_n261_), .C(men_men_n105_), .Y(men_men_n262_));
  AN2        u0234(.A(men_men_n262_), .B(men_men_n260_), .Y(men_men_n263_));
  NAi21      u0235(.An(h), .B(i), .Y(men_men_n264_));
  NA2        u0236(.A(men_men_n186_), .B(k), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA2        u0238(.A(men_men_n263_), .B(men_men_n256_), .Y(men_men_n267_));
  NOi21      u0239(.An(g), .B(e), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n269_));
  NA2        u0241(.A(men_men_n269_), .B(men_men_n268_), .Y(men_men_n270_));
  NOi32      u0242(.An(l), .Bn(j), .C(i), .Y(men_men_n271_));
  AOI210     u0243(.A0(men_men_n74_), .A1(men_men_n87_), .B0(men_men_n271_), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n264_), .B(men_men_n44_), .Y(men_men_n273_));
  NAi21      u0245(.An(f), .B(g), .Y(men_men_n274_));
  NO2        u0246(.A(men_men_n274_), .B(men_men_n63_), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n67_), .B(men_men_n119_), .Y(men_men_n276_));
  AOI220     u0248(.A0(men_men_n276_), .A1(men_men_n275_), .B0(men_men_n273_), .B1(men_men_n65_), .Y(men_men_n277_));
  OAI210     u0249(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n277_), .Y(men_men_n278_));
  NO3        u0250(.A(men_men_n135_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n279_));
  NOi41      u0251(.An(men_men_n253_), .B(men_men_n278_), .C(men_men_n267_), .D(men_men_n229_), .Y(men_men_n280_));
  NO4        u0252(.A(men_men_n210_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n281_));
  NO2        u0253(.A(men_men_n281_), .B(men_men_n113_), .Y(men_men_n282_));
  NA3        u0254(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n283_));
  NAi21      u0255(.An(h), .B(g), .Y(men_men_n284_));
  OR4        u0256(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n232_), .D(e), .Y(men_men_n285_));
  NO2        u0257(.A(men_men_n259_), .B(men_men_n274_), .Y(men_men_n286_));
  NAi31      u0258(.An(g), .B(k), .C(h), .Y(men_men_n287_));
  NO3        u0259(.A(men_men_n134_), .B(men_men_n287_), .C(l), .Y(men_men_n288_));
  NAi31      u0260(.An(e), .B(d), .C(a), .Y(men_men_n289_));
  NA2        u0261(.A(men_men_n288_), .B(men_men_n132_), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n290_), .B(men_men_n285_), .Y(men_men_n291_));
  NA4        u0263(.A(men_men_n164_), .B(men_men_n80_), .C(men_men_n76_), .D(men_men_n119_), .Y(men_men_n292_));
  BUFFER     u0264(.A(men_men_n292_), .Y(men_men_n293_));
  NA3        u0265(.A(e), .B(c), .C(b), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n60_), .B(men_men_n294_), .Y(men_men_n295_));
  NAi32      u0267(.An(k), .Bn(i), .C(j), .Y(men_men_n296_));
  INV        u0268(.A(men_men_n49_), .Y(men_men_n297_));
  OAI210     u0269(.A0(men_men_n275_), .A1(men_men_n295_), .B0(men_men_n297_), .Y(men_men_n298_));
  NAi21      u0270(.An(l), .B(k), .Y(men_men_n299_));
  NO2        u0271(.A(men_men_n299_), .B(men_men_n49_), .Y(men_men_n300_));
  NOi21      u0272(.An(l), .B(j), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n167_), .B(men_men_n301_), .Y(men_men_n302_));
  NA3        u0274(.A(men_men_n120_), .B(men_men_n119_), .C(g), .Y(men_men_n303_));
  OR3        u0275(.A(men_men_n71_), .B(men_men_n73_), .C(e), .Y(men_men_n304_));
  AOI210     u0276(.A0(men_men_n303_), .A1(men_men_n302_), .B0(men_men_n304_), .Y(men_men_n305_));
  INV        u0277(.A(men_men_n305_), .Y(men_men_n306_));
  NAi32      u0278(.An(j), .Bn(h), .C(i), .Y(men_men_n307_));
  NAi21      u0279(.An(m), .B(l), .Y(men_men_n308_));
  NO3        u0280(.A(men_men_n308_), .B(men_men_n307_), .C(men_men_n84_), .Y(men_men_n309_));
  NA2        u0281(.A(h), .B(g), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n173_), .B(men_men_n45_), .Y(men_men_n311_));
  NO2        u0283(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n312_));
  OAI210     u0284(.A0(men_men_n312_), .A1(men_men_n309_), .B0(men_men_n168_), .Y(men_men_n313_));
  NA4        u0285(.A(men_men_n313_), .B(men_men_n306_), .C(men_men_n298_), .D(men_men_n293_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n148_), .B(d), .Y(men_men_n315_));
  NA2        u0287(.A(men_men_n315_), .B(men_men_n53_), .Y(men_men_n316_));
  NAi32      u0288(.An(n), .Bn(m), .C(l), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n317_), .B(men_men_n307_), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n318_), .B(men_men_n190_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n124_), .B(men_men_n118_), .Y(men_men_n320_));
  NAi31      u0292(.An(k), .B(l), .C(j), .Y(men_men_n321_));
  OAI210     u0293(.A0(men_men_n299_), .A1(j), .B0(men_men_n321_), .Y(men_men_n322_));
  NOi21      u0294(.An(men_men_n322_), .B(men_men_n122_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n319_), .B(men_men_n316_), .Y(men_men_n324_));
  NO4        u0296(.A(men_men_n324_), .B(men_men_n314_), .C(men_men_n291_), .D(men_men_n282_), .Y(men_men_n325_));
  NA2        u0297(.A(men_men_n266_), .B(men_men_n200_), .Y(men_men_n326_));
  NAi21      u0298(.An(m), .B(k), .Y(men_men_n327_));
  NO2        u0299(.A(men_men_n235_), .B(men_men_n327_), .Y(men_men_n328_));
  NAi41      u0300(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n329_), .B(men_men_n154_), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n330_), .B(men_men_n328_), .Y(men_men_n331_));
  NAi31      u0303(.An(i), .B(l), .C(h), .Y(men_men_n332_));
  NO4        u0304(.A(men_men_n332_), .B(men_men_n154_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n333_));
  NA2        u0305(.A(e), .B(c), .Y(men_men_n334_));
  NO3        u0306(.A(men_men_n334_), .B(n), .C(d), .Y(men_men_n335_));
  NOi21      u0307(.An(f), .B(h), .Y(men_men_n336_));
  NA2        u0308(.A(men_men_n336_), .B(men_men_n120_), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n337_), .B(men_men_n223_), .Y(men_men_n338_));
  NAi31      u0310(.An(d), .B(e), .C(b), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n134_), .B(men_men_n339_), .Y(men_men_n340_));
  NAi31      u0312(.An(men_men_n333_), .B(men_men_n331_), .C(men_men_n326_), .Y(men_men_n341_));
  NO4        u0313(.A(men_men_n329_), .B(men_men_n79_), .C(men_men_n70_), .D(men_men_n223_), .Y(men_men_n342_));
  NA2        u0314(.A(men_men_n261_), .B(men_men_n105_), .Y(men_men_n343_));
  OR2        u0315(.A(men_men_n343_), .B(men_men_n212_), .Y(men_men_n344_));
  NOi31      u0316(.An(l), .B(n), .C(m), .Y(men_men_n345_));
  NA2        u0317(.A(men_men_n345_), .B(men_men_n224_), .Y(men_men_n346_));
  NO2        u0318(.A(men_men_n346_), .B(men_men_n201_), .Y(men_men_n347_));
  NAi32      u0319(.An(men_men_n347_), .Bn(men_men_n342_), .C(men_men_n344_), .Y(men_men_n348_));
  NAi32      u0320(.An(m), .Bn(j), .C(k), .Y(men_men_n349_));
  NAi41      u0321(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n350_));
  NA2        u0322(.A(men_men_n220_), .B(men_men_n350_), .Y(men_men_n351_));
  NOi31      u0323(.An(j), .B(m), .C(k), .Y(men_men_n352_));
  NO2        u0324(.A(men_men_n127_), .B(men_men_n352_), .Y(men_men_n353_));
  AN3        u0325(.A(h), .B(g), .C(f), .Y(men_men_n354_));
  NAi31      u0326(.An(men_men_n353_), .B(men_men_n354_), .C(men_men_n351_), .Y(men_men_n355_));
  NOi32      u0327(.An(m), .Bn(j), .C(l), .Y(men_men_n356_));
  NO2        u0328(.A(men_men_n356_), .B(men_men_n98_), .Y(men_men_n357_));
  NAi32      u0329(.An(men_men_n357_), .Bn(men_men_n209_), .C(men_men_n315_), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n308_), .B(men_men_n307_), .Y(men_men_n359_));
  NO2        u0331(.A(men_men_n226_), .B(g), .Y(men_men_n360_));
  NO2        u0332(.A(men_men_n160_), .B(men_men_n84_), .Y(men_men_n361_));
  AOI220     u0333(.A0(men_men_n361_), .A1(men_men_n360_), .B0(men_men_n258_), .B1(men_men_n359_), .Y(men_men_n362_));
  INV        u0334(.A(men_men_n243_), .Y(men_men_n363_));
  NA3        u0335(.A(men_men_n363_), .B(men_men_n354_), .C(men_men_n221_), .Y(men_men_n364_));
  NA4        u0336(.A(men_men_n364_), .B(men_men_n362_), .C(men_men_n358_), .D(men_men_n355_), .Y(men_men_n365_));
  NA3        u0337(.A(h), .B(g), .C(f), .Y(men_men_n366_));
  NO2        u0338(.A(men_men_n366_), .B(men_men_n75_), .Y(men_men_n367_));
  NA2        u0339(.A(men_men_n350_), .B(men_men_n220_), .Y(men_men_n368_));
  NA2        u0340(.A(men_men_n167_), .B(e), .Y(men_men_n369_));
  NO2        u0341(.A(men_men_n369_), .B(men_men_n41_), .Y(men_men_n370_));
  AOI220     u0342(.A0(men_men_n370_), .A1(men_men_n320_), .B0(men_men_n368_), .B1(men_men_n367_), .Y(men_men_n371_));
  NOi32      u0343(.An(j), .Bn(g), .C(i), .Y(men_men_n372_));
  NA3        u0344(.A(men_men_n372_), .B(men_men_n299_), .C(men_men_n115_), .Y(men_men_n373_));
  AO210      u0345(.A0(men_men_n113_), .A1(men_men_n32_), .B0(men_men_n373_), .Y(men_men_n374_));
  NOi32      u0346(.An(e), .Bn(b), .C(a), .Y(men_men_n375_));
  AN2        u0347(.A(l), .B(j), .Y(men_men_n376_));
  INV        u0348(.A(men_men_n327_), .Y(men_men_n377_));
  NO3        u0349(.A(men_men_n329_), .B(men_men_n70_), .C(men_men_n223_), .Y(men_men_n378_));
  NA3        u0350(.A(men_men_n217_), .B(men_men_n215_), .C(men_men_n35_), .Y(men_men_n379_));
  AOI220     u0351(.A0(men_men_n379_), .A1(men_men_n375_), .B0(men_men_n378_), .B1(men_men_n377_), .Y(men_men_n380_));
  NO2        u0352(.A(men_men_n339_), .B(n), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n216_), .B(k), .Y(men_men_n382_));
  NA3        u0354(.A(m), .B(men_men_n114_), .C(men_men_n222_), .Y(men_men_n383_));
  NA4        u0355(.A(men_men_n211_), .B(men_men_n87_), .C(g), .D(men_men_n222_), .Y(men_men_n384_));
  OAI210     u0356(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n384_), .Y(men_men_n385_));
  NAi41      u0357(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n51_), .B(men_men_n115_), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n388_));
  AOI220     u0360(.A0(men_men_n388_), .A1(b), .B0(men_men_n385_), .B1(men_men_n381_), .Y(men_men_n389_));
  NA4        u0361(.A(men_men_n389_), .B(men_men_n380_), .C(men_men_n374_), .D(men_men_n371_), .Y(men_men_n390_));
  NO4        u0362(.A(men_men_n390_), .B(men_men_n365_), .C(men_men_n348_), .D(men_men_n341_), .Y(men_men_n391_));
  NA4        u0363(.A(men_men_n391_), .B(men_men_n325_), .C(men_men_n280_), .D(men_men_n207_), .Y(men10));
  NA3        u0364(.A(m), .B(k), .C(i), .Y(men_men_n393_));
  NO3        u0365(.A(men_men_n393_), .B(j), .C(men_men_n223_), .Y(men_men_n394_));
  NOi21      u0366(.An(e), .B(f), .Y(men_men_n395_));
  NO4        u0367(.A(men_men_n155_), .B(men_men_n395_), .C(n), .D(men_men_n112_), .Y(men_men_n396_));
  NAi31      u0368(.An(b), .B(f), .C(c), .Y(men_men_n397_));
  INV        u0369(.A(men_men_n397_), .Y(men_men_n398_));
  NOi32      u0370(.An(k), .Bn(h), .C(j), .Y(men_men_n399_));
  NA2        u0371(.A(men_men_n399_), .B(men_men_n230_), .Y(men_men_n400_));
  NA2        u0372(.A(men_men_n165_), .B(men_men_n400_), .Y(men_men_n401_));
  AOI220     u0373(.A0(men_men_n401_), .A1(men_men_n398_), .B0(men_men_n396_), .B1(men_men_n394_), .Y(men_men_n402_));
  AN2        u0374(.A(j), .B(h), .Y(men_men_n403_));
  NO3        u0375(.A(n), .B(m), .C(k), .Y(men_men_n404_));
  NA2        u0376(.A(men_men_n404_), .B(men_men_n403_), .Y(men_men_n405_));
  NO3        u0377(.A(men_men_n405_), .B(men_men_n155_), .C(men_men_n222_), .Y(men_men_n406_));
  OR2        u0378(.A(m), .B(k), .Y(men_men_n407_));
  NO2        u0379(.A(men_men_n180_), .B(men_men_n407_), .Y(men_men_n408_));
  NA4        u0380(.A(n), .B(f), .C(c), .D(men_men_n118_), .Y(men_men_n409_));
  NOi21      u0381(.An(men_men_n408_), .B(men_men_n409_), .Y(men_men_n410_));
  NOi32      u0382(.An(d), .Bn(a), .C(c), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n411_), .B(men_men_n188_), .Y(men_men_n412_));
  NAi21      u0384(.An(i), .B(g), .Y(men_men_n413_));
  NAi31      u0385(.An(k), .B(m), .C(j), .Y(men_men_n414_));
  NO3        u0386(.A(men_men_n414_), .B(men_men_n413_), .C(n), .Y(men_men_n415_));
  NOi21      u0387(.An(men_men_n415_), .B(men_men_n412_), .Y(men_men_n416_));
  NO3        u0388(.A(men_men_n416_), .B(men_men_n410_), .C(men_men_n406_), .Y(men_men_n417_));
  NO2        u0389(.A(men_men_n409_), .B(men_men_n308_), .Y(men_men_n418_));
  NOi32      u0390(.An(f), .Bn(d), .C(c), .Y(men_men_n419_));
  AOI220     u0391(.A0(men_men_n419_), .A1(men_men_n318_), .B0(men_men_n418_), .B1(men_men_n224_), .Y(men_men_n420_));
  NA3        u0392(.A(men_men_n420_), .B(men_men_n417_), .C(men_men_n402_), .Y(men_men_n421_));
  NO2        u0393(.A(men_men_n59_), .B(men_men_n118_), .Y(men_men_n422_));
  NA2        u0394(.A(men_men_n261_), .B(men_men_n422_), .Y(men_men_n423_));
  INV        u0395(.A(e), .Y(men_men_n424_));
  NA2        u0396(.A(men_men_n46_), .B(e), .Y(men_men_n425_));
  OAI220     u0397(.A0(men_men_n425_), .A1(men_men_n208_), .B0(men_men_n212_), .B1(men_men_n424_), .Y(men_men_n426_));
  AN2        u0398(.A(g), .B(e), .Y(men_men_n427_));
  NA3        u0399(.A(men_men_n427_), .B(men_men_n211_), .C(i), .Y(men_men_n428_));
  OAI210     u0400(.A0(men_men_n89_), .A1(men_men_n424_), .B0(men_men_n428_), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n101_), .B(men_men_n424_), .Y(men_men_n430_));
  NO3        u0402(.A(men_men_n430_), .B(men_men_n429_), .C(men_men_n426_), .Y(men_men_n431_));
  NOi32      u0403(.An(h), .Bn(e), .C(g), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n432_), .B(men_men_n301_), .C(m), .Y(men_men_n433_));
  NOi21      u0405(.An(g), .B(h), .Y(men_men_n434_));
  AN3        u0406(.A(m), .B(l), .C(i), .Y(men_men_n435_));
  NA3        u0407(.A(men_men_n435_), .B(men_men_n434_), .C(e), .Y(men_men_n436_));
  AN3        u0408(.A(h), .B(g), .C(e), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n437_), .B(men_men_n98_), .Y(men_men_n438_));
  AN3        u0410(.A(men_men_n438_), .B(men_men_n436_), .C(men_men_n433_), .Y(men_men_n439_));
  AOI210     u0411(.A0(men_men_n439_), .A1(men_men_n431_), .B0(men_men_n423_), .Y(men_men_n440_));
  NA3        u0412(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n441_), .B(men_men_n423_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n411_), .B(men_men_n188_), .C(men_men_n84_), .Y(men_men_n443_));
  NAi31      u0415(.An(b), .B(c), .C(a), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n444_), .B(n), .Y(men_men_n445_));
  OAI210     u0417(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n446_), .B(men_men_n151_), .Y(men_men_n447_));
  NA2        u0419(.A(men_men_n447_), .B(men_men_n445_), .Y(men_men_n448_));
  INV        u0420(.A(men_men_n448_), .Y(men_men_n449_));
  NO4        u0421(.A(men_men_n449_), .B(men_men_n442_), .C(men_men_n440_), .D(men_men_n421_), .Y(men_men_n450_));
  NA2        u0422(.A(i), .B(g), .Y(men_men_n451_));
  NO3        u0423(.A(men_men_n289_), .B(men_men_n451_), .C(c), .Y(men_men_n452_));
  NOi21      u0424(.An(a), .B(n), .Y(men_men_n453_));
  NOi21      u0425(.An(d), .B(c), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  NA3        u0427(.A(i), .B(g), .C(f), .Y(men_men_n456_));
  OR2        u0428(.A(men_men_n456_), .B(men_men_n69_), .Y(men_men_n457_));
  NA3        u0429(.A(men_men_n435_), .B(men_men_n434_), .C(men_men_n188_), .Y(men_men_n458_));
  AOI210     u0430(.A0(men_men_n458_), .A1(men_men_n457_), .B0(men_men_n455_), .Y(men_men_n459_));
  AOI210     u0431(.A0(men_men_n452_), .A1(men_men_n300_), .B0(men_men_n459_), .Y(men_men_n460_));
  OR2        u0432(.A(n), .B(m), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n461_), .B(men_men_n156_), .Y(men_men_n462_));
  NO2        u0434(.A(men_men_n189_), .B(men_men_n151_), .Y(men_men_n463_));
  OAI210     u0435(.A0(men_men_n462_), .A1(men_men_n182_), .B0(men_men_n463_), .Y(men_men_n464_));
  INV        u0436(.A(men_men_n387_), .Y(men_men_n465_));
  NA3        u0437(.A(men_men_n465_), .B(men_men_n375_), .C(d), .Y(men_men_n466_));
  NO2        u0438(.A(men_men_n444_), .B(men_men_n49_), .Y(men_men_n467_));
  NO3        u0439(.A(men_men_n64_), .B(men_men_n114_), .C(e), .Y(men_men_n468_));
  NAi21      u0440(.An(k), .B(j), .Y(men_men_n469_));
  NA2        u0441(.A(men_men_n264_), .B(men_men_n469_), .Y(men_men_n470_));
  NA3        u0442(.A(men_men_n470_), .B(men_men_n468_), .C(men_men_n467_), .Y(men_men_n471_));
  NAi21      u0443(.An(e), .B(d), .Y(men_men_n472_));
  INV        u0444(.A(men_men_n472_), .Y(men_men_n473_));
  NO2        u0445(.A(men_men_n265_), .B(men_men_n222_), .Y(men_men_n474_));
  NA3        u0446(.A(men_men_n474_), .B(men_men_n473_), .C(men_men_n236_), .Y(men_men_n475_));
  NA4        u0447(.A(men_men_n475_), .B(men_men_n471_), .C(men_men_n466_), .D(men_men_n464_), .Y(men_men_n476_));
  NO2        u0448(.A(men_men_n346_), .B(men_men_n222_), .Y(men_men_n477_));
  NA2        u0449(.A(men_men_n477_), .B(men_men_n473_), .Y(men_men_n478_));
  NOi31      u0450(.An(n), .B(m), .C(k), .Y(men_men_n479_));
  AOI220     u0451(.A0(men_men_n479_), .A1(men_men_n403_), .B0(men_men_n230_), .B1(men_men_n50_), .Y(men_men_n480_));
  NAi31      u0452(.An(g), .B(f), .C(c), .Y(men_men_n481_));
  OR3        u0453(.A(men_men_n481_), .B(men_men_n480_), .C(e), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n482_), .B(men_men_n478_), .C(men_men_n319_), .Y(men_men_n483_));
  NOi41      u0455(.An(men_men_n460_), .B(men_men_n483_), .C(men_men_n476_), .D(men_men_n278_), .Y(men_men_n484_));
  NOi32      u0456(.An(c), .Bn(a), .C(b), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n485_), .B(men_men_n115_), .Y(men_men_n486_));
  INV        u0458(.A(men_men_n287_), .Y(men_men_n487_));
  AN2        u0459(.A(e), .B(d), .Y(men_men_n488_));
  NA2        u0460(.A(men_men_n488_), .B(men_men_n487_), .Y(men_men_n489_));
  INV        u0461(.A(men_men_n151_), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n133_), .B(men_men_n41_), .Y(men_men_n491_));
  NO2        u0463(.A(men_men_n64_), .B(e), .Y(men_men_n492_));
  NOi31      u0464(.An(j), .B(k), .C(i), .Y(men_men_n493_));
  NOi21      u0465(.An(men_men_n170_), .B(men_men_n493_), .Y(men_men_n494_));
  NA4        u0466(.A(men_men_n332_), .B(men_men_n494_), .C(men_men_n272_), .D(men_men_n121_), .Y(men_men_n495_));
  AOI220     u0467(.A0(men_men_n495_), .A1(men_men_n492_), .B0(men_men_n491_), .B1(men_men_n490_), .Y(men_men_n496_));
  AOI210     u0468(.A0(men_men_n496_), .A1(men_men_n489_), .B0(men_men_n486_), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n218_), .B(men_men_n213_), .Y(men_men_n498_));
  NOi21      u0470(.An(a), .B(b), .Y(men_men_n499_));
  NA3        u0471(.A(e), .B(d), .C(c), .Y(men_men_n500_));
  NAi21      u0472(.An(men_men_n500_), .B(men_men_n499_), .Y(men_men_n501_));
  NO2        u0473(.A(men_men_n443_), .B(men_men_n212_), .Y(men_men_n502_));
  NOi21      u0474(.An(men_men_n501_), .B(men_men_n502_), .Y(men_men_n503_));
  AOI210     u0475(.A0(men_men_n281_), .A1(men_men_n498_), .B0(men_men_n503_), .Y(men_men_n504_));
  NO4        u0476(.A(men_men_n195_), .B(men_men_n104_), .C(men_men_n56_), .D(b), .Y(men_men_n505_));
  OR2        u0477(.A(k), .B(j), .Y(men_men_n506_));
  NA2        u0478(.A(l), .B(k), .Y(men_men_n507_));
  OR3        u0479(.A(men_men_n1588_), .B(men_men_n147_), .C(men_men_n137_), .Y(men_men_n508_));
  NA3        u0480(.A(men_men_n292_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n411_), .B(men_men_n115_), .Y(men_men_n510_));
  NO4        u0482(.A(men_men_n510_), .B(men_men_n95_), .C(men_men_n114_), .D(e), .Y(men_men_n511_));
  NO3        u0483(.A(men_men_n443_), .B(men_men_n92_), .C(men_men_n133_), .Y(men_men_n512_));
  NO4        u0484(.A(men_men_n512_), .B(men_men_n511_), .C(men_men_n509_), .D(men_men_n333_), .Y(men_men_n513_));
  NA2        u0485(.A(men_men_n513_), .B(men_men_n508_), .Y(men_men_n514_));
  NO4        u0486(.A(men_men_n514_), .B(men_men_n505_), .C(men_men_n504_), .D(men_men_n497_), .Y(men_men_n515_));
  NA2        u0487(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n516_));
  NAi31      u0488(.An(j), .B(l), .C(i), .Y(men_men_n517_));
  OAI210     u0489(.A0(men_men_n517_), .A1(men_men_n134_), .B0(men_men_n104_), .Y(men_men_n518_));
  NO3        u0490(.A(men_men_n412_), .B(men_men_n357_), .C(men_men_n209_), .Y(men_men_n519_));
  NO2        u0491(.A(men_men_n412_), .B(men_men_n387_), .Y(men_men_n520_));
  NO3        u0492(.A(men_men_n520_), .B(men_men_n519_), .C(men_men_n191_), .Y(men_men_n521_));
  NA3        u0493(.A(men_men_n521_), .B(men_men_n516_), .C(men_men_n253_), .Y(men_men_n522_));
  OAI210     u0494(.A0(men_men_n129_), .A1(men_men_n127_), .B0(n), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n523_), .B(men_men_n133_), .Y(men_men_n524_));
  OR2        u0496(.A(men_men_n309_), .B(men_men_n255_), .Y(men_men_n525_));
  OA210      u0497(.A0(men_men_n525_), .A1(men_men_n524_), .B0(men_men_n200_), .Y(men_men_n526_));
  XO2        u0498(.A(i), .B(h), .Y(men_men_n527_));
  NA3        u0499(.A(men_men_n527_), .B(men_men_n164_), .C(n), .Y(men_men_n528_));
  NAi41      u0500(.An(men_men_n309_), .B(men_men_n528_), .C(men_men_n480_), .D(men_men_n400_), .Y(men_men_n529_));
  NOi32      u0501(.An(men_men_n529_), .Bn(men_men_n492_), .C(men_men_n283_), .Y(men_men_n530_));
  NAi31      u0502(.An(c), .B(f), .C(d), .Y(men_men_n531_));
  NO2        u0503(.A(men_men_n203_), .B(men_men_n531_), .Y(men_men_n532_));
  BUFFER     u0504(.A(men_men_n82_), .Y(men_men_n533_));
  NA3        u0505(.A(men_men_n396_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n534_));
  NA2        u0506(.A(men_men_n237_), .B(men_men_n110_), .Y(men_men_n535_));
  AOI210     u0507(.A0(men_men_n535_), .A1(men_men_n187_), .B0(men_men_n531_), .Y(men_men_n536_));
  AOI210     u0508(.A0(men_men_n373_), .A1(men_men_n35_), .B0(men_men_n501_), .Y(men_men_n537_));
  NOi31      u0509(.An(men_men_n534_), .B(men_men_n537_), .C(men_men_n536_), .Y(men_men_n538_));
  AO220      u0510(.A0(men_men_n297_), .A1(men_men_n275_), .B0(men_men_n171_), .B1(men_men_n65_), .Y(men_men_n539_));
  NA3        u0511(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n540_));
  NO2        u0512(.A(men_men_n540_), .B(men_men_n455_), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(men_men_n305_), .Y(men_men_n542_));
  NAi41      u0514(.An(men_men_n539_), .B(men_men_n542_), .C(men_men_n538_), .D(men_men_n533_), .Y(men_men_n543_));
  NO4        u0515(.A(men_men_n543_), .B(men_men_n530_), .C(men_men_n526_), .D(men_men_n522_), .Y(men_men_n544_));
  NA4        u0516(.A(men_men_n544_), .B(men_men_n515_), .C(men_men_n484_), .D(men_men_n450_), .Y(men11));
  NO2        u0517(.A(men_men_n71_), .B(f), .Y(men_men_n546_));
  NA2        u0518(.A(j), .B(g), .Y(men_men_n547_));
  NAi31      u0519(.An(i), .B(m), .C(l), .Y(men_men_n548_));
  NA3        u0520(.A(m), .B(k), .C(j), .Y(men_men_n549_));
  OAI220     u0521(.A0(men_men_n549_), .A1(men_men_n133_), .B0(men_men_n548_), .B1(men_men_n547_), .Y(men_men_n550_));
  NA2        u0522(.A(men_men_n550_), .B(men_men_n546_), .Y(men_men_n551_));
  NOi32      u0523(.An(e), .Bn(b), .C(f), .Y(men_men_n552_));
  NA2        u0524(.A(men_men_n271_), .B(men_men_n115_), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n46_), .B(j), .Y(men_men_n554_));
  NO2        u0526(.A(men_men_n554_), .B(men_men_n311_), .Y(men_men_n555_));
  NAi31      u0527(.An(d), .B(e), .C(a), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n556_), .B(n), .Y(men_men_n557_));
  AOI220     u0529(.A0(men_men_n557_), .A1(men_men_n102_), .B0(men_men_n555_), .B1(men_men_n552_), .Y(men_men_n558_));
  NAi41      u0530(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n559_));
  AN2        u0531(.A(men_men_n559_), .B(men_men_n386_), .Y(men_men_n560_));
  AOI210     u0532(.A0(men_men_n560_), .A1(men_men_n412_), .B0(men_men_n284_), .Y(men_men_n561_));
  NA2        u0533(.A(j), .B(i), .Y(men_men_n562_));
  NAi31      u0534(.An(n), .B(m), .C(k), .Y(men_men_n563_));
  NO3        u0535(.A(men_men_n563_), .B(men_men_n562_), .C(men_men_n114_), .Y(men_men_n564_));
  NO4        u0536(.A(n), .B(d), .C(men_men_n118_), .D(a), .Y(men_men_n565_));
  OR2        u0537(.A(n), .B(c), .Y(men_men_n566_));
  NO2        u0538(.A(men_men_n566_), .B(men_men_n153_), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(men_men_n565_), .Y(men_men_n568_));
  NOi32      u0540(.An(g), .Bn(f), .C(i), .Y(men_men_n569_));
  AOI220     u0541(.A0(men_men_n569_), .A1(men_men_n100_), .B0(men_men_n550_), .B1(f), .Y(men_men_n570_));
  NO2        u0542(.A(men_men_n287_), .B(men_men_n49_), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n570_), .B(men_men_n568_), .Y(men_men_n572_));
  AOI210     u0544(.A0(men_men_n564_), .A1(men_men_n561_), .B0(men_men_n572_), .Y(men_men_n573_));
  NA2        u0545(.A(men_men_n143_), .B(men_men_n34_), .Y(men_men_n574_));
  OAI220     u0546(.A0(men_men_n574_), .A1(m), .B0(men_men_n554_), .B1(men_men_n243_), .Y(men_men_n575_));
  NOi41      u0547(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n576_));
  NAi32      u0548(.An(e), .Bn(b), .C(c), .Y(men_men_n577_));
  OR2        u0549(.A(men_men_n577_), .B(men_men_n84_), .Y(men_men_n578_));
  AN2        u0550(.A(men_men_n350_), .B(men_men_n329_), .Y(men_men_n579_));
  NA2        u0551(.A(men_men_n579_), .B(men_men_n578_), .Y(men_men_n580_));
  OA210      u0552(.A0(men_men_n580_), .A1(men_men_n576_), .B0(men_men_n575_), .Y(men_men_n581_));
  OAI220     u0553(.A0(men_men_n414_), .A1(men_men_n413_), .B0(men_men_n548_), .B1(men_men_n547_), .Y(men_men_n582_));
  NAi31      u0554(.An(d), .B(c), .C(a), .Y(men_men_n583_));
  NO2        u0555(.A(men_men_n583_), .B(n), .Y(men_men_n584_));
  NA3        u0556(.A(men_men_n584_), .B(men_men_n582_), .C(e), .Y(men_men_n585_));
  NO3        u0557(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n223_), .Y(men_men_n586_));
  NO2        u0558(.A(men_men_n240_), .B(men_men_n112_), .Y(men_men_n587_));
  OAI210     u0559(.A0(men_men_n586_), .A1(men_men_n415_), .B0(men_men_n587_), .Y(men_men_n588_));
  NA2        u0560(.A(men_men_n588_), .B(men_men_n585_), .Y(men_men_n589_));
  NO2        u0561(.A(men_men_n289_), .B(n), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n445_), .B(men_men_n590_), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n582_), .B(f), .Y(men_men_n592_));
  NAi32      u0564(.An(d), .Bn(a), .C(b), .Y(men_men_n593_));
  NO2        u0565(.A(men_men_n593_), .B(men_men_n49_), .Y(men_men_n594_));
  NA2        u0566(.A(h), .B(f), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n595_), .B(men_men_n95_), .Y(men_men_n596_));
  NO3        u0568(.A(men_men_n183_), .B(men_men_n180_), .C(g), .Y(men_men_n597_));
  AOI220     u0569(.A0(men_men_n597_), .A1(men_men_n58_), .B0(men_men_n596_), .B1(men_men_n594_), .Y(men_men_n598_));
  OAI210     u0570(.A0(men_men_n592_), .A1(men_men_n591_), .B0(men_men_n598_), .Y(men_men_n599_));
  AN3        u0571(.A(j), .B(h), .C(g), .Y(men_men_n600_));
  NO2        u0572(.A(men_men_n150_), .B(c), .Y(men_men_n601_));
  NA3        u0573(.A(men_men_n601_), .B(men_men_n600_), .C(men_men_n479_), .Y(men_men_n602_));
  NA3        u0574(.A(f), .B(d), .C(b), .Y(men_men_n603_));
  NO4        u0575(.A(men_men_n603_), .B(men_men_n183_), .C(men_men_n180_), .D(g), .Y(men_men_n604_));
  NAi21      u0576(.An(men_men_n604_), .B(men_men_n602_), .Y(men_men_n605_));
  NO4        u0577(.A(men_men_n605_), .B(men_men_n599_), .C(men_men_n589_), .D(men_men_n581_), .Y(men_men_n606_));
  AN4        u0578(.A(men_men_n606_), .B(men_men_n573_), .C(men_men_n558_), .D(men_men_n551_), .Y(men_men_n607_));
  INV        u0579(.A(k), .Y(men_men_n608_));
  NA3        u0580(.A(l), .B(men_men_n608_), .C(i), .Y(men_men_n609_));
  INV        u0581(.A(men_men_n609_), .Y(men_men_n610_));
  NA4        u0582(.A(men_men_n411_), .B(men_men_n434_), .C(men_men_n188_), .D(men_men_n115_), .Y(men_men_n611_));
  NAi32      u0583(.An(h), .Bn(f), .C(g), .Y(men_men_n612_));
  NAi41      u0584(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n613_));
  OAI210     u0585(.A0(men_men_n556_), .A1(n), .B0(men_men_n613_), .Y(men_men_n614_));
  NA2        u0586(.A(men_men_n614_), .B(m), .Y(men_men_n615_));
  NAi31      u0587(.An(h), .B(g), .C(f), .Y(men_men_n616_));
  OR3        u0588(.A(men_men_n616_), .B(men_men_n289_), .C(men_men_n49_), .Y(men_men_n617_));
  NA4        u0589(.A(men_men_n434_), .B(men_men_n123_), .C(men_men_n115_), .D(e), .Y(men_men_n618_));
  AN2        u0590(.A(men_men_n618_), .B(men_men_n617_), .Y(men_men_n619_));
  OA210      u0591(.A0(men_men_n615_), .A1(men_men_n612_), .B0(men_men_n619_), .Y(men_men_n620_));
  NO3        u0592(.A(men_men_n612_), .B(men_men_n71_), .C(men_men_n73_), .Y(men_men_n621_));
  NO4        u0593(.A(men_men_n616_), .B(men_men_n566_), .C(men_men_n153_), .D(men_men_n73_), .Y(men_men_n622_));
  OR2        u0594(.A(men_men_n622_), .B(men_men_n621_), .Y(men_men_n623_));
  NAi31      u0595(.An(men_men_n623_), .B(men_men_n620_), .C(men_men_n611_), .Y(men_men_n624_));
  NAi31      u0596(.An(f), .B(h), .C(g), .Y(men_men_n625_));
  NO4        u0597(.A(men_men_n321_), .B(men_men_n625_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n626_));
  NOi32      u0598(.An(b), .Bn(a), .C(c), .Y(men_men_n627_));
  NOi41      u0599(.An(men_men_n627_), .B(men_men_n366_), .C(men_men_n67_), .D(men_men_n119_), .Y(men_men_n628_));
  OR2        u0600(.A(men_men_n628_), .B(men_men_n626_), .Y(men_men_n629_));
  NOi32      u0601(.An(d), .Bn(a), .C(e), .Y(men_men_n630_));
  NA2        u0602(.A(men_men_n630_), .B(men_men_n115_), .Y(men_men_n631_));
  NO2        u0603(.A(n), .B(c), .Y(men_men_n632_));
  NA3        u0604(.A(men_men_n632_), .B(men_men_n29_), .C(m), .Y(men_men_n633_));
  NAi32      u0605(.An(n), .Bn(f), .C(m), .Y(men_men_n634_));
  NA3        u0606(.A(men_men_n634_), .B(men_men_n633_), .C(men_men_n631_), .Y(men_men_n635_));
  NOi32      u0607(.An(e), .Bn(a), .C(d), .Y(men_men_n636_));
  AOI210     u0608(.A0(men_men_n29_), .A1(d), .B0(men_men_n636_), .Y(men_men_n637_));
  AOI210     u0609(.A0(men_men_n637_), .A1(men_men_n222_), .B0(men_men_n574_), .Y(men_men_n638_));
  AOI210     u0610(.A0(men_men_n638_), .A1(men_men_n635_), .B0(men_men_n629_), .Y(men_men_n639_));
  OAI210     u0611(.A0(men_men_n260_), .A1(men_men_n87_), .B0(men_men_n639_), .Y(men_men_n640_));
  AOI210     u0612(.A0(men_men_n624_), .A1(men_men_n610_), .B0(men_men_n640_), .Y(men_men_n641_));
  NA3        u0613(.A(men_men_n531_), .B(men_men_n178_), .C(men_men_n177_), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n481_), .B(men_men_n240_), .Y(men_men_n643_));
  NA2        u0615(.A(men_men_n74_), .B(men_men_n115_), .Y(men_men_n644_));
  NO2        u0616(.A(men_men_n644_), .B(men_men_n45_), .Y(men_men_n645_));
  NA2        u0617(.A(men_men_n645_), .B(men_men_n561_), .Y(men_men_n646_));
  NO2        u0618(.A(men_men_n646_), .B(men_men_n87_), .Y(men_men_n647_));
  NA3        u0619(.A(men_men_n576_), .B(men_men_n352_), .C(men_men_n46_), .Y(men_men_n648_));
  NOi32      u0620(.An(e), .Bn(c), .C(f), .Y(men_men_n649_));
  NOi21      u0621(.An(f), .B(g), .Y(men_men_n650_));
  NO2        u0622(.A(men_men_n650_), .B(men_men_n220_), .Y(men_men_n651_));
  AOI220     u0623(.A0(men_men_n651_), .A1(men_men_n408_), .B0(men_men_n649_), .B1(men_men_n182_), .Y(men_men_n652_));
  NA3        u0624(.A(men_men_n652_), .B(men_men_n648_), .C(men_men_n185_), .Y(men_men_n653_));
  AOI210     u0625(.A0(men_men_n560_), .A1(men_men_n412_), .B0(men_men_n310_), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n654_), .B(men_men_n276_), .Y(men_men_n655_));
  NOi21      u0627(.An(j), .B(l), .Y(men_men_n656_));
  NAi21      u0628(.An(k), .B(h), .Y(men_men_n657_));
  NO2        u0629(.A(men_men_n657_), .B(men_men_n274_), .Y(men_men_n658_));
  NA2        u0630(.A(men_men_n658_), .B(men_men_n656_), .Y(men_men_n659_));
  OR2        u0631(.A(men_men_n659_), .B(men_men_n615_), .Y(men_men_n660_));
  NOi31      u0632(.An(m), .B(n), .C(k), .Y(men_men_n661_));
  NA2        u0633(.A(men_men_n656_), .B(men_men_n661_), .Y(men_men_n662_));
  AOI210     u0634(.A0(men_men_n412_), .A1(men_men_n386_), .B0(men_men_n310_), .Y(men_men_n663_));
  NAi21      u0635(.An(men_men_n662_), .B(men_men_n663_), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n289_), .B(men_men_n49_), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n321_), .B(men_men_n625_), .Y(men_men_n666_));
  NO2        u0638(.A(men_men_n556_), .B(men_men_n49_), .Y(men_men_n667_));
  AOI220     u0639(.A0(men_men_n667_), .A1(men_men_n666_), .B0(men_men_n665_), .B1(men_men_n596_), .Y(men_men_n668_));
  NA4        u0640(.A(men_men_n668_), .B(men_men_n664_), .C(men_men_n660_), .D(men_men_n655_), .Y(men_men_n669_));
  NA2        u0641(.A(men_men_n110_), .B(men_men_n36_), .Y(men_men_n670_));
  NO2        u0642(.A(k), .B(men_men_n223_), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n552_), .B(men_men_n375_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n672_), .B(n), .Y(men_men_n673_));
  NAi31      u0645(.An(men_men_n670_), .B(men_men_n673_), .C(men_men_n671_), .Y(men_men_n674_));
  NO2        u0646(.A(men_men_n554_), .B(men_men_n183_), .Y(men_men_n675_));
  NA3        u0647(.A(men_men_n577_), .B(men_men_n283_), .C(men_men_n148_), .Y(men_men_n676_));
  NA2        u0648(.A(men_men_n527_), .B(men_men_n164_), .Y(men_men_n677_));
  NO3        u0649(.A(men_men_n409_), .B(men_men_n677_), .C(men_men_n87_), .Y(men_men_n678_));
  AOI210     u0650(.A0(men_men_n676_), .A1(men_men_n675_), .B0(men_men_n678_), .Y(men_men_n679_));
  AN3        u0651(.A(f), .B(d), .C(b), .Y(men_men_n680_));
  OAI210     u0652(.A0(men_men_n680_), .A1(men_men_n132_), .B0(n), .Y(men_men_n681_));
  NA3        u0653(.A(men_men_n527_), .B(men_men_n164_), .C(men_men_n223_), .Y(men_men_n682_));
  AOI210     u0654(.A0(men_men_n681_), .A1(men_men_n242_), .B0(men_men_n682_), .Y(men_men_n683_));
  NAi31      u0655(.An(m), .B(n), .C(k), .Y(men_men_n684_));
  OR2        u0656(.A(men_men_n137_), .B(men_men_n61_), .Y(men_men_n685_));
  OAI210     u0657(.A0(men_men_n685_), .A1(men_men_n684_), .B0(men_men_n262_), .Y(men_men_n686_));
  OAI210     u0658(.A0(men_men_n686_), .A1(men_men_n683_), .B0(j), .Y(men_men_n687_));
  NA3        u0659(.A(men_men_n687_), .B(men_men_n679_), .C(men_men_n674_), .Y(men_men_n688_));
  NO4        u0660(.A(men_men_n688_), .B(men_men_n669_), .C(men_men_n653_), .D(men_men_n647_), .Y(men_men_n689_));
  NA2        u0661(.A(men_men_n396_), .B(men_men_n167_), .Y(men_men_n690_));
  NAi31      u0662(.An(g), .B(h), .C(f), .Y(men_men_n691_));
  OR3        u0663(.A(men_men_n691_), .B(men_men_n289_), .C(n), .Y(men_men_n692_));
  OA210      u0664(.A0(men_men_n556_), .A1(n), .B0(men_men_n613_), .Y(men_men_n693_));
  NA3        u0665(.A(men_men_n432_), .B(men_men_n123_), .C(men_men_n84_), .Y(men_men_n694_));
  OAI210     u0666(.A0(men_men_n693_), .A1(men_men_n91_), .B0(men_men_n694_), .Y(men_men_n695_));
  NOi21      u0667(.An(men_men_n692_), .B(men_men_n695_), .Y(men_men_n696_));
  AOI210     u0668(.A0(men_men_n696_), .A1(men_men_n690_), .B0(men_men_n549_), .Y(men_men_n697_));
  NAi21      u0669(.An(h), .B(j), .Y(men_men_n698_));
  OR2        u0670(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n699_));
  NA2        u0671(.A(men_men_n627_), .B(men_men_n354_), .Y(men_men_n700_));
  OA220      u0672(.A0(men_men_n662_), .A1(men_men_n700_), .B0(men_men_n659_), .B1(men_men_n699_), .Y(men_men_n701_));
  NA3        u0673(.A(men_men_n546_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n702_));
  NA2        u0674(.A(h), .B(men_men_n37_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n100_), .B(men_men_n46_), .Y(men_men_n704_));
  OAI220     u0676(.A0(men_men_n704_), .A1(men_men_n343_), .B0(men_men_n703_), .B1(men_men_n486_), .Y(men_men_n705_));
  AOI210     u0677(.A0(men_men_n593_), .A1(men_men_n444_), .B0(men_men_n49_), .Y(men_men_n706_));
  OAI220     u0678(.A0(men_men_n616_), .A1(men_men_n609_), .B0(men_men_n337_), .B1(men_men_n547_), .Y(men_men_n707_));
  AOI210     u0679(.A0(men_men_n707_), .A1(men_men_n706_), .B0(men_men_n705_), .Y(men_men_n708_));
  NA3        u0680(.A(men_men_n708_), .B(men_men_n702_), .C(men_men_n701_), .Y(men_men_n709_));
  NO2        u0681(.A(men_men_n264_), .B(f), .Y(men_men_n710_));
  NA2        u0682(.A(men_men_n340_), .B(men_men_n143_), .Y(men_men_n711_));
  NA2        u0683(.A(men_men_n134_), .B(men_men_n49_), .Y(men_men_n712_));
  AOI220     u0684(.A0(men_men_n712_), .A1(men_men_n552_), .B0(men_men_n375_), .B1(men_men_n115_), .Y(men_men_n713_));
  OA220      u0685(.A0(men_men_n713_), .A1(men_men_n574_), .B0(men_men_n373_), .B1(men_men_n113_), .Y(men_men_n714_));
  OAI210     u0686(.A0(men_men_n711_), .A1(men_men_n264_), .B0(men_men_n714_), .Y(men_men_n715_));
  NO3        u0687(.A(men_men_n419_), .B(men_men_n200_), .C(men_men_n199_), .Y(men_men_n716_));
  NA2        u0688(.A(men_men_n716_), .B(men_men_n240_), .Y(men_men_n717_));
  NA3        u0689(.A(men_men_n717_), .B(men_men_n266_), .C(j), .Y(men_men_n718_));
  NO3        u0690(.A(men_men_n481_), .B(men_men_n180_), .C(i), .Y(men_men_n719_));
  NA2        u0691(.A(men_men_n485_), .B(men_men_n84_), .Y(men_men_n720_));
  NO4        u0692(.A(men_men_n549_), .B(men_men_n720_), .C(men_men_n133_), .D(men_men_n222_), .Y(men_men_n721_));
  INV        u0693(.A(men_men_n721_), .Y(men_men_n722_));
  NA4        u0694(.A(men_men_n722_), .B(men_men_n718_), .C(men_men_n534_), .D(men_men_n417_), .Y(men_men_n723_));
  NO4        u0695(.A(men_men_n723_), .B(men_men_n715_), .C(men_men_n709_), .D(men_men_n697_), .Y(men_men_n724_));
  NA4        u0696(.A(men_men_n724_), .B(men_men_n689_), .C(men_men_n641_), .D(men_men_n607_), .Y(men08));
  NO2        u0697(.A(k), .B(h), .Y(men_men_n726_));
  AO210      u0698(.A0(men_men_n264_), .A1(men_men_n469_), .B0(men_men_n726_), .Y(men_men_n727_));
  NO2        u0699(.A(men_men_n727_), .B(men_men_n308_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n649_), .B(men_men_n84_), .Y(men_men_n729_));
  INV        u0701(.A(men_men_n729_), .Y(men_men_n730_));
  AOI210     u0702(.A0(men_men_n730_), .A1(men_men_n728_), .B0(men_men_n512_), .Y(men_men_n731_));
  NA2        u0703(.A(men_men_n84_), .B(men_men_n112_), .Y(men_men_n732_));
  NO2        u0704(.A(men_men_n732_), .B(men_men_n57_), .Y(men_men_n733_));
  NO4        u0705(.A(men_men_n393_), .B(men_men_n114_), .C(j), .D(men_men_n223_), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n603_), .B(men_men_n242_), .Y(men_men_n735_));
  AOI220     u0707(.A0(men_men_n735_), .A1(men_men_n360_), .B0(men_men_n734_), .B1(men_men_n733_), .Y(men_men_n736_));
  AOI210     u0708(.A0(men_men_n603_), .A1(men_men_n160_), .B0(men_men_n84_), .Y(men_men_n737_));
  NA4        u0709(.A(men_men_n225_), .B(men_men_n143_), .C(men_men_n45_), .D(h), .Y(men_men_n738_));
  AN2        u0710(.A(l), .B(k), .Y(men_men_n739_));
  NA4        u0711(.A(men_men_n739_), .B(men_men_n110_), .C(men_men_n73_), .D(men_men_n223_), .Y(men_men_n740_));
  OAI210     u0712(.A0(men_men_n738_), .A1(g), .B0(men_men_n740_), .Y(men_men_n741_));
  NA2        u0713(.A(men_men_n741_), .B(men_men_n737_), .Y(men_men_n742_));
  NA4        u0714(.A(men_men_n742_), .B(men_men_n736_), .C(men_men_n731_), .D(men_men_n362_), .Y(men_men_n743_));
  AN2        u0715(.A(men_men_n557_), .B(men_men_n96_), .Y(men_men_n744_));
  NO4        u0716(.A(men_men_n180_), .B(men_men_n407_), .C(men_men_n114_), .D(g), .Y(men_men_n745_));
  AOI210     u0717(.A0(men_men_n745_), .A1(men_men_n735_), .B0(men_men_n541_), .Y(men_men_n746_));
  NO2        u0718(.A(men_men_n38_), .B(men_men_n222_), .Y(men_men_n747_));
  AOI220     u0719(.A0(men_men_n651_), .A1(men_men_n359_), .B0(men_men_n747_), .B1(men_men_n590_), .Y(men_men_n748_));
  NAi31      u0720(.An(men_men_n744_), .B(men_men_n748_), .C(men_men_n746_), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n560_), .B(men_men_n35_), .Y(men_men_n750_));
  OAI210     u0722(.A0(men_men_n577_), .A1(men_men_n47_), .B0(men_men_n685_), .Y(men_men_n751_));
  NO2        u0723(.A(men_men_n507_), .B(men_men_n134_), .Y(men_men_n752_));
  AOI210     u0724(.A0(men_men_n752_), .A1(men_men_n751_), .B0(men_men_n750_), .Y(men_men_n753_));
  NO3        u0725(.A(men_men_n327_), .B(men_men_n133_), .C(men_men_n41_), .Y(men_men_n754_));
  NAi21      u0726(.An(men_men_n754_), .B(men_men_n740_), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n727_), .B(men_men_n138_), .Y(men_men_n756_));
  AOI220     u0728(.A0(men_men_n756_), .A1(men_men_n418_), .B0(men_men_n755_), .B1(men_men_n76_), .Y(men_men_n757_));
  OAI210     u0729(.A0(men_men_n753_), .A1(men_men_n87_), .B0(men_men_n757_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n375_), .B(men_men_n43_), .Y(men_men_n759_));
  NA3        u0731(.A(men_men_n717_), .B(men_men_n345_), .C(men_men_n399_), .Y(men_men_n760_));
  NA2        u0732(.A(men_men_n739_), .B(men_men_n230_), .Y(men_men_n761_));
  NO2        u0733(.A(men_men_n761_), .B(men_men_n339_), .Y(men_men_n762_));
  AOI210     u0734(.A0(men_men_n762_), .A1(men_men_n710_), .B0(men_men_n511_), .Y(men_men_n763_));
  NA3        u0735(.A(m), .B(l), .C(k), .Y(men_men_n764_));
  AOI210     u0736(.A0(men_men_n694_), .A1(men_men_n692_), .B0(men_men_n764_), .Y(men_men_n765_));
  NO2        u0737(.A(men_men_n559_), .B(men_men_n284_), .Y(men_men_n766_));
  NOi21      u0738(.An(men_men_n766_), .B(men_men_n553_), .Y(men_men_n767_));
  NA4        u0739(.A(men_men_n115_), .B(l), .C(k), .D(men_men_n87_), .Y(men_men_n768_));
  NA3        u0740(.A(men_men_n123_), .B(men_men_n427_), .C(i), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n769_), .B(men_men_n768_), .Y(men_men_n770_));
  NO3        u0742(.A(men_men_n770_), .B(men_men_n767_), .C(men_men_n765_), .Y(men_men_n771_));
  NA4        u0743(.A(men_men_n771_), .B(men_men_n763_), .C(men_men_n760_), .D(men_men_n759_), .Y(men_men_n772_));
  NO4        u0744(.A(men_men_n772_), .B(men_men_n758_), .C(men_men_n749_), .D(men_men_n743_), .Y(men_men_n773_));
  NA2        u0745(.A(men_men_n651_), .B(men_men_n408_), .Y(men_men_n774_));
  NOi31      u0746(.An(g), .B(h), .C(f), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n667_), .B(men_men_n775_), .Y(men_men_n776_));
  AO210      u0748(.A0(men_men_n776_), .A1(men_men_n617_), .B0(men_men_n562_), .Y(men_men_n777_));
  NO3        u0749(.A(men_men_n412_), .B(men_men_n547_), .C(h), .Y(men_men_n778_));
  AOI210     u0750(.A0(men_men_n778_), .A1(men_men_n115_), .B0(men_men_n520_), .Y(men_men_n779_));
  NA4        u0751(.A(men_men_n779_), .B(men_men_n777_), .C(men_men_n774_), .D(men_men_n263_), .Y(men_men_n780_));
  NA2        u0752(.A(men_men_n739_), .B(men_men_n73_), .Y(men_men_n781_));
  NOi21      u0753(.An(h), .B(j), .Y(men_men_n782_));
  NA2        u0754(.A(men_men_n782_), .B(f), .Y(men_men_n783_));
  NO2        u0755(.A(men_men_n783_), .B(men_men_n257_), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n784_), .B(men_men_n719_), .Y(men_men_n785_));
  OAI220     u0757(.A0(men_men_n785_), .A1(men_men_n781_), .B0(men_men_n619_), .B1(men_men_n62_), .Y(men_men_n786_));
  AOI210     u0758(.A0(men_men_n780_), .A1(l), .B0(men_men_n786_), .Y(men_men_n787_));
  NO2        u0759(.A(j), .B(i), .Y(men_men_n788_));
  NA3        u0760(.A(men_men_n788_), .B(men_men_n80_), .C(l), .Y(men_men_n789_));
  NA2        u0761(.A(men_men_n788_), .B(men_men_n33_), .Y(men_men_n790_));
  NA2        u0762(.A(men_men_n437_), .B(men_men_n123_), .Y(men_men_n791_));
  OA220      u0763(.A0(men_men_n791_), .A1(men_men_n790_), .B0(men_men_n789_), .B1(men_men_n615_), .Y(men_men_n792_));
  NO3        u0764(.A(men_men_n155_), .B(men_men_n49_), .C(men_men_n112_), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n566_), .B(men_men_n153_), .C(men_men_n73_), .Y(men_men_n794_));
  NO3        u0766(.A(men_men_n507_), .B(men_men_n456_), .C(j), .Y(men_men_n795_));
  OAI210     u0767(.A0(men_men_n794_), .A1(men_men_n793_), .B0(men_men_n795_), .Y(men_men_n796_));
  OAI210     u0768(.A0(men_men_n776_), .A1(men_men_n62_), .B0(men_men_n796_), .Y(men_men_n797_));
  NA2        u0769(.A(k), .B(j), .Y(men_men_n798_));
  NO3        u0770(.A(men_men_n308_), .B(men_men_n798_), .C(men_men_n40_), .Y(men_men_n799_));
  AOI210     u0771(.A0(men_men_n552_), .A1(n), .B0(men_men_n576_), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n800_), .B(men_men_n579_), .Y(men_men_n801_));
  AN3        u0773(.A(men_men_n801_), .B(men_men_n799_), .C(men_men_n99_), .Y(men_men_n802_));
  NO3        u0774(.A(men_men_n180_), .B(men_men_n407_), .C(men_men_n114_), .Y(men_men_n803_));
  AOI220     u0775(.A0(men_men_n803_), .A1(men_men_n258_), .B0(men_men_n643_), .B1(men_men_n318_), .Y(men_men_n804_));
  NAi31      u0776(.An(men_men_n637_), .B(men_men_n93_), .C(men_men_n84_), .Y(men_men_n805_));
  NA2        u0777(.A(men_men_n805_), .B(men_men_n804_), .Y(men_men_n806_));
  NO2        u0778(.A(men_men_n308_), .B(men_men_n138_), .Y(men_men_n807_));
  AOI220     u0779(.A0(men_men_n807_), .A1(men_men_n651_), .B0(men_men_n754_), .B1(men_men_n737_), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n764_), .B(men_men_n91_), .Y(men_men_n809_));
  NA2        u0781(.A(men_men_n809_), .B(men_men_n614_), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n616_), .B(men_men_n119_), .Y(men_men_n811_));
  OAI210     u0783(.A0(men_men_n811_), .A1(men_men_n795_), .B0(men_men_n706_), .Y(men_men_n812_));
  NA3        u0784(.A(men_men_n812_), .B(men_men_n810_), .C(men_men_n808_), .Y(men_men_n813_));
  OR4        u0785(.A(men_men_n813_), .B(men_men_n806_), .C(men_men_n802_), .D(men_men_n797_), .Y(men_men_n814_));
  NA3        u0786(.A(men_men_n800_), .B(men_men_n579_), .C(men_men_n578_), .Y(men_men_n815_));
  NA4        u0787(.A(men_men_n815_), .B(men_men_n225_), .C(men_men_n469_), .D(men_men_n34_), .Y(men_men_n816_));
  NO4        u0788(.A(men_men_n507_), .B(men_men_n451_), .C(j), .D(f), .Y(men_men_n817_));
  NA2        u0789(.A(men_men_n817_), .B(men_men_n269_), .Y(men_men_n818_));
  NA3        u0790(.A(men_men_n569_), .B(men_men_n301_), .C(h), .Y(men_men_n819_));
  NOi21      u0791(.An(men_men_n706_), .B(men_men_n819_), .Y(men_men_n820_));
  NO2        u0792(.A(men_men_n92_), .B(men_men_n47_), .Y(men_men_n821_));
  OAI220     u0793(.A0(men_men_n819_), .A1(men_men_n633_), .B0(men_men_n789_), .B1(men_men_n699_), .Y(men_men_n822_));
  AOI210     u0794(.A0(men_men_n821_), .A1(men_men_n673_), .B0(men_men_n822_), .Y(men_men_n823_));
  NAi41      u0795(.An(men_men_n820_), .B(men_men_n823_), .C(men_men_n818_), .D(men_men_n816_), .Y(men_men_n824_));
  OR2        u0796(.A(men_men_n809_), .B(men_men_n96_), .Y(men_men_n825_));
  AOI220     u0797(.A0(men_men_n825_), .A1(men_men_n248_), .B0(men_men_n795_), .B1(men_men_n665_), .Y(men_men_n826_));
  NO2        u0798(.A(men_men_n693_), .B(men_men_n73_), .Y(men_men_n827_));
  AOI210     u0799(.A0(men_men_n817_), .A1(men_men_n827_), .B0(men_men_n347_), .Y(men_men_n828_));
  OAI210     u0800(.A0(men_men_n764_), .A1(men_men_n691_), .B0(men_men_n540_), .Y(men_men_n829_));
  NA3        u0801(.A(men_men_n261_), .B(men_men_n59_), .C(b), .Y(men_men_n830_));
  AOI220     u0802(.A0(men_men_n632_), .A1(men_men_n29_), .B0(men_men_n485_), .B1(men_men_n84_), .Y(men_men_n831_));
  NA2        u0803(.A(men_men_n831_), .B(men_men_n830_), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n819_), .B(men_men_n510_), .Y(men_men_n833_));
  AOI210     u0805(.A0(men_men_n832_), .A1(men_men_n829_), .B0(men_men_n833_), .Y(men_men_n834_));
  NA3        u0806(.A(men_men_n834_), .B(men_men_n828_), .C(men_men_n826_), .Y(men_men_n835_));
  NOi41      u0807(.An(men_men_n792_), .B(men_men_n835_), .C(men_men_n824_), .D(men_men_n814_), .Y(men_men_n836_));
  OR3        u0808(.A(men_men_n738_), .B(men_men_n242_), .C(g), .Y(men_men_n837_));
  NO3        u0809(.A(men_men_n353_), .B(men_men_n310_), .C(men_men_n114_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n838_), .B(men_men_n801_), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n840_));
  NO3        u0812(.A(men_men_n840_), .B(men_men_n790_), .C(men_men_n289_), .Y(men_men_n841_));
  NO3        u0813(.A(men_men_n547_), .B(men_men_n94_), .C(h), .Y(men_men_n842_));
  AOI210     u0814(.A0(men_men_n842_), .A1(men_men_n733_), .B0(men_men_n841_), .Y(men_men_n843_));
  NA4        u0815(.A(men_men_n843_), .B(men_men_n839_), .C(men_men_n837_), .D(men_men_n420_), .Y(men_men_n844_));
  OR2        u0816(.A(men_men_n691_), .B(men_men_n92_), .Y(men_men_n845_));
  NOi31      u0817(.An(b), .B(d), .C(a), .Y(men_men_n846_));
  NO2        u0818(.A(men_men_n846_), .B(men_men_n630_), .Y(men_men_n847_));
  NO2        u0819(.A(men_men_n847_), .B(n), .Y(men_men_n848_));
  NOi21      u0820(.An(men_men_n831_), .B(men_men_n848_), .Y(men_men_n849_));
  OAI220     u0821(.A0(men_men_n849_), .A1(men_men_n845_), .B0(men_men_n819_), .B1(men_men_n631_), .Y(men_men_n850_));
  NO2        u0822(.A(men_men_n577_), .B(men_men_n84_), .Y(men_men_n851_));
  NO3        u0823(.A(men_men_n650_), .B(men_men_n339_), .C(men_men_n119_), .Y(men_men_n852_));
  NOi21      u0824(.An(men_men_n852_), .B(men_men_n165_), .Y(men_men_n853_));
  AOI210     u0825(.A0(men_men_n838_), .A1(men_men_n851_), .B0(men_men_n853_), .Y(men_men_n854_));
  OAI210     u0826(.A0(men_men_n738_), .A1(men_men_n409_), .B0(men_men_n854_), .Y(men_men_n855_));
  NO2        u0827(.A(men_men_n716_), .B(n), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n856_), .B(men_men_n728_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n334_), .B(men_men_n247_), .Y(men_men_n858_));
  OAI210     u0830(.A0(men_men_n96_), .A1(men_men_n93_), .B0(men_men_n858_), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n123_), .B(men_men_n84_), .Y(men_men_n860_));
  AOI210     u0832(.A0(men_men_n441_), .A1(men_men_n433_), .B0(men_men_n860_), .Y(men_men_n861_));
  NAi21      u0833(.An(men_men_n861_), .B(men_men_n859_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n762_), .B(men_men_n34_), .Y(men_men_n863_));
  NAi21      u0835(.An(men_men_n768_), .B(men_men_n452_), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n284_), .B(i), .Y(men_men_n865_));
  NA2        u0837(.A(men_men_n745_), .B(men_men_n361_), .Y(men_men_n866_));
  OAI210     u0838(.A0(men_men_n622_), .A1(men_men_n621_), .B0(men_men_n376_), .Y(men_men_n867_));
  AN3        u0839(.A(men_men_n867_), .B(men_men_n866_), .C(men_men_n864_), .Y(men_men_n868_));
  NAi41      u0840(.An(men_men_n862_), .B(men_men_n868_), .C(men_men_n863_), .D(men_men_n857_), .Y(men_men_n869_));
  NO4        u0841(.A(men_men_n869_), .B(men_men_n855_), .C(men_men_n850_), .D(men_men_n844_), .Y(men_men_n870_));
  NA4        u0842(.A(men_men_n870_), .B(men_men_n836_), .C(men_men_n787_), .D(men_men_n773_), .Y(men09));
  INV        u0843(.A(men_men_n124_), .Y(men_men_n872_));
  NA2        u0844(.A(f), .B(e), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n235_), .B(men_men_n114_), .Y(men_men_n874_));
  NA2        u0846(.A(men_men_n874_), .B(g), .Y(men_men_n875_));
  NA4        u0847(.A(men_men_n321_), .B(men_men_n494_), .C(men_men_n272_), .D(men_men_n121_), .Y(men_men_n876_));
  AOI210     u0848(.A0(men_men_n876_), .A1(g), .B0(men_men_n491_), .Y(men_men_n877_));
  AOI210     u0849(.A0(men_men_n877_), .A1(men_men_n875_), .B0(men_men_n873_), .Y(men_men_n878_));
  NA2        u0850(.A(men_men_n462_), .B(e), .Y(men_men_n879_));
  NO2        u0851(.A(men_men_n879_), .B(men_men_n531_), .Y(men_men_n880_));
  AOI210     u0852(.A0(men_men_n878_), .A1(men_men_n872_), .B0(men_men_n880_), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n212_), .B(men_men_n222_), .Y(men_men_n882_));
  NA3        u0854(.A(m), .B(l), .C(i), .Y(men_men_n883_));
  OAI220     u0855(.A0(men_men_n616_), .A1(men_men_n883_), .B0(men_men_n366_), .B1(men_men_n548_), .Y(men_men_n884_));
  NA4        u0856(.A(men_men_n88_), .B(men_men_n87_), .C(g), .D(f), .Y(men_men_n885_));
  NAi31      u0857(.An(men_men_n884_), .B(men_men_n885_), .C(men_men_n457_), .Y(men_men_n886_));
  OR2        u0858(.A(men_men_n886_), .B(men_men_n882_), .Y(men_men_n887_));
  NA3        u0859(.A(men_men_n845_), .B(men_men_n592_), .C(men_men_n540_), .Y(men_men_n888_));
  OA210      u0860(.A0(men_men_n888_), .A1(men_men_n887_), .B0(men_men_n848_), .Y(men_men_n889_));
  INV        u0861(.A(men_men_n350_), .Y(men_men_n890_));
  NOi31      u0862(.An(k), .B(m), .C(l), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n352_), .B(men_men_n891_), .Y(men_men_n892_));
  NO2        u0864(.A(men_men_n892_), .B(men_men_n625_), .Y(men_men_n893_));
  NA2        u0865(.A(men_men_n830_), .B(men_men_n343_), .Y(men_men_n894_));
  NA2        u0866(.A(men_men_n354_), .B(men_men_n356_), .Y(men_men_n895_));
  OAI210     u0867(.A0(men_men_n212_), .A1(men_men_n222_), .B0(men_men_n895_), .Y(men_men_n896_));
  AOI220     u0868(.A0(men_men_n896_), .A1(men_men_n894_), .B0(men_men_n893_), .B1(men_men_n890_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n174_), .B(men_men_n116_), .Y(men_men_n898_));
  NA3        u0870(.A(men_men_n898_), .B(men_men_n727_), .C(men_men_n138_), .Y(men_men_n899_));
  NA3        u0871(.A(men_men_n899_), .B(men_men_n197_), .C(men_men_n31_), .Y(men_men_n900_));
  NA4        u0872(.A(men_men_n900_), .B(men_men_n897_), .C(men_men_n652_), .D(men_men_n82_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n612_), .B(men_men_n517_), .Y(men_men_n902_));
  NA2        u0874(.A(men_men_n902_), .B(men_men_n197_), .Y(men_men_n903_));
  NOi21      u0875(.An(f), .B(d), .Y(men_men_n904_));
  NA2        u0876(.A(men_men_n904_), .B(m), .Y(men_men_n905_));
  NO2        u0877(.A(men_men_n905_), .B(men_men_n52_), .Y(men_men_n906_));
  NOi32      u0878(.An(g), .Bn(f), .C(d), .Y(men_men_n907_));
  NA4        u0879(.A(men_men_n907_), .B(men_men_n632_), .C(men_men_n29_), .D(m), .Y(men_men_n908_));
  NOi21      u0880(.An(men_men_n322_), .B(men_men_n908_), .Y(men_men_n909_));
  AOI210     u0881(.A0(men_men_n906_), .A1(men_men_n567_), .B0(men_men_n909_), .Y(men_men_n910_));
  NA3        u0882(.A(men_men_n321_), .B(men_men_n272_), .C(men_men_n121_), .Y(men_men_n911_));
  AN2        u0883(.A(f), .B(d), .Y(men_men_n912_));
  NA3        u0884(.A(men_men_n499_), .B(men_men_n912_), .C(men_men_n84_), .Y(men_men_n913_));
  NO3        u0885(.A(men_men_n913_), .B(men_men_n73_), .C(men_men_n223_), .Y(men_men_n914_));
  INV        u0886(.A(men_men_n296_), .Y(men_men_n915_));
  NA2        u0887(.A(men_men_n911_), .B(men_men_n914_), .Y(men_men_n916_));
  NAi41      u0888(.An(men_men_n509_), .B(men_men_n916_), .C(men_men_n910_), .D(men_men_n903_), .Y(men_men_n917_));
  NO4        u0889(.A(men_men_n650_), .B(men_men_n134_), .C(men_men_n339_), .D(men_men_n156_), .Y(men_men_n918_));
  NO2        u0890(.A(men_men_n684_), .B(men_men_n339_), .Y(men_men_n919_));
  AN2        u0891(.A(men_men_n919_), .B(men_men_n710_), .Y(men_men_n920_));
  NO3        u0892(.A(men_men_n920_), .B(men_men_n918_), .C(men_men_n244_), .Y(men_men_n921_));
  NA2        u0893(.A(men_men_n630_), .B(men_men_n84_), .Y(men_men_n922_));
  NO2        u0894(.A(men_men_n895_), .B(men_men_n922_), .Y(men_men_n923_));
  NA3        u0895(.A(men_men_n164_), .B(men_men_n110_), .C(men_men_n109_), .Y(men_men_n924_));
  OAI220     u0896(.A0(men_men_n913_), .A1(men_men_n446_), .B0(men_men_n350_), .B1(men_men_n924_), .Y(men_men_n925_));
  NOi31      u0897(.An(men_men_n233_), .B(men_men_n925_), .C(men_men_n923_), .Y(men_men_n926_));
  NA2        u0898(.A(c), .B(men_men_n118_), .Y(men_men_n927_));
  NO2        u0899(.A(men_men_n927_), .B(men_men_n424_), .Y(men_men_n928_));
  NA3        u0900(.A(men_men_n928_), .B(men_men_n529_), .C(f), .Y(men_men_n929_));
  OR2        u0901(.A(men_men_n691_), .B(men_men_n563_), .Y(men_men_n930_));
  INV        u0902(.A(men_men_n930_), .Y(men_men_n931_));
  NA2        u0903(.A(men_men_n847_), .B(men_men_n113_), .Y(men_men_n932_));
  NA2        u0904(.A(men_men_n932_), .B(men_men_n931_), .Y(men_men_n933_));
  NA4        u0905(.A(men_men_n933_), .B(men_men_n929_), .C(men_men_n926_), .D(men_men_n921_), .Y(men_men_n934_));
  NO4        u0906(.A(men_men_n934_), .B(men_men_n917_), .C(men_men_n901_), .D(men_men_n889_), .Y(men_men_n935_));
  OR2        u0907(.A(men_men_n913_), .B(men_men_n73_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n874_), .B(g), .Y(men_men_n937_));
  AOI210     u0909(.A0(men_men_n937_), .A1(men_men_n302_), .B0(men_men_n936_), .Y(men_men_n938_));
  NO2        u0910(.A(men_men_n343_), .B(men_men_n885_), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n940_));
  NO2        u0912(.A(men_men_n240_), .B(men_men_n234_), .Y(men_men_n941_));
  AOI220     u0913(.A0(men_men_n941_), .A1(men_men_n237_), .B0(men_men_n315_), .B1(men_men_n940_), .Y(men_men_n942_));
  NO2        u0914(.A(men_men_n446_), .B(men_men_n873_), .Y(men_men_n943_));
  NA2        u0915(.A(men_men_n943_), .B(men_men_n584_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n944_), .B(men_men_n942_), .Y(men_men_n945_));
  NA2        u0917(.A(e), .B(d), .Y(men_men_n946_));
  OAI220     u0918(.A0(men_men_n946_), .A1(c), .B0(men_men_n334_), .B1(d), .Y(men_men_n947_));
  NA3        u0919(.A(men_men_n947_), .B(men_men_n474_), .C(men_men_n527_), .Y(men_men_n948_));
  AOI210     u0920(.A0(men_men_n535_), .A1(men_men_n187_), .B0(men_men_n240_), .Y(men_men_n949_));
  AOI210     u0921(.A0(men_men_n651_), .A1(men_men_n359_), .B0(men_men_n949_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n296_), .B(men_men_n170_), .Y(men_men_n951_));
  NA2        u0923(.A(men_men_n914_), .B(men_men_n951_), .Y(men_men_n952_));
  NA3        u0924(.A(men_men_n952_), .B(men_men_n950_), .C(men_men_n948_), .Y(men_men_n953_));
  NO4        u0925(.A(men_men_n953_), .B(men_men_n945_), .C(men_men_n939_), .D(men_men_n938_), .Y(men_men_n954_));
  NA2        u0926(.A(men_men_n890_), .B(men_men_n31_), .Y(men_men_n955_));
  AO210      u0927(.A0(men_men_n955_), .A1(men_men_n729_), .B0(men_men_n226_), .Y(men_men_n956_));
  NO2        u0928(.A(men_men_n310_), .B(j), .Y(men_men_n957_));
  NA2        u0929(.A(men_men_n957_), .B(men_men_n919_), .Y(men_men_n958_));
  OAI210     u0930(.A0(men_men_n879_), .A1(men_men_n177_), .B0(men_men_n958_), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n874_), .A1(men_men_n951_), .B0(men_men_n907_), .Y(men_men_n960_));
  NO2        u0932(.A(men_men_n960_), .B(men_men_n633_), .Y(men_men_n961_));
  AOI210     u0933(.A0(men_men_n120_), .A1(men_men_n119_), .B0(men_men_n271_), .Y(men_men_n962_));
  NO2        u0934(.A(men_men_n962_), .B(men_men_n908_), .Y(men_men_n963_));
  AO210      u0935(.A0(men_men_n894_), .A1(men_men_n884_), .B0(men_men_n963_), .Y(men_men_n964_));
  NOi31      u0936(.An(men_men_n567_), .B(men_men_n905_), .C(men_men_n302_), .Y(men_men_n965_));
  NO4        u0937(.A(men_men_n965_), .B(men_men_n964_), .C(men_men_n961_), .D(men_men_n959_), .Y(men_men_n966_));
  AN2        u0938(.A(men_men_n182_), .B(f), .Y(men_men_n967_));
  OAI210     u0939(.A0(men_men_n967_), .A1(men_men_n477_), .B0(men_men_n947_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n456_), .B(men_men_n69_), .Y(men_men_n969_));
  OAI210     u0941(.A0(men_men_n888_), .A1(men_men_n969_), .B0(men_men_n733_), .Y(men_men_n970_));
  AN4        u0942(.A(men_men_n970_), .B(men_men_n968_), .C(men_men_n966_), .D(men_men_n956_), .Y(men_men_n971_));
  NA4        u0943(.A(men_men_n971_), .B(men_men_n954_), .C(men_men_n935_), .D(men_men_n881_), .Y(men12));
  NO2        u0944(.A(men_men_n472_), .B(c), .Y(men_men_n973_));
  NO4        u0945(.A(men_men_n461_), .B(men_men_n264_), .C(men_men_n608_), .D(men_men_n223_), .Y(men_men_n974_));
  NA2        u0946(.A(men_men_n974_), .B(men_men_n973_), .Y(men_men_n975_));
  NA2        u0947(.A(men_men_n567_), .B(men_men_n969_), .Y(men_men_n976_));
  NO2        u0948(.A(men_men_n472_), .B(men_men_n118_), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n691_), .B(men_men_n393_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n978_), .B(men_men_n565_), .Y(men_men_n979_));
  NA4        u0951(.A(men_men_n979_), .B(men_men_n976_), .C(men_men_n975_), .D(men_men_n460_), .Y(men_men_n980_));
  AOI210     u0952(.A0(men_men_n243_), .A1(men_men_n349_), .B0(men_men_n209_), .Y(men_men_n981_));
  BUFFER     u0953(.A(men_men_n974_), .Y(men_men_n982_));
  AOI210     u0954(.A0(men_men_n346_), .A1(men_men_n405_), .B0(men_men_n223_), .Y(men_men_n983_));
  OAI210     u0955(.A0(men_men_n983_), .A1(men_men_n982_), .B0(men_men_n419_), .Y(men_men_n984_));
  NO2        u0956(.A(men_men_n670_), .B(men_men_n274_), .Y(men_men_n985_));
  NO2        u0957(.A(men_men_n616_), .B(men_men_n883_), .Y(men_men_n986_));
  AOI220     u0958(.A0(men_men_n986_), .A1(men_men_n590_), .B0(men_men_n858_), .B1(men_men_n985_), .Y(men_men_n987_));
  NO2        u0959(.A(men_men_n155_), .B(men_men_n247_), .Y(men_men_n988_));
  NA3        u0960(.A(men_men_n988_), .B(men_men_n250_), .C(i), .Y(men_men_n989_));
  NA3        u0961(.A(men_men_n989_), .B(men_men_n987_), .C(men_men_n984_), .Y(men_men_n990_));
  OR2        u0962(.A(men_men_n335_), .B(men_men_n977_), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n991_), .B(men_men_n367_), .Y(men_men_n992_));
  NO3        u0964(.A(men_men_n134_), .B(men_men_n156_), .C(men_men_n223_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n993_), .B(men_men_n552_), .Y(men_men_n994_));
  NA4        u0966(.A(men_men_n462_), .B(men_men_n454_), .C(men_men_n188_), .D(g), .Y(men_men_n995_));
  NA3        u0967(.A(men_men_n995_), .B(men_men_n994_), .C(men_men_n992_), .Y(men_men_n996_));
  NO3        u0968(.A(men_men_n696_), .B(men_men_n92_), .C(men_men_n45_), .Y(men_men_n997_));
  NO4        u0969(.A(men_men_n997_), .B(men_men_n996_), .C(men_men_n990_), .D(men_men_n980_), .Y(men_men_n998_));
  NO2        u0970(.A(men_men_n383_), .B(men_men_n382_), .Y(men_men_n999_));
  NA2        u0971(.A(men_men_n613_), .B(men_men_n71_), .Y(men_men_n1000_));
  NOi21      u0972(.An(men_men_n34_), .B(men_men_n684_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n1000_), .B(men_men_n999_), .Y(men_men_n1002_));
  OAI210     u0974(.A0(men_men_n262_), .A1(men_men_n45_), .B0(men_men_n1002_), .Y(men_men_n1003_));
  NA2        u0975(.A(men_men_n452_), .B(men_men_n276_), .Y(men_men_n1004_));
  NO3        u0976(.A(men_men_n860_), .B(men_men_n89_), .C(men_men_n424_), .Y(men_men_n1005_));
  NAi31      u0977(.An(men_men_n1005_), .B(men_men_n1004_), .C(men_men_n331_), .Y(men_men_n1006_));
  NO2        u0978(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1007_));
  NO2        u0979(.A(men_men_n523_), .B(men_men_n310_), .Y(men_men_n1008_));
  INV        u0980(.A(men_men_n661_), .Y(men_men_n1009_));
  OAI210     u0981(.A0(men_men_n769_), .A1(men_men_n1009_), .B0(men_men_n380_), .Y(men_men_n1010_));
  NO3        u0982(.A(men_men_n1010_), .B(men_men_n1006_), .C(men_men_n1003_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n359_), .B(g), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n167_), .B(i), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n46_), .B(i), .Y(men_men_n1014_));
  OAI220     u0986(.A0(men_men_n1014_), .A1(men_men_n208_), .B0(men_men_n1013_), .B1(men_men_n92_), .Y(men_men_n1015_));
  AOI210     u0987(.A0(men_men_n435_), .A1(men_men_n37_), .B0(men_men_n1015_), .Y(men_men_n1016_));
  NO2        u0988(.A(men_men_n148_), .B(men_men_n84_), .Y(men_men_n1017_));
  OR2        u0989(.A(men_men_n1017_), .B(men_men_n576_), .Y(men_men_n1018_));
  INV        u0990(.A(men_men_n1018_), .Y(men_men_n1019_));
  OAI220     u0991(.A0(men_men_n1019_), .A1(men_men_n1012_), .B0(men_men_n1016_), .B1(men_men_n343_), .Y(men_men_n1020_));
  NO2        u0992(.A(men_men_n691_), .B(men_men_n517_), .Y(men_men_n1021_));
  NA3        u0993(.A(men_men_n354_), .B(men_men_n656_), .C(i), .Y(men_men_n1022_));
  OAI210     u0994(.A0(men_men_n456_), .A1(men_men_n321_), .B0(men_men_n1022_), .Y(men_men_n1023_));
  OAI220     u0995(.A0(men_men_n1023_), .A1(men_men_n1021_), .B0(men_men_n706_), .B1(men_men_n794_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n636_), .B(men_men_n115_), .Y(men_men_n1025_));
  OR3        u0997(.A(men_men_n321_), .B(men_men_n451_), .C(f), .Y(men_men_n1026_));
  NA3        u0998(.A(men_men_n656_), .B(men_men_n80_), .C(i), .Y(men_men_n1027_));
  OA220      u0999(.A0(men_men_n1027_), .A1(men_men_n1025_), .B0(men_men_n1026_), .B1(men_men_n615_), .Y(men_men_n1028_));
  NA2        u1000(.A(men_men_n720_), .B(men_men_n922_), .Y(men_men_n1029_));
  NA2        u1001(.A(men_men_n885_), .B(men_men_n457_), .Y(men_men_n1030_));
  NA2        u1002(.A(men_men_n231_), .B(men_men_n77_), .Y(men_men_n1031_));
  NA3        u1003(.A(men_men_n1031_), .B(men_men_n1027_), .C(men_men_n1026_), .Y(men_men_n1032_));
  AOI220     u1004(.A0(men_men_n1032_), .A1(men_men_n269_), .B0(men_men_n1030_), .B1(men_men_n1029_), .Y(men_men_n1033_));
  NA3        u1005(.A(men_men_n1033_), .B(men_men_n1028_), .C(men_men_n1024_), .Y(men_men_n1034_));
  NO2        u1006(.A(men_men_n393_), .B(men_men_n91_), .Y(men_men_n1035_));
  OAI210     u1007(.A0(men_men_n1035_), .A1(men_men_n985_), .B0(men_men_n248_), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n695_), .B(men_men_n88_), .Y(men_men_n1037_));
  NO2        u1009(.A(men_men_n480_), .B(men_men_n223_), .Y(men_men_n1038_));
  AOI220     u1010(.A0(men_men_n1038_), .A1(men_men_n398_), .B0(men_men_n991_), .B1(men_men_n227_), .Y(men_men_n1039_));
  AOI220     u1011(.A0(men_men_n978_), .A1(men_men_n988_), .B0(men_men_n614_), .B1(men_men_n90_), .Y(men_men_n1040_));
  NA4        u1012(.A(men_men_n1040_), .B(men_men_n1039_), .C(men_men_n1037_), .D(men_men_n1036_), .Y(men_men_n1041_));
  OAI210     u1013(.A0(men_men_n1030_), .A1(men_men_n986_), .B0(men_men_n565_), .Y(men_men_n1042_));
  AOI210     u1014(.A0(men_men_n436_), .A1(men_men_n428_), .B0(men_men_n860_), .Y(men_men_n1043_));
  OAI210     u1015(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n111_), .Y(men_men_n1044_));
  AOI210     u1016(.A0(men_men_n1044_), .A1(men_men_n557_), .B0(men_men_n1043_), .Y(men_men_n1045_));
  NO3        u1017(.A(l), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1046_));
  AOI220     u1018(.A0(men_men_n1046_), .A1(men_men_n654_), .B0(men_men_n675_), .B1(men_men_n552_), .Y(men_men_n1047_));
  NA3        u1019(.A(men_men_n1047_), .B(men_men_n1045_), .C(men_men_n1042_), .Y(men_men_n1048_));
  NO4        u1020(.A(men_men_n1048_), .B(men_men_n1041_), .C(men_men_n1034_), .D(men_men_n1020_), .Y(men_men_n1049_));
  NAi31      u1021(.An(men_men_n144_), .B(men_men_n437_), .C(n), .Y(men_men_n1050_));
  NO3        u1022(.A(men_men_n127_), .B(men_men_n352_), .C(men_men_n891_), .Y(men_men_n1051_));
  NO2        u1023(.A(men_men_n1051_), .B(men_men_n1050_), .Y(men_men_n1052_));
  NO3        u1024(.A(men_men_n284_), .B(men_men_n144_), .C(men_men_n424_), .Y(men_men_n1053_));
  AOI210     u1025(.A0(men_men_n1053_), .A1(men_men_n518_), .B0(men_men_n1052_), .Y(men_men_n1054_));
  NA2        u1026(.A(men_men_n512_), .B(i), .Y(men_men_n1055_));
  NA2        u1027(.A(men_men_n1055_), .B(men_men_n1054_), .Y(men_men_n1056_));
  NA2        u1028(.A(men_men_n240_), .B(men_men_n178_), .Y(men_men_n1057_));
  NO3        u1029(.A(men_men_n318_), .B(men_men_n462_), .C(men_men_n182_), .Y(men_men_n1058_));
  NOi31      u1030(.An(men_men_n1057_), .B(men_men_n1058_), .C(men_men_n223_), .Y(men_men_n1059_));
  NAi21      u1031(.An(men_men_n577_), .B(men_men_n1038_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n455_), .B(men_men_n922_), .Y(men_men_n1061_));
  NO2        u1033(.A(men_men_n456_), .B(men_men_n321_), .Y(men_men_n1062_));
  AOI220     u1034(.A0(men_men_n1062_), .A1(men_men_n1061_), .B0(men_men_n505_), .B1(g), .Y(men_men_n1063_));
  NA2        u1035(.A(men_men_n1063_), .B(men_men_n1060_), .Y(men_men_n1064_));
  OAI220     u1036(.A0(men_men_n1050_), .A1(men_men_n243_), .B0(men_men_n1022_), .B1(men_men_n631_), .Y(men_men_n1065_));
  NO2        u1037(.A(men_men_n692_), .B(men_men_n393_), .Y(men_men_n1066_));
  NA2        u1038(.A(men_men_n981_), .B(men_men_n973_), .Y(men_men_n1067_));
  NO3        u1039(.A(men_men_n566_), .B(men_men_n153_), .C(men_men_n222_), .Y(men_men_n1068_));
  OAI210     u1040(.A0(men_men_n1068_), .A1(men_men_n546_), .B0(men_men_n394_), .Y(men_men_n1069_));
  OAI220     u1041(.A0(men_men_n978_), .A1(men_men_n986_), .B0(men_men_n567_), .B1(men_men_n445_), .Y(men_men_n1070_));
  NA4        u1042(.A(men_men_n1070_), .B(men_men_n1069_), .C(men_men_n1067_), .D(men_men_n648_), .Y(men_men_n1071_));
  OAI210     u1043(.A0(men_men_n981_), .A1(men_men_n974_), .B0(men_men_n1057_), .Y(men_men_n1072_));
  AOI210     u1044(.A0(men_men_n396_), .A1(men_men_n394_), .B0(men_men_n342_), .Y(men_men_n1073_));
  NA3        u1045(.A(men_men_n1073_), .B(men_men_n1072_), .C(men_men_n285_), .Y(men_men_n1074_));
  OR4        u1046(.A(men_men_n1074_), .B(men_men_n1071_), .C(men_men_n1066_), .D(men_men_n1065_), .Y(men_men_n1075_));
  NO4        u1047(.A(men_men_n1075_), .B(men_men_n1064_), .C(men_men_n1059_), .D(men_men_n1056_), .Y(men_men_n1076_));
  NA4        u1048(.A(men_men_n1076_), .B(men_men_n1049_), .C(men_men_n1011_), .D(men_men_n998_), .Y(men13));
  NA2        u1049(.A(men_men_n46_), .B(men_men_n87_), .Y(men_men_n1078_));
  AN2        u1050(.A(c), .B(b), .Y(men_men_n1079_));
  NA3        u1051(.A(men_men_n261_), .B(men_men_n1079_), .C(m), .Y(men_men_n1080_));
  NO4        u1052(.A(e), .B(men_men_n1080_), .C(men_men_n1078_), .D(men_men_n609_), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n276_), .B(men_men_n1079_), .Y(men_men_n1082_));
  NO4        u1054(.A(men_men_n1082_), .B(e), .C(men_men_n1013_), .D(a), .Y(men_men_n1083_));
  NAi32      u1055(.An(d), .Bn(c), .C(e), .Y(men_men_n1084_));
  NA2        u1056(.A(men_men_n143_), .B(men_men_n45_), .Y(men_men_n1085_));
  NO4        u1057(.A(men_men_n1085_), .B(men_men_n1084_), .C(men_men_n616_), .D(men_men_n317_), .Y(men_men_n1086_));
  NA2        u1058(.A(men_men_n698_), .B(men_men_n234_), .Y(men_men_n1087_));
  NA2        u1059(.A(men_men_n427_), .B(men_men_n222_), .Y(men_men_n1088_));
  AN2        u1060(.A(d), .B(c), .Y(men_men_n1089_));
  NA2        u1061(.A(men_men_n1089_), .B(men_men_n118_), .Y(men_men_n1090_));
  NO4        u1062(.A(men_men_n1090_), .B(men_men_n1088_), .C(men_men_n183_), .D(men_men_n174_), .Y(men_men_n1091_));
  NA2        u1063(.A(d), .B(c), .Y(men_men_n1092_));
  NO4        u1064(.A(men_men_n1085_), .B(men_men_n612_), .C(men_men_n1092_), .D(men_men_n317_), .Y(men_men_n1093_));
  AO210      u1065(.A0(men_men_n1091_), .A1(men_men_n1087_), .B0(men_men_n1093_), .Y(men_men_n1094_));
  OR4        u1066(.A(men_men_n1094_), .B(men_men_n1086_), .C(men_men_n1083_), .D(men_men_n1081_), .Y(men_men_n1095_));
  NAi32      u1067(.An(f), .Bn(e), .C(c), .Y(men_men_n1096_));
  NO2        u1068(.A(men_men_n1096_), .B(men_men_n150_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n1097_), .B(g), .Y(men_men_n1098_));
  OR3        u1070(.A(men_men_n234_), .B(men_men_n183_), .C(men_men_n174_), .Y(men_men_n1099_));
  NO2        u1071(.A(men_men_n1099_), .B(men_men_n1098_), .Y(men_men_n1100_));
  NO2        u1072(.A(men_men_n1092_), .B(men_men_n317_), .Y(men_men_n1101_));
  NO2        u1073(.A(j), .B(men_men_n45_), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n658_), .B(men_men_n1102_), .Y(men_men_n1103_));
  NOi21      u1075(.An(men_men_n1101_), .B(men_men_n1103_), .Y(men_men_n1104_));
  NO2        u1076(.A(men_men_n798_), .B(men_men_n114_), .Y(men_men_n1105_));
  NOi41      u1077(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1106_));
  NA2        u1078(.A(men_men_n1106_), .B(men_men_n1105_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n1107_), .B(men_men_n1098_), .Y(men_men_n1108_));
  OR3        u1080(.A(e), .B(d), .C(c), .Y(men_men_n1109_));
  NA3        u1081(.A(k), .B(j), .C(i), .Y(men_men_n1110_));
  NO3        u1082(.A(men_men_n1110_), .B(men_men_n317_), .C(men_men_n91_), .Y(men_men_n1111_));
  NOi21      u1083(.An(men_men_n1111_), .B(men_men_n1109_), .Y(men_men_n1112_));
  OR4        u1084(.A(men_men_n1112_), .B(men_men_n1108_), .C(men_men_n1104_), .D(men_men_n1100_), .Y(men_men_n1113_));
  NA3        u1085(.A(men_men_n488_), .B(men_men_n345_), .C(men_men_n56_), .Y(men_men_n1114_));
  NO2        u1086(.A(men_men_n1114_), .B(men_men_n1103_), .Y(men_men_n1115_));
  NO4        u1087(.A(men_men_n1114_), .B(men_men_n612_), .C(men_men_n469_), .D(men_men_n45_), .Y(men_men_n1116_));
  NO2        u1088(.A(f), .B(c), .Y(men_men_n1117_));
  NOi21      u1089(.An(men_men_n1117_), .B(men_men_n461_), .Y(men_men_n1118_));
  NA2        u1090(.A(men_men_n1118_), .B(men_men_n59_), .Y(men_men_n1119_));
  NO3        u1091(.A(k), .B(men_men_n254_), .C(l), .Y(men_men_n1120_));
  NOi31      u1092(.An(men_men_n1120_), .B(men_men_n1119_), .C(j), .Y(men_men_n1121_));
  OR3        u1093(.A(men_men_n1121_), .B(men_men_n1116_), .C(men_men_n1115_), .Y(men_men_n1122_));
  OR3        u1094(.A(men_men_n1122_), .B(men_men_n1113_), .C(men_men_n1095_), .Y(men02));
  OR2        u1095(.A(l), .B(k), .Y(men_men_n1124_));
  OR3        u1096(.A(h), .B(g), .C(f), .Y(men_men_n1125_));
  OR3        u1097(.A(n), .B(m), .C(i), .Y(men_men_n1126_));
  NO4        u1098(.A(men_men_n1126_), .B(men_men_n1125_), .C(men_men_n1124_), .D(men_men_n1109_), .Y(men_men_n1127_));
  NOi31      u1099(.An(e), .B(d), .C(c), .Y(men_men_n1128_));
  AOI210     u1100(.A0(men_men_n1111_), .A1(men_men_n1128_), .B0(men_men_n1086_), .Y(men_men_n1129_));
  AN3        u1101(.A(g), .B(f), .C(c), .Y(men_men_n1130_));
  NA3        u1102(.A(men_men_n1130_), .B(men_men_n488_), .C(h), .Y(men_men_n1131_));
  OR2        u1103(.A(men_men_n1110_), .B(men_men_n1131_), .Y(men_men_n1132_));
  NO3        u1104(.A(men_men_n1114_), .B(men_men_n1085_), .C(men_men_n612_), .Y(men_men_n1133_));
  NO2        u1105(.A(men_men_n1133_), .B(men_men_n1100_), .Y(men_men_n1134_));
  NA3        u1106(.A(l), .B(k), .C(j), .Y(men_men_n1135_));
  NA2        u1107(.A(i), .B(h), .Y(men_men_n1136_));
  NO3        u1108(.A(men_men_n1136_), .B(men_men_n1135_), .C(men_men_n134_), .Y(men_men_n1137_));
  NO3        u1109(.A(men_men_n145_), .B(men_men_n294_), .C(men_men_n223_), .Y(men_men_n1138_));
  INV        u1110(.A(men_men_n1104_), .Y(men_men_n1139_));
  NA3        u1111(.A(c), .B(b), .C(a), .Y(men_men_n1140_));
  NO3        u1112(.A(men_men_n1140_), .B(men_men_n946_), .C(men_men_n222_), .Y(men_men_n1141_));
  INV        u1113(.A(men_men_n1115_), .Y(men_men_n1142_));
  AN4        u1114(.A(men_men_n1142_), .B(men_men_n1139_), .C(men_men_n1134_), .D(men_men_n1132_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n1090_), .B(men_men_n1088_), .Y(men_men_n1144_));
  NA2        u1116(.A(men_men_n1107_), .B(men_men_n1099_), .Y(men_men_n1145_));
  AOI210     u1117(.A0(men_men_n1145_), .A1(men_men_n1144_), .B0(men_men_n1081_), .Y(men_men_n1146_));
  NAi41      u1118(.An(men_men_n1127_), .B(men_men_n1146_), .C(men_men_n1143_), .D(men_men_n1129_), .Y(men03));
  NO2        u1119(.A(men_men_n548_), .B(men_men_n625_), .Y(men_men_n1148_));
  NA4        u1120(.A(men_men_n88_), .B(men_men_n87_), .C(g), .D(men_men_n222_), .Y(men_men_n1149_));
  NA4        u1121(.A(men_men_n600_), .B(m), .C(men_men_n114_), .D(men_men_n222_), .Y(men_men_n1150_));
  NA3        u1122(.A(men_men_n1150_), .B(men_men_n384_), .C(men_men_n1149_), .Y(men_men_n1151_));
  NO3        u1123(.A(men_men_n1151_), .B(men_men_n1148_), .C(men_men_n1044_), .Y(men_men_n1152_));
  NOi41      u1124(.An(men_men_n845_), .B(men_men_n896_), .C(men_men_n886_), .D(men_men_n747_), .Y(men_men_n1153_));
  OAI220     u1125(.A0(men_men_n1153_), .A1(men_men_n720_), .B0(men_men_n1152_), .B1(men_men_n613_), .Y(men_men_n1154_));
  NOi31      u1126(.An(i), .B(k), .C(j), .Y(men_men_n1155_));
  NA4        u1127(.A(men_men_n1155_), .B(men_men_n1128_), .C(men_men_n354_), .D(men_men_n345_), .Y(men_men_n1156_));
  OAI210     u1128(.A0(men_men_n860_), .A1(men_men_n438_), .B0(men_men_n1156_), .Y(men_men_n1157_));
  NOi31      u1129(.An(m), .B(n), .C(f), .Y(men_men_n1158_));
  NA2        u1130(.A(men_men_n1158_), .B(men_men_n51_), .Y(men_men_n1159_));
  AN2        u1131(.A(e), .B(c), .Y(men_men_n1160_));
  NA2        u1132(.A(men_men_n1160_), .B(a), .Y(men_men_n1161_));
  OAI220     u1133(.A0(men_men_n1161_), .A1(men_men_n1159_), .B0(men_men_n930_), .B1(men_men_n444_), .Y(men_men_n1162_));
  NA2        u1134(.A(men_men_n527_), .B(l), .Y(men_men_n1163_));
  NOi31      u1135(.An(men_men_n907_), .B(men_men_n1080_), .C(men_men_n1163_), .Y(men_men_n1164_));
  NO4        u1136(.A(men_men_n1164_), .B(men_men_n1162_), .C(men_men_n1157_), .D(men_men_n1043_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n294_), .B(a), .Y(men_men_n1166_));
  INV        u1138(.A(men_men_n1086_), .Y(men_men_n1167_));
  NO2        u1139(.A(men_men_n1136_), .B(men_men_n507_), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n87_), .B(g), .Y(men_men_n1169_));
  AOI210     u1141(.A0(men_men_n1169_), .A1(men_men_n1168_), .B0(men_men_n1120_), .Y(men_men_n1170_));
  OR2        u1142(.A(men_men_n1170_), .B(men_men_n1119_), .Y(men_men_n1171_));
  NA3        u1143(.A(men_men_n1171_), .B(men_men_n1167_), .C(men_men_n1165_), .Y(men_men_n1172_));
  NO4        u1144(.A(men_men_n1172_), .B(men_men_n1154_), .C(men_men_n862_), .D(men_men_n589_), .Y(men_men_n1173_));
  NA2        u1145(.A(c), .B(b), .Y(men_men_n1174_));
  NO2        u1146(.A(men_men_n732_), .B(men_men_n1174_), .Y(men_men_n1175_));
  OAI210     u1147(.A0(men_men_n905_), .A1(men_men_n877_), .B0(men_men_n431_), .Y(men_men_n1176_));
  OAI210     u1148(.A0(men_men_n1176_), .A1(men_men_n906_), .B0(men_men_n1175_), .Y(men_men_n1177_));
  NAi21      u1149(.An(men_men_n439_), .B(men_men_n1175_), .Y(men_men_n1178_));
  NA2        u1150(.A(men_men_n445_), .B(men_men_n582_), .Y(men_men_n1179_));
  OAI210     u1151(.A0(men_men_n571_), .A1(men_men_n39_), .B0(men_men_n1166_), .Y(men_men_n1180_));
  NA3        u1152(.A(men_men_n1180_), .B(men_men_n1179_), .C(men_men_n1178_), .Y(men_men_n1181_));
  INV        u1153(.A(g), .Y(men_men_n1182_));
  NAi21      u1154(.An(f), .B(d), .Y(men_men_n1183_));
  NO2        u1155(.A(men_men_n1183_), .B(men_men_n1140_), .Y(men_men_n1184_));
  INV        u1156(.A(men_men_n1184_), .Y(men_men_n1185_));
  AOI210     u1157(.A0(men_men_n1182_), .A1(men_men_n302_), .B0(men_men_n1185_), .Y(men_men_n1186_));
  AOI210     u1158(.A0(men_men_n1186_), .A1(men_men_n115_), .B0(men_men_n1181_), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n491_), .B(men_men_n490_), .Y(men_men_n1188_));
  NO2        u1160(.A(men_men_n189_), .B(men_men_n247_), .Y(men_men_n1189_));
  NA2        u1161(.A(men_men_n1189_), .B(m), .Y(men_men_n1190_));
  NA3        u1162(.A(men_men_n962_), .B(men_men_n1163_), .C(men_men_n494_), .Y(men_men_n1191_));
  OAI210     u1163(.A0(men_men_n1191_), .A1(men_men_n322_), .B0(men_men_n492_), .Y(men_men_n1192_));
  AOI210     u1164(.A0(men_men_n1192_), .A1(men_men_n1188_), .B0(men_men_n1190_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n584_), .B(men_men_n426_), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n465_), .B(men_men_n1184_), .Y(men_men_n1195_));
  NO2        u1167(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n1196_));
  AOI210     u1168(.A0(men_men_n1189_), .A1(men_men_n447_), .B0(men_men_n1005_), .Y(men_men_n1197_));
  NAi41      u1169(.An(men_men_n1196_), .B(men_men_n1197_), .C(men_men_n1195_), .D(men_men_n1194_), .Y(men_men_n1198_));
  NO2        u1170(.A(men_men_n1198_), .B(men_men_n1193_), .Y(men_men_n1199_));
  NA4        u1171(.A(men_men_n1199_), .B(men_men_n1187_), .C(men_men_n1177_), .D(men_men_n1173_), .Y(men00));
  NO2        u1172(.A(men_men_n309_), .B(men_men_n288_), .Y(men_men_n1201_));
  NO2        u1173(.A(men_men_n1201_), .B(men_men_n603_), .Y(men_men_n1202_));
  AOI210     u1174(.A0(men_men_n943_), .A1(men_men_n988_), .B0(men_men_n1157_), .Y(men_men_n1203_));
  NO3        u1175(.A(men_men_n1133_), .B(men_men_n1005_), .C(men_men_n744_), .Y(men_men_n1204_));
  NA3        u1176(.A(men_men_n1204_), .B(men_men_n1203_), .C(men_men_n1045_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n529_), .B(f), .Y(men_men_n1206_));
  OAI210     u1178(.A0(men_men_n1051_), .A1(men_men_n40_), .B0(men_men_n677_), .Y(men_men_n1207_));
  NA3        u1179(.A(men_men_n1207_), .B(men_men_n268_), .C(n), .Y(men_men_n1208_));
  AOI210     u1180(.A0(men_men_n1208_), .A1(men_men_n1206_), .B0(men_men_n1090_), .Y(men_men_n1209_));
  NO4        u1181(.A(men_men_n1209_), .B(men_men_n1205_), .C(men_men_n1202_), .D(men_men_n1113_), .Y(men_men_n1210_));
  NA3        u1182(.A(men_men_n173_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1211_));
  NA3        u1183(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1212_));
  NOi31      u1184(.An(n), .B(m), .C(i), .Y(men_men_n1213_));
  NA3        u1185(.A(men_men_n1213_), .B(men_men_n680_), .C(men_men_n51_), .Y(men_men_n1214_));
  OAI210     u1186(.A0(men_men_n1212_), .A1(men_men_n1211_), .B0(men_men_n1214_), .Y(men_men_n1215_));
  INV        u1187(.A(men_men_n602_), .Y(men_men_n1216_));
  NO4        u1188(.A(men_men_n1216_), .B(men_men_n1215_), .C(men_men_n1196_), .D(men_men_n965_), .Y(men_men_n1217_));
  NA3        u1189(.A(men_men_n399_), .B(men_men_n230_), .C(g), .Y(men_men_n1218_));
  OA220      u1190(.A0(men_men_n1218_), .A1(men_men_n1212_), .B0(men_men_n400_), .B1(men_men_n137_), .Y(men_men_n1219_));
  NO2        u1191(.A(h), .B(g), .Y(men_men_n1220_));
  NA4        u1192(.A(men_men_n518_), .B(men_men_n488_), .C(men_men_n1220_), .D(men_men_n1079_), .Y(men_men_n1221_));
  OAI220     u1193(.A0(men_men_n548_), .A1(men_men_n625_), .B0(men_men_n92_), .B1(men_men_n91_), .Y(men_men_n1222_));
  AOI220     u1194(.A0(men_men_n1222_), .A1(men_men_n557_), .B0(men_men_n993_), .B1(men_men_n601_), .Y(men_men_n1223_));
  AOI220     u1195(.A0(men_men_n328_), .A1(men_men_n258_), .B0(men_men_n184_), .B1(men_men_n152_), .Y(men_men_n1224_));
  NA4        u1196(.A(men_men_n1224_), .B(men_men_n1223_), .C(men_men_n1221_), .D(men_men_n1219_), .Y(men_men_n1225_));
  NO2        u1197(.A(men_men_n1225_), .B(men_men_n278_), .Y(men_men_n1226_));
  INV        u1198(.A(men_men_n333_), .Y(men_men_n1227_));
  AOI210     u1199(.A0(men_men_n258_), .A1(men_men_n359_), .B0(men_men_n604_), .Y(men_men_n1228_));
  NA3        u1200(.A(men_men_n1228_), .B(men_men_n1227_), .C(men_men_n158_), .Y(men_men_n1229_));
  NO2        u1201(.A(men_men_n249_), .B(men_men_n188_), .Y(men_men_n1230_));
  NA2        u1202(.A(men_men_n1230_), .B(men_men_n445_), .Y(men_men_n1231_));
  NA3        u1203(.A(men_men_n186_), .B(men_men_n114_), .C(g), .Y(men_men_n1232_));
  NA3        u1204(.A(men_men_n488_), .B(men_men_n40_), .C(f), .Y(men_men_n1233_));
  NOi31      u1205(.An(men_men_n915_), .B(men_men_n1233_), .C(men_men_n1232_), .Y(men_men_n1234_));
  NAi31      u1206(.An(men_men_n193_), .B(men_men_n902_), .C(men_men_n488_), .Y(men_men_n1235_));
  NAi31      u1207(.An(men_men_n1234_), .B(men_men_n1235_), .C(men_men_n1231_), .Y(men_men_n1236_));
  NO2        u1208(.A(men_men_n287_), .B(men_men_n73_), .Y(men_men_n1237_));
  NO3        u1209(.A(men_men_n444_), .B(men_men_n873_), .C(n), .Y(men_men_n1238_));
  AOI210     u1210(.A0(men_men_n1238_), .A1(men_men_n1237_), .B0(men_men_n1127_), .Y(men_men_n1239_));
  NAi31      u1211(.An(men_men_n1093_), .B(men_men_n1239_), .C(men_men_n72_), .Y(men_men_n1240_));
  NO4        u1212(.A(men_men_n1240_), .B(men_men_n1236_), .C(men_men_n1229_), .D(men_men_n539_), .Y(men_men_n1241_));
  AN3        u1213(.A(men_men_n1241_), .B(men_men_n1226_), .C(men_men_n1217_), .Y(men_men_n1242_));
  NA2        u1214(.A(men_men_n557_), .B(men_men_n102_), .Y(men_men_n1243_));
  NA3        u1215(.A(men_men_n1158_), .B(men_men_n636_), .C(men_men_n487_), .Y(men_men_n1244_));
  NA4        u1216(.A(men_men_n1244_), .B(men_men_n585_), .C(men_men_n1243_), .D(men_men_n252_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n1151_), .B(men_men_n557_), .Y(men_men_n1246_));
  NA4        u1218(.A(men_men_n680_), .B(men_men_n214_), .C(men_men_n230_), .D(men_men_n167_), .Y(men_men_n1247_));
  NA3        u1219(.A(men_men_n1247_), .B(men_men_n1246_), .C(men_men_n306_), .Y(men_men_n1248_));
  OAI210     u1220(.A0(men_men_n486_), .A1(men_men_n122_), .B0(men_men_n908_), .Y(men_men_n1249_));
  AOI220     u1221(.A0(men_men_n1249_), .A1(men_men_n1191_), .B0(men_men_n584_), .B1(men_men_n426_), .Y(men_men_n1250_));
  OR4        u1222(.A(men_men_n1090_), .B(men_men_n284_), .C(men_men_n232_), .D(e), .Y(men_men_n1251_));
  NO2        u1223(.A(men_men_n226_), .B(men_men_n223_), .Y(men_men_n1252_));
  NA2        u1224(.A(n), .B(e), .Y(men_men_n1253_));
  NO2        u1225(.A(men_men_n1253_), .B(men_men_n150_), .Y(men_men_n1254_));
  AOI220     u1226(.A0(men_men_n1254_), .A1(men_men_n286_), .B0(men_men_n890_), .B1(men_men_n1252_), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n370_), .A1(men_men_n323_), .B0(men_men_n467_), .Y(men_men_n1256_));
  NA4        u1228(.A(men_men_n1256_), .B(men_men_n1255_), .C(men_men_n1251_), .D(men_men_n1250_), .Y(men_men_n1257_));
  AOI210     u1229(.A0(men_men_n1254_), .A1(men_men_n893_), .B0(men_men_n861_), .Y(men_men_n1258_));
  AOI220     u1230(.A0(men_men_n1001_), .A1(men_men_n601_), .B0(men_men_n680_), .B1(men_men_n255_), .Y(men_men_n1259_));
  NO2        u1231(.A(men_men_n66_), .B(h), .Y(men_men_n1260_));
  NO3        u1232(.A(men_men_n1090_), .B(men_men_n1088_), .C(men_men_n761_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n1124_), .B(men_men_n134_), .Y(men_men_n1262_));
  AN2        u1234(.A(men_men_n1262_), .B(men_men_n1138_), .Y(men_men_n1263_));
  OAI210     u1235(.A0(men_men_n1263_), .A1(men_men_n1261_), .B0(men_men_n1260_), .Y(men_men_n1264_));
  NA4        u1236(.A(men_men_n1264_), .B(men_men_n1259_), .C(men_men_n1258_), .D(men_men_n910_), .Y(men_men_n1265_));
  NO4        u1237(.A(men_men_n1265_), .B(men_men_n1257_), .C(men_men_n1248_), .D(men_men_n1245_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n878_), .B(men_men_n793_), .Y(men_men_n1267_));
  NA4        u1239(.A(men_men_n1267_), .B(men_men_n1266_), .C(men_men_n1242_), .D(men_men_n1210_), .Y(men01));
  AN2        u1240(.A(men_men_n1069_), .B(men_men_n1067_), .Y(men_men_n1269_));
  NO3        u1241(.A(men_men_n841_), .B(men_men_n833_), .C(men_men_n502_), .Y(men_men_n1270_));
  NO2        u1242(.A(men_men_n618_), .B(men_men_n299_), .Y(men_men_n1271_));
  OAI210     u1243(.A0(men_men_n1271_), .A1(men_men_n410_), .B0(i), .Y(men_men_n1272_));
  NA3        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n1269_), .Y(men_men_n1273_));
  NA2        u1245(.A(men_men_n614_), .B(men_men_n90_), .Y(men_men_n1274_));
  NA2        u1246(.A(men_men_n577_), .B(men_men_n283_), .Y(men_men_n1275_));
  NA2        u1247(.A(men_men_n1008_), .B(men_men_n1275_), .Y(men_men_n1276_));
  NA4        u1248(.A(men_men_n1276_), .B(men_men_n1274_), .C(men_men_n958_), .D(men_men_n344_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n739_), .B(men_men_n97_), .Y(men_men_n1278_));
  NO2        u1250(.A(men_men_n1278_), .B(i), .Y(men_men_n1279_));
  OAI210     u1251(.A0(men_men_n819_), .A1(men_men_n631_), .B0(men_men_n1247_), .Y(men_men_n1280_));
  AOI210     u1252(.A0(men_men_n1279_), .A1(men_men_n665_), .B0(men_men_n1280_), .Y(men_men_n1281_));
  NA2        u1253(.A(men_men_n120_), .B(l), .Y(men_men_n1282_));
  OA220      u1254(.A0(men_men_n1282_), .A1(men_men_n611_), .B0(men_men_n693_), .B1(men_men_n384_), .Y(men_men_n1283_));
  NAi41      u1255(.An(men_men_n166_), .B(men_men_n1283_), .C(men_men_n1281_), .D(men_men_n942_), .Y(men_men_n1284_));
  NO3        u1256(.A(men_men_n820_), .B(men_men_n705_), .C(men_men_n532_), .Y(men_men_n1285_));
  NA3        u1257(.A(men_men_n739_), .B(men_men_n97_), .C(men_men_n222_), .Y(men_men_n1286_));
  OR2        u1258(.A(men_men_n203_), .B(men_men_n201_), .Y(men_men_n1287_));
  NA3        u1259(.A(men_men_n1287_), .B(men_men_n1285_), .C(men_men_n140_), .Y(men_men_n1288_));
  NO4        u1260(.A(men_men_n1288_), .B(men_men_n1284_), .C(men_men_n1277_), .D(men_men_n1273_), .Y(men_men_n1289_));
  NA2        u1261(.A(men_men_n1218_), .B(men_men_n215_), .Y(men_men_n1290_));
  OAI210     u1262(.A0(men_men_n1290_), .A1(men_men_n312_), .B0(men_men_n552_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n560_), .B(men_men_n412_), .Y(men_men_n1292_));
  NA2        u1264(.A(men_men_n74_), .B(i), .Y(men_men_n1293_));
  AOI210     u1265(.A0(men_men_n617_), .A1(men_men_n611_), .B0(men_men_n1293_), .Y(men_men_n1294_));
  AOI210     u1266(.A0(men_men_n586_), .A1(men_men_n1292_), .B0(men_men_n1294_), .Y(men_men_n1295_));
  AOI210     u1267(.A0(men_men_n212_), .A1(men_men_n89_), .B0(men_men_n222_), .Y(men_men_n1296_));
  OAI210     u1268(.A0(men_men_n848_), .A1(men_men_n445_), .B0(men_men_n1296_), .Y(men_men_n1297_));
  AN3        u1269(.A(m), .B(l), .C(k), .Y(men_men_n1298_));
  OAI210     u1270(.A0(men_men_n372_), .A1(men_men_n34_), .B0(men_men_n1298_), .Y(men_men_n1299_));
  NA2        u1271(.A(men_men_n211_), .B(men_men_n34_), .Y(men_men_n1300_));
  AO210      u1272(.A0(men_men_n1300_), .A1(men_men_n1299_), .B0(men_men_n343_), .Y(men_men_n1301_));
  NA4        u1273(.A(men_men_n1301_), .B(men_men_n1297_), .C(men_men_n1295_), .D(men_men_n1291_), .Y(men_men_n1302_));
  AOI210     u1274(.A0(men_men_n623_), .A1(men_men_n120_), .B0(men_men_n629_), .Y(men_men_n1303_));
  OAI210     u1275(.A0(men_men_n1282_), .A1(men_men_n620_), .B0(men_men_n1303_), .Y(men_men_n1304_));
  NO3        u1276(.A(men_men_n860_), .B(men_men_n212_), .C(men_men_n424_), .Y(men_men_n1305_));
  NO2        u1277(.A(men_men_n1305_), .B(men_men_n1005_), .Y(men_men_n1306_));
  OAI210     u1278(.A0(men_men_n1279_), .A1(men_men_n338_), .B0(men_men_n706_), .Y(men_men_n1307_));
  NA3        u1279(.A(men_men_n1307_), .B(men_men_n1306_), .C(men_men_n823_), .Y(men_men_n1308_));
  NO3        u1280(.A(men_men_n1308_), .B(men_men_n1304_), .C(men_men_n1302_), .Y(men_men_n1309_));
  NA3        u1281(.A(men_men_n632_), .B(men_men_n29_), .C(f), .Y(men_men_n1310_));
  NO2        u1282(.A(men_men_n1310_), .B(men_men_n212_), .Y(men_men_n1311_));
  AOI210     u1283(.A0(men_men_n524_), .A1(men_men_n58_), .B0(men_men_n1311_), .Y(men_men_n1312_));
  OR3        u1284(.A(men_men_n1278_), .B(men_men_n633_), .C(i), .Y(men_men_n1313_));
  NA3        u1285(.A(men_men_n775_), .B(men_men_n74_), .C(i), .Y(men_men_n1314_));
  AOI210     u1286(.A0(men_men_n1314_), .A1(men_men_n1286_), .B0(men_men_n1025_), .Y(men_men_n1315_));
  NO2        u1287(.A(men_men_n215_), .B(men_men_n113_), .Y(men_men_n1316_));
  NO3        u1288(.A(men_men_n1316_), .B(men_men_n1315_), .C(men_men_n1215_), .Y(men_men_n1317_));
  NA4        u1289(.A(men_men_n1317_), .B(men_men_n1313_), .C(men_men_n1312_), .D(men_men_n792_), .Y(men_men_n1318_));
  NO2        u1290(.A(men_men_n1013_), .B(men_men_n242_), .Y(men_men_n1319_));
  NO2        u1291(.A(men_men_n1014_), .B(men_men_n579_), .Y(men_men_n1320_));
  OAI210     u1292(.A0(men_men_n1320_), .A1(men_men_n1319_), .B0(men_men_n352_), .Y(men_men_n1321_));
  NA2        u1293(.A(men_men_n596_), .B(men_men_n594_), .Y(men_men_n1322_));
  NO3        u1294(.A(men_men_n79_), .B(men_men_n310_), .C(men_men_n45_), .Y(men_men_n1323_));
  NA2        u1295(.A(men_men_n1323_), .B(men_men_n576_), .Y(men_men_n1324_));
  NA3        u1296(.A(men_men_n1324_), .B(men_men_n1322_), .C(men_men_n701_), .Y(men_men_n1325_));
  OR2        u1297(.A(men_men_n1218_), .B(men_men_n1212_), .Y(men_men_n1326_));
  NO2        u1298(.A(men_men_n384_), .B(men_men_n71_), .Y(men_men_n1327_));
  AOI210     u1299(.A0(men_men_n766_), .A1(men_men_n645_), .B0(men_men_n1327_), .Y(men_men_n1328_));
  NA2        u1300(.A(men_men_n1323_), .B(men_men_n851_), .Y(men_men_n1329_));
  NA4        u1301(.A(men_men_n1329_), .B(men_men_n1328_), .C(men_men_n1326_), .D(men_men_n402_), .Y(men_men_n1330_));
  NOi41      u1302(.An(men_men_n1321_), .B(men_men_n1330_), .C(men_men_n1325_), .D(men_men_n1318_), .Y(men_men_n1331_));
  NO2        u1303(.A(men_men_n133_), .B(men_men_n45_), .Y(men_men_n1332_));
  NO2        u1304(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1333_));
  AO220      u1305(.A0(men_men_n1333_), .A1(men_men_n651_), .B0(men_men_n1332_), .B1(men_men_n737_), .Y(men_men_n1334_));
  NA2        u1306(.A(men_men_n1334_), .B(men_men_n352_), .Y(men_men_n1335_));
  INV        u1307(.A(men_men_n137_), .Y(men_men_n1336_));
  NO3        u1308(.A(men_men_n1136_), .B(men_men_n183_), .C(men_men_n87_), .Y(men_men_n1337_));
  AOI220     u1309(.A0(men_men_n1337_), .A1(men_men_n1336_), .B0(men_men_n1323_), .B1(men_men_n1017_), .Y(men_men_n1338_));
  NA2        u1310(.A(men_men_n1338_), .B(men_men_n1335_), .Y(men_men_n1339_));
  NO2        u1311(.A(men_men_n643_), .B(men_men_n642_), .Y(men_men_n1340_));
  NO4        u1312(.A(men_men_n1136_), .B(men_men_n1340_), .C(men_men_n181_), .D(men_men_n87_), .Y(men_men_n1341_));
  NO3        u1313(.A(men_men_n1341_), .B(men_men_n1339_), .C(men_men_n669_), .Y(men_men_n1342_));
  NA4        u1314(.A(men_men_n1342_), .B(men_men_n1331_), .C(men_men_n1309_), .D(men_men_n1289_), .Y(men06));
  NO2        u1315(.A(men_men_n425_), .B(men_men_n583_), .Y(men_men_n1344_));
  NA2        u1316(.A(men_men_n279_), .B(men_men_n1344_), .Y(men_men_n1345_));
  NO2        u1317(.A(men_men_n234_), .B(men_men_n104_), .Y(men_men_n1346_));
  OAI210     u1318(.A0(men_men_n1346_), .A1(men_men_n1337_), .B0(men_men_n398_), .Y(men_men_n1347_));
  NO3        u1319(.A(men_men_n627_), .B(men_men_n846_), .C(men_men_n630_), .Y(men_men_n1348_));
  OR2        u1320(.A(men_men_n1348_), .B(men_men_n930_), .Y(men_men_n1349_));
  NA4        u1321(.A(men_men_n1349_), .B(men_men_n1347_), .C(men_men_n1345_), .D(men_men_n1321_), .Y(men_men_n1350_));
  NO3        u1322(.A(men_men_n1350_), .B(men_men_n1325_), .C(men_men_n267_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n310_), .B(men_men_n45_), .Y(men_men_n1352_));
  NA2        u1324(.A(men_men_n1352_), .B(men_men_n1018_), .Y(men_men_n1353_));
  AOI210     u1325(.A0(men_men_n1352_), .A1(men_men_n580_), .B0(men_men_n1334_), .Y(men_men_n1354_));
  AOI210     u1326(.A0(men_men_n1354_), .A1(men_men_n1353_), .B0(men_men_n349_), .Y(men_men_n1355_));
  OAI210     u1327(.A0(men_men_n89_), .A1(men_men_n40_), .B0(men_men_n704_), .Y(men_men_n1356_));
  NA2        u1328(.A(men_men_n1356_), .B(men_men_n673_), .Y(men_men_n1357_));
  NO2        u1329(.A(men_men_n535_), .B(men_men_n178_), .Y(men_men_n1358_));
  NO2        u1330(.A(men_men_n637_), .B(men_men_n1159_), .Y(men_men_n1359_));
  NO3        u1331(.A(men_men_n1359_), .B(men_men_n139_), .C(men_men_n1358_), .Y(men_men_n1360_));
  OR2        u1332(.A(men_men_n628_), .B(men_men_n626_), .Y(men_men_n1361_));
  NO2        u1333(.A(men_men_n383_), .B(men_men_n138_), .Y(men_men_n1362_));
  AOI210     u1334(.A0(men_men_n1362_), .A1(men_men_n614_), .B0(men_men_n1361_), .Y(men_men_n1363_));
  NA3        u1335(.A(men_men_n1363_), .B(men_men_n1360_), .C(men_men_n1357_), .Y(men_men_n1364_));
  NO2        u1336(.A(men_men_n783_), .B(men_men_n382_), .Y(men_men_n1365_));
  NO3        u1337(.A(men_men_n706_), .B(men_men_n794_), .C(men_men_n665_), .Y(men_men_n1366_));
  NOi21      u1338(.An(men_men_n1365_), .B(men_men_n1366_), .Y(men_men_n1367_));
  AN2        u1339(.A(men_men_n1001_), .B(men_men_n676_), .Y(men_men_n1368_));
  NO4        u1340(.A(men_men_n1368_), .B(men_men_n1367_), .C(men_men_n1364_), .D(men_men_n1355_), .Y(men_men_n1369_));
  NO2        u1341(.A(men_men_n840_), .B(men_men_n289_), .Y(men_men_n1370_));
  OAI220     u1342(.A0(men_men_n768_), .A1(men_men_n47_), .B0(men_men_n234_), .B1(men_men_n644_), .Y(men_men_n1371_));
  OAI210     u1343(.A0(men_men_n289_), .A1(c), .B0(men_men_n672_), .Y(men_men_n1372_));
  AOI220     u1344(.A0(men_men_n1372_), .A1(men_men_n1371_), .B0(men_men_n1370_), .B1(men_men_n279_), .Y(men_men_n1373_));
  NO3        u1345(.A(men_men_n254_), .B(men_men_n104_), .C(men_men_n294_), .Y(men_men_n1374_));
  OAI220     u1346(.A0(men_men_n729_), .A1(men_men_n259_), .B0(men_men_n531_), .B1(men_men_n535_), .Y(men_men_n1375_));
  OAI210     u1347(.A0(l), .A1(i), .B0(k), .Y(men_men_n1376_));
  NO3        u1348(.A(men_men_n1376_), .B(men_men_n625_), .C(j), .Y(men_men_n1377_));
  NOi21      u1349(.An(men_men_n1377_), .B(men_men_n699_), .Y(men_men_n1378_));
  NO4        u1350(.A(men_men_n1378_), .B(men_men_n1375_), .C(men_men_n1374_), .D(men_men_n1162_), .Y(men_men_n1379_));
  NA4        u1351(.A(men_men_n831_), .B(men_men_n830_), .C(men_men_n455_), .D(men_men_n922_), .Y(men_men_n1380_));
  NAi31      u1352(.An(men_men_n783_), .B(men_men_n1380_), .C(men_men_n211_), .Y(men_men_n1381_));
  NA4        u1353(.A(men_men_n1381_), .B(men_men_n1379_), .C(men_men_n1373_), .D(men_men_n1259_), .Y(men_men_n1382_));
  OR2        u1354(.A(men_men_n819_), .B(men_men_n563_), .Y(men_men_n1383_));
  OR3        u1355(.A(men_men_n386_), .B(men_men_n234_), .C(men_men_n644_), .Y(men_men_n1384_));
  AOI210     u1356(.A0(men_men_n596_), .A1(men_men_n467_), .B0(men_men_n388_), .Y(men_men_n1385_));
  NA2        u1357(.A(men_men_n1377_), .B(men_men_n827_), .Y(men_men_n1386_));
  NA4        u1358(.A(men_men_n1386_), .B(men_men_n1385_), .C(men_men_n1384_), .D(men_men_n1383_), .Y(men_men_n1387_));
  AOI220     u1359(.A0(men_men_n1365_), .A1(men_men_n793_), .B0(men_men_n1362_), .B1(men_men_n248_), .Y(men_men_n1388_));
  AN2        u1360(.A(men_men_n974_), .B(men_men_n973_), .Y(men_men_n1389_));
  NO4        u1361(.A(men_men_n1389_), .B(men_men_n920_), .C(men_men_n520_), .D(men_men_n505_), .Y(men_men_n1390_));
  NA3        u1362(.A(men_men_n1390_), .B(men_men_n1388_), .C(men_men_n1329_), .Y(men_men_n1391_));
  NAi21      u1363(.An(j), .B(i), .Y(men_men_n1392_));
  NO4        u1364(.A(men_men_n1340_), .B(men_men_n1392_), .C(men_men_n461_), .D(men_men_n245_), .Y(men_men_n1393_));
  NO4        u1365(.A(men_men_n1393_), .B(men_men_n1391_), .C(men_men_n1387_), .D(men_men_n1382_), .Y(men_men_n1394_));
  NA4        u1366(.A(men_men_n1394_), .B(men_men_n1369_), .C(men_men_n1351_), .D(men_men_n1342_), .Y(men07));
  NOi21      u1367(.An(j), .B(k), .Y(men_men_n1396_));
  NAi32      u1368(.An(m), .Bn(b), .C(n), .Y(men_men_n1397_));
  NO3        u1369(.A(men_men_n1397_), .B(g), .C(f), .Y(men_men_n1398_));
  OAI210     u1370(.A0(men_men_n332_), .A1(men_men_n506_), .B0(men_men_n1398_), .Y(men_men_n1399_));
  NAi21      u1371(.An(f), .B(c), .Y(men_men_n1400_));
  NOi31      u1372(.An(n), .B(m), .C(b), .Y(men_men_n1401_));
  INV        u1373(.A(men_men_n1399_), .Y(men_men_n1402_));
  NOi41      u1374(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1403_), .B(men_men_n912_), .C(men_men_n427_), .Y(men_men_n1404_));
  NO2        u1376(.A(men_men_n1404_), .B(men_men_n56_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1138_), .B(men_men_n230_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1406_), .B(men_men_n61_), .Y(men_men_n1407_));
  NA2        u1379(.A(men_men_n87_), .B(men_men_n45_), .Y(men_men_n1408_));
  NO2        u1380(.A(men_men_n1096_), .B(men_men_n461_), .Y(men_men_n1409_));
  NA3        u1381(.A(men_men_n1409_), .B(men_men_n1408_), .C(men_men_n223_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1110_), .B(men_men_n317_), .Y(men_men_n1411_));
  NA2        u1383(.A(men_men_n1260_), .B(men_men_n300_), .Y(men_men_n1412_));
  NA2        u1384(.A(men_men_n1412_), .B(men_men_n1410_), .Y(men_men_n1413_));
  NO4        u1385(.A(men_men_n1413_), .B(men_men_n1407_), .C(men_men_n1405_), .D(men_men_n1402_), .Y(men_men_n1414_));
  NO3        u1386(.A(e), .B(d), .C(c), .Y(men_men_n1415_));
  OAI210     u1387(.A0(men_men_n134_), .A1(men_men_n223_), .B0(men_men_n634_), .Y(men_men_n1416_));
  NA2        u1388(.A(men_men_n1416_), .B(men_men_n1415_), .Y(men_men_n1417_));
  INV        u1389(.A(men_men_n1417_), .Y(men_men_n1418_));
  OR2        u1390(.A(h), .B(f), .Y(men_men_n1419_));
  NO3        u1391(.A(n), .B(m), .C(i), .Y(men_men_n1420_));
  OAI210     u1392(.A0(men_men_n1160_), .A1(men_men_n161_), .B0(men_men_n1420_), .Y(men_men_n1421_));
  NO2        u1393(.A(i), .B(g), .Y(men_men_n1422_));
  OR3        u1394(.A(men_men_n1422_), .B(men_men_n1397_), .C(men_men_n70_), .Y(men_men_n1423_));
  OAI220     u1395(.A0(men_men_n1423_), .A1(men_men_n506_), .B0(men_men_n1421_), .B1(men_men_n1419_), .Y(men_men_n1424_));
  NA3        u1396(.A(men_men_n726_), .B(men_men_n712_), .C(men_men_n114_), .Y(men_men_n1425_));
  NA3        u1397(.A(men_men_n1401_), .B(men_men_n1105_), .C(h), .Y(men_men_n1426_));
  AOI210     u1398(.A0(men_men_n1426_), .A1(men_men_n1425_), .B0(men_men_n45_), .Y(men_men_n1427_));
  NA2        u1399(.A(men_men_n1420_), .B(men_men_n671_), .Y(men_men_n1428_));
  NO2        u1400(.A(l), .B(k), .Y(men_men_n1429_));
  NO3        u1401(.A(men_men_n461_), .B(d), .C(c), .Y(men_men_n1430_));
  NO3        u1402(.A(men_men_n1427_), .B(men_men_n1424_), .C(men_men_n1418_), .Y(men_men_n1431_));
  NO2        u1403(.A(men_men_n151_), .B(h), .Y(men_men_n1432_));
  NO2        u1404(.A(g), .B(c), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n472_), .B(a), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1434_), .B(men_men_n1586_), .C(men_men_n115_), .Y(men_men_n1435_));
  NO2        u1407(.A(i), .B(h), .Y(men_men_n1436_));
  NA2        u1408(.A(men_men_n1436_), .B(men_men_n230_), .Y(men_men_n1437_));
  AOI210     u1409(.A0(men_men_n1183_), .A1(h), .B0(men_men_n432_), .Y(men_men_n1438_));
  NA2        u1410(.A(men_men_n141_), .B(men_men_n230_), .Y(men_men_n1439_));
  AOI210     u1411(.A0(men_men_n268_), .A1(men_men_n118_), .B0(men_men_n552_), .Y(men_men_n1440_));
  OAI220     u1412(.A0(men_men_n1440_), .A1(men_men_n1437_), .B0(men_men_n1439_), .B1(men_men_n1438_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n790_), .B(men_men_n195_), .Y(men_men_n1442_));
  NOi31      u1414(.An(m), .B(n), .C(b), .Y(men_men_n1443_));
  NOi31      u1415(.An(f), .B(d), .C(c), .Y(men_men_n1444_));
  NA2        u1416(.A(men_men_n1444_), .B(men_men_n1443_), .Y(men_men_n1445_));
  INV        u1417(.A(men_men_n1445_), .Y(men_men_n1446_));
  NO3        u1418(.A(men_men_n1446_), .B(men_men_n1442_), .C(men_men_n1441_), .Y(men_men_n1447_));
  NA2        u1419(.A(men_men_n1130_), .B(men_men_n488_), .Y(men_men_n1448_));
  OAI210     u1420(.A0(men_men_n189_), .A1(men_men_n547_), .B0(men_men_n1106_), .Y(men_men_n1449_));
  AN3        u1421(.A(men_men_n1449_), .B(men_men_n1447_), .C(men_men_n1435_), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1401_), .B(men_men_n395_), .Y(men_men_n1451_));
  NO2        u1423(.A(men_men_n1451_), .B(men_men_n1087_), .Y(men_men_n1452_));
  NO2        u1424(.A(men_men_n195_), .B(b), .Y(men_men_n1453_));
  AOI220     u1425(.A0(men_men_n1213_), .A1(men_men_n1453_), .B0(men_men_n1137_), .B1(men_men_n1448_), .Y(men_men_n1454_));
  NO2        u1426(.A(i), .B(men_men_n222_), .Y(men_men_n1455_));
  NA4        u1427(.A(men_men_n1189_), .B(men_men_n1455_), .C(men_men_n105_), .D(m), .Y(men_men_n1456_));
  NAi31      u1428(.An(men_men_n1452_), .B(men_men_n1456_), .C(men_men_n1454_), .Y(men_men_n1457_));
  NO4        u1429(.A(men_men_n134_), .B(g), .C(f), .D(e), .Y(men_men_n1458_));
  NA2        u1430(.A(men_men_n301_), .B(h), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n202_), .B(men_men_n99_), .Y(men_men_n1460_));
  NA2        u1432(.A(men_men_n30_), .B(h), .Y(men_men_n1461_));
  NO2        u1433(.A(men_men_n1461_), .B(men_men_n1126_), .Y(men_men_n1462_));
  NOi41      u1434(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n1463_), .B(men_men_n115_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n1403_), .B(men_men_n1429_), .Y(men_men_n1465_));
  NA2        u1437(.A(men_men_n1465_), .B(men_men_n1464_), .Y(men_men_n1466_));
  OR3        u1438(.A(men_men_n563_), .B(men_men_n562_), .C(men_men_n114_), .Y(men_men_n1467_));
  NA2        u1439(.A(men_men_n1158_), .B(men_men_n424_), .Y(men_men_n1468_));
  OAI220     u1440(.A0(men_men_n1468_), .A1(men_men_n454_), .B0(men_men_n1467_), .B1(men_men_n310_), .Y(men_men_n1469_));
  AO210      u1441(.A0(men_men_n1469_), .A1(men_men_n118_), .B0(men_men_n1466_), .Y(men_men_n1470_));
  NO3        u1442(.A(men_men_n1470_), .B(men_men_n1462_), .C(men_men_n1457_), .Y(men_men_n1471_));
  NA4        u1443(.A(men_men_n1471_), .B(men_men_n1450_), .C(men_men_n1431_), .D(men_men_n1414_), .Y(men_men_n1472_));
  NO2        u1444(.A(men_men_n1174_), .B(men_men_n112_), .Y(men_men_n1473_));
  NA2        u1445(.A(men_men_n395_), .B(men_men_n56_), .Y(men_men_n1474_));
  AOI210     u1446(.A0(men_men_n1474_), .A1(men_men_n1096_), .B0(men_men_n1428_), .Y(men_men_n1475_));
  NA2        u1447(.A(men_men_n224_), .B(men_men_n186_), .Y(men_men_n1476_));
  AOI210     u1448(.A0(men_men_n1476_), .A1(men_men_n1232_), .B0(men_men_n1474_), .Y(men_men_n1477_));
  NO2        u1449(.A(men_men_n1131_), .B(men_men_n1126_), .Y(men_men_n1478_));
  NO3        u1450(.A(men_men_n1478_), .B(men_men_n1477_), .C(men_men_n1475_), .Y(men_men_n1479_));
  NO2        u1451(.A(men_men_n407_), .B(j), .Y(men_men_n1480_));
  NA3        u1452(.A(g), .B(men_men_n1480_), .C(men_men_n163_), .Y(men_men_n1481_));
  INV        u1453(.A(men_men_n1481_), .Y(men_men_n1482_));
  NO3        u1454(.A(men_men_n783_), .B(men_men_n181_), .C(men_men_n427_), .Y(men_men_n1483_));
  NO2        u1455(.A(men_men_n1483_), .B(men_men_n1482_), .Y(men_men_n1484_));
  NO3        u1456(.A(men_men_n1126_), .B(men_men_n608_), .C(g), .Y(men_men_n1485_));
  NOi21      u1457(.An(men_men_n1476_), .B(men_men_n1485_), .Y(men_men_n1486_));
  AOI210     u1458(.A0(men_men_n1486_), .A1(men_men_n1460_), .B0(men_men_n1096_), .Y(men_men_n1487_));
  INV        u1459(.A(men_men_n49_), .Y(men_men_n1488_));
  AOI220     u1460(.A0(men_men_n1488_), .A1(men_men_n1220_), .B0(men_men_n865_), .B1(men_men_n202_), .Y(men_men_n1489_));
  INV        u1461(.A(men_men_n1489_), .Y(men_men_n1490_));
  OAI220     u1462(.A0(men_men_n698_), .A1(g), .B0(men_men_n234_), .B1(c), .Y(men_men_n1491_));
  AOI210     u1463(.A0(men_men_n1453_), .A1(men_men_n41_), .B0(men_men_n1491_), .Y(men_men_n1492_));
  NO2        u1464(.A(men_men_n1492_), .B(men_men_n183_), .Y(men_men_n1493_));
  NO3        u1465(.A(men_men_n1467_), .B(men_men_n488_), .C(men_men_n366_), .Y(men_men_n1494_));
  NO4        u1466(.A(men_men_n1494_), .B(men_men_n1493_), .C(men_men_n1490_), .D(men_men_n1487_), .Y(men_men_n1495_));
  NA2        u1467(.A(men_men_n1141_), .B(men_men_n1587_), .Y(men_men_n1496_));
  NO2        u1468(.A(men_men_n1126_), .B(h), .Y(men_men_n1497_));
  NA3        u1469(.A(men_men_n1497_), .B(d), .C(men_men_n1088_), .Y(men_men_n1498_));
  OAI220     u1470(.A0(men_men_n1498_), .A1(c), .B0(men_men_n1496_), .B1(j), .Y(men_men_n1499_));
  NA3        u1471(.A(men_men_n1473_), .B(men_men_n488_), .C(f), .Y(men_men_n1500_));
  NO2        u1472(.A(men_men_n1396_), .B(men_men_n42_), .Y(men_men_n1501_));
  AOI210     u1473(.A0(men_men_n115_), .A1(men_men_n40_), .B0(men_men_n1501_), .Y(men_men_n1502_));
  NO2        u1474(.A(men_men_n1502_), .B(men_men_n1500_), .Y(men_men_n1503_));
  AOI210     u1475(.A0(men_men_n547_), .A1(h), .B0(men_men_n67_), .Y(men_men_n1504_));
  NA2        u1476(.A(men_men_n1504_), .B(men_men_n1434_), .Y(men_men_n1505_));
  NO2        u1477(.A(men_men_n1392_), .B(men_men_n181_), .Y(men_men_n1506_));
  NOi21      u1478(.An(d), .B(f), .Y(men_men_n1507_));
  NO3        u1479(.A(men_men_n1444_), .B(men_men_n1507_), .C(men_men_n40_), .Y(men_men_n1508_));
  NA2        u1480(.A(men_men_n1508_), .B(men_men_n1506_), .Y(men_men_n1509_));
  NA2        u1481(.A(men_men_n1434_), .B(men_men_n1501_), .Y(men_men_n1510_));
  NO2        u1482(.A(men_men_n310_), .B(c), .Y(men_men_n1511_));
  NA2        u1483(.A(men_men_n1511_), .B(men_men_n564_), .Y(men_men_n1512_));
  NA4        u1484(.A(men_men_n1512_), .B(men_men_n1510_), .C(men_men_n1509_), .D(men_men_n1505_), .Y(men_men_n1513_));
  NO3        u1485(.A(men_men_n1513_), .B(men_men_n1503_), .C(men_men_n1499_), .Y(men_men_n1514_));
  NA4        u1486(.A(men_men_n1514_), .B(men_men_n1495_), .C(men_men_n1484_), .D(men_men_n1479_), .Y(men_men_n1515_));
  NO3        u1487(.A(men_men_n1130_), .B(men_men_n1117_), .C(men_men_n40_), .Y(men_men_n1516_));
  NA2        u1488(.A(men_men_n1516_), .B(men_men_n1411_), .Y(men_men_n1517_));
  OAI210     u1489(.A0(men_men_n1458_), .A1(men_men_n1401_), .B0(men_men_n927_), .Y(men_men_n1518_));
  OAI220     u1490(.A0(men_men_n1084_), .A1(men_men_n134_), .B0(men_men_n698_), .B1(men_men_n181_), .Y(men_men_n1519_));
  NA2        u1491(.A(men_men_n1519_), .B(men_men_n650_), .Y(men_men_n1520_));
  NA3        u1492(.A(men_men_n1520_), .B(men_men_n1518_), .C(men_men_n1517_), .Y(men_men_n1521_));
  NA2        u1493(.A(men_men_n1433_), .B(men_men_n1507_), .Y(men_men_n1522_));
  NO2        u1494(.A(men_men_n1522_), .B(m), .Y(men_men_n1523_));
  NA3        u1495(.A(men_men_n1138_), .B(men_men_n110_), .C(men_men_n230_), .Y(men_men_n1524_));
  OAI220     u1496(.A0(men_men_n155_), .A1(men_men_n188_), .B0(men_men_n469_), .B1(g), .Y(men_men_n1525_));
  OAI210     u1497(.A0(men_men_n1525_), .A1(men_men_n112_), .B0(men_men_n1443_), .Y(men_men_n1526_));
  NA2        u1498(.A(men_men_n1526_), .B(men_men_n1524_), .Y(men_men_n1527_));
  NO3        u1499(.A(men_men_n1527_), .B(men_men_n1523_), .C(men_men_n1521_), .Y(men_men_n1528_));
  NO2        u1500(.A(men_men_n1400_), .B(e), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1169_), .B(men_men_n661_), .Y(men_men_n1530_));
  NO2        u1502(.A(men_men_n1530_), .B(men_men_n463_), .Y(men_men_n1531_));
  NO3        u1503(.A(men_men_n1467_), .B(men_men_n366_), .C(a), .Y(men_men_n1532_));
  NO2        u1504(.A(men_men_n1532_), .B(men_men_n1531_), .Y(men_men_n1533_));
  NO2        u1505(.A(men_men_n188_), .B(c), .Y(men_men_n1534_));
  OAI210     u1506(.A0(men_men_n1534_), .A1(men_men_n1529_), .B0(men_men_n186_), .Y(men_men_n1535_));
  AOI220     u1507(.A0(men_men_n1535_), .A1(men_men_n1119_), .B0(men_men_n554_), .B1(men_men_n382_), .Y(men_men_n1536_));
  NA2        u1508(.A(men_men_n562_), .B(g), .Y(men_men_n1537_));
  NA2        u1509(.A(men_men_n1537_), .B(men_men_n1430_), .Y(men_men_n1538_));
  NA2        u1510(.A(men_men_n1169_), .B(a), .Y(men_men_n1539_));
  OAI220     u1511(.A0(men_men_n1539_), .A1(men_men_n67_), .B0(men_men_n1538_), .B1(men_men_n222_), .Y(men_men_n1540_));
  AOI210     u1512(.A0(men_men_n946_), .A1(men_men_n434_), .B0(men_men_n106_), .Y(men_men_n1541_));
  OR2        u1513(.A(men_men_n1541_), .B(men_men_n562_), .Y(men_men_n1542_));
  NO2        u1514(.A(men_men_n1542_), .B(men_men_n181_), .Y(men_men_n1543_));
  NO2        u1515(.A(men_men_n49_), .B(l), .Y(men_men_n1544_));
  INV        u1516(.A(men_men_n506_), .Y(men_men_n1545_));
  NA2        u1517(.A(men_men_n1545_), .B(men_men_n1544_), .Y(men_men_n1546_));
  NO2        u1518(.A(men_men_n264_), .B(g), .Y(men_men_n1547_));
  NO2        u1519(.A(m), .B(i), .Y(men_men_n1548_));
  AOI220     u1520(.A0(men_men_n1548_), .A1(men_men_n1432_), .B0(men_men_n1118_), .B1(men_men_n1547_), .Y(men_men_n1549_));
  NA2        u1521(.A(men_men_n1549_), .B(men_men_n1546_), .Y(men_men_n1550_));
  NO4        u1522(.A(men_men_n1550_), .B(men_men_n1543_), .C(men_men_n1540_), .D(men_men_n1536_), .Y(men_men_n1551_));
  NA3        u1523(.A(men_men_n1551_), .B(men_men_n1533_), .C(men_men_n1528_), .Y(men_men_n1552_));
  NA3        u1524(.A(men_men_n1007_), .B(men_men_n141_), .C(men_men_n46_), .Y(men_men_n1553_));
  AOI210     u1525(.A0(men_men_n152_), .A1(c), .B0(men_men_n1553_), .Y(men_men_n1554_));
  OAI210     u1526(.A0(men_men_n608_), .A1(g), .B0(men_men_n192_), .Y(men_men_n1555_));
  NA2        u1527(.A(men_men_n1555_), .B(men_men_n1497_), .Y(men_men_n1556_));
  AO210      u1528(.A0(men_men_n135_), .A1(l), .B0(men_men_n1451_), .Y(men_men_n1557_));
  NO2        u1529(.A(men_men_n70_), .B(c), .Y(men_men_n1558_));
  NO4        u1530(.A(men_men_n1419_), .B(men_men_n193_), .C(men_men_n469_), .D(men_men_n45_), .Y(men_men_n1559_));
  AOI210     u1531(.A0(men_men_n1506_), .A1(men_men_n1558_), .B0(men_men_n1559_), .Y(men_men_n1560_));
  NA3        u1532(.A(men_men_n1560_), .B(men_men_n1557_), .C(men_men_n1556_), .Y(men_men_n1561_));
  NO2        u1533(.A(men_men_n1561_), .B(men_men_n1554_), .Y(men_men_n1562_));
  NO4        u1534(.A(men_men_n234_), .B(men_men_n193_), .C(men_men_n268_), .D(k), .Y(men_men_n1563_));
  NO2        u1535(.A(men_men_n1553_), .B(men_men_n112_), .Y(men_men_n1564_));
  NO2        u1536(.A(men_men_n1564_), .B(men_men_n1563_), .Y(men_men_n1565_));
  AN2        u1537(.A(men_men_n1138_), .B(men_men_n1124_), .Y(men_men_n1566_));
  AOI220     u1538(.A0(men_men_n1548_), .A1(men_men_n671_), .B0(men_men_n1102_), .B1(men_men_n164_), .Y(men_men_n1567_));
  NOi31      u1539(.An(men_men_n30_), .B(men_men_n1567_), .C(n), .Y(men_men_n1568_));
  AOI210     u1540(.A0(men_men_n1566_), .A1(men_men_n1213_), .B0(men_men_n1568_), .Y(men_men_n1569_));
  NO2        u1541(.A(men_men_n1500_), .B(men_men_n67_), .Y(men_men_n1570_));
  NA2        u1542(.A(men_men_n59_), .B(a), .Y(men_men_n1571_));
  NO2        u1543(.A(men_men_n1468_), .B(men_men_n1571_), .Y(men_men_n1572_));
  NO2        u1544(.A(men_men_n1572_), .B(men_men_n1570_), .Y(men_men_n1573_));
  NA4        u1545(.A(men_men_n1573_), .B(men_men_n1569_), .C(men_men_n1565_), .D(men_men_n1562_), .Y(men_men_n1574_));
  OR4        u1546(.A(men_men_n1574_), .B(men_men_n1552_), .C(men_men_n1515_), .D(men_men_n1472_), .Y(men04));
  NOi31      u1547(.An(men_men_n1458_), .B(men_men_n1459_), .C(men_men_n1090_), .Y(men_men_n1576_));
  NO4        u1548(.A(men_men_n284_), .B(men_men_n1080_), .C(men_men_n507_), .D(j), .Y(men_men_n1577_));
  OR3        u1549(.A(men_men_n1577_), .B(men_men_n1576_), .C(men_men_n1108_), .Y(men_men_n1578_));
  NO3        u1550(.A(men_men_n1408_), .B(men_men_n91_), .C(k), .Y(men_men_n1579_));
  AOI210     u1551(.A0(men_men_n1579_), .A1(men_men_n1101_), .B0(men_men_n1234_), .Y(men_men_n1580_));
  NA2        u1552(.A(men_men_n1580_), .B(men_men_n1264_), .Y(men_men_n1581_));
  NO4        u1553(.A(men_men_n1581_), .B(men_men_n1578_), .C(men_men_n1116_), .D(men_men_n1095_), .Y(men_men_n1582_));
  NA4        u1554(.A(men_men_n1582_), .B(men_men_n1171_), .C(men_men_n1156_), .D(men_men_n1143_), .Y(men05));
  INV        u1555(.A(i), .Y(men_men_n1586_));
  INV        u1556(.A(n), .Y(men_men_n1587_));
  INV        u1557(.A(men_men_n230_), .Y(men_men_n1588_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule