//Benchmark atmr_intb_466_0.5

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n246_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n286_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n339_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n409_, men_men_n410_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  INV        o004(.A(ori_ori_n26_), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  INV        o017(.A(x05), .Y(ori_ori_n40_));
  NO2        o018(.A(x09), .B(x02), .Y(ori_ori_n41_));
  NO2        o019(.A(ori_ori_n39_), .B(ori_ori_n34_), .Y(ori00));
  INV        o020(.A(x01), .Y(ori_ori_n43_));
  INV        o021(.A(x06), .Y(ori_ori_n44_));
  NA2        o022(.A(ori_ori_n44_), .B(ori_ori_n28_), .Y(ori_ori_n45_));
  INV        o023(.A(x09), .Y(ori_ori_n46_));
  NO2        o024(.A(x10), .B(x02), .Y(ori_ori_n47_));
  NOi21      o025(.An(x01), .B(x09), .Y(ori_ori_n48_));
  INV        o026(.A(x00), .Y(ori_ori_n49_));
  NO2        o027(.A(ori_ori_n46_), .B(ori_ori_n49_), .Y(ori_ori_n50_));
  NO2        o028(.A(ori_ori_n50_), .B(ori_ori_n48_), .Y(ori_ori_n51_));
  NA2        o029(.A(x09), .B(ori_ori_n49_), .Y(ori_ori_n52_));
  INV        o030(.A(x07), .Y(ori_ori_n53_));
  INV        o031(.A(ori_ori_n51_), .Y(ori_ori_n54_));
  NA2        o032(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n55_), .B(ori_ori_n24_), .Y(ori_ori_n56_));
  NO2        o034(.A(ori_ori_n56_), .B(ori_ori_n54_), .Y(ori_ori_n57_));
  NA2        o035(.A(ori_ori_n53_), .B(ori_ori_n44_), .Y(ori_ori_n58_));
  OAI210     o036(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n58_), .Y(ori_ori_n59_));
  AOI220     o037(.A0(ori_ori_n59_), .A1(ori_ori_n51_), .B0(ori_ori_n57_), .B1(ori_ori_n31_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n61_));
  NO2        o039(.A(ori_ori_n53_), .B(ori_ori_n23_), .Y(ori_ori_n62_));
  NA2        o040(.A(x09), .B(x05), .Y(ori_ori_n63_));
  NA2        o041(.A(x10), .B(x06), .Y(ori_ori_n64_));
  INV        o042(.A(ori_ori_n64_), .Y(ori_ori_n65_));
  OAI210     o043(.A0(ori_ori_n65_), .A1(ori_ori_n62_), .B0(x03), .Y(ori_ori_n66_));
  NOi31      o044(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n67_));
  INV        o045(.A(x07), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n68_), .B(ori_ori_n24_), .Y(ori_ori_n69_));
  NO2        o047(.A(x09), .B(ori_ori_n40_), .Y(ori_ori_n70_));
  INV        o048(.A(ori_ori_n70_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n70_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n72_));
  AOI210     o050(.A0(ori_ori_n71_), .A1(ori_ori_n44_), .B0(ori_ori_n72_), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n74_));
  NO2        o052(.A(x08), .B(x01), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n35_), .Y(ori_ori_n76_));
  NO3        o054(.A(ori_ori_n76_), .B(ori_ori_n73_), .C(ori_ori_n69_), .Y(ori_ori_n77_));
  AN2        o055(.A(ori_ori_n77_), .B(ori_ori_n66_), .Y(ori_ori_n78_));
  INV        o056(.A(ori_ori_n76_), .Y(ori_ori_n79_));
  NA2        o057(.A(x11), .B(x00), .Y(ori_ori_n80_));
  NO2        o058(.A(x11), .B(ori_ori_n43_), .Y(ori_ori_n81_));
  NOi21      o059(.An(ori_ori_n80_), .B(ori_ori_n81_), .Y(ori_ori_n82_));
  INV        o060(.A(ori_ori_n82_), .Y(ori_ori_n83_));
  NOi21      o061(.An(x01), .B(x10), .Y(ori_ori_n84_));
  NO2        o062(.A(ori_ori_n29_), .B(ori_ori_n49_), .Y(ori_ori_n85_));
  NO2        o063(.A(ori_ori_n83_), .B(x07), .Y(ori_ori_n86_));
  NO3        o064(.A(ori_ori_n86_), .B(ori_ori_n78_), .C(ori_ori_n61_), .Y(ori01));
  INV        o065(.A(x12), .Y(ori_ori_n88_));
  INV        o066(.A(x13), .Y(ori_ori_n89_));
  NO2        o067(.A(x10), .B(x01), .Y(ori_ori_n90_));
  NO2        o068(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n91_));
  NO2        o069(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n48_), .B(x05), .Y(ori_ori_n93_));
  NOi21      o071(.An(ori_ori_n93_), .B(ori_ori_n50_), .Y(ori_ori_n94_));
  NA2        o072(.A(ori_ori_n29_), .B(ori_ori_n43_), .Y(ori_ori_n95_));
  NA2        o073(.A(x10), .B(ori_ori_n49_), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n96_), .B(ori_ori_n95_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n46_), .B(x05), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n99_));
  NO3        o077(.A(ori_ori_n95_), .B(x06), .C(x03), .Y(ori_ori_n100_));
  INV        o078(.A(ori_ori_n100_), .Y(ori_ori_n101_));
  OAI210     o079(.A0(ori_ori_n75_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n102_), .B(ori_ori_n267_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n46_), .B(ori_ori_n40_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n105_));
  AOI210     o083(.A0(ori_ori_n105_), .A1(ori_ori_n45_), .B0(ori_ori_n104_), .Y(ori_ori_n106_));
  NO2        o084(.A(x09), .B(x05), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n107_), .B(ori_ori_n43_), .Y(ori_ori_n108_));
  NA2        o086(.A(x09), .B(x00), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n93_), .B(ori_ori_n109_), .Y(ori_ori_n110_));
  NO2        o088(.A(x03), .B(x02), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n76_), .B(ori_ori_n89_), .Y(ori_ori_n112_));
  OAI210     o090(.A0(ori_ori_n112_), .A1(ori_ori_n94_), .B0(ori_ori_n111_), .Y(ori_ori_n113_));
  OA210      o091(.A0(ori_ori_n268_), .A1(x11), .B0(ori_ori_n113_), .Y(ori_ori_n114_));
  OAI210     o092(.A0(ori_ori_n101_), .A1(ori_ori_n23_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  INV        o093(.A(ori_ori_n92_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n40_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n89_), .B(x01), .Y(ori_ori_n119_));
  AOI210     o097(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n117_), .B(ori_ori_n120_), .Y(ori_ori_n121_));
  NA2        o099(.A(x04), .B(x02), .Y(ori_ori_n122_));
  NA2        o100(.A(x10), .B(x05), .Y(ori_ori_n123_));
  NO2        o101(.A(x09), .B(x01), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n93_), .B(x08), .Y(ori_ori_n125_));
  NO2        o103(.A(ori_ori_n85_), .B(x06), .Y(ori_ori_n126_));
  NOi21      o104(.An(x09), .B(x00), .Y(ori_ori_n127_));
  NO3        o105(.A(ori_ori_n74_), .B(ori_ori_n127_), .C(ori_ori_n43_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n96_), .Y(ori_ori_n129_));
  NA2        o107(.A(x06), .B(x05), .Y(ori_ori_n130_));
  OAI210     o108(.A0(ori_ori_n130_), .A1(ori_ori_n35_), .B0(ori_ori_n88_), .Y(ori_ori_n131_));
  AOI210     o109(.A0(x10), .A1(ori_ori_n50_), .B0(ori_ori_n131_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n129_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n89_), .B(x12), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n135_), .B(ori_ori_n133_), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n137_), .B(ori_ori_n121_), .Y(ori_ori_n138_));
  AOI210     o116(.A0(ori_ori_n115_), .A1(ori_ori_n88_), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n28_), .B(ori_ori_n103_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n46_), .B(ori_ori_n43_), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n140_), .B(x12), .Y(ori_ori_n142_));
  NO2        o120(.A(ori_ori_n84_), .B(x06), .Y(ori_ori_n143_));
  AOI210     o121(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n46_), .Y(ori_ori_n144_));
  NO3        o122(.A(ori_ori_n144_), .B(ori_ori_n143_), .C(ori_ori_n40_), .Y(ori_ori_n145_));
  INV        o123(.A(ori_ori_n105_), .Y(ori_ori_n146_));
  OAI210     o124(.A0(ori_ori_n146_), .A1(ori_ori_n145_), .B0(x02), .Y(ori_ori_n147_));
  AOI210     o125(.A0(ori_ori_n147_), .A1(ori_ori_n49_), .B0(ori_ori_n23_), .Y(ori_ori_n148_));
  OAI210     o126(.A0(ori_ori_n142_), .A1(ori_ori_n49_), .B0(ori_ori_n148_), .Y(ori_ori_n149_));
  INV        o127(.A(ori_ori_n105_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n46_), .B(x03), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n152_));
  NOi21      o130(.An(x13), .B(x04), .Y(ori_ori_n153_));
  NO3        o131(.A(ori_ori_n153_), .B(ori_ori_n67_), .C(ori_ori_n127_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n154_), .B(x05), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n155_), .B(ori_ori_n152_), .Y(ori_ori_n156_));
  INV        o134(.A(ori_ori_n156_), .Y(ori_ori_n157_));
  INV        o135(.A(ori_ori_n81_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n158_), .B(x12), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n23_), .B(ori_ori_n43_), .Y(ori_ori_n160_));
  INV        o138(.A(x00), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n29_), .B(ori_ori_n44_), .Y(ori_ori_n162_));
  NA2        o140(.A(x13), .B(ori_ori_n88_), .Y(ori_ori_n163_));
  NA3        o141(.A(ori_ori_n163_), .B(ori_ori_n131_), .C(ori_ori_n82_), .Y(ori_ori_n164_));
  INV        o142(.A(ori_ori_n164_), .Y(ori_ori_n165_));
  AOI210     o143(.A0(ori_ori_n159_), .A1(ori_ori_n157_), .B0(ori_ori_n165_), .Y(ori_ori_n166_));
  AOI210     o144(.A0(ori_ori_n166_), .A1(ori_ori_n149_), .B0(x07), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n63_), .B(ori_ori_n29_), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n168_), .Y(ori_ori_n169_));
  NO2        o147(.A(x12), .B(x02), .Y(ori_ori_n170_));
  INV        o148(.A(ori_ori_n170_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n171_), .B(ori_ori_n158_), .Y(ori_ori_n172_));
  OA210      o150(.A0(ori_ori_n67_), .A1(ori_ori_n169_), .B0(ori_ori_n172_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n46_), .B(ori_ori_n40_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n174_), .B(x01), .Y(ori_ori_n175_));
  NO3        o153(.A(ori_ori_n80_), .B(x12), .C(x03), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n175_), .B(ori_ori_n176_), .Y(ori_ori_n177_));
  NOi21      o155(.An(ori_ori_n168_), .B(ori_ori_n143_), .Y(ori_ori_n178_));
  INV        o156(.A(ori_ori_n25_), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n178_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n181_));
  NO3        o159(.A(ori_ori_n181_), .B(ori_ori_n144_), .C(ori_ori_n126_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n160_), .B(ori_ori_n28_), .Y(ori_ori_n183_));
  OAI210     o161(.A0(ori_ori_n182_), .A1(ori_ori_n150_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  NA3        o162(.A(ori_ori_n184_), .B(ori_ori_n180_), .C(ori_ori_n177_), .Y(ori_ori_n185_));
  NO3        o163(.A(ori_ori_n185_), .B(ori_ori_n173_), .C(ori_ori_n167_), .Y(ori_ori_n186_));
  OAI210     o164(.A0(ori_ori_n139_), .A1(ori_ori_n53_), .B0(ori_ori_n186_), .Y(ori02));
  INV        o165(.A(ori_ori_n98_), .Y(ori_ori_n188_));
  NOi21      o166(.An(ori_ori_n154_), .B(ori_ori_n124_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n189_), .B(ori_ori_n32_), .Y(ori_ori_n190_));
  OAI210     o168(.A0(ori_ori_n190_), .A1(ori_ori_n188_), .B0(ori_ori_n123_), .Y(ori_ori_n191_));
  INV        o169(.A(ori_ori_n123_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n76_), .B(ori_ori_n46_), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  AOI210     o172(.A0(ori_ori_n194_), .A1(ori_ori_n191_), .B0(ori_ori_n44_), .Y(ori_ori_n195_));
  NO2        o173(.A(x05), .B(x02), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n196_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n197_), .B(ori_ori_n105_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n162_), .B(ori_ori_n43_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n199_), .B(ori_ori_n155_), .Y(ori_ori_n200_));
  BUFFER     o178(.A(ori_ori_n108_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(x06), .Y(ori_ori_n202_));
  NA2        o180(.A(ori_ori_n202_), .B(ori_ori_n85_), .Y(ori_ori_n203_));
  INV        o181(.A(ori_ori_n111_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(ori_ori_n97_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n205_), .B(x13), .Y(ori_ori_n206_));
  NA3        o184(.A(ori_ori_n206_), .B(ori_ori_n203_), .C(ori_ori_n200_), .Y(ori_ori_n207_));
  NO3        o185(.A(ori_ori_n207_), .B(ori_ori_n198_), .C(ori_ori_n195_), .Y(ori_ori_n208_));
  INV        o186(.A(x03), .Y(ori_ori_n209_));
  NA2        o187(.A(x08), .B(ori_ori_n90_), .Y(ori_ori_n210_));
  NA2        o188(.A(ori_ori_n122_), .B(ori_ori_n119_), .Y(ori_ori_n211_));
  AN2        o189(.A(ori_ori_n211_), .B(ori_ori_n125_), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n212_), .B(ori_ori_n91_), .Y(ori_ori_n213_));
  NA3        o191(.A(ori_ori_n213_), .B(ori_ori_n210_), .C(ori_ori_n44_), .Y(ori_ori_n214_));
  INV        o192(.A(ori_ori_n136_), .Y(ori_ori_n215_));
  INV        o193(.A(x05), .Y(ori_ori_n216_));
  OAI220     o194(.A0(ori_ori_n216_), .A1(ori_ori_n31_), .B0(ori_ori_n215_), .B1(ori_ori_n51_), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n217_), .B(x02), .Y(ori_ori_n218_));
  NO3        o196(.A(ori_ori_n134_), .B(ori_ori_n118_), .C(ori_ori_n47_), .Y(ori_ori_n219_));
  OAI210     o197(.A0(ori_ori_n109_), .A1(ori_ori_n36_), .B0(ori_ori_n88_), .Y(ori_ori_n220_));
  OAI210     o198(.A0(ori_ori_n220_), .A1(ori_ori_n128_), .B0(ori_ori_n219_), .Y(ori_ori_n221_));
  NA3        o199(.A(ori_ori_n221_), .B(ori_ori_n218_), .C(x06), .Y(ori_ori_n222_));
  NA2        o200(.A(x09), .B(x03), .Y(ori_ori_n223_));
  OAI220     o201(.A0(ori_ori_n223_), .A1(ori_ori_n96_), .B0(ori_ori_n141_), .B1(ori_ori_n55_), .Y(ori_ori_n224_));
  NO3        o202(.A(ori_ori_n181_), .B(ori_ori_n95_), .C(x08), .Y(ori_ori_n225_));
  INV        o203(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n44_), .B(ori_ori_n40_), .Y(ori_ori_n227_));
  NO3        o205(.A(ori_ori_n93_), .B(ori_ori_n96_), .C(ori_ori_n38_), .Y(ori_ori_n228_));
  AOI210     o206(.A0(ori_ori_n219_), .A1(ori_ori_n227_), .B0(ori_ori_n228_), .Y(ori_ori_n229_));
  OAI210     o207(.A0(ori_ori_n226_), .A1(ori_ori_n28_), .B0(ori_ori_n229_), .Y(ori_ori_n230_));
  AO220      o208(.A0(ori_ori_n230_), .A1(x04), .B0(ori_ori_n224_), .B1(x05), .Y(ori_ori_n231_));
  AOI210     o209(.A0(ori_ori_n222_), .A1(ori_ori_n214_), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  OAI210     o210(.A0(ori_ori_n208_), .A1(x12), .B0(ori_ori_n232_), .Y(ori03));
  OR2        o211(.A(ori_ori_n41_), .B(ori_ori_n151_), .Y(ori_ori_n234_));
  AOI210     o212(.A0(ori_ori_n112_), .A1(ori_ori_n88_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n134_), .B(ori_ori_n111_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  OAI210     o215(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(x05), .Y(ori_ori_n238_));
  AOI210     o216(.A0(ori_ori_n108_), .A1(ori_ori_n52_), .B0(ori_ori_n38_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n124_), .B(ori_ori_n99_), .Y(ori_ori_n240_));
  OAI220     o218(.A0(ori_ori_n240_), .A1(ori_ori_n37_), .B0(ori_ori_n110_), .B1(x13), .Y(ori_ori_n241_));
  OAI210     o219(.A0(ori_ori_n241_), .A1(ori_ori_n239_), .B0(x04), .Y(ori_ori_n242_));
  NO3        o220(.A(x05), .B(ori_ori_n76_), .C(ori_ori_n51_), .Y(ori_ori_n243_));
  INV        o221(.A(ori_ori_n243_), .Y(ori_ori_n244_));
  NA3        o222(.A(ori_ori_n244_), .B(ori_ori_n242_), .C(ori_ori_n238_), .Y(ori04));
  NO2        o223(.A(ori_ori_n79_), .B(ori_ori_n39_), .Y(ori_ori_n246_));
  XO2        o224(.A(ori_ori_n246_), .B(ori_ori_n163_), .Y(ori05));
  NA2        o225(.A(ori_ori_n161_), .B(ori_ori_n158_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n33_), .B(ori_ori_n88_), .Y(ori_ori_n249_));
  AOI210     o227(.A0(ori_ori_n249_), .A1(ori_ori_n81_), .B0(x07), .Y(ori_ori_n250_));
  AOI210     o228(.A0(ori_ori_n250_), .A1(ori_ori_n248_), .B0(x07), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n43_), .B(x04), .Y(ori_ori_n252_));
  NO4        o230(.A(ori_ori_n252_), .B(ori_ori_n269_), .C(ori_ori_n134_), .D(x08), .Y(ori_ori_n253_));
  BUFFER     o231(.A(ori_ori_n163_), .Y(ori_ori_n254_));
  NA4        o232(.A(ori_ori_n254_), .B(x04), .C(x03), .D(x08), .Y(ori_ori_n255_));
  INV        o233(.A(ori_ori_n255_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n253_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  NA2        o235(.A(x09), .B(ori_ori_n209_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n119_), .B(x07), .C(ori_ori_n49_), .Y(ori_ori_n259_));
  INV        o237(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n260_), .B(ori_ori_n258_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n249_), .B(ori_ori_n53_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n262_), .B(x05), .Y(ori_ori_n263_));
  NO4        o241(.A(ori_ori_n263_), .B(ori_ori_n261_), .C(ori_ori_n257_), .D(ori_ori_n251_), .Y(ori06));
  INV        o242(.A(x13), .Y(ori_ori_n267_));
  INV        o243(.A(ori_ori_n106_), .Y(ori_ori_n268_));
  INV        o244(.A(x02), .Y(ori_ori_n269_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NO2        m030(.A(x09), .B(x07), .Y(mai_mai_n53_));
  OAI210     m031(.A0(mai_mai_n53_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n54_));
  NOi21      m032(.An(x01), .B(x09), .Y(mai_mai_n55_));
  INV        m033(.A(x00), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n51_), .B(mai_mai_n56_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(x09), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m037(.A(x07), .Y(mai_mai_n60_));
  AOI220     m038(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n60_), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n58_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n63_), .B(mai_mai_n24_), .Y(mai_mai_n64_));
  OAI220     m042(.A0(mai_mai_n64_), .A1(mai_mai_n62_), .B0(mai_mai_n61_), .B1(mai_mai_n59_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n65_), .B(mai_mai_n31_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(mai_mai_n66_), .A1(mai_mai_n54_), .B0(x05), .Y(mai_mai_n67_));
  NA2        m045(.A(x09), .B(x05), .Y(mai_mai_n68_));
  NA2        m046(.A(x10), .B(x06), .Y(mai_mai_n69_));
  NO2        m047(.A(mai_mai_n60_), .B(mai_mai_n41_), .Y(mai_mai_n70_));
  NOi31      m048(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n71_));
  NO2        m049(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n72_));
  OAI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n74_));
  NO2        m052(.A(x08), .B(x01), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n35_), .Y(mai_mai_n76_));
  INV        m054(.A(mai_mai_n76_), .Y(mai_mai_n77_));
  NO2        m055(.A(x06), .B(x05), .Y(mai_mai_n78_));
  NA2        m056(.A(x11), .B(x00), .Y(mai_mai_n79_));
  NO2        m057(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n80_));
  NOi21      m058(.An(mai_mai_n79_), .B(mai_mai_n80_), .Y(mai_mai_n81_));
  AOI210     m059(.A0(mai_mai_n78_), .A1(mai_mai_n77_), .B0(mai_mai_n81_), .Y(mai_mai_n82_));
  NOi21      m060(.An(x01), .B(x10), .Y(mai_mai_n83_));
  NO2        m061(.A(mai_mai_n29_), .B(mai_mai_n56_), .Y(mai_mai_n84_));
  NO3        m062(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(x06), .Y(mai_mai_n85_));
  NA2        m063(.A(mai_mai_n85_), .B(mai_mai_n27_), .Y(mai_mai_n86_));
  OAI210     m064(.A0(mai_mai_n82_), .A1(x07), .B0(mai_mai_n86_), .Y(mai_mai_n87_));
  NO2        m065(.A(mai_mai_n87_), .B(mai_mai_n67_), .Y(mai01));
  INV        m066(.A(x12), .Y(mai_mai_n89_));
  INV        m067(.A(x13), .Y(mai_mai_n90_));
  NA2        m068(.A(x08), .B(x04), .Y(mai_mai_n91_));
  NA2        m069(.A(mai_mai_n83_), .B(mai_mai_n28_), .Y(mai_mai_n92_));
  NO2        m070(.A(x10), .B(x01), .Y(mai_mai_n93_));
  NO2        m071(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n95_));
  NO3        m073(.A(mai_mai_n342_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n96_));
  NO2        m074(.A(mai_mai_n55_), .B(x05), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n98_));
  NA3        m076(.A(x08), .B(mai_mai_n98_), .C(x06), .Y(mai_mai_n99_));
  INV        m077(.A(mai_mai_n99_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n75_), .B(x13), .Y(mai_mai_n101_));
  AOI210     m079(.A0(x00), .A1(mai_mai_n101_), .B0(mai_mai_n69_), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n103_));
  NA2        m081(.A(x10), .B(mai_mai_n56_), .Y(mai_mai_n104_));
  NA2        m082(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n106_));
  INV        m084(.A(x13), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n59_), .B(x05), .Y(mai_mai_n108_));
  NO3        m086(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n109_));
  NO4        m087(.A(mai_mai_n109_), .B(mai_mai_n102_), .C(mai_mai_n100_), .D(mai_mai_n96_), .Y(mai_mai_n110_));
  OAI210     m088(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n112_));
  NA2        m090(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n113_));
  NO2        m091(.A(x09), .B(x05), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n114_), .B(mai_mai_n47_), .Y(mai_mai_n115_));
  AOI210     m093(.A0(mai_mai_n115_), .A1(mai_mai_n95_), .B0(mai_mai_n49_), .Y(mai_mai_n116_));
  NA2        m094(.A(x09), .B(x00), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n97_), .B(mai_mai_n117_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n71_), .B(mai_mai_n51_), .Y(mai_mai_n119_));
  AOI210     m097(.A0(mai_mai_n119_), .A1(mai_mai_n118_), .B0(mai_mai_n113_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(mai_mai_n116_), .Y(mai_mai_n121_));
  NO2        m099(.A(x03), .B(x02), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n76_), .B(mai_mai_n90_), .Y(mai_mai_n123_));
  OR2        m101(.A(mai_mai_n121_), .B(x11), .Y(mai_mai_n124_));
  OAI210     m102(.A0(mai_mai_n110_), .A1(mai_mai_n23_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n95_), .B(mai_mai_n40_), .Y(mai_mai_n126_));
  NAi21      m104(.An(x06), .B(x10), .Y(mai_mai_n127_));
  NOi21      m105(.An(x01), .B(x13), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n129_));
  OR2        m107(.A(mai_mai_n129_), .B(x08), .Y(mai_mai_n130_));
  AOI210     m108(.A0(mai_mai_n130_), .A1(mai_mai_n126_), .B0(mai_mai_n41_), .Y(mai_mai_n131_));
  NO2        m109(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n90_), .B(x01), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n133_), .B(x08), .Y(mai_mai_n134_));
  OAI210     m112(.A0(x05), .A1(mai_mai_n134_), .B0(mai_mai_n51_), .Y(mai_mai_n135_));
  AOI210     m113(.A0(mai_mai_n135_), .A1(mai_mai_n132_), .B0(mai_mai_n48_), .Y(mai_mai_n136_));
  AOI210     m114(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n137_));
  OAI210     m115(.A0(mai_mai_n136_), .A1(mai_mai_n131_), .B0(mai_mai_n137_), .Y(mai_mai_n138_));
  NA2        m116(.A(x04), .B(x02), .Y(mai_mai_n139_));
  NA2        m117(.A(x10), .B(x05), .Y(mai_mai_n140_));
  NO2        m118(.A(mai_mai_n97_), .B(x08), .Y(mai_mai_n141_));
  AOI210     m119(.A0(mai_mai_n141_), .A1(x06), .B0(mai_mai_n128_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n142_), .B(x11), .Y(mai_mai_n143_));
  NAi21      m121(.An(mai_mai_n139_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  INV        m122(.A(mai_mai_n25_), .Y(mai_mai_n145_));
  NAi21      m123(.An(x13), .B(x00), .Y(mai_mai_n146_));
  AOI210     m124(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n146_), .Y(mai_mai_n147_));
  AN2        m125(.A(x04), .B(mai_mai_n147_), .Y(mai_mai_n148_));
  BUFFER     m126(.A(mai_mai_n68_), .Y(mai_mai_n149_));
  NO2        m127(.A(mai_mai_n146_), .B(mai_mai_n36_), .Y(mai_mai_n150_));
  INV        m128(.A(mai_mai_n150_), .Y(mai_mai_n151_));
  OAI210     m129(.A0(mai_mai_n56_), .A1(mai_mai_n149_), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  OAI210     m130(.A0(mai_mai_n152_), .A1(mai_mai_n148_), .B0(mai_mai_n145_), .Y(mai_mai_n153_));
  NOi21      m131(.An(x09), .B(x00), .Y(mai_mai_n154_));
  NA2        m132(.A(x06), .B(x05), .Y(mai_mai_n155_));
  NO2        m133(.A(mai_mai_n90_), .B(x12), .Y(mai_mai_n156_));
  NA2        m134(.A(mai_mai_n83_), .B(mai_mai_n51_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(x02), .Y(mai_mai_n159_));
  NO2        m137(.A(mai_mai_n159_), .B(mai_mai_n157_), .Y(mai_mai_n160_));
  INV        m138(.A(mai_mai_n160_), .Y(mai_mai_n161_));
  NA4        m139(.A(mai_mai_n161_), .B(mai_mai_n153_), .C(mai_mai_n144_), .D(mai_mai_n138_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n125_), .A1(mai_mai_n89_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  NA2        m141(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n164_));
  NA2        m142(.A(mai_mai_n164_), .B(mai_mai_n111_), .Y(mai_mai_n165_));
  AOI210     m143(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n103_), .B(x06), .Y(mai_mai_n167_));
  AOI210     m145(.A0(mai_mai_n166_), .A1(mai_mai_n165_), .B0(mai_mai_n167_), .Y(mai_mai_n168_));
  NO2        m146(.A(mai_mai_n168_), .B(x12), .Y(mai_mai_n169_));
  INV        m147(.A(mai_mai_n71_), .Y(mai_mai_n170_));
  NA2        m148(.A(mai_mai_n129_), .B(mai_mai_n56_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NA4        m150(.A(mai_mai_n127_), .B(mai_mai_n55_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(mai_mai_n113_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n174_), .B(x02), .Y(mai_mai_n175_));
  AOI210     m153(.A0(mai_mai_n175_), .A1(mai_mai_n172_), .B0(mai_mai_n23_), .Y(mai_mai_n176_));
  OAI210     m154(.A0(mai_mai_n169_), .A1(mai_mai_n56_), .B0(mai_mai_n176_), .Y(mai_mai_n177_));
  INV        m155(.A(mai_mai_n113_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n90_), .B(x03), .Y(mai_mai_n179_));
  AOI210     m157(.A0(mai_mai_n71_), .A1(mai_mai_n346_), .B0(mai_mai_n179_), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n181_));
  INV        m159(.A(mai_mai_n127_), .Y(mai_mai_n182_));
  NOi21      m160(.An(x13), .B(x04), .Y(mai_mai_n183_));
  NO3        m161(.A(mai_mai_n183_), .B(mai_mai_n71_), .C(mai_mai_n154_), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n184_), .B(x05), .Y(mai_mai_n185_));
  AOI220     m163(.A0(mai_mai_n185_), .A1(mai_mai_n181_), .B0(mai_mai_n182_), .B1(mai_mai_n56_), .Y(mai_mai_n186_));
  OAI210     m164(.A0(mai_mai_n180_), .A1(mai_mai_n178_), .B0(mai_mai_n186_), .Y(mai_mai_n187_));
  INV        m165(.A(mai_mai_n80_), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n188_), .B(x12), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n190_));
  INV        m168(.A(mai_mai_n147_), .Y(mai_mai_n191_));
  AOI210     m169(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n192_));
  NO2        m170(.A(x06), .B(x00), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(x03), .Y(mai_mai_n195_));
  OA210      m173(.A0(mai_mai_n195_), .A1(mai_mai_n193_), .B0(mai_mai_n191_), .Y(mai_mai_n196_));
  NA2        m174(.A(x13), .B(mai_mai_n89_), .Y(mai_mai_n197_));
  NA2        m175(.A(x12), .B(mai_mai_n81_), .Y(mai_mai_n198_));
  OAI210     m176(.A0(mai_mai_n196_), .A1(mai_mai_n190_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  AOI210     m177(.A0(mai_mai_n189_), .A1(mai_mai_n187_), .B0(mai_mai_n199_), .Y(mai_mai_n200_));
  AOI210     m178(.A0(mai_mai_n200_), .A1(mai_mai_n177_), .B0(x07), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n68_), .B(mai_mai_n29_), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n183_), .B(mai_mai_n154_), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n203_), .A1(mai_mai_n119_), .B0(mai_mai_n202_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n90_), .B(x06), .Y(mai_mai_n205_));
  INV        m183(.A(mai_mai_n205_), .Y(mai_mai_n206_));
  NO2        m184(.A(x08), .B(x05), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n207_), .B(mai_mai_n192_), .Y(mai_mai_n208_));
  NA2        m186(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n209_));
  OAI210     m187(.A0(mai_mai_n208_), .A1(mai_mai_n206_), .B0(mai_mai_n209_), .Y(mai_mai_n210_));
  NO2        m188(.A(x12), .B(x02), .Y(mai_mai_n211_));
  INV        m189(.A(mai_mai_n211_), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n212_), .B(mai_mai_n188_), .Y(mai_mai_n213_));
  OA210      m191(.A0(mai_mai_n210_), .A1(mai_mai_n204_), .B0(mai_mai_n213_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n215_), .B(x01), .Y(mai_mai_n216_));
  BUFFER     m194(.A(mai_mai_n75_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  AOI210     m196(.A0(mai_mai_n218_), .A1(mai_mai_n107_), .B0(mai_mai_n29_), .Y(mai_mai_n219_));
  INV        m197(.A(mai_mai_n205_), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n90_), .B(x04), .Y(mai_mai_n221_));
  OAI210     m199(.A0(x02), .A1(mai_mai_n101_), .B0(mai_mai_n220_), .Y(mai_mai_n222_));
  NO3        m200(.A(mai_mai_n79_), .B(x12), .C(x03), .Y(mai_mai_n223_));
  OAI210     m201(.A0(mai_mai_n222_), .A1(mai_mai_n219_), .B0(mai_mai_n223_), .Y(mai_mai_n224_));
  AOI210     m202(.A0(mai_mai_n157_), .A1(mai_mai_n155_), .B0(mai_mai_n91_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n225_), .B(mai_mai_n226_), .Y(mai_mai_n227_));
  NA2        m205(.A(mai_mai_n227_), .B(mai_mai_n224_), .Y(mai_mai_n228_));
  NO3        m206(.A(mai_mai_n228_), .B(mai_mai_n214_), .C(mai_mai_n201_), .Y(mai_mai_n229_));
  OAI210     m207(.A0(mai_mai_n163_), .A1(mai_mai_n60_), .B0(mai_mai_n229_), .Y(mai02));
  NO2        m208(.A(mai_mai_n90_), .B(mai_mai_n35_), .Y(mai_mai_n231_));
  INV        m209(.A(mai_mai_n140_), .Y(mai_mai_n232_));
  AOI220     m210(.A0(x13), .A1(mai_mai_n232_), .B0(mai_mai_n123_), .B1(mai_mai_n122_), .Y(mai_mai_n233_));
  AOI210     m211(.A0(mai_mai_n233_), .A1(mai_mai_n32_), .B0(mai_mai_n48_), .Y(mai_mai_n234_));
  NO2        m212(.A(x05), .B(x02), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n165_), .B(mai_mai_n235_), .Y(mai_mai_n236_));
  AOI220     m214(.A0(mai_mai_n207_), .A1(mai_mai_n57_), .B0(mai_mai_n55_), .B1(mai_mai_n36_), .Y(mai_mai_n237_));
  NOi21      m215(.An(mai_mai_n231_), .B(mai_mai_n237_), .Y(mai_mai_n238_));
  AOI210     m216(.A0(mai_mai_n183_), .A1(mai_mai_n72_), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  AOI210     m217(.A0(mai_mai_n239_), .A1(mai_mai_n236_), .B0(mai_mai_n113_), .Y(mai_mai_n240_));
  NO2        m218(.A(mai_mai_n194_), .B(mai_mai_n47_), .Y(mai_mai_n241_));
  OAI210     m219(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n242_));
  INV        m220(.A(mai_mai_n242_), .Y(mai_mai_n243_));
  OAI210     m221(.A0(mai_mai_n243_), .A1(mai_mai_n179_), .B0(mai_mai_n84_), .Y(mai_mai_n244_));
  NA2        m222(.A(mai_mai_n84_), .B(mai_mai_n75_), .Y(mai_mai_n245_));
  NA3        m223(.A(mai_mai_n83_), .B(mai_mai_n74_), .C(mai_mai_n42_), .Y(mai_mai_n246_));
  AOI210     m224(.A0(mai_mai_n246_), .A1(mai_mai_n245_), .B0(x04), .Y(mai_mai_n247_));
  INV        m225(.A(mai_mai_n247_), .Y(mai_mai_n248_));
  NA3        m226(.A(mai_mai_n248_), .B(mai_mai_n244_), .C(mai_mai_n343_), .Y(mai_mai_n249_));
  NO3        m227(.A(mai_mai_n249_), .B(mai_mai_n240_), .C(mai_mai_n234_), .Y(mai_mai_n250_));
  NA2        m228(.A(mai_mai_n112_), .B(x03), .Y(mai_mai_n251_));
  OAI210     m229(.A0(mai_mai_n146_), .A1(mai_mai_n51_), .B0(mai_mai_n251_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n252_), .B(mai_mai_n93_), .Y(mai_mai_n253_));
  OAI220     m231(.A0(mai_mai_n221_), .A1(x09), .B0(mai_mai_n106_), .B1(mai_mai_n28_), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n254_), .B(mai_mai_n94_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n221_), .B(mai_mai_n89_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n89_), .B(mai_mai_n41_), .Y(mai_mai_n257_));
  NA3        m235(.A(mai_mai_n257_), .B(mai_mai_n256_), .C(mai_mai_n105_), .Y(mai_mai_n258_));
  NA4        m236(.A(mai_mai_n258_), .B(mai_mai_n255_), .C(mai_mai_n253_), .D(mai_mai_n48_), .Y(mai_mai_n259_));
  INV        m237(.A(mai_mai_n158_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n134_), .B(mai_mai_n40_), .Y(mai_mai_n261_));
  OAI220     m239(.A0(mai_mai_n344_), .A1(mai_mai_n261_), .B0(mai_mai_n260_), .B1(mai_mai_n58_), .Y(mai_mai_n262_));
  NA2        m240(.A(mai_mai_n262_), .B(x02), .Y(mai_mai_n263_));
  OAI210     m241(.A0(mai_mai_n345_), .A1(x04), .B0(mai_mai_n84_), .Y(mai_mai_n264_));
  NO3        m242(.A(mai_mai_n156_), .B(mai_mai_n132_), .C(mai_mai_n52_), .Y(mai_mai_n265_));
  OAI210     m243(.A0(mai_mai_n117_), .A1(mai_mai_n36_), .B0(mai_mai_n89_), .Y(mai_mai_n266_));
  NA2        m244(.A(mai_mai_n266_), .B(mai_mai_n265_), .Y(mai_mai_n267_));
  NA4        m245(.A(mai_mai_n267_), .B(mai_mai_n264_), .C(mai_mai_n263_), .D(x06), .Y(mai_mai_n268_));
  NA2        m246(.A(x09), .B(x03), .Y(mai_mai_n269_));
  OAI220     m247(.A0(mai_mai_n269_), .A1(mai_mai_n104_), .B0(mai_mai_n164_), .B1(mai_mai_n63_), .Y(mai_mai_n270_));
  OAI220     m248(.A0(mai_mai_n133_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n271_), .B(mai_mai_n178_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n273_));
  NA2        m251(.A(mai_mai_n265_), .B(mai_mai_n273_), .Y(mai_mai_n274_));
  OAI210     m252(.A0(mai_mai_n272_), .A1(mai_mai_n28_), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  AO220      m253(.A0(mai_mai_n275_), .A1(x04), .B0(mai_mai_n270_), .B1(x05), .Y(mai_mai_n276_));
  AOI210     m254(.A0(mai_mai_n268_), .A1(mai_mai_n259_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  OAI210     m255(.A0(mai_mai_n250_), .A1(x12), .B0(mai_mai_n277_), .Y(mai03));
  NO2        m256(.A(mai_mai_n90_), .B(mai_mai_n58_), .Y(mai_mai_n279_));
  OAI210     m257(.A0(mai_mai_n279_), .A1(x05), .B0(mai_mai_n89_), .Y(mai_mai_n280_));
  NO3        m258(.A(mai_mai_n257_), .B(mai_mai_n76_), .C(mai_mai_n58_), .Y(mai_mai_n281_));
  AOI210     m259(.A0(mai_mai_n151_), .A1(mai_mai_n89_), .B0(mai_mai_n115_), .Y(mai_mai_n282_));
  OA210      m260(.A0(mai_mai_n134_), .A1(x12), .B0(mai_mai_n108_), .Y(mai_mai_n283_));
  NO3        m261(.A(mai_mai_n283_), .B(mai_mai_n282_), .C(mai_mai_n281_), .Y(mai_mai_n284_));
  NA2        m262(.A(mai_mai_n284_), .B(mai_mai_n280_), .Y(mai04));
  NO2        m263(.A(mai_mai_n77_), .B(mai_mai_n39_), .Y(mai_mai_n286_));
  XO2        m264(.A(mai_mai_n286_), .B(mai_mai_n197_), .Y(mai05));
  NO2        m265(.A(mai_mai_n52_), .B(mai_mai_n167_), .Y(mai_mai_n288_));
  AOI210     m266(.A0(mai_mai_n288_), .A1(mai_mai_n242_), .B0(mai_mai_n25_), .Y(mai_mai_n289_));
  NA2        m267(.A(mai_mai_n113_), .B(mai_mai_n31_), .Y(mai_mai_n290_));
  AOI210     m268(.A0(x06), .A1(mai_mai_n290_), .B0(mai_mai_n24_), .Y(mai_mai_n291_));
  OAI210     m269(.A0(mai_mai_n291_), .A1(mai_mai_n289_), .B0(mai_mai_n89_), .Y(mai_mai_n292_));
  NA2        m270(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n293_));
  NA2        m271(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n294_));
  NA2        m272(.A(mai_mai_n202_), .B(x03), .Y(mai_mai_n295_));
  OAI220     m273(.A0(mai_mai_n295_), .A1(mai_mai_n294_), .B0(mai_mai_n293_), .B1(mai_mai_n73_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n26_), .A1(mai_mai_n89_), .B0(x07), .Y(mai_mai_n297_));
  AOI210     m275(.A0(mai_mai_n296_), .A1(x06), .B0(mai_mai_n297_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n128_), .B(x05), .Y(mai_mai_n299_));
  NA3        m277(.A(mai_mai_n299_), .B(mai_mai_n193_), .C(mai_mai_n188_), .Y(mai_mai_n300_));
  NO2        m278(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n301_));
  OAI210     m279(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n302_));
  OR3        m280(.A(mai_mai_n302_), .B(mai_mai_n301_), .C(mai_mai_n44_), .Y(mai_mai_n303_));
  NA2        m281(.A(mai_mai_n303_), .B(mai_mai_n300_), .Y(mai_mai_n304_));
  NA2        m282(.A(mai_mai_n304_), .B(mai_mai_n89_), .Y(mai_mai_n305_));
  NA2        m283(.A(mai_mai_n33_), .B(mai_mai_n89_), .Y(mai_mai_n306_));
  AOI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n80_), .B0(x07), .Y(mai_mai_n307_));
  AOI220     m285(.A0(mai_mai_n307_), .A1(mai_mai_n305_), .B0(mai_mai_n298_), .B1(mai_mai_n292_), .Y(mai_mai_n308_));
  NO2        m286(.A(mai_mai_n70_), .B(mai_mai_n112_), .Y(mai_mai_n309_));
  OR2        m287(.A(mai_mai_n309_), .B(x03), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n273_), .B(mai_mai_n60_), .Y(mai_mai_n311_));
  NO2        m289(.A(mai_mai_n311_), .B(x11), .Y(mai_mai_n312_));
  NO3        m290(.A(mai_mai_n312_), .B(mai_mai_n114_), .C(mai_mai_n28_), .Y(mai_mai_n313_));
  AOI210     m291(.A0(mai_mai_n313_), .A1(mai_mai_n310_), .B0(mai_mai_n47_), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n314_), .B(mai_mai_n90_), .Y(mai_mai_n315_));
  NOi21      m293(.An(mai_mai_n251_), .B(mai_mai_n108_), .Y(mai_mai_n316_));
  NO2        m294(.A(mai_mai_n316_), .B(mai_mai_n212_), .Y(mai_mai_n317_));
  OAI210     m295(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n318_));
  AOI210     m296(.A0(mai_mai_n197_), .A1(mai_mai_n47_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  NO3        m297(.A(mai_mai_n319_), .B(mai_mai_n317_), .C(x08), .Y(mai_mai_n320_));
  NO2        m298(.A(mai_mai_n106_), .B(mai_mai_n28_), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n321_), .B(mai_mai_n216_), .Y(mai_mai_n322_));
  AOI210     m300(.A0(mai_mai_n320_), .A1(mai_mai_n315_), .B0(x08), .Y(mai_mai_n323_));
  OAI210     m301(.A0(mai_mai_n311_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n232_), .B(x07), .Y(mai_mai_n325_));
  OAI220     m303(.A0(mai_mai_n325_), .A1(mai_mai_n294_), .B0(mai_mai_n114_), .B1(mai_mai_n43_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n326_), .A1(mai_mai_n324_), .B0(mai_mai_n150_), .Y(mai_mai_n327_));
  NA3        m305(.A(mai_mai_n322_), .B(mai_mai_n316_), .C(mai_mai_n256_), .Y(mai_mai_n328_));
  INV        m306(.A(x14), .Y(mai_mai_n329_));
  NO3        m307(.A(mai_mai_n251_), .B(mai_mai_n92_), .C(x11), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n330_), .B(mai_mai_n329_), .Y(mai_mai_n331_));
  NA3        m309(.A(mai_mai_n331_), .B(mai_mai_n328_), .C(mai_mai_n327_), .Y(mai_mai_n332_));
  AOI220     m310(.A0(mai_mai_n306_), .A1(mai_mai_n60_), .B0(mai_mai_n321_), .B1(mai_mai_n132_), .Y(mai_mai_n333_));
  NOi21      m311(.An(mai_mai_n221_), .B(mai_mai_n118_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n226_), .B(mai_mai_n182_), .Y(mai_mai_n335_));
  OAI210     m313(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n335_), .Y(mai_mai_n336_));
  OAI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n334_), .B0(mai_mai_n89_), .Y(mai_mai_n337_));
  OAI210     m315(.A0(mai_mai_n333_), .A1(mai_mai_n79_), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  NO4        m316(.A(mai_mai_n338_), .B(mai_mai_n332_), .C(mai_mai_n323_), .D(mai_mai_n308_), .Y(mai06));
  INV        m317(.A(x04), .Y(mai_mai_n342_));
  INV        m318(.A(mai_mai_n241_), .Y(mai_mai_n343_));
  INV        m319(.A(x05), .Y(mai_mai_n344_));
  INV        m320(.A(x13), .Y(mai_mai_n345_));
  INV        m321(.A(x03), .Y(mai_mai_n346_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  INV        u004(.A(x02), .Y(men_men_n27_));
  INV        u005(.A(x10), .Y(men_men_n28_));
  NA2        u006(.A(men_men_n28_), .B(men_men_n27_), .Y(men_men_n29_));
  INV        u007(.A(x03), .Y(men_men_n30_));
  NA2        u008(.A(x10), .B(men_men_n30_), .Y(men_men_n31_));
  INV        u009(.A(x04), .Y(men_men_n32_));
  INV        u010(.A(x08), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(x02), .Y(men_men_n34_));
  NA2        u012(.A(x08), .B(x03), .Y(men_men_n35_));
  AOI210     u013(.A0(men_men_n35_), .A1(men_men_n34_), .B0(men_men_n32_), .Y(men_men_n36_));
  NA2        u014(.A(x09), .B(men_men_n30_), .Y(men_men_n37_));
  INV        u015(.A(x05), .Y(men_men_n38_));
  NO2        u016(.A(x09), .B(x02), .Y(men_men_n39_));
  NO2        u017(.A(men_men_n39_), .B(men_men_n38_), .Y(men_men_n40_));
  NA2        u018(.A(men_men_n40_), .B(men_men_n37_), .Y(men_men_n41_));
  INV        u019(.A(men_men_n41_), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n36_), .Y(men00));
  INV        u021(.A(x01), .Y(men_men_n44_));
  INV        u022(.A(x06), .Y(men_men_n45_));
  NA2        u023(.A(men_men_n45_), .B(men_men_n27_), .Y(men_men_n46_));
  INV        u024(.A(x09), .Y(men_men_n47_));
  NO2        u025(.A(x10), .B(x02), .Y(men_men_n48_));
  NOi21      u026(.An(x01), .B(x09), .Y(men_men_n49_));
  INV        u027(.A(x00), .Y(men_men_n50_));
  NO2        u028(.A(men_men_n47_), .B(men_men_n50_), .Y(men_men_n51_));
  NA2        u029(.A(x09), .B(men_men_n50_), .Y(men_men_n52_));
  INV        u030(.A(x07), .Y(men_men_n53_));
  NA2        u031(.A(men_men_n53_), .B(men_men_n45_), .Y(men_men_n54_));
  INV        u032(.A(men_men_n29_), .Y(men_men_n55_));
  NO2        u033(.A(men_men_n55_), .B(men_men_n50_), .Y(men_men_n56_));
  AOI210     u034(.A0(men_men_n56_), .A1(men_men_n46_), .B0(x05), .Y(men_men_n57_));
  NA2        u035(.A(x10), .B(x09), .Y(men_men_n58_));
  NA2        u036(.A(x09), .B(x05), .Y(men_men_n59_));
  NA2        u037(.A(x10), .B(x06), .Y(men_men_n60_));
  NA3        u038(.A(men_men_n60_), .B(men_men_n59_), .C(men_men_n27_), .Y(men_men_n61_));
  NO2        u039(.A(men_men_n53_), .B(men_men_n38_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n61_), .B(x03), .Y(men_men_n63_));
  NOi31      u041(.An(x08), .B(x04), .C(x00), .Y(men_men_n64_));
  NO2        u042(.A(x09), .B(men_men_n38_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n65_), .B(men_men_n33_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n65_), .A1(men_men_n28_), .B0(x02), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n45_), .B(men_men_n67_), .Y(men_men_n68_));
  NO2        u046(.A(men_men_n33_), .B(x00), .Y(men_men_n69_));
  NO2        u047(.A(x08), .B(x01), .Y(men_men_n70_));
  OAI210     u048(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n32_), .Y(men_men_n71_));
  NA2        u049(.A(men_men_n47_), .B(men_men_n33_), .Y(men_men_n72_));
  NO2        u050(.A(men_men_n71_), .B(men_men_n68_), .Y(men_men_n73_));
  AN2        u051(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n74_));
  INV        u052(.A(men_men_n71_), .Y(men_men_n75_));
  NO2        u053(.A(x06), .B(x05), .Y(men_men_n76_));
  NA2        u054(.A(x11), .B(x00), .Y(men_men_n77_));
  NO2        u055(.A(x11), .B(men_men_n44_), .Y(men_men_n78_));
  NOi21      u056(.An(men_men_n77_), .B(men_men_n78_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n76_), .B(men_men_n79_), .Y(men_men_n80_));
  NOi21      u058(.An(x01), .B(x10), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n28_), .B(men_men_n50_), .Y(men_men_n82_));
  NO3        u060(.A(men_men_n82_), .B(men_men_n81_), .C(x06), .Y(men_men_n83_));
  INV        u061(.A(men_men_n83_), .Y(men_men_n84_));
  OAI210     u062(.A0(men_men_n80_), .A1(x07), .B0(men_men_n84_), .Y(men_men_n85_));
  NO3        u063(.A(men_men_n85_), .B(men_men_n74_), .C(men_men_n57_), .Y(men01));
  INV        u064(.A(x12), .Y(men_men_n87_));
  INV        u065(.A(x13), .Y(men_men_n88_));
  NA2        u066(.A(x08), .B(x04), .Y(men_men_n89_));
  NO2        u067(.A(men_men_n89_), .B(men_men_n50_), .Y(men_men_n90_));
  NA2        u068(.A(men_men_n90_), .B(men_men_n76_), .Y(men_men_n91_));
  NA2        u069(.A(men_men_n81_), .B(men_men_n27_), .Y(men_men_n92_));
  NO2        u070(.A(x10), .B(x01), .Y(men_men_n93_));
  NO2        u071(.A(men_men_n28_), .B(x00), .Y(men_men_n94_));
  NO2        u072(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u073(.A(x04), .B(men_men_n27_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n33_), .C(men_men_n38_), .Y(men_men_n97_));
  NA2        u075(.A(men_men_n97_), .B(men_men_n95_), .Y(men_men_n98_));
  AOI210     u076(.A0(men_men_n98_), .A1(men_men_n91_), .B0(men_men_n88_), .Y(men_men_n99_));
  NO2        u077(.A(men_men_n49_), .B(x05), .Y(men_men_n100_));
  NOi21      u078(.An(men_men_n100_), .B(men_men_n51_), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n32_), .B(x02), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n88_), .B(men_men_n33_), .Y(men_men_n103_));
  NA3        u081(.A(men_men_n103_), .B(men_men_n102_), .C(x06), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n101_), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n70_), .B(x13), .Y(men_men_n106_));
  NA2        u084(.A(x09), .B(men_men_n32_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NA2        u086(.A(x13), .B(men_men_n32_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(x05), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n110_), .B(men_men_n108_), .Y(men_men_n111_));
  NA2        u089(.A(men_men_n32_), .B(men_men_n50_), .Y(men_men_n112_));
  NA2        u090(.A(men_men_n112_), .B(men_men_n88_), .Y(men_men_n113_));
  AOI210     u091(.A0(men_men_n113_), .A1(men_men_n66_), .B0(men_men_n101_), .Y(men_men_n114_));
  AOI210     u092(.A0(men_men_n114_), .A1(men_men_n111_), .B0(men_men_n60_), .Y(men_men_n115_));
  NA2        u093(.A(men_men_n28_), .B(men_men_n44_), .Y(men_men_n116_));
  NA2        u094(.A(x10), .B(men_men_n50_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n47_), .B(x05), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n33_), .B(x04), .Y(men_men_n120_));
  NA3        u098(.A(men_men_n120_), .B(men_men_n119_), .C(x13), .Y(men_men_n121_));
  NO3        u099(.A(men_men_n112_), .B(men_men_n65_), .C(men_men_n33_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n52_), .B(x05), .Y(men_men_n123_));
  NOi41      u101(.An(men_men_n121_), .B(men_men_n123_), .C(men_men_n122_), .D(men_men_n118_), .Y(men_men_n124_));
  NO3        u102(.A(men_men_n124_), .B(x06), .C(x03), .Y(men_men_n125_));
  NO4        u103(.A(men_men_n125_), .B(men_men_n115_), .C(men_men_n105_), .D(men_men_n99_), .Y(men_men_n126_));
  NA2        u104(.A(x13), .B(men_men_n33_), .Y(men_men_n127_));
  OAI210     u105(.A0(men_men_n70_), .A1(x13), .B0(men_men_n32_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n129_));
  BUFFER     u107(.A(x04), .Y(men_men_n130_));
  NO2        u108(.A(men_men_n47_), .B(men_men_n38_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n28_), .B(x06), .Y(men_men_n132_));
  AOI210     u110(.A0(men_men_n132_), .A1(men_men_n46_), .B0(men_men_n131_), .Y(men_men_n133_));
  OA210      u111(.A0(men_men_n133_), .A1(men_men_n130_), .B0(men_men_n129_), .Y(men_men_n134_));
  NO2        u112(.A(x09), .B(x05), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(men_men_n44_), .Y(men_men_n136_));
  AOI210     u114(.A0(men_men_n136_), .A1(men_men_n95_), .B0(men_men_n46_), .Y(men_men_n137_));
  NA2        u115(.A(x09), .B(x00), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n100_), .B(men_men_n138_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n64_), .B(men_men_n47_), .Y(men_men_n140_));
  AOI210     u118(.A0(men_men_n140_), .A1(men_men_n139_), .B0(men_men_n132_), .Y(men_men_n141_));
  NO3        u119(.A(men_men_n141_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n142_));
  NO2        u120(.A(x03), .B(x02), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n71_), .B(men_men_n88_), .Y(men_men_n144_));
  OAI210     u122(.A0(men_men_n144_), .A1(men_men_n101_), .B0(men_men_n143_), .Y(men_men_n145_));
  OA210      u123(.A0(men_men_n142_), .A1(x11), .B0(men_men_n145_), .Y(men_men_n146_));
  OAI210     u124(.A0(men_men_n126_), .A1(men_men_n23_), .B0(men_men_n146_), .Y(men_men_n147_));
  NAi21      u125(.An(x06), .B(x10), .Y(men_men_n148_));
  NOi21      u126(.An(x01), .B(x13), .Y(men_men_n149_));
  NA2        u127(.A(men_men_n149_), .B(men_men_n148_), .Y(men_men_n150_));
  OR2        u128(.A(men_men_n150_), .B(x08), .Y(men_men_n151_));
  NO2        u129(.A(men_men_n151_), .B(men_men_n38_), .Y(men_men_n152_));
  NO2        u130(.A(men_men_n28_), .B(x03), .Y(men_men_n153_));
  NA2        u131(.A(men_men_n88_), .B(x01), .Y(men_men_n154_));
  OAI210     u132(.A0(x05), .A1(men_men_n88_), .B0(men_men_n47_), .Y(men_men_n155_));
  AOI210     u133(.A0(men_men_n155_), .A1(men_men_n153_), .B0(men_men_n45_), .Y(men_men_n156_));
  AOI210     u134(.A0(x11), .A1(men_men_n30_), .B0(men_men_n27_), .Y(men_men_n157_));
  OAI210     u135(.A0(men_men_n156_), .A1(men_men_n152_), .B0(men_men_n157_), .Y(men_men_n158_));
  NA2        u136(.A(x04), .B(x02), .Y(men_men_n159_));
  NA2        u137(.A(x10), .B(x05), .Y(men_men_n160_));
  NA2        u138(.A(x09), .B(x06), .Y(men_men_n161_));
  NO2        u139(.A(x09), .B(x01), .Y(men_men_n162_));
  NO3        u140(.A(men_men_n162_), .B(men_men_n93_), .C(men_men_n30_), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n163_), .B(x00), .Y(men_men_n164_));
  NA3        u142(.A(men_men_n149_), .B(men_men_n148_), .C(men_men_n47_), .Y(men_men_n165_));
  OAI210     u143(.A0(men_men_n165_), .A1(x11), .B0(men_men_n164_), .Y(men_men_n166_));
  NAi21      u144(.An(men_men_n159_), .B(men_men_n166_), .Y(men_men_n167_));
  INV        u145(.A(men_men_n25_), .Y(men_men_n168_));
  NAi21      u146(.An(x13), .B(x00), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n28_), .A1(men_men_n45_), .B0(men_men_n169_), .Y(men_men_n170_));
  AOI220     u148(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n160_), .A1(men_men_n32_), .B0(men_men_n171_), .Y(men_men_n172_));
  AN2        u150(.A(men_men_n172_), .B(men_men_n170_), .Y(men_men_n173_));
  AN2        u151(.A(men_men_n60_), .B(men_men_n59_), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n82_), .B(x06), .Y(men_men_n175_));
  NO2        u153(.A(men_men_n169_), .B(men_men_n33_), .Y(men_men_n176_));
  OAI220     u154(.A0(men_men_n169_), .A1(men_men_n161_), .B0(men_men_n175_), .B1(men_men_n174_), .Y(men_men_n177_));
  OAI210     u155(.A0(men_men_n177_), .A1(men_men_n173_), .B0(men_men_n168_), .Y(men_men_n178_));
  NOi21      u156(.An(x09), .B(x00), .Y(men_men_n179_));
  NO3        u157(.A(men_men_n69_), .B(men_men_n179_), .C(men_men_n44_), .Y(men_men_n180_));
  NA2        u158(.A(men_men_n180_), .B(men_men_n117_), .Y(men_men_n181_));
  NA2        u159(.A(x10), .B(x08), .Y(men_men_n182_));
  INV        u160(.A(men_men_n182_), .Y(men_men_n183_));
  NA2        u161(.A(x06), .B(x05), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(men_men_n32_), .B0(men_men_n87_), .Y(men_men_n185_));
  AOI210     u163(.A0(men_men_n183_), .A1(men_men_n51_), .B0(men_men_n185_), .Y(men_men_n186_));
  NA2        u164(.A(men_men_n186_), .B(men_men_n181_), .Y(men_men_n187_));
  NO2        u165(.A(men_men_n88_), .B(x12), .Y(men_men_n188_));
  AOI210     u166(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n188_), .Y(men_men_n189_));
  NA2        u167(.A(men_men_n81_), .B(men_men_n47_), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n32_), .B(men_men_n30_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n191_), .B(x02), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n192_), .B(men_men_n190_), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n189_), .A1(men_men_n187_), .B0(men_men_n193_), .Y(men_men_n194_));
  NA4        u172(.A(men_men_n194_), .B(men_men_n178_), .C(men_men_n167_), .D(men_men_n158_), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n147_), .A1(men_men_n87_), .B0(men_men_n195_), .Y(men_men_n196_));
  INV        u174(.A(men_men_n61_), .Y(men_men_n197_));
  NA2        u175(.A(men_men_n197_), .B(men_men_n129_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n199_));
  NA2        u177(.A(men_men_n199_), .B(men_men_n128_), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n29_), .A1(x06), .B0(x05), .Y(men_men_n201_));
  NO2        u179(.A(men_men_n116_), .B(x06), .Y(men_men_n202_));
  AOI210     u180(.A0(men_men_n201_), .A1(men_men_n200_), .B0(men_men_n202_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n203_), .A1(men_men_n198_), .B0(x12), .Y(men_men_n204_));
  INV        u182(.A(men_men_n64_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n182_), .A1(x05), .B0(men_men_n47_), .Y(men_men_n206_));
  OAI210     u184(.A0(men_men_n206_), .A1(men_men_n150_), .B0(men_men_n50_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(men_men_n205_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n81_), .B(x06), .Y(men_men_n209_));
  AOI210     u187(.A0(men_men_n33_), .A1(x04), .B0(men_men_n47_), .Y(men_men_n210_));
  NO2        u188(.A(men_men_n210_), .B(men_men_n38_), .Y(men_men_n211_));
  OAI210     u189(.A0(men_men_n49_), .A1(men_men_n211_), .B0(x02), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n212_), .A1(men_men_n208_), .B0(men_men_n23_), .Y(men_men_n213_));
  OAI210     u191(.A0(men_men_n204_), .A1(men_men_n50_), .B0(men_men_n213_), .Y(men_men_n214_));
  INV        u192(.A(men_men_n132_), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n47_), .B(x03), .Y(men_men_n216_));
  OAI210     u194(.A0(men_men_n65_), .A1(men_men_n33_), .B0(men_men_n107_), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n88_), .B(x03), .Y(men_men_n218_));
  AOI220     u196(.A0(men_men_n218_), .A1(men_men_n217_), .B0(men_men_n64_), .B1(men_men_n216_), .Y(men_men_n219_));
  INV        u197(.A(men_men_n148_), .Y(men_men_n220_));
  NOi21      u198(.An(x13), .B(x04), .Y(men_men_n221_));
  NO3        u199(.A(men_men_n221_), .B(men_men_n64_), .C(men_men_n179_), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n220_), .B(men_men_n50_), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n219_), .B(men_men_n223_), .Y(men_men_n224_));
  INV        u202(.A(men_men_n78_), .Y(men_men_n225_));
  NA2        u203(.A(men_men_n23_), .B(men_men_n44_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n47_), .B(men_men_n33_), .Y(men_men_n227_));
  OAI210     u205(.A0(men_men_n227_), .A1(men_men_n172_), .B0(men_men_n170_), .Y(men_men_n228_));
  AOI210     u206(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n229_), .B(men_men_n38_), .Y(men_men_n230_));
  OAI210     u208(.A0(men_men_n89_), .A1(men_men_n138_), .B0(men_men_n60_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  INV        u210(.A(x03), .Y(men_men_n233_));
  OA210      u211(.A0(men_men_n233_), .A1(men_men_n232_), .B0(men_men_n228_), .Y(men_men_n234_));
  NA2        u212(.A(x13), .B(men_men_n87_), .Y(men_men_n235_));
  NA3        u213(.A(men_men_n235_), .B(men_men_n185_), .C(men_men_n79_), .Y(men_men_n236_));
  OAI210     u214(.A0(men_men_n234_), .A1(men_men_n226_), .B0(men_men_n236_), .Y(men_men_n237_));
  AOI210     u215(.A0(men_men_n78_), .A1(men_men_n224_), .B0(men_men_n237_), .Y(men_men_n238_));
  AOI210     u216(.A0(men_men_n238_), .A1(men_men_n214_), .B0(x07), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n59_), .B(men_men_n28_), .Y(men_men_n240_));
  AOI210     u218(.A0(men_men_n127_), .A1(men_men_n140_), .B0(men_men_n240_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n88_), .B(x06), .Y(men_men_n242_));
  INV        u220(.A(men_men_n242_), .Y(men_men_n243_));
  NO2        u221(.A(x08), .B(x05), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n244_), .B(men_men_n229_), .Y(men_men_n245_));
  OAI210     u223(.A0(men_men_n64_), .A1(x13), .B0(men_men_n30_), .Y(men_men_n246_));
  OAI210     u224(.A0(men_men_n245_), .A1(men_men_n243_), .B0(men_men_n246_), .Y(men_men_n247_));
  NO2        u225(.A(x12), .B(x02), .Y(men_men_n248_));
  INV        u226(.A(men_men_n248_), .Y(men_men_n249_));
  NO2        u227(.A(men_men_n249_), .B(men_men_n225_), .Y(men_men_n250_));
  OA210      u228(.A0(men_men_n247_), .A1(men_men_n241_), .B0(men_men_n250_), .Y(men_men_n251_));
  NA2        u229(.A(men_men_n47_), .B(men_men_n38_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(x01), .Y(men_men_n253_));
  AOI210     u231(.A0(men_men_n107_), .A1(men_men_n121_), .B0(men_men_n28_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n242_), .B(men_men_n217_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n88_), .B(x04), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n256_), .B(men_men_n27_), .Y(men_men_n257_));
  NA2        u235(.A(men_men_n257_), .B(men_men_n255_), .Y(men_men_n258_));
  NO3        u236(.A(men_men_n77_), .B(x12), .C(x03), .Y(men_men_n259_));
  OAI210     u237(.A0(men_men_n258_), .A1(men_men_n254_), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n190_), .A1(men_men_n184_), .B0(men_men_n89_), .Y(men_men_n261_));
  NOi21      u239(.An(men_men_n240_), .B(men_men_n209_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n25_), .B(x00), .Y(men_men_n263_));
  OAI210     u241(.A0(men_men_n262_), .A1(men_men_n261_), .B0(men_men_n263_), .Y(men_men_n264_));
  NO2        u242(.A(men_men_n51_), .B(x05), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n265_), .B(men_men_n210_), .Y(men_men_n266_));
  NO2        u244(.A(men_men_n226_), .B(men_men_n27_), .Y(men_men_n267_));
  OAI210     u245(.A0(men_men_n266_), .A1(men_men_n215_), .B0(men_men_n267_), .Y(men_men_n268_));
  NA3        u246(.A(men_men_n268_), .B(men_men_n264_), .C(men_men_n260_), .Y(men_men_n269_));
  NO3        u247(.A(men_men_n269_), .B(men_men_n251_), .C(men_men_n239_), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n196_), .A1(men_men_n53_), .B0(men_men_n270_), .Y(men02));
  AOI210     u249(.A0(men_men_n127_), .A1(men_men_n71_), .B0(men_men_n119_), .Y(men_men_n272_));
  BUFFER     u250(.A(men_men_n222_), .Y(men_men_n273_));
  NA3        u251(.A(x13), .B(men_men_n183_), .C(men_men_n49_), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n273_), .A1(men_men_n31_), .B0(men_men_n274_), .Y(men_men_n275_));
  OAI210     u253(.A0(men_men_n275_), .A1(men_men_n272_), .B0(men_men_n160_), .Y(men_men_n276_));
  INV        u254(.A(men_men_n160_), .Y(men_men_n277_));
  AOI210     u255(.A0(men_men_n102_), .A1(men_men_n72_), .B0(men_men_n210_), .Y(men_men_n278_));
  OAI220     u256(.A0(men_men_n278_), .A1(men_men_n88_), .B0(men_men_n71_), .B1(men_men_n47_), .Y(men_men_n279_));
  AOI220     u257(.A0(men_men_n279_), .A1(men_men_n277_), .B0(men_men_n144_), .B1(men_men_n143_), .Y(men_men_n280_));
  AOI210     u258(.A0(men_men_n280_), .A1(men_men_n276_), .B0(men_men_n45_), .Y(men_men_n281_));
  NOi21      u259(.An(x13), .B(men_men_n409_), .Y(men_men_n282_));
  NO2        u260(.A(men_men_n221_), .B(men_men_n282_), .Y(men_men_n283_));
  AOI210     u261(.A0(men_men_n283_), .A1(men_men_n410_), .B0(men_men_n132_), .Y(men_men_n284_));
  INV        u262(.A(men_men_n219_), .Y(men_men_n285_));
  NA2        u263(.A(x01), .B(men_men_n285_), .Y(men_men_n286_));
  AN2        u264(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n287_));
  OAI210     u265(.A0(men_men_n39_), .A1(men_men_n38_), .B0(men_men_n45_), .Y(men_men_n288_));
  NA2        u266(.A(x13), .B(men_men_n27_), .Y(men_men_n289_));
  OA210      u267(.A0(men_men_n289_), .A1(x08), .B0(men_men_n136_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n290_), .A1(men_men_n128_), .B0(men_men_n288_), .Y(men_men_n291_));
  OAI210     u269(.A0(men_men_n291_), .A1(men_men_n287_), .B0(men_men_n82_), .Y(men_men_n292_));
  NA3        u270(.A(men_men_n82_), .B(men_men_n70_), .C(men_men_n216_), .Y(men_men_n293_));
  NA3        u271(.A(men_men_n81_), .B(men_men_n69_), .C(men_men_n39_), .Y(men_men_n294_));
  AOI210     u272(.A0(men_men_n294_), .A1(men_men_n293_), .B0(x04), .Y(men_men_n295_));
  NO2        u273(.A(men_men_n245_), .B(men_men_n92_), .Y(men_men_n296_));
  AOI210     u274(.A0(men_men_n296_), .A1(x13), .B0(men_men_n295_), .Y(men_men_n297_));
  NA3        u275(.A(men_men_n297_), .B(men_men_n292_), .C(men_men_n286_), .Y(men_men_n298_));
  NO3        u276(.A(men_men_n298_), .B(men_men_n284_), .C(men_men_n281_), .Y(men_men_n299_));
  NA2        u277(.A(men_men_n131_), .B(x03), .Y(men_men_n300_));
  INV        u278(.A(men_men_n169_), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n47_), .A1(men_men_n32_), .B0(men_men_n33_), .Y(men_men_n302_));
  AOI220     u280(.A0(men_men_n302_), .A1(men_men_n301_), .B0(men_men_n191_), .B1(x08), .Y(men_men_n303_));
  OAI210     u281(.A0(men_men_n303_), .A1(men_men_n265_), .B0(men_men_n300_), .Y(men_men_n304_));
  NA2        u282(.A(men_men_n304_), .B(men_men_n93_), .Y(men_men_n305_));
  OAI210     u283(.A0(men_men_n49_), .A1(x05), .B0(men_men_n94_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n256_), .B(men_men_n87_), .Y(men_men_n307_));
  NA2        u285(.A(men_men_n87_), .B(men_men_n38_), .Y(men_men_n308_));
  NA3        u286(.A(men_men_n308_), .B(men_men_n307_), .C(men_men_n118_), .Y(men_men_n309_));
  NA4        u287(.A(men_men_n309_), .B(men_men_n306_), .C(men_men_n305_), .D(men_men_n45_), .Y(men_men_n310_));
  INV        u288(.A(men_men_n191_), .Y(men_men_n311_));
  INV        u289(.A(men_men_n227_), .Y(men_men_n312_));
  NA2        u290(.A(men_men_n188_), .B(x04), .Y(men_men_n313_));
  NO2        u291(.A(men_men_n313_), .B(men_men_n312_), .Y(men_men_n314_));
  NO3        u292(.A(men_men_n171_), .B(x13), .C(men_men_n30_), .Y(men_men_n315_));
  OAI210     u293(.A0(men_men_n315_), .A1(men_men_n314_), .B0(men_men_n82_), .Y(men_men_n316_));
  NO3        u294(.A(men_men_n188_), .B(men_men_n153_), .C(men_men_n48_), .Y(men_men_n317_));
  OAI210     u295(.A0(x12), .A1(men_men_n180_), .B0(men_men_n317_), .Y(men_men_n318_));
  NA3        u296(.A(men_men_n318_), .B(men_men_n316_), .C(x06), .Y(men_men_n319_));
  NO3        u297(.A(men_men_n265_), .B(men_men_n116_), .C(x08), .Y(men_men_n320_));
  AOI210     u298(.A0(x01), .A1(men_men_n215_), .B0(men_men_n320_), .Y(men_men_n321_));
  NO3        u299(.A(men_men_n100_), .B(men_men_n117_), .C(men_men_n35_), .Y(men_men_n322_));
  INV        u300(.A(men_men_n322_), .Y(men_men_n323_));
  OAI210     u301(.A0(men_men_n321_), .A1(men_men_n27_), .B0(men_men_n323_), .Y(men_men_n324_));
  AN2        u302(.A(men_men_n324_), .B(x04), .Y(men_men_n325_));
  AOI210     u303(.A0(men_men_n319_), .A1(men_men_n310_), .B0(men_men_n325_), .Y(men_men_n326_));
  OAI210     u304(.A0(men_men_n299_), .A1(x12), .B0(men_men_n326_), .Y(men03));
  OR2        u305(.A(men_men_n39_), .B(men_men_n216_), .Y(men_men_n328_));
  NO2        u306(.A(men_men_n87_), .B(men_men_n328_), .Y(men_men_n329_));
  AO210      u307(.A0(men_men_n312_), .A1(men_men_n72_), .B0(men_men_n313_), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(men_men_n192_), .Y(men_men_n331_));
  OAI210     u309(.A0(men_men_n331_), .A1(men_men_n329_), .B0(x05), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n328_), .B(x05), .Y(men_men_n333_));
  AOI210     u311(.A0(men_men_n128_), .A1(men_men_n205_), .B0(men_men_n333_), .Y(men_men_n334_));
  AOI210     u312(.A0(men_men_n218_), .A1(men_men_n66_), .B0(men_men_n110_), .Y(men_men_n335_));
  OAI210     u313(.A0(men_men_n289_), .A1(men_men_n409_), .B0(men_men_n335_), .Y(men_men_n336_));
  OAI210     u314(.A0(men_men_n336_), .A1(men_men_n334_), .B0(men_men_n87_), .Y(men_men_n337_));
  NA3        u315(.A(men_men_n139_), .B(men_men_n337_), .C(men_men_n332_), .Y(men04));
  NO2        u316(.A(men_men_n75_), .B(men_men_n36_), .Y(men_men_n339_));
  XO2        u317(.A(men_men_n339_), .B(men_men_n235_), .Y(men05));
  AOI210     u318(.A0(men_men_n59_), .A1(men_men_n48_), .B0(men_men_n202_), .Y(men_men_n341_));
  AOI210     u319(.A0(men_men_n341_), .A1(men_men_n288_), .B0(men_men_n25_), .Y(men_men_n342_));
  NA3        u320(.A(men_men_n132_), .B(men_men_n119_), .C(men_men_n30_), .Y(men_men_n343_));
  AOI210     u321(.A0(men_men_n220_), .A1(men_men_n50_), .B0(men_men_n76_), .Y(men_men_n344_));
  AOI210     u322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n24_), .Y(men_men_n345_));
  OAI210     u323(.A0(men_men_n345_), .A1(men_men_n342_), .B0(men_men_n87_), .Y(men_men_n346_));
  NA2        u324(.A(x11), .B(men_men_n30_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n23_), .B(men_men_n27_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n240_), .B(x03), .Y(men_men_n349_));
  OAI220     u327(.A0(men_men_n349_), .A1(men_men_n348_), .B0(men_men_n347_), .B1(men_men_n67_), .Y(men_men_n350_));
  OAI210     u328(.A0(men_men_n26_), .A1(men_men_n87_), .B0(x07), .Y(men_men_n351_));
  AOI210     u329(.A0(men_men_n350_), .A1(x06), .B0(men_men_n351_), .Y(men_men_n352_));
  AOI220     u330(.A0(men_men_n67_), .A1(men_men_n30_), .B0(men_men_n48_), .B1(men_men_n47_), .Y(men_men_n353_));
  NO3        u331(.A(men_men_n353_), .B(men_men_n23_), .C(x00), .Y(men_men_n354_));
  NA2        u332(.A(men_men_n58_), .B(x02), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n355_), .A1(men_men_n349_), .B0(men_men_n242_), .Y(men_men_n356_));
  OR2        u334(.A(men_men_n356_), .B(men_men_n226_), .Y(men_men_n357_));
  NO2        u335(.A(men_men_n23_), .B(x10), .Y(men_men_n358_));
  OAI210     u336(.A0(x11), .A1(men_men_n28_), .B0(men_men_n45_), .Y(men_men_n359_));
  OR3        u337(.A(men_men_n359_), .B(men_men_n358_), .C(men_men_n41_), .Y(men_men_n360_));
  NA2        u338(.A(men_men_n360_), .B(men_men_n357_), .Y(men_men_n361_));
  OAI210     u339(.A0(men_men_n361_), .A1(men_men_n354_), .B0(men_men_n87_), .Y(men_men_n362_));
  INV        u340(.A(x07), .Y(men_men_n363_));
  AOI220     u341(.A0(men_men_n363_), .A1(men_men_n362_), .B0(men_men_n352_), .B1(men_men_n346_), .Y(men_men_n364_));
  NA3        u342(.A(men_men_n23_), .B(men_men_n53_), .C(men_men_n45_), .Y(men_men_n365_));
  AO210      u343(.A0(men_men_n365_), .A1(men_men_n252_), .B0(men_men_n249_), .Y(men_men_n366_));
  AOI210     u344(.A0(men_men_n358_), .A1(men_men_n62_), .B0(men_men_n131_), .Y(men_men_n367_));
  OR2        u345(.A(men_men_n367_), .B(x03), .Y(men_men_n368_));
  NA2        u346(.A(x05), .B(men_men_n53_), .Y(men_men_n369_));
  NO2        u347(.A(men_men_n369_), .B(x11), .Y(men_men_n370_));
  NO3        u348(.A(men_men_n370_), .B(men_men_n135_), .C(men_men_n27_), .Y(men_men_n371_));
  AOI220     u349(.A0(men_men_n371_), .A1(men_men_n368_), .B0(men_men_n366_), .B1(men_men_n44_), .Y(men_men_n372_));
  NO4        u350(.A(men_men_n308_), .B(men_men_n31_), .C(x11), .D(x09), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n88_), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n313_), .A1(men_men_n96_), .B0(men_men_n248_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n375_), .B(x08), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n358_), .A1(men_men_n27_), .B0(men_men_n30_), .Y(men_men_n377_));
  NA2        u355(.A(x09), .B(men_men_n38_), .Y(men_men_n378_));
  OAI220     u356(.A0(men_men_n378_), .A1(men_men_n377_), .B0(men_men_n347_), .B1(men_men_n54_), .Y(men_men_n379_));
  NO2        u357(.A(x13), .B(x12), .Y(men_men_n380_));
  NO2        u358(.A(men_men_n119_), .B(men_men_n27_), .Y(men_men_n381_));
  NO2        u359(.A(men_men_n381_), .B(men_men_n253_), .Y(men_men_n382_));
  OR3        u360(.A(men_men_n382_), .B(x12), .C(x03), .Y(men_men_n383_));
  NA3        u361(.A(men_men_n311_), .B(men_men_n112_), .C(x12), .Y(men_men_n384_));
  AO210      u362(.A0(men_men_n311_), .A1(men_men_n112_), .B0(men_men_n235_), .Y(men_men_n385_));
  NA4        u363(.A(men_men_n385_), .B(men_men_n384_), .C(men_men_n383_), .D(x08), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n380_), .A1(men_men_n379_), .B0(men_men_n386_), .Y(men_men_n387_));
  AOI210     u365(.A0(men_men_n376_), .A1(men_men_n374_), .B0(men_men_n387_), .Y(men_men_n388_));
  OAI210     u366(.A0(men_men_n369_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n389_));
  NA2        u367(.A(men_men_n277_), .B(x07), .Y(men_men_n390_));
  OAI220     u368(.A0(men_men_n390_), .A1(men_men_n348_), .B0(men_men_n135_), .B1(men_men_n40_), .Y(men_men_n391_));
  OAI210     u369(.A0(men_men_n391_), .A1(men_men_n389_), .B0(men_men_n176_), .Y(men_men_n392_));
  NA3        u370(.A(men_men_n382_), .B(men_men_n47_), .C(men_men_n307_), .Y(men_men_n393_));
  INV        u371(.A(x14), .Y(men_men_n394_));
  NO3        u372(.A(men_men_n300_), .B(men_men_n92_), .C(x11), .Y(men_men_n395_));
  NO3        u373(.A(men_men_n154_), .B(men_men_n62_), .C(men_men_n50_), .Y(men_men_n396_));
  NO3        u374(.A(men_men_n365_), .B(men_men_n308_), .C(men_men_n169_), .Y(men_men_n397_));
  NO4        u375(.A(men_men_n397_), .B(men_men_n396_), .C(men_men_n395_), .D(men_men_n394_), .Y(men_men_n398_));
  NA3        u376(.A(men_men_n398_), .B(men_men_n393_), .C(men_men_n392_), .Y(men_men_n399_));
  INV        u377(.A(men_men_n381_), .Y(men_men_n400_));
  NO3        u378(.A(men_men_n116_), .B(men_men_n24_), .C(x06), .Y(men_men_n401_));
  AOI210     u379(.A0(men_men_n263_), .A1(men_men_n220_), .B0(men_men_n401_), .Y(men_men_n402_));
  OAI210     u380(.A0(men_men_n41_), .A1(x04), .B0(men_men_n402_), .Y(men_men_n403_));
  NA2        u381(.A(men_men_n403_), .B(men_men_n87_), .Y(men_men_n404_));
  OAI210     u382(.A0(men_men_n400_), .A1(men_men_n77_), .B0(men_men_n404_), .Y(men_men_n405_));
  NO4        u383(.A(men_men_n405_), .B(men_men_n399_), .C(men_men_n388_), .D(men_men_n364_), .Y(men06));
  INV        u384(.A(men_men_n244_), .Y(men_men_n409_));
  INV        u385(.A(men_men_n179_), .Y(men_men_n410_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule