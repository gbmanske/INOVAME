// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n42_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n108_, new_new_n109_, new_new_n110_, new_new_n112_,
    new_new_n113_, new_new_n114_, new_new_n115_, new_new_n116_,
    new_new_n117_, new_new_n118_, new_new_n119_, new_new_n120_,
    new_new_n121_, new_new_n122_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n258_, new_new_n259_, new_new_n260_, new_new_n261_,
    new_new_n262_, new_new_n263_, new_new_n264_, new_new_n265_,
    new_new_n266_, new_new_n267_, new_new_n268_, new_new_n269_,
    new_new_n270_, new_new_n271_, new_new_n272_, new_new_n273_,
    new_new_n274_, new_new_n275_, new_new_n276_, new_new_n277_,
    new_new_n278_, new_new_n279_, new_new_n280_, new_new_n281_,
    new_new_n282_, new_new_n283_, new_new_n284_, new_new_n285_,
    new_new_n286_, new_new_n287_, new_new_n288_, new_new_n289_,
    new_new_n290_, new_new_n291_, new_new_n292_, new_new_n293_,
    new_new_n294_, new_new_n295_, new_new_n296_, new_new_n297_,
    new_new_n298_, new_new_n299_, new_new_n300_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n314_, new_new_n315_, new_new_n316_, new_new_n317_,
    new_new_n318_, new_new_n319_, new_new_n320_, new_new_n321_,
    new_new_n322_, new_new_n323_, new_new_n324_, new_new_n325_,
    new_new_n326_, new_new_n327_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n337_, new_new_n338_,
    new_new_n339_, new_new_n340_, new_new_n341_, new_new_n342_,
    new_new_n343_, new_new_n344_, new_new_n345_, new_new_n346_,
    new_new_n347_, new_new_n348_, new_new_n349_, new_new_n350_,
    new_new_n351_, new_new_n352_, new_new_n353_, new_new_n354_,
    new_new_n355_, new_new_n357_, new_new_n358_, new_new_n359_,
    new_new_n360_, new_new_n361_, new_new_n362_, new_new_n363_,
    new_new_n364_, new_new_n365_, new_new_n366_, new_new_n367_,
    new_new_n368_, new_new_n369_, new_new_n370_, new_new_n371_,
    new_new_n372_, new_new_n373_, new_new_n374_, new_new_n375_,
    new_new_n376_, new_new_n377_, new_new_n378_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n452_, new_new_n453_, new_new_n454_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  AO210      g008(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n31_));
  OR2        g009(.A(new_new_n31_), .B(i_11_), .Y(new_new_n32_));
  NA2        g010(.A(new_new_n32_), .B(new_new_n30_), .Y(new_new_n33_));
  XO2        g011(.A(new_new_n33_), .B(new_new_n23_), .Y(new_new_n34_));
  INV        g012(.A(i_4_), .Y(new_new_n35_));
  INV        g013(.A(i_10_), .Y(new_new_n36_));
  NAi21      g014(.An(i_11_), .B(i_9_), .Y(new_new_n37_));
  NO3        g015(.A(new_new_n37_), .B(i_12_), .C(new_new_n36_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n34_), .Y(ori1));
  INV        g019(.A(i_11_), .Y(new_new_n42_));
  NO2        g020(.A(new_new_n42_), .B(i_6_), .Y(new_new_n43_));
  INV        g021(.A(i_2_), .Y(new_new_n44_));
  INV        g022(.A(i_5_), .Y(new_new_n45_));
  NO2        g023(.A(i_7_), .B(i_10_), .Y(new_new_n46_));
  AOI210     g024(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n46_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_2_), .Y(new_new_n48_));
  NA2        g026(.A(i_7_), .B(i_9_), .Y(new_new_n49_));
  NO2        g027(.A(new_new_n49_), .B(new_new_n48_), .Y(new_new_n50_));
  NO2        g028(.A(i_1_), .B(i_6_), .Y(new_new_n51_));
  NA2        g029(.A(i_8_), .B(i_7_), .Y(new_new_n52_));
  NAi21      g030(.An(i_2_), .B(i_7_), .Y(new_new_n53_));
  INV        g031(.A(i_1_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n54_), .B(i_6_), .Y(new_new_n55_));
  INV        g033(.A(i_10_), .Y(new_new_n56_));
  NO2        g034(.A(new_new_n56_), .B(i_6_), .Y(new_new_n57_));
  NAi21      g035(.An(new_new_n57_), .B(new_new_n52_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n47_), .B(i_2_), .Y(new_new_n59_));
  AOI210     g037(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(i_1_), .B(i_6_), .Y(new_new_n61_));
  NO2        g039(.A(new_new_n61_), .B(new_new_n25_), .Y(new_new_n62_));
  INV        g040(.A(i_0_), .Y(new_new_n63_));
  NA2        g041(.A(i_5_), .B(i_9_), .Y(new_new_n64_));
  INV        g042(.A(new_new_n62_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n59_), .B(new_new_n65_), .Y(new_new_n66_));
  OAI210     g044(.A0(new_new_n66_), .A1(new_new_n58_), .B0(i_0_), .Y(new_new_n67_));
  NA2        g045(.A(i_12_), .B(i_5_), .Y(new_new_n68_));
  NO2        g046(.A(i_3_), .B(i_9_), .Y(new_new_n69_));
  NO2        g047(.A(i_3_), .B(i_7_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n69_), .B(new_new_n54_), .Y(new_new_n71_));
  INV        g049(.A(i_6_), .Y(new_new_n72_));
  NO2        g050(.A(i_2_), .B(i_7_), .Y(new_new_n73_));
  INV        g051(.A(new_new_n73_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n71_), .A1(i_8_), .B0(new_new_n74_), .Y(new_new_n75_));
  NAi21      g053(.An(i_6_), .B(i_10_), .Y(new_new_n76_));
  NA2        g054(.A(i_6_), .B(i_9_), .Y(new_new_n77_));
  AOI210     g055(.A0(new_new_n77_), .A1(new_new_n76_), .B0(new_new_n54_), .Y(new_new_n78_));
  NA2        g056(.A(i_2_), .B(i_6_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n79_), .B(new_new_n25_), .Y(new_new_n80_));
  NO2        g058(.A(new_new_n80_), .B(new_new_n78_), .Y(new_new_n81_));
  AOI210     g059(.A0(new_new_n81_), .A1(new_new_n75_), .B0(new_new_n68_), .Y(new_new_n82_));
  AN3        g060(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_11_), .Y(new_new_n84_));
  INV        g062(.A(i_7_), .Y(new_new_n85_));
  NA2        g063(.A(new_new_n44_), .B(new_new_n85_), .Y(new_new_n86_));
  NO2        g064(.A(i_0_), .B(i_5_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n87_), .B(new_new_n72_), .Y(new_new_n88_));
  NA2        g066(.A(i_12_), .B(i_3_), .Y(new_new_n89_));
  INV        g067(.A(new_new_n89_), .Y(new_new_n90_));
  NA3        g068(.A(new_new_n90_), .B(new_new_n88_), .C(new_new_n86_), .Y(new_new_n91_));
  NAi21      g069(.An(i_7_), .B(i_11_), .Y(new_new_n92_));
  AN2        g070(.A(i_2_), .B(i_10_), .Y(new_new_n93_));
  BUFFER     g071(.A(new_new_n68_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n54_), .B(new_new_n26_), .Y(new_new_n95_));
  NA2        g073(.A(i_11_), .B(i_12_), .Y(new_new_n96_));
  INV        g074(.A(new_new_n91_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n85_), .B(new_new_n36_), .Y(new_new_n98_));
  NA2        g076(.A(i_7_), .B(new_new_n25_), .Y(new_new_n99_));
  NA2        g077(.A(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n100_), .B(new_new_n44_), .Y(new_new_n101_));
  NA2        g079(.A(new_new_n77_), .B(new_new_n76_), .Y(new_new_n102_));
  NAi21      g080(.An(i_3_), .B(i_8_), .Y(new_new_n103_));
  NO2        g081(.A(i_1_), .B(new_new_n72_), .Y(new_new_n104_));
  NO2        g082(.A(i_6_), .B(i_5_), .Y(new_new_n105_));
  NO3        g083(.A(i_11_), .B(new_new_n97_), .C(new_new_n82_), .Y(new_new_n106_));
  NA2        g084(.A(new_new_n106_), .B(new_new_n67_), .Y(ori2));
  NO2        g085(.A(new_new_n54_), .B(new_new_n36_), .Y(new_new_n108_));
  INV        g086(.A(i_6_), .Y(new_new_n109_));
  NA2        g087(.A(new_new_n109_), .B(new_new_n108_), .Y(new_new_n110_));
  NA4        g088(.A(new_new_n110_), .B(new_new_n65_), .C(new_new_n59_), .D(new_new_n30_), .Y(ori0));
  AN2        g089(.A(i_8_), .B(i_7_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(i_6_), .Y(new_new_n113_));
  NO2        g091(.A(i_12_), .B(i_13_), .Y(new_new_n114_));
  NAi21      g092(.An(i_5_), .B(i_11_), .Y(new_new_n115_));
  NO2        g093(.A(i_0_), .B(i_1_), .Y(new_new_n116_));
  AN2        g094(.A(new_new_n114_), .B(new_new_n69_), .Y(new_new_n117_));
  NA2        g095(.A(i_1_), .B(i_5_), .Y(new_new_n118_));
  OR2        g096(.A(i_0_), .B(i_1_), .Y(new_new_n119_));
  NOi21      g097(.An(i_4_), .B(i_10_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(new_new_n39_), .Y(new_new_n121_));
  NOi21      g099(.An(i_4_), .B(i_9_), .Y(new_new_n122_));
  NOi21      g100(.An(i_11_), .B(i_13_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n63_), .B(new_new_n54_), .Y(new_new_n124_));
  NO2        g102(.A(new_new_n63_), .B(i_5_), .Y(new_new_n125_));
  NO2        g103(.A(i_2_), .B(i_1_), .Y(new_new_n126_));
  NAi21      g104(.An(i_4_), .B(i_12_), .Y(new_new_n127_));
  INV        g105(.A(i_8_), .Y(new_new_n128_));
  NO2        g106(.A(i_3_), .B(i_8_), .Y(new_new_n129_));
  NO3        g107(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n130_));
  NO2        g108(.A(new_new_n87_), .B(new_new_n51_), .Y(new_new_n131_));
  NO2        g109(.A(i_13_), .B(i_9_), .Y(new_new_n132_));
  NO2        g110(.A(new_new_n42_), .B(i_5_), .Y(new_new_n133_));
  NA2        g111(.A(i_0_), .B(i_5_), .Y(new_new_n134_));
  NAi31      g112(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n135_));
  INV        g113(.A(i_13_), .Y(new_new_n136_));
  NO2        g114(.A(i_12_), .B(new_new_n136_), .Y(new_new_n137_));
  INV        g115(.A(i_12_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n42_), .B(new_new_n138_), .Y(new_new_n139_));
  NO3        g117(.A(new_new_n35_), .B(i_8_), .C(i_10_), .Y(new_new_n140_));
  NA2        g118(.A(i_2_), .B(i_1_), .Y(new_new_n141_));
  NO3        g119(.A(i_11_), .B(i_7_), .C(new_new_n36_), .Y(new_new_n142_));
  NAi21      g120(.An(i_4_), .B(i_3_), .Y(new_new_n143_));
  NOi41      g121(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n144_));
  NO2        g122(.A(i_11_), .B(new_new_n136_), .Y(new_new_n145_));
  NOi21      g123(.An(i_1_), .B(i_6_), .Y(new_new_n146_));
  NAi21      g124(.An(i_3_), .B(i_7_), .Y(new_new_n147_));
  NA2        g125(.A(new_new_n138_), .B(i_9_), .Y(new_new_n148_));
  OR4        g126(.A(new_new_n148_), .B(new_new_n147_), .C(new_new_n146_), .D(new_new_n125_), .Y(new_new_n149_));
  NA2        g127(.A(new_new_n63_), .B(i_5_), .Y(new_new_n150_));
  NA2        g128(.A(i_3_), .B(i_9_), .Y(new_new_n151_));
  NAi21      g129(.An(i_7_), .B(i_10_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n152_), .B(new_new_n151_), .Y(new_new_n153_));
  NA3        g131(.A(new_new_n153_), .B(new_new_n150_), .C(new_new_n55_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n154_), .B(new_new_n149_), .Y(new_new_n155_));
  INV        g133(.A(new_new_n113_), .Y(new_new_n156_));
  NA2        g134(.A(new_new_n138_), .B(i_13_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(new_new_n64_), .Y(new_new_n158_));
  AOI220     g136(.A0(new_new_n158_), .A1(new_new_n156_), .B0(new_new_n155_), .B1(new_new_n145_), .Y(new_new_n159_));
  NA2        g137(.A(i_12_), .B(i_6_), .Y(new_new_n160_));
  OR2        g138(.A(i_13_), .B(i_9_), .Y(new_new_n161_));
  NO2        g139(.A(new_new_n143_), .B(i_2_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n145_), .B(i_9_), .Y(new_new_n163_));
  NO3        g141(.A(i_12_), .B(new_new_n136_), .C(new_new_n36_), .Y(new_new_n164_));
  AN2        g142(.A(i_3_), .B(i_10_), .Y(new_new_n165_));
  NO2        g143(.A(i_5_), .B(new_new_n36_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n44_), .B(new_new_n26_), .Y(new_new_n167_));
  NO3        g145(.A(new_new_n42_), .B(i_13_), .C(i_9_), .Y(new_new_n168_));
  NO2        g146(.A(i_2_), .B(i_3_), .Y(new_new_n169_));
  NO2        g147(.A(i_12_), .B(i_10_), .Y(new_new_n170_));
  NO2        g148(.A(i_1_), .B(i_7_), .Y(new_new_n171_));
  NOi21      g149(.An(new_new_n118_), .B(new_new_n88_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n172_), .B(new_new_n99_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(i_3_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n128_), .B(i_9_), .Y(new_new_n175_));
  NA2        g153(.A(new_new_n175_), .B(new_new_n131_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n176_), .B(new_new_n44_), .Y(new_new_n177_));
  INV        g155(.A(new_new_n177_), .Y(new_new_n178_));
  AOI210     g156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(new_new_n121_), .Y(new_new_n179_));
  INV        g157(.A(new_new_n179_), .Y(new_new_n180_));
  NOi32      g158(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n181_));
  INV        g159(.A(new_new_n181_), .Y(new_new_n182_));
  NOi32      g160(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n183_));
  NO2        g161(.A(i_1_), .B(new_new_n85_), .Y(new_new_n184_));
  NAi21      g162(.An(i_3_), .B(i_4_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(i_9_), .Y(new_new_n186_));
  AN2        g164(.A(i_6_), .B(i_7_), .Y(new_new_n187_));
  OAI210     g165(.A0(new_new_n187_), .A1(new_new_n184_), .B0(new_new_n186_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n185_), .B(i_10_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n188_), .B(new_new_n125_), .Y(new_new_n190_));
  AOI220     g168(.A0(new_new_n189_), .A1(new_new_n171_), .B0(new_new_n140_), .B1(new_new_n126_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n191_), .B(i_5_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n192_), .B(new_new_n190_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n193_), .B(new_new_n182_), .Y(new_new_n194_));
  AN2        g172(.A(i_12_), .B(i_5_), .Y(new_new_n195_));
  NO2        g173(.A(i_11_), .B(i_6_), .Y(new_new_n196_));
  NO2        g174(.A(i_5_), .B(i_10_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n36_), .B(new_new_n25_), .Y(new_new_n198_));
  NO3        g176(.A(i_1_), .B(i_12_), .C(new_new_n72_), .Y(new_new_n199_));
  NO2        g177(.A(i_0_), .B(i_11_), .Y(new_new_n200_));
  BUFFER     g178(.A(i_6_), .Y(new_new_n201_));
  NAi21      g179(.An(i_9_), .B(i_4_), .Y(new_new_n202_));
  OR2        g180(.A(i_13_), .B(i_10_), .Y(new_new_n203_));
  NO3        g181(.A(new_new_n203_), .B(new_new_n96_), .C(new_new_n202_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n205_));
  NA2        g183(.A(new_new_n164_), .B(new_new_n205_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n206_), .B(new_new_n172_), .Y(new_new_n207_));
  NA2        g185(.A(new_new_n128_), .B(i_10_), .Y(new_new_n208_));
  NA3        g186(.A(new_new_n150_), .B(new_new_n55_), .C(i_2_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n210_));
  INV        g188(.A(new_new_n210_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(new_new_n163_), .Y(new_new_n212_));
  NO3        g190(.A(new_new_n212_), .B(new_new_n207_), .C(new_new_n194_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n63_), .B(i_13_), .Y(new_new_n214_));
  NO3        g192(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n215_));
  NA2        g193(.A(new_new_n160_), .B(new_new_n84_), .Y(new_new_n216_));
  NA2        g194(.A(i_8_), .B(i_9_), .Y(new_new_n217_));
  NO2        g195(.A(i_7_), .B(i_2_), .Y(new_new_n218_));
  OR2        g196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n164_), .B(new_new_n131_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  NA2        g199(.A(new_new_n145_), .B(new_new_n166_), .Y(new_new_n222_));
  NO3        g200(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n223_));
  INV        g201(.A(new_new_n223_), .Y(new_new_n224_));
  NA3        g202(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n225_));
  NA4        g203(.A(new_new_n115_), .B(new_new_n95_), .C(new_new_n68_), .D(new_new_n23_), .Y(new_new_n226_));
  OAI220     g204(.A0(new_new_n226_), .A1(new_new_n225_), .B0(new_new_n224_), .B1(new_new_n222_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n221_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n83_), .B(i_13_), .Y(new_new_n229_));
  NO2        g207(.A(i_11_), .B(i_1_), .Y(new_new_n230_));
  NA3        g208(.A(new_new_n144_), .B(new_new_n123_), .C(new_new_n105_), .Y(new_new_n231_));
  NA2        g209(.A(new_new_n44_), .B(new_new_n42_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n119_), .B(i_3_), .Y(new_new_n233_));
  NAi31      g211(.An(new_new_n232_), .B(new_new_n233_), .C(new_new_n137_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n234_), .B(new_new_n231_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n235_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n215_), .B(new_new_n195_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n223_), .B(new_new_n197_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n27_), .B(i_10_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n168_), .B(new_new_n140_), .Y(new_new_n240_));
  OAI220     g218(.A0(new_new_n240_), .A1(new_new_n209_), .B0(new_new_n239_), .B1(new_new_n229_), .Y(new_new_n241_));
  INV        g219(.A(new_new_n241_), .Y(new_new_n242_));
  NA3        g220(.A(new_new_n242_), .B(new_new_n236_), .C(new_new_n228_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n195_), .B(new_new_n136_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n187_), .B(new_new_n183_), .Y(new_new_n245_));
  OR2        g223(.A(new_new_n244_), .B(new_new_n245_), .Y(new_new_n246_));
  AOI210     g224(.A0(new_new_n38_), .A1(i_13_), .B0(new_new_n204_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n247_), .B(new_new_n246_), .Y(new_new_n248_));
  NA3        g226(.A(new_new_n134_), .B(new_new_n61_), .C(new_new_n42_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n164_), .B(new_new_n70_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n249_), .B(new_new_n250_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n203_), .B(i_1_), .Y(new_new_n252_));
  NOi31      g230(.An(new_new_n252_), .B(new_new_n216_), .C(new_new_n63_), .Y(new_new_n253_));
  NOi21      g231(.An(i_10_), .B(i_6_), .Y(new_new_n254_));
  OR2        g232(.A(i_2_), .B(i_5_), .Y(new_new_n255_));
  NO3        g233(.A(new_new_n251_), .B(new_new_n248_), .C(new_new_n243_), .Y(new_new_n256_));
  NA4        g234(.A(new_new_n256_), .B(new_new_n213_), .C(new_new_n180_), .D(new_new_n159_), .Y(ori7));
  NO2        g235(.A(new_new_n79_), .B(new_new_n49_), .Y(new_new_n258_));
  INV        g236(.A(i_11_), .Y(new_new_n259_));
  NA3        g237(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n138_), .B(i_4_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n261_), .B(i_8_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n89_), .B(new_new_n260_), .Y(new_new_n263_));
  NA2        g241(.A(i_2_), .B(new_new_n72_), .Y(new_new_n264_));
  OAI210     g242(.A0(new_new_n73_), .A1(new_new_n129_), .B0(new_new_n130_), .Y(new_new_n265_));
  INV        g243(.A(new_new_n165_), .Y(new_new_n266_));
  OAI220     g244(.A0(new_new_n266_), .A1(new_new_n264_), .B0(new_new_n265_), .B1(i_13_), .Y(new_new_n267_));
  NO3        g245(.A(new_new_n267_), .B(new_new_n263_), .C(new_new_n258_), .Y(new_new_n268_));
  AOI210     g246(.A0(new_new_n103_), .A1(new_new_n53_), .B0(i_10_), .Y(new_new_n269_));
  AOI210     g247(.A0(new_new_n269_), .A1(new_new_n138_), .B0(new_new_n120_), .Y(new_new_n270_));
  OR2        g248(.A(i_6_), .B(i_10_), .Y(new_new_n271_));
  OR3        g249(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n272_));
  OR2        g250(.A(new_new_n270_), .B(new_new_n161_), .Y(new_new_n273_));
  AOI210     g251(.A0(new_new_n273_), .A1(new_new_n268_), .B0(new_new_n54_), .Y(new_new_n274_));
  NOi21      g252(.An(i_11_), .B(i_7_), .Y(new_new_n275_));
  AO210      g253(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(new_new_n275_), .Y(new_new_n277_));
  NA2        g255(.A(new_new_n277_), .B(new_new_n132_), .Y(new_new_n278_));
  NA3        g256(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n278_), .B(new_new_n54_), .Y(new_new_n280_));
  OR2        g258(.A(new_new_n191_), .B(new_new_n40_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n137_), .B(new_new_n54_), .Y(new_new_n282_));
  NO2        g260(.A(i_1_), .B(i_12_), .Y(new_new_n283_));
  NA2        g261(.A(new_new_n282_), .B(new_new_n281_), .Y(new_new_n284_));
  OAI210     g262(.A0(new_new_n284_), .A1(new_new_n280_), .B0(i_6_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n279_), .B(new_new_n92_), .Y(new_new_n286_));
  NO3        g264(.A(new_new_n271_), .B(i_7_), .C(new_new_n23_), .Y(new_new_n287_));
  AOI210     g265(.A0(i_1_), .A1(new_new_n153_), .B0(new_new_n287_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n288_), .B(new_new_n42_), .Y(new_new_n289_));
  INV        g267(.A(i_2_), .Y(new_new_n290_));
  NA2        g268(.A(new_new_n108_), .B(i_9_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n291_), .B(new_new_n290_), .Y(new_new_n292_));
  AOI210     g270(.A0(new_new_n230_), .A1(new_new_n205_), .B0(new_new_n142_), .Y(new_new_n293_));
  NO2        g271(.A(new_new_n293_), .B(new_new_n264_), .Y(new_new_n294_));
  OR2        g272(.A(new_new_n294_), .B(new_new_n292_), .Y(new_new_n295_));
  NO3        g273(.A(new_new_n295_), .B(new_new_n289_), .C(new_new_n286_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n138_), .B(new_new_n85_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n297_), .B(new_new_n275_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n298_), .B(i_1_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n299_), .B(new_new_n272_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n202_), .B(new_new_n72_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n300_), .B(new_new_n44_), .Y(new_new_n302_));
  NO2        g280(.A(i_7_), .B(new_new_n42_), .Y(new_new_n303_));
  NO3        g281(.A(new_new_n303_), .B(new_new_n167_), .C(new_new_n139_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n96_), .B(new_new_n36_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n305_), .B(i_6_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n72_), .B(i_9_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n307_), .B(new_new_n54_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n308_), .B(new_new_n283_), .Y(new_new_n309_));
  NO4        g287(.A(new_new_n309_), .B(new_new_n306_), .C(new_new_n304_), .D(i_4_), .Y(new_new_n310_));
  INV        g288(.A(new_new_n310_), .Y(new_new_n311_));
  NA4        g289(.A(new_new_n311_), .B(new_new_n302_), .C(new_new_n296_), .D(new_new_n285_), .Y(new_new_n312_));
  INV        g290(.A(i_1_), .Y(new_new_n313_));
  OR2        g291(.A(i_11_), .B(i_7_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n49_), .B(i_12_), .Y(new_new_n315_));
  INV        g293(.A(new_new_n315_), .Y(new_new_n316_));
  NA2        g294(.A(i_7_), .B(new_new_n301_), .Y(new_new_n317_));
  OAI220     g295(.A0(new_new_n317_), .A1(new_new_n40_), .B0(new_new_n316_), .B1(new_new_n79_), .Y(new_new_n318_));
  INV        g296(.A(new_new_n318_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n102_), .B(i_13_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(new_new_n313_), .Y(new_new_n321_));
  INV        g299(.A(i_7_), .Y(new_new_n322_));
  AOI220     g300(.A0(new_new_n196_), .A1(new_new_n454_), .B0(new_new_n78_), .B1(new_new_n86_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n323_), .B(new_new_n262_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n324_), .B(new_new_n321_), .Y(new_new_n325_));
  OR2        g303(.A(i_11_), .B(i_6_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n261_), .B(i_7_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(new_new_n326_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n328_), .B(new_new_n54_), .Y(new_new_n329_));
  NO2        g307(.A(i_2_), .B(i_12_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n184_), .B(new_new_n330_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n186_), .B(new_new_n184_), .Y(new_new_n332_));
  NA2        g310(.A(new_new_n332_), .B(new_new_n331_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n333_), .B(new_new_n43_), .Y(new_new_n334_));
  NA4        g312(.A(new_new_n334_), .B(new_new_n329_), .C(new_new_n325_), .D(new_new_n319_), .Y(new_new_n335_));
  OR3        g313(.A(new_new_n335_), .B(new_new_n312_), .C(new_new_n274_), .Y(ori5));
  NA2        g314(.A(new_new_n298_), .B(new_new_n162_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n24_), .B(new_new_n330_), .C(new_new_n92_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n262_), .B(i_11_), .Y(new_new_n339_));
  NA2        g317(.A(new_new_n73_), .B(new_new_n339_), .Y(new_new_n340_));
  NA3        g318(.A(new_new_n340_), .B(new_new_n338_), .C(new_new_n337_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n99_), .B(new_new_n23_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  INV        g321(.A(new_new_n123_), .Y(new_new_n344_));
  INV        g322(.A(new_new_n144_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n345_), .B(new_new_n344_), .Y(new_new_n346_));
  INV        g324(.A(new_new_n346_), .Y(new_new_n347_));
  NO3        g325(.A(new_new_n276_), .B(new_new_n37_), .C(new_new_n26_), .Y(new_new_n348_));
  OA210      g326(.A0(new_new_n277_), .A1(new_new_n101_), .B0(i_13_), .Y(new_new_n349_));
  NA3        g327(.A(i_2_), .B(new_new_n165_), .C(new_new_n99_), .Y(new_new_n350_));
  NO4        g328(.A(new_new_n453_), .B(new_new_n117_), .C(new_new_n349_), .D(new_new_n348_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n53_), .B(i_12_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n352_), .B(new_new_n101_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n353_), .B(new_new_n259_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n354_), .B(new_new_n35_), .Y(new_new_n355_));
  NA4        g333(.A(new_new_n355_), .B(new_new_n351_), .C(new_new_n347_), .D(new_new_n343_), .Y(ori6));
  NO2        g334(.A(new_new_n135_), .B(new_new_n232_), .Y(new_new_n357_));
  INV        g335(.A(new_new_n170_), .Y(new_new_n358_));
  NA2        g336(.A(new_new_n64_), .B(new_new_n104_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n146_), .B(i_9_), .Y(new_new_n361_));
  NA2        g339(.A(new_new_n361_), .B(new_new_n352_), .Y(new_new_n362_));
  AOI210     g340(.A0(new_new_n362_), .A1(new_new_n245_), .B0(new_new_n125_), .Y(new_new_n363_));
  NAi32      g341(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n326_), .B(new_new_n364_), .Y(new_new_n365_));
  OR3        g343(.A(new_new_n365_), .B(new_new_n363_), .C(new_new_n360_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n314_), .B(i_2_), .Y(new_new_n367_));
  BUFFER     g345(.A(new_new_n277_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n368_), .B(new_new_n116_), .Y(new_new_n369_));
  OR2        g347(.A(new_new_n238_), .B(new_new_n35_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n370_), .B(new_new_n369_), .Y(new_new_n371_));
  NA2        g349(.A(new_new_n357_), .B(new_new_n322_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n372_), .B(new_new_n265_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n271_), .B(new_new_n86_), .Y(new_new_n374_));
  OAI210     g352(.A0(new_new_n374_), .A1(new_new_n94_), .B0(new_new_n200_), .Y(new_new_n375_));
  NA3        g353(.A(new_new_n452_), .B(new_new_n170_), .C(i_7_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n377_));
  NO4        g355(.A(new_new_n377_), .B(new_new_n373_), .C(new_new_n371_), .D(new_new_n366_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n378_), .B(new_new_n193_), .Y(ori3));
  NA2        g357(.A(i_12_), .B(i_10_), .Y(new_new_n380_));
  NO2        g358(.A(i_11_), .B(new_new_n138_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n265_), .B(new_new_n188_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n382_), .B(new_new_n39_), .Y(new_new_n383_));
  NOi21      g361(.An(new_new_n83_), .B(new_new_n25_), .Y(new_new_n384_));
  AN2        g362(.A(new_new_n216_), .B(new_new_n50_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n386_));
  AOI210     g364(.A0(new_new_n386_), .A1(new_new_n383_), .B0(new_new_n45_), .Y(new_new_n387_));
  NO3        g365(.A(new_new_n195_), .B(new_new_n37_), .C(i_0_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n125_), .B(new_new_n254_), .Y(new_new_n389_));
  NOi21      g367(.An(new_new_n389_), .B(new_new_n388_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n54_), .Y(new_new_n391_));
  NOi21      g369(.An(i_5_), .B(i_9_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n392_), .B(new_new_n214_), .Y(new_new_n393_));
  BUFFER     g371(.A(new_new_n160_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n394_), .B(new_new_n230_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n395_), .B(new_new_n393_), .Y(new_new_n396_));
  NO3        g374(.A(new_new_n396_), .B(new_new_n391_), .C(new_new_n387_), .Y(new_new_n397_));
  NO4        g375(.A(new_new_n255_), .B(i_12_), .C(new_new_n203_), .D(new_new_n201_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n398_), .B(i_11_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n148_), .B(new_new_n118_), .Y(new_new_n400_));
  NA2        g378(.A(i_0_), .B(i_10_), .Y(new_new_n401_));
  AN2        g379(.A(new_new_n400_), .B(i_6_), .Y(new_new_n402_));
  INV        g380(.A(new_new_n402_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n403_), .B(new_new_n399_), .Y(new_new_n404_));
  NA2        g382(.A(i_11_), .B(i_9_), .Y(new_new_n405_));
  NO3        g383(.A(i_12_), .B(new_new_n405_), .C(new_new_n264_), .Y(new_new_n406_));
  AN2        g384(.A(new_new_n406_), .B(i_5_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n198_), .B(new_new_n124_), .Y(new_new_n408_));
  INV        g386(.A(new_new_n408_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n405_), .B(new_new_n63_), .Y(new_new_n410_));
  INV        g388(.A(new_new_n199_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(new_new_n393_), .Y(new_new_n412_));
  NO3        g390(.A(new_new_n412_), .B(new_new_n409_), .C(new_new_n407_), .Y(new_new_n413_));
  INV        g391(.A(new_new_n413_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n380_), .B(new_new_n169_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(new_new_n410_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n246_), .B(new_new_n416_), .Y(new_new_n417_));
  NO3        g395(.A(new_new_n417_), .B(new_new_n414_), .C(new_new_n404_), .Y(new_new_n418_));
  NO3        g396(.A(new_new_n401_), .B(new_new_n392_), .C(new_new_n127_), .Y(new_new_n419_));
  AOI220     g397(.A0(new_new_n419_), .A1(i_11_), .B0(new_new_n253_), .B1(new_new_n64_), .Y(new_new_n420_));
  NO3        g398(.A(new_new_n133_), .B(new_new_n195_), .C(i_0_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n421_), .B(i_13_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n422_), .B(new_new_n420_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n237_), .B(new_new_n231_), .Y(new_new_n424_));
  INV        g402(.A(new_new_n424_), .Y(new_new_n425_));
  NA3        g403(.A(new_new_n197_), .B(new_new_n123_), .C(new_new_n122_), .Y(new_new_n426_));
  INV        g404(.A(new_new_n426_), .Y(new_new_n427_));
  NO3        g405(.A(new_new_n405_), .B(new_new_n134_), .C(new_new_n127_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n428_), .B(new_new_n427_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n425_), .Y(new_new_n430_));
  NO2        g408(.A(new_new_n72_), .B(i_5_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n381_), .B(new_new_n93_), .Y(new_new_n432_));
  INV        g410(.A(new_new_n432_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n433_), .B(new_new_n431_), .Y(new_new_n434_));
  NAi21      g412(.An(new_new_n142_), .B(new_new_n143_), .Y(new_new_n435_));
  NO4        g413(.A(new_new_n141_), .B(new_new_n133_), .C(i_0_), .D(i_12_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n436_), .B(new_new_n435_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n437_), .B(new_new_n434_), .Y(new_new_n438_));
  NO3        g416(.A(new_new_n438_), .B(new_new_n430_), .C(new_new_n423_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n367_), .B(new_new_n36_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n270_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n441_), .B(new_new_n132_), .Y(new_new_n442_));
  NA2        g420(.A(i_2_), .B(i_10_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n60_), .B(new_new_n443_), .Y(new_new_n444_));
  AOI210     g422(.A0(new_new_n444_), .A1(new_new_n45_), .B0(new_new_n398_), .Y(new_new_n445_));
  AOI210     g423(.A0(new_new_n445_), .A1(new_new_n442_), .B0(new_new_n63_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n191_), .B(new_new_n344_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n447_), .B(new_new_n446_), .Y(new_new_n448_));
  NA4        g426(.A(new_new_n448_), .B(new_new_n439_), .C(new_new_n418_), .D(new_new_n397_), .Y(ori4));
  INV        g427(.A(new_new_n255_), .Y(new_new_n452_));
  INV        g428(.A(new_new_n350_), .Y(new_new_n453_));
  INV        g429(.A(i_1_), .Y(new_new_n454_));
endmodule


