//Benchmark atmr_misex3_1774_0.0625

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1468_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  NA3        o0002(.A(e), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n31_));
  NOi32      o0003(.An(m), .Bn(l), .C(n), .Y(ori_ori_n32_));
  NOi32      o0004(.An(i), .Bn(g), .C(h), .Y(ori_ori_n33_));
  NA2        o0005(.A(ori_ori_n33_), .B(ori_ori_n32_), .Y(ori_ori_n34_));
  AN2        o0006(.A(m), .B(l), .Y(ori_ori_n35_));
  NOi32      o0007(.An(j), .Bn(g), .C(k), .Y(ori_ori_n36_));
  NA2        o0008(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n37_));
  NO2        o0009(.A(ori_ori_n37_), .B(n), .Y(ori_ori_n38_));
  INV        o0010(.A(h), .Y(ori_ori_n39_));
  NAi21      o0011(.An(j), .B(l), .Y(ori_ori_n40_));
  NAi31      o0012(.An(n), .B(m), .C(l), .Y(ori_ori_n41_));
  INV        o0013(.A(i), .Y(ori_ori_n42_));
  AN2        o0014(.A(h), .B(g), .Y(ori_ori_n43_));
  NA2        o0015(.A(ori_ori_n43_), .B(ori_ori_n42_), .Y(ori_ori_n44_));
  NO2        o0016(.A(ori_ori_n44_), .B(ori_ori_n41_), .Y(ori_ori_n45_));
  NAi21      o0017(.An(n), .B(m), .Y(ori_ori_n46_));
  NOi32      o0018(.An(k), .Bn(h), .C(l), .Y(ori_ori_n47_));
  NOi32      o0019(.An(k), .Bn(h), .C(g), .Y(ori_ori_n48_));
  INV        o0020(.A(ori_ori_n48_), .Y(ori_ori_n49_));
  NO2        o0021(.A(ori_ori_n49_), .B(ori_ori_n46_), .Y(ori_ori_n50_));
  NO3        o0022(.A(ori_ori_n50_), .B(ori_ori_n45_), .C(ori_ori_n38_), .Y(ori_ori_n51_));
  AOI210     o0023(.A0(ori_ori_n51_), .A1(ori_ori_n34_), .B0(ori_ori_n31_), .Y(ori_ori_n52_));
  INV        o0024(.A(c), .Y(ori_ori_n53_));
  NA2        o0025(.A(e), .B(b), .Y(ori_ori_n54_));
  NO2        o0026(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  INV        o0027(.A(d), .Y(ori_ori_n56_));
  NA2        o0028(.A(g), .B(ori_ori_n56_), .Y(ori_ori_n57_));
  NAi21      o0029(.An(i), .B(h), .Y(ori_ori_n58_));
  NAi31      o0030(.An(i), .B(l), .C(j), .Y(ori_ori_n59_));
  NAi41      o0031(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n60_));
  NA2        o0032(.A(g), .B(f), .Y(ori_ori_n61_));
  NO2        o0033(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n62_));
  NAi32      o0034(.An(n), .Bn(k), .C(m), .Y(ori_ori_n63_));
  NAi31      o0035(.An(l), .B(m), .C(k), .Y(ori_ori_n64_));
  NAi21      o0036(.An(e), .B(h), .Y(ori_ori_n65_));
  NAi41      o0037(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n66_));
  INV        o0038(.A(m), .Y(ori_ori_n67_));
  NOi21      o0039(.An(k), .B(l), .Y(ori_ori_n68_));
  NA2        o0040(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  AN4        o0041(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n70_));
  NOi31      o0042(.An(h), .B(g), .C(f), .Y(ori_ori_n71_));
  NA2        o0043(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n72_));
  NAi32      o0044(.An(m), .Bn(k), .C(j), .Y(ori_ori_n73_));
  NOi32      o0045(.An(h), .Bn(g), .C(f), .Y(ori_ori_n74_));
  NA2        o0046(.A(ori_ori_n74_), .B(ori_ori_n70_), .Y(ori_ori_n75_));
  OA220      o0047(.A0(ori_ori_n75_), .A1(ori_ori_n73_), .B0(ori_ori_n72_), .B1(ori_ori_n69_), .Y(ori_ori_n76_));
  INV        o0048(.A(ori_ori_n76_), .Y(ori_ori_n77_));
  INV        o0049(.A(n), .Y(ori_ori_n78_));
  NOi32      o0050(.An(e), .Bn(b), .C(d), .Y(ori_ori_n79_));
  NA2        o0051(.A(ori_ori_n79_), .B(ori_ori_n78_), .Y(ori_ori_n80_));
  INV        o0052(.A(j), .Y(ori_ori_n81_));
  AN3        o0053(.A(m), .B(k), .C(i), .Y(ori_ori_n82_));
  NA3        o0054(.A(ori_ori_n82_), .B(ori_ori_n81_), .C(g), .Y(ori_ori_n83_));
  NO2        o0055(.A(ori_ori_n83_), .B(f), .Y(ori_ori_n84_));
  NAi32      o0056(.An(g), .Bn(f), .C(h), .Y(ori_ori_n85_));
  NAi31      o0057(.An(j), .B(m), .C(l), .Y(ori_ori_n86_));
  NO2        o0058(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n87_));
  NA2        o0059(.A(m), .B(l), .Y(ori_ori_n88_));
  NAi31      o0060(.An(k), .B(j), .C(g), .Y(ori_ori_n89_));
  NO3        o0061(.A(ori_ori_n89_), .B(ori_ori_n88_), .C(f), .Y(ori_ori_n90_));
  AN2        o0062(.A(j), .B(g), .Y(ori_ori_n91_));
  NOi32      o0063(.An(m), .Bn(l), .C(i), .Y(ori_ori_n92_));
  NOi21      o0064(.An(g), .B(i), .Y(ori_ori_n93_));
  NOi32      o0065(.An(m), .Bn(j), .C(k), .Y(ori_ori_n94_));
  AOI220     o0066(.A0(ori_ori_n94_), .A1(ori_ori_n93_), .B0(ori_ori_n92_), .B1(ori_ori_n91_), .Y(ori_ori_n95_));
  NO2        o0067(.A(ori_ori_n95_), .B(f), .Y(ori_ori_n96_));
  NAi41      o0068(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n97_));
  AN2        o0069(.A(e), .B(b), .Y(ori_ori_n98_));
  NOi31      o0070(.An(c), .B(h), .C(f), .Y(ori_ori_n99_));
  NA2        o0071(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  NO2        o0072(.A(ori_ori_n100_), .B(ori_ori_n97_), .Y(ori_ori_n101_));
  NOi21      o0073(.An(g), .B(f), .Y(ori_ori_n102_));
  NOi21      o0074(.An(i), .B(h), .Y(ori_ori_n103_));
  NA3        o0075(.A(ori_ori_n103_), .B(ori_ori_n102_), .C(ori_ori_n35_), .Y(ori_ori_n104_));
  INV        o0076(.A(a), .Y(ori_ori_n105_));
  NA2        o0077(.A(ori_ori_n98_), .B(ori_ori_n105_), .Y(ori_ori_n106_));
  INV        o0078(.A(l), .Y(ori_ori_n107_));
  NOi21      o0079(.An(m), .B(n), .Y(ori_ori_n108_));
  AN2        o0080(.A(k), .B(h), .Y(ori_ori_n109_));
  INV        o0081(.A(b), .Y(ori_ori_n110_));
  NA2        o0082(.A(l), .B(j), .Y(ori_ori_n111_));
  AN2        o0083(.A(k), .B(i), .Y(ori_ori_n112_));
  NA2        o0084(.A(g), .B(e), .Y(ori_ori_n113_));
  NOi32      o0085(.An(c), .Bn(a), .C(d), .Y(ori_ori_n114_));
  NA2        o0086(.A(ori_ori_n114_), .B(ori_ori_n108_), .Y(ori_ori_n115_));
  INV        o0087(.A(ori_ori_n101_), .Y(ori_ori_n116_));
  OAI210     o0088(.A0(ori_ori_n1224_), .A1(ori_ori_n80_), .B0(ori_ori_n116_), .Y(ori_ori_n117_));
  NOi31      o0089(.An(k), .B(m), .C(j), .Y(ori_ori_n118_));
  NA3        o0090(.A(ori_ori_n118_), .B(ori_ori_n71_), .C(ori_ori_n70_), .Y(ori_ori_n119_));
  NOi31      o0091(.An(k), .B(m), .C(i), .Y(ori_ori_n120_));
  NA3        o0092(.A(ori_ori_n120_), .B(ori_ori_n74_), .C(ori_ori_n70_), .Y(ori_ori_n121_));
  NA2        o0093(.A(ori_ori_n121_), .B(ori_ori_n119_), .Y(ori_ori_n122_));
  NAi21      o0094(.An(g), .B(h), .Y(ori_ori_n123_));
  NAi21      o0095(.An(m), .B(n), .Y(ori_ori_n124_));
  NAi41      o0096(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n125_));
  NAi31      o0097(.An(j), .B(k), .C(h), .Y(ori_ori_n126_));
  NO3        o0098(.A(ori_ori_n126_), .B(ori_ori_n125_), .C(ori_ori_n124_), .Y(ori_ori_n127_));
  INV        o0099(.A(ori_ori_n127_), .Y(ori_ori_n128_));
  NO2        o0100(.A(k), .B(j), .Y(ori_ori_n129_));
  NO2        o0101(.A(ori_ori_n129_), .B(ori_ori_n124_), .Y(ori_ori_n130_));
  AN2        o0102(.A(k), .B(j), .Y(ori_ori_n131_));
  NAi21      o0103(.An(c), .B(b), .Y(ori_ori_n132_));
  NA2        o0104(.A(f), .B(d), .Y(ori_ori_n133_));
  NO4        o0105(.A(ori_ori_n133_), .B(ori_ori_n132_), .C(ori_ori_n131_), .D(ori_ori_n123_), .Y(ori_ori_n134_));
  NA2        o0106(.A(h), .B(c), .Y(ori_ori_n135_));
  NAi31      o0107(.An(f), .B(e), .C(b), .Y(ori_ori_n136_));
  NA2        o0108(.A(ori_ori_n134_), .B(ori_ori_n130_), .Y(ori_ori_n137_));
  NA2        o0109(.A(d), .B(b), .Y(ori_ori_n138_));
  NAi21      o0110(.An(e), .B(f), .Y(ori_ori_n139_));
  NO2        o0111(.A(ori_ori_n139_), .B(ori_ori_n138_), .Y(ori_ori_n140_));
  NA2        o0112(.A(b), .B(a), .Y(ori_ori_n141_));
  NAi21      o0113(.An(e), .B(g), .Y(ori_ori_n142_));
  NAi21      o0114(.An(c), .B(d), .Y(ori_ori_n143_));
  NAi31      o0115(.An(l), .B(k), .C(h), .Y(ori_ori_n144_));
  NO2        o0116(.A(ori_ori_n124_), .B(ori_ori_n144_), .Y(ori_ori_n145_));
  NA2        o0117(.A(ori_ori_n145_), .B(ori_ori_n140_), .Y(ori_ori_n146_));
  NAi41      o0118(.An(ori_ori_n122_), .B(ori_ori_n146_), .C(ori_ori_n137_), .D(ori_ori_n128_), .Y(ori_ori_n147_));
  NAi31      o0119(.An(e), .B(f), .C(b), .Y(ori_ori_n148_));
  NOi21      o0120(.An(g), .B(d), .Y(ori_ori_n149_));
  NO2        o0121(.A(ori_ori_n149_), .B(ori_ori_n148_), .Y(ori_ori_n150_));
  NOi21      o0122(.An(h), .B(i), .Y(ori_ori_n151_));
  NOi21      o0123(.An(k), .B(m), .Y(ori_ori_n152_));
  NA3        o0124(.A(ori_ori_n152_), .B(ori_ori_n151_), .C(n), .Y(ori_ori_n153_));
  NOi21      o0125(.An(ori_ori_n150_), .B(ori_ori_n153_), .Y(ori_ori_n154_));
  NOi21      o0126(.An(h), .B(g), .Y(ori_ori_n155_));
  NO2        o0127(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n156_));
  NAi31      o0128(.An(l), .B(j), .C(h), .Y(ori_ori_n157_));
  INV        o0129(.A(ori_ori_n46_), .Y(ori_ori_n158_));
  NA2        o0130(.A(ori_ori_n158_), .B(ori_ori_n62_), .Y(ori_ori_n159_));
  NOi32      o0131(.An(n), .Bn(k), .C(m), .Y(ori_ori_n160_));
  INV        o0132(.A(ori_ori_n159_), .Y(ori_ori_n161_));
  NAi31      o0133(.An(d), .B(f), .C(c), .Y(ori_ori_n162_));
  NAi31      o0134(.An(e), .B(f), .C(c), .Y(ori_ori_n163_));
  NA2        o0135(.A(ori_ori_n163_), .B(ori_ori_n162_), .Y(ori_ori_n164_));
  NA2        o0136(.A(j), .B(h), .Y(ori_ori_n165_));
  OR3        o0137(.A(n), .B(m), .C(k), .Y(ori_ori_n166_));
  NO2        o0138(.A(ori_ori_n166_), .B(ori_ori_n165_), .Y(ori_ori_n167_));
  NAi32      o0139(.An(m), .Bn(k), .C(n), .Y(ori_ori_n168_));
  NO2        o0140(.A(ori_ori_n168_), .B(ori_ori_n165_), .Y(ori_ori_n169_));
  AOI220     o0141(.A0(ori_ori_n169_), .A1(ori_ori_n150_), .B0(ori_ori_n167_), .B1(ori_ori_n164_), .Y(ori_ori_n170_));
  NO2        o0142(.A(n), .B(m), .Y(ori_ori_n171_));
  NA2        o0143(.A(ori_ori_n171_), .B(ori_ori_n47_), .Y(ori_ori_n172_));
  NAi21      o0144(.An(f), .B(e), .Y(ori_ori_n173_));
  NA2        o0145(.A(d), .B(c), .Y(ori_ori_n174_));
  NO2        o0146(.A(ori_ori_n174_), .B(ori_ori_n173_), .Y(ori_ori_n175_));
  NOi21      o0147(.An(ori_ori_n175_), .B(ori_ori_n172_), .Y(ori_ori_n176_));
  NAi21      o0148(.An(h), .B(f), .Y(ori_ori_n177_));
  NOi32      o0149(.An(f), .Bn(c), .C(d), .Y(ori_ori_n178_));
  NOi32      o0150(.An(f), .Bn(c), .C(e), .Y(ori_ori_n179_));
  NO2        o0151(.A(ori_ori_n179_), .B(ori_ori_n178_), .Y(ori_ori_n180_));
  NO3        o0152(.A(n), .B(m), .C(j), .Y(ori_ori_n181_));
  NA2        o0153(.A(ori_ori_n181_), .B(ori_ori_n109_), .Y(ori_ori_n182_));
  AO210      o0154(.A0(ori_ori_n182_), .A1(ori_ori_n172_), .B0(ori_ori_n180_), .Y(ori_ori_n183_));
  NAi31      o0155(.An(ori_ori_n176_), .B(ori_ori_n183_), .C(ori_ori_n170_), .Y(ori_ori_n184_));
  OR4        o0156(.A(ori_ori_n184_), .B(ori_ori_n161_), .C(ori_ori_n154_), .D(ori_ori_n147_), .Y(ori_ori_n185_));
  NO4        o0157(.A(ori_ori_n185_), .B(ori_ori_n117_), .C(ori_ori_n77_), .D(ori_ori_n52_), .Y(ori_ori_n186_));
  NA3        o0158(.A(m), .B(ori_ori_n107_), .C(j), .Y(ori_ori_n187_));
  NAi31      o0159(.An(n), .B(h), .C(g), .Y(ori_ori_n188_));
  NO2        o0160(.A(ori_ori_n188_), .B(ori_ori_n187_), .Y(ori_ori_n189_));
  NOi32      o0161(.An(m), .Bn(k), .C(l), .Y(ori_ori_n190_));
  NA3        o0162(.A(ori_ori_n190_), .B(ori_ori_n81_), .C(g), .Y(ori_ori_n191_));
  NOi21      o0163(.An(k), .B(j), .Y(ori_ori_n192_));
  NA4        o0164(.A(ori_ori_n192_), .B(ori_ori_n108_), .C(i), .D(g), .Y(ori_ori_n193_));
  NA3        o0165(.A(ori_ori_n68_), .B(g), .C(ori_ori_n108_), .Y(ori_ori_n194_));
  NA2        o0166(.A(ori_ori_n194_), .B(ori_ori_n193_), .Y(ori_ori_n195_));
  NO2        o0167(.A(ori_ori_n195_), .B(ori_ori_n189_), .Y(ori_ori_n196_));
  NAi41      o0168(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n197_));
  INV        o0169(.A(ori_ori_n197_), .Y(ori_ori_n198_));
  INV        o0170(.A(f), .Y(ori_ori_n199_));
  INV        o0171(.A(g), .Y(ori_ori_n200_));
  NOi31      o0172(.An(i), .B(j), .C(h), .Y(ori_ori_n201_));
  NOi21      o0173(.An(l), .B(m), .Y(ori_ori_n202_));
  NA2        o0174(.A(ori_ori_n202_), .B(ori_ori_n201_), .Y(ori_ori_n203_));
  NO3        o0175(.A(ori_ori_n203_), .B(ori_ori_n200_), .C(ori_ori_n199_), .Y(ori_ori_n204_));
  NA2        o0176(.A(ori_ori_n204_), .B(ori_ori_n198_), .Y(ori_ori_n205_));
  OAI210     o0177(.A0(ori_ori_n196_), .A1(ori_ori_n31_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  NOi21      o0178(.An(n), .B(m), .Y(ori_ori_n207_));
  NOi32      o0179(.An(l), .Bn(i), .C(j), .Y(ori_ori_n208_));
  NA2        o0180(.A(ori_ori_n208_), .B(ori_ori_n207_), .Y(ori_ori_n209_));
  OA220      o0181(.A0(ori_ori_n209_), .A1(ori_ori_n100_), .B0(ori_ori_n73_), .B1(ori_ori_n72_), .Y(ori_ori_n210_));
  NAi21      o0182(.An(j), .B(h), .Y(ori_ori_n211_));
  XN2        o0183(.A(i), .B(h), .Y(ori_ori_n212_));
  NA2        o0184(.A(ori_ori_n212_), .B(ori_ori_n211_), .Y(ori_ori_n213_));
  NOi31      o0185(.An(k), .B(n), .C(m), .Y(ori_ori_n214_));
  NOi31      o0186(.An(ori_ori_n214_), .B(ori_ori_n174_), .C(ori_ori_n173_), .Y(ori_ori_n215_));
  NA2        o0187(.A(ori_ori_n215_), .B(ori_ori_n213_), .Y(ori_ori_n216_));
  NAi31      o0188(.An(f), .B(e), .C(c), .Y(ori_ori_n217_));
  NO4        o0189(.A(ori_ori_n217_), .B(ori_ori_n166_), .C(ori_ori_n165_), .D(ori_ori_n56_), .Y(ori_ori_n218_));
  NA4        o0190(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n219_));
  NAi32      o0191(.An(m), .Bn(i), .C(k), .Y(ori_ori_n220_));
  INV        o0192(.A(k), .Y(ori_ori_n221_));
  INV        o0193(.A(ori_ori_n218_), .Y(ori_ori_n222_));
  NAi21      o0194(.An(n), .B(a), .Y(ori_ori_n223_));
  NO2        o0195(.A(ori_ori_n223_), .B(ori_ori_n138_), .Y(ori_ori_n224_));
  NAi41      o0196(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n225_));
  NO2        o0197(.A(ori_ori_n225_), .B(e), .Y(ori_ori_n226_));
  NA2        o0198(.A(ori_ori_n226_), .B(ori_ori_n224_), .Y(ori_ori_n227_));
  AN4        o0199(.A(ori_ori_n227_), .B(ori_ori_n222_), .C(ori_ori_n216_), .D(ori_ori_n210_), .Y(ori_ori_n228_));
  NAi41      o0200(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n229_));
  NO2        o0201(.A(ori_ori_n229_), .B(ori_ori_n199_), .Y(ori_ori_n230_));
  NA2        o0202(.A(ori_ori_n152_), .B(ori_ori_n103_), .Y(ori_ori_n231_));
  NAi21      o0203(.An(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NO2        o0204(.A(n), .B(a), .Y(ori_ori_n233_));
  NAi31      o0205(.An(ori_ori_n225_), .B(ori_ori_n233_), .C(ori_ori_n98_), .Y(ori_ori_n234_));
  AN2        o0206(.A(ori_ori_n234_), .B(ori_ori_n232_), .Y(ori_ori_n235_));
  NAi21      o0207(.An(h), .B(i), .Y(ori_ori_n236_));
  NA2        o0208(.A(ori_ori_n171_), .B(k), .Y(ori_ori_n237_));
  NO2        o0209(.A(ori_ori_n237_), .B(ori_ori_n236_), .Y(ori_ori_n238_));
  NA2        o0210(.A(ori_ori_n238_), .B(ori_ori_n178_), .Y(ori_ori_n239_));
  NA2        o0211(.A(ori_ori_n239_), .B(ori_ori_n235_), .Y(ori_ori_n240_));
  NOi21      o0212(.An(g), .B(e), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n66_), .B(ori_ori_n67_), .Y(ori_ori_n242_));
  NOi32      o0214(.An(l), .Bn(j), .C(i), .Y(ori_ori_n243_));
  AOI210     o0215(.A0(ori_ori_n68_), .A1(ori_ori_n81_), .B0(ori_ori_n243_), .Y(ori_ori_n244_));
  NAi21      o0216(.An(f), .B(g), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(ori_ori_n60_), .Y(ori_ori_n246_));
  NOi31      o0218(.An(ori_ori_n228_), .B(ori_ori_n240_), .C(ori_ori_n206_), .Y(ori_ori_n247_));
  NA3        o0219(.A(ori_ori_n56_), .B(c), .C(b), .Y(ori_ori_n248_));
  NAi21      o0220(.An(h), .B(g), .Y(ori_ori_n249_));
  OR4        o0221(.A(ori_ori_n249_), .B(ori_ori_n248_), .C(ori_ori_n209_), .D(e), .Y(ori_ori_n250_));
  INV        o0222(.A(ori_ori_n231_), .Y(ori_ori_n251_));
  NAi31      o0223(.An(e), .B(d), .C(a), .Y(ori_ori_n252_));
  INV        o0224(.A(ori_ori_n250_), .Y(ori_ori_n253_));
  NA4        o0225(.A(ori_ori_n152_), .B(ori_ori_n74_), .C(ori_ori_n70_), .D(ori_ori_n111_), .Y(ori_ori_n254_));
  NA3        o0226(.A(ori_ori_n152_), .B(ori_ori_n151_), .C(ori_ori_n78_), .Y(ori_ori_n255_));
  NO2        o0227(.A(ori_ori_n255_), .B(ori_ori_n180_), .Y(ori_ori_n256_));
  NOi21      o0228(.An(ori_ori_n254_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  NA3        o0229(.A(e), .B(c), .C(b), .Y(ori_ori_n258_));
  NO2        o0230(.A(ori_ori_n57_), .B(ori_ori_n258_), .Y(ori_ori_n259_));
  NAi32      o0231(.An(k), .Bn(i), .C(j), .Y(ori_ori_n260_));
  NAi31      o0232(.An(h), .B(l), .C(i), .Y(ori_ori_n261_));
  NA3        o0233(.A(ori_ori_n261_), .B(ori_ori_n260_), .C(ori_ori_n157_), .Y(ori_ori_n262_));
  NOi21      o0234(.An(ori_ori_n262_), .B(ori_ori_n46_), .Y(ori_ori_n263_));
  OAI210     o0235(.A0(ori_ori_n246_), .A1(ori_ori_n259_), .B0(ori_ori_n263_), .Y(ori_ori_n264_));
  NAi21      o0236(.An(l), .B(k), .Y(ori_ori_n265_));
  NOi21      o0237(.An(l), .B(j), .Y(ori_ori_n266_));
  NAi32      o0238(.An(j), .Bn(h), .C(i), .Y(ori_ori_n267_));
  NAi21      o0239(.An(m), .B(l), .Y(ori_ori_n268_));
  NA2        o0240(.A(h), .B(g), .Y(ori_ori_n269_));
  NA2        o0241(.A(ori_ori_n160_), .B(ori_ori_n42_), .Y(ori_ori_n270_));
  NO2        o0242(.A(ori_ori_n270_), .B(ori_ori_n269_), .Y(ori_ori_n271_));
  NA2        o0243(.A(ori_ori_n271_), .B(ori_ori_n156_), .Y(ori_ori_n272_));
  NA3        o0244(.A(ori_ori_n272_), .B(ori_ori_n264_), .C(ori_ori_n257_), .Y(ori_ori_n273_));
  NO2        o0245(.A(ori_ori_n100_), .B(ori_ori_n97_), .Y(ori_ori_n274_));
  NAi32      o0246(.An(n), .Bn(m), .C(l), .Y(ori_ori_n275_));
  NO2        o0247(.A(ori_ori_n275_), .B(ori_ori_n267_), .Y(ori_ori_n276_));
  NA2        o0248(.A(ori_ori_n276_), .B(ori_ori_n175_), .Y(ori_ori_n277_));
  NAi31      o0249(.An(k), .B(l), .C(j), .Y(ori_ori_n278_));
  OAI210     o0250(.A0(ori_ori_n265_), .A1(j), .B0(ori_ori_n278_), .Y(ori_ori_n279_));
  NOi21      o0251(.An(ori_ori_n279_), .B(ori_ori_n113_), .Y(ori_ori_n280_));
  NO3        o0252(.A(ori_ori_n1223_), .B(ori_ori_n273_), .C(ori_ori_n253_), .Y(ori_ori_n281_));
  NA2        o0253(.A(ori_ori_n238_), .B(ori_ori_n179_), .Y(ori_ori_n282_));
  NAi21      o0254(.An(m), .B(k), .Y(ori_ori_n283_));
  NO2        o0255(.A(ori_ori_n212_), .B(ori_ori_n283_), .Y(ori_ori_n284_));
  NAi41      o0256(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n285_));
  NO2        o0257(.A(ori_ori_n285_), .B(ori_ori_n142_), .Y(ori_ori_n286_));
  NA2        o0258(.A(ori_ori_n286_), .B(ori_ori_n284_), .Y(ori_ori_n287_));
  NO4        o0259(.A(i), .B(ori_ori_n142_), .C(ori_ori_n66_), .D(ori_ori_n67_), .Y(ori_ori_n288_));
  NA2        o0260(.A(e), .B(c), .Y(ori_ori_n289_));
  NO3        o0261(.A(ori_ori_n289_), .B(n), .C(d), .Y(ori_ori_n290_));
  NOi21      o0262(.An(f), .B(h), .Y(ori_ori_n291_));
  NAi31      o0263(.An(d), .B(e), .C(b), .Y(ori_ori_n292_));
  NAi31      o0264(.An(ori_ori_n288_), .B(ori_ori_n287_), .C(ori_ori_n282_), .Y(ori_ori_n293_));
  NO4        o0265(.A(ori_ori_n285_), .B(ori_ori_n73_), .C(ori_ori_n65_), .D(ori_ori_n200_), .Y(ori_ori_n294_));
  NA2        o0266(.A(ori_ori_n233_), .B(ori_ori_n98_), .Y(ori_ori_n295_));
  NOi31      o0267(.An(l), .B(n), .C(m), .Y(ori_ori_n296_));
  NA2        o0268(.A(ori_ori_n296_), .B(ori_ori_n201_), .Y(ori_ori_n297_));
  NO2        o0269(.A(ori_ori_n297_), .B(ori_ori_n180_), .Y(ori_ori_n298_));
  OR2        o0270(.A(ori_ori_n298_), .B(ori_ori_n294_), .Y(ori_ori_n299_));
  NAi32      o0271(.An(m), .Bn(j), .C(k), .Y(ori_ori_n300_));
  NAi41      o0272(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n301_));
  NOi31      o0273(.An(j), .B(m), .C(k), .Y(ori_ori_n302_));
  NO2        o0274(.A(ori_ori_n118_), .B(ori_ori_n302_), .Y(ori_ori_n303_));
  AN3        o0275(.A(h), .B(g), .C(f), .Y(ori_ori_n304_));
  NOi32      o0276(.An(m), .Bn(j), .C(l), .Y(ori_ori_n305_));
  NO2        o0277(.A(ori_ori_n268_), .B(ori_ori_n267_), .Y(ori_ori_n306_));
  NA2        o0278(.A(ori_ori_n230_), .B(ori_ori_n306_), .Y(ori_ori_n307_));
  INV        o0279(.A(ori_ori_n220_), .Y(ori_ori_n308_));
  NA3        o0280(.A(ori_ori_n308_), .B(ori_ori_n304_), .C(ori_ori_n198_), .Y(ori_ori_n309_));
  NA2        o0281(.A(ori_ori_n309_), .B(ori_ori_n307_), .Y(ori_ori_n310_));
  NA3        o0282(.A(h), .B(g), .C(f), .Y(ori_ori_n311_));
  NO2        o0283(.A(ori_ori_n311_), .B(ori_ori_n69_), .Y(ori_ori_n312_));
  NA2        o0284(.A(ori_ori_n301_), .B(ori_ori_n197_), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n155_), .B(e), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n314_), .B(ori_ori_n40_), .Y(ori_ori_n315_));
  NA2        o0287(.A(ori_ori_n313_), .B(ori_ori_n312_), .Y(ori_ori_n316_));
  NOi32      o0288(.An(j), .Bn(g), .C(i), .Y(ori_ori_n317_));
  NA2        o0289(.A(ori_ori_n317_), .B(ori_ori_n108_), .Y(ori_ori_n318_));
  AO210      o0290(.A0(ori_ori_n106_), .A1(ori_ori_n31_), .B0(ori_ori_n318_), .Y(ori_ori_n319_));
  NOi32      o0291(.An(e), .Bn(b), .C(a), .Y(ori_ori_n320_));
  AN2        o0292(.A(l), .B(j), .Y(ori_ori_n321_));
  NO2        o0293(.A(ori_ori_n283_), .B(ori_ori_n321_), .Y(ori_ori_n322_));
  NO3        o0294(.A(ori_ori_n285_), .B(ori_ori_n65_), .C(ori_ori_n200_), .Y(ori_ori_n323_));
  NA3        o0295(.A(ori_ori_n194_), .B(ori_ori_n193_), .C(ori_ori_n34_), .Y(ori_ori_n324_));
  AOI220     o0296(.A0(ori_ori_n324_), .A1(ori_ori_n320_), .B0(ori_ori_n323_), .B1(ori_ori_n322_), .Y(ori_ori_n325_));
  NA2        o0297(.A(g), .B(k), .Y(ori_ori_n326_));
  NA3        o0298(.A(m), .B(ori_ori_n107_), .C(ori_ori_n199_), .Y(ori_ori_n327_));
  NA4        o0299(.A(ori_ori_n190_), .B(ori_ori_n81_), .C(g), .D(ori_ori_n199_), .Y(ori_ori_n328_));
  NAi41      o0300(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n329_));
  NA2        o0301(.A(ori_ori_n48_), .B(ori_ori_n108_), .Y(ori_ori_n330_));
  NO2        o0302(.A(ori_ori_n330_), .B(ori_ori_n329_), .Y(ori_ori_n331_));
  NA2        o0303(.A(ori_ori_n331_), .B(b), .Y(ori_ori_n332_));
  NA4        o0304(.A(ori_ori_n332_), .B(ori_ori_n325_), .C(ori_ori_n319_), .D(ori_ori_n316_), .Y(ori_ori_n333_));
  NO4        o0305(.A(ori_ori_n333_), .B(ori_ori_n310_), .C(ori_ori_n299_), .D(ori_ori_n293_), .Y(ori_ori_n334_));
  NA4        o0306(.A(ori_ori_n334_), .B(ori_ori_n281_), .C(ori_ori_n247_), .D(ori_ori_n186_), .Y(ori10));
  NA3        o0307(.A(m), .B(k), .C(i), .Y(ori_ori_n336_));
  NOi21      o0308(.An(e), .B(f), .Y(ori_ori_n337_));
  NO4        o0309(.A(ori_ori_n143_), .B(ori_ori_n337_), .C(n), .D(ori_ori_n105_), .Y(ori_ori_n338_));
  NAi31      o0310(.An(b), .B(f), .C(c), .Y(ori_ori_n339_));
  INV        o0311(.A(ori_ori_n339_), .Y(ori_ori_n340_));
  NOi32      o0312(.An(k), .Bn(h), .C(j), .Y(ori_ori_n341_));
  NA2        o0313(.A(ori_ori_n341_), .B(ori_ori_n207_), .Y(ori_ori_n342_));
  NA2        o0314(.A(ori_ori_n153_), .B(ori_ori_n342_), .Y(ori_ori_n343_));
  NA2        o0315(.A(ori_ori_n343_), .B(ori_ori_n340_), .Y(ori_ori_n344_));
  AN2        o0316(.A(j), .B(h), .Y(ori_ori_n345_));
  NO3        o0317(.A(n), .B(m), .C(k), .Y(ori_ori_n346_));
  NA2        o0318(.A(ori_ori_n346_), .B(ori_ori_n345_), .Y(ori_ori_n347_));
  NO3        o0319(.A(ori_ori_n347_), .B(ori_ori_n143_), .C(ori_ori_n199_), .Y(ori_ori_n348_));
  OR2        o0320(.A(m), .B(k), .Y(ori_ori_n349_));
  NO2        o0321(.A(ori_ori_n165_), .B(ori_ori_n349_), .Y(ori_ori_n350_));
  NA4        o0322(.A(n), .B(f), .C(c), .D(ori_ori_n110_), .Y(ori_ori_n351_));
  NOi21      o0323(.An(ori_ori_n350_), .B(ori_ori_n351_), .Y(ori_ori_n352_));
  NOi32      o0324(.An(d), .Bn(a), .C(c), .Y(ori_ori_n353_));
  NA2        o0325(.A(ori_ori_n353_), .B(ori_ori_n173_), .Y(ori_ori_n354_));
  NAi21      o0326(.An(i), .B(g), .Y(ori_ori_n355_));
  NAi31      o0327(.An(k), .B(m), .C(j), .Y(ori_ori_n356_));
  NO3        o0328(.A(ori_ori_n356_), .B(ori_ori_n355_), .C(n), .Y(ori_ori_n357_));
  NOi21      o0329(.An(ori_ori_n357_), .B(ori_ori_n354_), .Y(ori_ori_n358_));
  NO3        o0330(.A(ori_ori_n358_), .B(ori_ori_n352_), .C(ori_ori_n348_), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n351_), .B(ori_ori_n268_), .Y(ori_ori_n360_));
  NOi32      o0332(.An(f), .Bn(d), .C(c), .Y(ori_ori_n361_));
  AOI220     o0333(.A0(ori_ori_n361_), .A1(ori_ori_n276_), .B0(ori_ori_n360_), .B1(ori_ori_n201_), .Y(ori_ori_n362_));
  NA3        o0334(.A(ori_ori_n362_), .B(ori_ori_n359_), .C(ori_ori_n344_), .Y(ori_ori_n363_));
  NO2        o0335(.A(ori_ori_n56_), .B(ori_ori_n110_), .Y(ori_ori_n364_));
  NA2        o0336(.A(ori_ori_n233_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  INV        o0337(.A(e), .Y(ori_ori_n366_));
  AN2        o0338(.A(g), .B(e), .Y(ori_ori_n367_));
  NA3        o0339(.A(ori_ori_n367_), .B(ori_ori_n190_), .C(i), .Y(ori_ori_n368_));
  OAI210     o0340(.A0(ori_ori_n83_), .A1(ori_ori_n366_), .B0(ori_ori_n368_), .Y(ori_ori_n369_));
  NO2        o0341(.A(ori_ori_n95_), .B(ori_ori_n366_), .Y(ori_ori_n370_));
  NO2        o0342(.A(ori_ori_n370_), .B(ori_ori_n369_), .Y(ori_ori_n371_));
  NOi32      o0343(.An(h), .Bn(e), .C(g), .Y(ori_ori_n372_));
  NOi21      o0344(.An(g), .B(h), .Y(ori_ori_n373_));
  AN3        o0345(.A(m), .B(l), .C(i), .Y(ori_ori_n374_));
  NA3        o0346(.A(ori_ori_n374_), .B(ori_ori_n373_), .C(e), .Y(ori_ori_n375_));
  AN3        o0347(.A(h), .B(g), .C(e), .Y(ori_ori_n376_));
  AOI210     o0348(.A0(ori_ori_n375_), .A1(ori_ori_n371_), .B0(ori_ori_n365_), .Y(ori_ori_n377_));
  NAi31      o0349(.An(b), .B(c), .C(a), .Y(ori_ori_n378_));
  NO2        o0350(.A(ori_ori_n378_), .B(n), .Y(ori_ori_n379_));
  NA2        o0351(.A(ori_ori_n48_), .B(m), .Y(ori_ori_n380_));
  NO2        o0352(.A(ori_ori_n380_), .B(ori_ori_n139_), .Y(ori_ori_n381_));
  NO2        o0353(.A(ori_ori_n377_), .B(ori_ori_n363_), .Y(ori_ori_n382_));
  INV        o0354(.A(g), .Y(ori_ori_n383_));
  NOi21      o0355(.An(a), .B(n), .Y(ori_ori_n384_));
  NOi21      o0356(.An(d), .B(c), .Y(ori_ori_n385_));
  NA2        o0357(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n386_));
  NA3        o0358(.A(i), .B(g), .C(f), .Y(ori_ori_n387_));
  OR2        o0359(.A(ori_ori_n387_), .B(ori_ori_n64_), .Y(ori_ori_n388_));
  NA3        o0360(.A(ori_ori_n374_), .B(ori_ori_n373_), .C(ori_ori_n173_), .Y(ori_ori_n389_));
  AOI210     o0361(.A0(ori_ori_n389_), .A1(ori_ori_n388_), .B0(ori_ori_n386_), .Y(ori_ori_n390_));
  INV        o0362(.A(ori_ori_n390_), .Y(ori_ori_n391_));
  OR2        o0363(.A(n), .B(m), .Y(ori_ori_n392_));
  NO2        o0364(.A(ori_ori_n392_), .B(ori_ori_n144_), .Y(ori_ori_n393_));
  NO2        o0365(.A(ori_ori_n174_), .B(ori_ori_n139_), .Y(ori_ori_n394_));
  OAI210     o0366(.A0(ori_ori_n393_), .A1(ori_ori_n167_), .B0(ori_ori_n394_), .Y(ori_ori_n395_));
  INV        o0367(.A(ori_ori_n330_), .Y(ori_ori_n396_));
  NA3        o0368(.A(ori_ori_n396_), .B(ori_ori_n320_), .C(d), .Y(ori_ori_n397_));
  NO2        o0369(.A(ori_ori_n378_), .B(ori_ori_n46_), .Y(ori_ori_n398_));
  NAi21      o0370(.An(k), .B(j), .Y(ori_ori_n399_));
  NAi21      o0371(.An(e), .B(d), .Y(ori_ori_n400_));
  INV        o0372(.A(ori_ori_n400_), .Y(ori_ori_n401_));
  NO2        o0373(.A(ori_ori_n237_), .B(ori_ori_n199_), .Y(ori_ori_n402_));
  NA3        o0374(.A(ori_ori_n402_), .B(ori_ori_n401_), .C(ori_ori_n213_), .Y(ori_ori_n403_));
  NA3        o0375(.A(ori_ori_n403_), .B(ori_ori_n397_), .C(ori_ori_n395_), .Y(ori_ori_n404_));
  NO2        o0376(.A(ori_ori_n297_), .B(ori_ori_n199_), .Y(ori_ori_n405_));
  NA2        o0377(.A(ori_ori_n405_), .B(ori_ori_n401_), .Y(ori_ori_n406_));
  NOi31      o0378(.An(n), .B(m), .C(k), .Y(ori_ori_n407_));
  AOI220     o0379(.A0(ori_ori_n407_), .A1(ori_ori_n345_), .B0(ori_ori_n207_), .B1(ori_ori_n47_), .Y(ori_ori_n408_));
  NAi31      o0380(.An(g), .B(f), .C(c), .Y(ori_ori_n409_));
  NA2        o0381(.A(ori_ori_n406_), .B(ori_ori_n277_), .Y(ori_ori_n410_));
  NOi31      o0382(.An(ori_ori_n391_), .B(ori_ori_n410_), .C(ori_ori_n404_), .Y(ori_ori_n411_));
  NOi32      o0383(.An(c), .Bn(a), .C(b), .Y(ori_ori_n412_));
  NA2        o0384(.A(ori_ori_n412_), .B(ori_ori_n108_), .Y(ori_ori_n413_));
  AN2        o0385(.A(e), .B(d), .Y(ori_ori_n414_));
  INV        o0386(.A(ori_ori_n139_), .Y(ori_ori_n415_));
  NO2        o0387(.A(ori_ori_n123_), .B(ori_ori_n40_), .Y(ori_ori_n416_));
  NO2        o0388(.A(ori_ori_n61_), .B(e), .Y(ori_ori_n417_));
  AOI210     o0389(.A0(ori_ori_n416_), .A1(ori_ori_n415_), .B0(ori_ori_n417_), .Y(ori_ori_n418_));
  NO2        o0390(.A(ori_ori_n418_), .B(ori_ori_n413_), .Y(ori_ori_n419_));
  INV        o0391(.A(ori_ori_n195_), .Y(ori_ori_n420_));
  NOi21      o0392(.An(a), .B(b), .Y(ori_ori_n421_));
  NA3        o0393(.A(e), .B(d), .C(c), .Y(ori_ori_n422_));
  NAi21      o0394(.An(ori_ori_n422_), .B(ori_ori_n421_), .Y(ori_ori_n423_));
  NO2        o0395(.A(ori_ori_n420_), .B(ori_ori_n423_), .Y(ori_ori_n424_));
  NA2        o0396(.A(ori_ori_n340_), .B(ori_ori_n145_), .Y(ori_ori_n425_));
  OR2        o0397(.A(k), .B(j), .Y(ori_ori_n426_));
  NA2        o0398(.A(l), .B(k), .Y(ori_ori_n427_));
  NA3        o0399(.A(ori_ori_n427_), .B(ori_ori_n426_), .C(ori_ori_n207_), .Y(ori_ori_n428_));
  AOI210     o0400(.A0(ori_ori_n220_), .A1(ori_ori_n300_), .B0(ori_ori_n78_), .Y(ori_ori_n429_));
  NOi21      o0401(.An(ori_ori_n428_), .B(ori_ori_n429_), .Y(ori_ori_n430_));
  OR3        o0402(.A(ori_ori_n430_), .B(ori_ori_n135_), .C(ori_ori_n125_), .Y(ori_ori_n431_));
  NA3        o0403(.A(ori_ori_n254_), .B(ori_ori_n121_), .C(ori_ori_n119_), .Y(ori_ori_n432_));
  NO2        o0404(.A(ori_ori_n432_), .B(ori_ori_n288_), .Y(ori_ori_n433_));
  NA3        o0405(.A(ori_ori_n433_), .B(ori_ori_n431_), .C(ori_ori_n425_), .Y(ori_ori_n434_));
  NO3        o0406(.A(ori_ori_n434_), .B(ori_ori_n424_), .C(ori_ori_n419_), .Y(ori_ori_n435_));
  INV        o0407(.A(e), .Y(ori_ori_n436_));
  NO2        o0408(.A(ori_ori_n177_), .B(ori_ori_n53_), .Y(ori_ori_n437_));
  NAi31      o0409(.An(j), .B(l), .C(i), .Y(ori_ori_n438_));
  OAI210     o0410(.A0(ori_ori_n438_), .A1(ori_ori_n124_), .B0(ori_ori_n97_), .Y(ori_ori_n439_));
  NA3        o0411(.A(ori_ori_n439_), .B(ori_ori_n437_), .C(ori_ori_n436_), .Y(ori_ori_n440_));
  NO2        o0412(.A(ori_ori_n354_), .B(ori_ori_n330_), .Y(ori_ori_n441_));
  NO3        o0413(.A(ori_ori_n441_), .B(ori_ori_n176_), .C(ori_ori_n274_), .Y(ori_ori_n442_));
  NA3        o0414(.A(ori_ori_n442_), .B(ori_ori_n440_), .C(ori_ori_n228_), .Y(ori_ori_n443_));
  OAI210     o0415(.A0(ori_ori_n120_), .A1(ori_ori_n118_), .B0(n), .Y(ori_ori_n444_));
  NO2        o0416(.A(ori_ori_n444_), .B(ori_ori_n123_), .Y(ori_ori_n445_));
  XO2        o0417(.A(i), .B(h), .Y(ori_ori_n446_));
  NA3        o0418(.A(ori_ori_n446_), .B(ori_ori_n152_), .C(n), .Y(ori_ori_n447_));
  NA3        o0419(.A(ori_ori_n447_), .B(ori_ori_n408_), .C(ori_ori_n342_), .Y(ori_ori_n448_));
  NOi32      o0420(.An(ori_ori_n448_), .Bn(ori_ori_n417_), .C(ori_ori_n248_), .Y(ori_ori_n449_));
  NAi31      o0421(.An(c), .B(f), .C(d), .Y(ori_ori_n450_));
  AOI210     o0422(.A0(ori_ori_n255_), .A1(ori_ori_n182_), .B0(ori_ori_n450_), .Y(ori_ori_n451_));
  NOi21      o0423(.An(ori_ori_n76_), .B(ori_ori_n451_), .Y(ori_ori_n452_));
  NA3        o0424(.A(ori_ori_n338_), .B(ori_ori_n92_), .C(ori_ori_n91_), .Y(ori_ori_n453_));
  NA2        o0425(.A(ori_ori_n214_), .B(ori_ori_n103_), .Y(ori_ori_n454_));
  AOI210     o0426(.A0(ori_ori_n454_), .A1(ori_ori_n172_), .B0(ori_ori_n450_), .Y(ori_ori_n455_));
  AOI210     o0427(.A0(ori_ori_n318_), .A1(ori_ori_n34_), .B0(ori_ori_n423_), .Y(ori_ori_n456_));
  NOi31      o0428(.An(ori_ori_n453_), .B(ori_ori_n456_), .C(ori_ori_n455_), .Y(ori_ori_n457_));
  AO220      o0429(.A0(ori_ori_n263_), .A1(ori_ori_n246_), .B0(ori_ori_n158_), .B1(ori_ori_n62_), .Y(ori_ori_n458_));
  NA3        o0430(.A(ori_ori_n36_), .B(ori_ori_n35_), .C(f), .Y(ori_ori_n459_));
  NAi31      o0431(.An(ori_ori_n458_), .B(ori_ori_n457_), .C(ori_ori_n452_), .Y(ori_ori_n460_));
  NO3        o0432(.A(ori_ori_n460_), .B(ori_ori_n449_), .C(ori_ori_n443_), .Y(ori_ori_n461_));
  NA4        o0433(.A(ori_ori_n461_), .B(ori_ori_n435_), .C(ori_ori_n411_), .D(ori_ori_n382_), .Y(ori11));
  NO2        o0434(.A(ori_ori_n66_), .B(f), .Y(ori_ori_n463_));
  NA2        o0435(.A(j), .B(g), .Y(ori_ori_n464_));
  NAi31      o0436(.An(i), .B(m), .C(l), .Y(ori_ori_n465_));
  NA3        o0437(.A(m), .B(k), .C(j), .Y(ori_ori_n466_));
  OAI220     o0438(.A0(ori_ori_n466_), .A1(ori_ori_n123_), .B0(ori_ori_n465_), .B1(ori_ori_n464_), .Y(ori_ori_n467_));
  NA2        o0439(.A(ori_ori_n467_), .B(ori_ori_n463_), .Y(ori_ori_n468_));
  NOi32      o0440(.An(e), .Bn(b), .C(f), .Y(ori_ori_n469_));
  NA2        o0441(.A(ori_ori_n43_), .B(j), .Y(ori_ori_n470_));
  NO2        o0442(.A(ori_ori_n470_), .B(ori_ori_n270_), .Y(ori_ori_n471_));
  NAi31      o0443(.An(d), .B(e), .C(a), .Y(ori_ori_n472_));
  NO2        o0444(.A(ori_ori_n472_), .B(n), .Y(ori_ori_n473_));
  AOI220     o0445(.A0(ori_ori_n473_), .A1(ori_ori_n96_), .B0(ori_ori_n471_), .B1(ori_ori_n469_), .Y(ori_ori_n474_));
  NAi41      o0446(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n475_));
  AN2        o0447(.A(ori_ori_n475_), .B(ori_ori_n329_), .Y(ori_ori_n476_));
  AOI210     o0448(.A0(ori_ori_n476_), .A1(ori_ori_n354_), .B0(ori_ori_n249_), .Y(ori_ori_n477_));
  NA2        o0449(.A(j), .B(i), .Y(ori_ori_n478_));
  NAi31      o0450(.An(n), .B(m), .C(k), .Y(ori_ori_n479_));
  NO3        o0451(.A(ori_ori_n479_), .B(ori_ori_n478_), .C(ori_ori_n107_), .Y(ori_ori_n480_));
  NO4        o0452(.A(n), .B(d), .C(ori_ori_n110_), .D(a), .Y(ori_ori_n481_));
  OR2        o0453(.A(n), .B(c), .Y(ori_ori_n482_));
  NO2        o0454(.A(ori_ori_n482_), .B(ori_ori_n141_), .Y(ori_ori_n483_));
  NO2        o0455(.A(ori_ori_n483_), .B(ori_ori_n481_), .Y(ori_ori_n484_));
  NOi32      o0456(.An(g), .Bn(f), .C(i), .Y(ori_ori_n485_));
  AOI220     o0457(.A0(ori_ori_n485_), .A1(ori_ori_n94_), .B0(ori_ori_n467_), .B1(f), .Y(ori_ori_n486_));
  NO2        o0458(.A(ori_ori_n486_), .B(ori_ori_n484_), .Y(ori_ori_n487_));
  AOI210     o0459(.A0(ori_ori_n480_), .A1(ori_ori_n477_), .B0(ori_ori_n487_), .Y(ori_ori_n488_));
  NA2        o0460(.A(ori_ori_n131_), .B(ori_ori_n33_), .Y(ori_ori_n489_));
  OAI220     o0461(.A0(ori_ori_n489_), .A1(m), .B0(ori_ori_n470_), .B1(ori_ori_n220_), .Y(ori_ori_n490_));
  NOi41      o0462(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n491_));
  NAi32      o0463(.An(e), .Bn(b), .C(c), .Y(ori_ori_n492_));
  OR2        o0464(.A(ori_ori_n492_), .B(ori_ori_n78_), .Y(ori_ori_n493_));
  AN2        o0465(.A(ori_ori_n301_), .B(ori_ori_n285_), .Y(ori_ori_n494_));
  NA2        o0466(.A(ori_ori_n494_), .B(ori_ori_n493_), .Y(ori_ori_n495_));
  OA210      o0467(.A0(ori_ori_n495_), .A1(ori_ori_n491_), .B0(ori_ori_n490_), .Y(ori_ori_n496_));
  OAI220     o0468(.A0(ori_ori_n356_), .A1(ori_ori_n355_), .B0(ori_ori_n465_), .B1(ori_ori_n464_), .Y(ori_ori_n497_));
  NO3        o0469(.A(ori_ori_n59_), .B(ori_ori_n46_), .C(ori_ori_n200_), .Y(ori_ori_n498_));
  NO2        o0470(.A(ori_ori_n217_), .B(ori_ori_n105_), .Y(ori_ori_n499_));
  OAI210     o0471(.A0(ori_ori_n498_), .A1(ori_ori_n357_), .B0(ori_ori_n499_), .Y(ori_ori_n500_));
  INV        o0472(.A(ori_ori_n500_), .Y(ori_ori_n501_));
  NO2        o0473(.A(ori_ori_n252_), .B(n), .Y(ori_ori_n502_));
  NO2        o0474(.A(ori_ori_n379_), .B(ori_ori_n502_), .Y(ori_ori_n503_));
  NA2        o0475(.A(ori_ori_n497_), .B(f), .Y(ori_ori_n504_));
  NAi32      o0476(.An(d), .Bn(a), .C(b), .Y(ori_ori_n505_));
  NO2        o0477(.A(ori_ori_n505_), .B(ori_ori_n46_), .Y(ori_ori_n506_));
  NA2        o0478(.A(h), .B(f), .Y(ori_ori_n507_));
  NO2        o0479(.A(ori_ori_n507_), .B(ori_ori_n89_), .Y(ori_ori_n508_));
  NO3        o0480(.A(ori_ori_n168_), .B(ori_ori_n165_), .C(g), .Y(ori_ori_n509_));
  AOI220     o0481(.A0(ori_ori_n509_), .A1(ori_ori_n55_), .B0(ori_ori_n508_), .B1(ori_ori_n506_), .Y(ori_ori_n510_));
  OAI210     o0482(.A0(ori_ori_n504_), .A1(ori_ori_n503_), .B0(ori_ori_n510_), .Y(ori_ori_n511_));
  AN3        o0483(.A(j), .B(h), .C(g), .Y(ori_ori_n512_));
  NO2        o0484(.A(ori_ori_n138_), .B(c), .Y(ori_ori_n513_));
  NA3        o0485(.A(ori_ori_n513_), .B(ori_ori_n512_), .C(ori_ori_n407_), .Y(ori_ori_n514_));
  NA3        o0486(.A(f), .B(d), .C(b), .Y(ori_ori_n515_));
  NO4        o0487(.A(ori_ori_n515_), .B(ori_ori_n168_), .C(ori_ori_n165_), .D(g), .Y(ori_ori_n516_));
  NAi21      o0488(.An(ori_ori_n516_), .B(ori_ori_n514_), .Y(ori_ori_n517_));
  NO4        o0489(.A(ori_ori_n517_), .B(ori_ori_n511_), .C(ori_ori_n501_), .D(ori_ori_n496_), .Y(ori_ori_n518_));
  AN4        o0490(.A(ori_ori_n518_), .B(ori_ori_n488_), .C(ori_ori_n474_), .D(ori_ori_n468_), .Y(ori_ori_n519_));
  INV        o0491(.A(k), .Y(ori_ori_n520_));
  NA3        o0492(.A(l), .B(ori_ori_n520_), .C(i), .Y(ori_ori_n521_));
  INV        o0493(.A(ori_ori_n521_), .Y(ori_ori_n522_));
  NA4        o0494(.A(ori_ori_n353_), .B(ori_ori_n373_), .C(ori_ori_n173_), .D(ori_ori_n108_), .Y(ori_ori_n523_));
  NAi32      o0495(.An(h), .Bn(f), .C(g), .Y(ori_ori_n524_));
  NAi41      o0496(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n525_));
  OAI210     o0497(.A0(ori_ori_n472_), .A1(n), .B0(ori_ori_n525_), .Y(ori_ori_n526_));
  NA2        o0498(.A(ori_ori_n526_), .B(m), .Y(ori_ori_n527_));
  NAi31      o0499(.An(h), .B(g), .C(f), .Y(ori_ori_n528_));
  OR3        o0500(.A(ori_ori_n528_), .B(ori_ori_n252_), .C(ori_ori_n46_), .Y(ori_ori_n529_));
  NA4        o0501(.A(ori_ori_n373_), .B(ori_ori_n114_), .C(ori_ori_n108_), .D(e), .Y(ori_ori_n530_));
  AN2        o0502(.A(ori_ori_n530_), .B(ori_ori_n529_), .Y(ori_ori_n531_));
  OA210      o0503(.A0(ori_ori_n527_), .A1(ori_ori_n524_), .B0(ori_ori_n531_), .Y(ori_ori_n532_));
  NO3        o0504(.A(ori_ori_n524_), .B(ori_ori_n66_), .C(ori_ori_n67_), .Y(ori_ori_n533_));
  NO4        o0505(.A(ori_ori_n528_), .B(ori_ori_n482_), .C(ori_ori_n141_), .D(ori_ori_n67_), .Y(ori_ori_n534_));
  OR2        o0506(.A(ori_ori_n534_), .B(ori_ori_n533_), .Y(ori_ori_n535_));
  NAi31      o0507(.An(ori_ori_n535_), .B(ori_ori_n532_), .C(ori_ori_n523_), .Y(ori_ori_n536_));
  NAi31      o0508(.An(f), .B(h), .C(g), .Y(ori_ori_n537_));
  NOi32      o0509(.An(b), .Bn(a), .C(c), .Y(ori_ori_n538_));
  NOi41      o0510(.An(ori_ori_n538_), .B(ori_ori_n311_), .C(ori_ori_n63_), .D(ori_ori_n111_), .Y(ori_ori_n539_));
  NOi32      o0511(.An(d), .Bn(a), .C(e), .Y(ori_ori_n540_));
  NA2        o0512(.A(ori_ori_n540_), .B(ori_ori_n108_), .Y(ori_ori_n541_));
  NO2        o0513(.A(n), .B(c), .Y(ori_ori_n542_));
  NA3        o0514(.A(ori_ori_n542_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n543_));
  NAi32      o0515(.An(n), .Bn(f), .C(m), .Y(ori_ori_n544_));
  NA3        o0516(.A(ori_ori_n544_), .B(ori_ori_n543_), .C(ori_ori_n541_), .Y(ori_ori_n545_));
  NOi32      o0517(.An(e), .Bn(a), .C(d), .Y(ori_ori_n546_));
  AOI210     o0518(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n546_), .Y(ori_ori_n547_));
  AOI210     o0519(.A0(ori_ori_n547_), .A1(ori_ori_n199_), .B0(ori_ori_n489_), .Y(ori_ori_n548_));
  AOI210     o0520(.A0(ori_ori_n548_), .A1(ori_ori_n545_), .B0(ori_ori_n539_), .Y(ori_ori_n549_));
  OAI210     o0521(.A0(ori_ori_n232_), .A1(ori_ori_n81_), .B0(ori_ori_n549_), .Y(ori_ori_n550_));
  AOI210     o0522(.A0(ori_ori_n536_), .A1(ori_ori_n522_), .B0(ori_ori_n550_), .Y(ori_ori_n551_));
  NO3        o0523(.A(ori_ori_n283_), .B(ori_ori_n58_), .C(n), .Y(ori_ori_n552_));
  NA3        o0524(.A(ori_ori_n450_), .B(ori_ori_n163_), .C(ori_ori_n162_), .Y(ori_ori_n553_));
  NA2        o0525(.A(ori_ori_n409_), .B(ori_ori_n217_), .Y(ori_ori_n554_));
  OR2        o0526(.A(ori_ori_n554_), .B(ori_ori_n553_), .Y(ori_ori_n555_));
  NA2        o0527(.A(ori_ori_n555_), .B(ori_ori_n552_), .Y(ori_ori_n556_));
  NO2        o0528(.A(ori_ori_n556_), .B(ori_ori_n81_), .Y(ori_ori_n557_));
  NA3        o0529(.A(ori_ori_n491_), .B(ori_ori_n302_), .C(ori_ori_n43_), .Y(ori_ori_n558_));
  NOi32      o0530(.An(e), .Bn(c), .C(f), .Y(ori_ori_n559_));
  NOi21      o0531(.An(f), .B(g), .Y(ori_ori_n560_));
  NO2        o0532(.A(ori_ori_n560_), .B(ori_ori_n197_), .Y(ori_ori_n561_));
  AOI220     o0533(.A0(ori_ori_n561_), .A1(ori_ori_n350_), .B0(ori_ori_n559_), .B1(ori_ori_n167_), .Y(ori_ori_n562_));
  NA3        o0534(.A(ori_ori_n562_), .B(ori_ori_n558_), .C(ori_ori_n170_), .Y(ori_ori_n563_));
  AOI210     o0535(.A0(ori_ori_n476_), .A1(ori_ori_n354_), .B0(ori_ori_n269_), .Y(ori_ori_n564_));
  NOi21      o0536(.An(j), .B(l), .Y(ori_ori_n565_));
  NAi21      o0537(.An(k), .B(h), .Y(ori_ori_n566_));
  NO2        o0538(.A(ori_ori_n566_), .B(ori_ori_n245_), .Y(ori_ori_n567_));
  NA2        o0539(.A(ori_ori_n567_), .B(ori_ori_n565_), .Y(ori_ori_n568_));
  OR2        o0540(.A(ori_ori_n568_), .B(ori_ori_n527_), .Y(ori_ori_n569_));
  NOi31      o0541(.An(m), .B(n), .C(k), .Y(ori_ori_n570_));
  NA2        o0542(.A(ori_ori_n565_), .B(ori_ori_n570_), .Y(ori_ori_n571_));
  AOI210     o0543(.A0(ori_ori_n354_), .A1(ori_ori_n329_), .B0(ori_ori_n269_), .Y(ori_ori_n572_));
  NAi21      o0544(.An(ori_ori_n571_), .B(ori_ori_n572_), .Y(ori_ori_n573_));
  NO2        o0545(.A(ori_ori_n472_), .B(ori_ori_n46_), .Y(ori_ori_n574_));
  NA2        o0546(.A(ori_ori_n573_), .B(ori_ori_n569_), .Y(ori_ori_n575_));
  NA2        o0547(.A(ori_ori_n103_), .B(ori_ori_n35_), .Y(ori_ori_n576_));
  NO2        o0548(.A(k), .B(ori_ori_n200_), .Y(ori_ori_n577_));
  INV        o0549(.A(ori_ori_n320_), .Y(ori_ori_n578_));
  NO2        o0550(.A(ori_ori_n578_), .B(n), .Y(ori_ori_n579_));
  NAi31      o0551(.An(ori_ori_n576_), .B(ori_ori_n579_), .C(ori_ori_n577_), .Y(ori_ori_n580_));
  NO2        o0552(.A(ori_ori_n470_), .B(ori_ori_n168_), .Y(ori_ori_n581_));
  NA3        o0553(.A(ori_ori_n492_), .B(ori_ori_n248_), .C(ori_ori_n136_), .Y(ori_ori_n582_));
  NA2        o0554(.A(ori_ori_n446_), .B(ori_ori_n152_), .Y(ori_ori_n583_));
  NO3        o0555(.A(ori_ori_n351_), .B(ori_ori_n583_), .C(ori_ori_n81_), .Y(ori_ori_n584_));
  AOI210     o0556(.A0(ori_ori_n582_), .A1(ori_ori_n581_), .B0(ori_ori_n584_), .Y(ori_ori_n585_));
  AN3        o0557(.A(f), .B(d), .C(b), .Y(ori_ori_n586_));
  NA3        o0558(.A(ori_ori_n446_), .B(ori_ori_n152_), .C(ori_ori_n200_), .Y(ori_ori_n587_));
  NO2        o0559(.A(ori_ori_n219_), .B(ori_ori_n587_), .Y(ori_ori_n588_));
  NAi31      o0560(.An(m), .B(n), .C(k), .Y(ori_ori_n589_));
  OR2        o0561(.A(ori_ori_n125_), .B(ori_ori_n58_), .Y(ori_ori_n590_));
  OAI210     o0562(.A0(ori_ori_n590_), .A1(ori_ori_n589_), .B0(ori_ori_n234_), .Y(ori_ori_n591_));
  OAI210     o0563(.A0(ori_ori_n591_), .A1(ori_ori_n588_), .B0(j), .Y(ori_ori_n592_));
  NA3        o0564(.A(ori_ori_n592_), .B(ori_ori_n585_), .C(ori_ori_n580_), .Y(ori_ori_n593_));
  NO4        o0565(.A(ori_ori_n593_), .B(ori_ori_n575_), .C(ori_ori_n563_), .D(ori_ori_n557_), .Y(ori_ori_n594_));
  NA2        o0566(.A(ori_ori_n338_), .B(ori_ori_n155_), .Y(ori_ori_n595_));
  NAi31      o0567(.An(g), .B(h), .C(f), .Y(ori_ori_n596_));
  OR3        o0568(.A(ori_ori_n596_), .B(ori_ori_n252_), .C(n), .Y(ori_ori_n597_));
  OA210      o0569(.A0(ori_ori_n472_), .A1(n), .B0(ori_ori_n525_), .Y(ori_ori_n598_));
  NA3        o0570(.A(ori_ori_n372_), .B(ori_ori_n114_), .C(ori_ori_n78_), .Y(ori_ori_n599_));
  OAI210     o0571(.A0(ori_ori_n598_), .A1(ori_ori_n85_), .B0(ori_ori_n599_), .Y(ori_ori_n600_));
  NOi21      o0572(.An(ori_ori_n597_), .B(ori_ori_n600_), .Y(ori_ori_n601_));
  AOI210     o0573(.A0(ori_ori_n601_), .A1(ori_ori_n595_), .B0(ori_ori_n466_), .Y(ori_ori_n602_));
  NO3        o0574(.A(g), .B(ori_ori_n199_), .C(ori_ori_n53_), .Y(ori_ori_n603_));
  NO2        o0575(.A(ori_ori_n454_), .B(ori_ori_n81_), .Y(ori_ori_n604_));
  OAI210     o0576(.A0(ori_ori_n604_), .A1(ori_ori_n350_), .B0(ori_ori_n603_), .Y(ori_ori_n605_));
  OR2        o0577(.A(ori_ori_n66_), .B(ori_ori_n67_), .Y(ori_ori_n606_));
  NA2        o0578(.A(ori_ori_n538_), .B(ori_ori_n304_), .Y(ori_ori_n607_));
  OA220      o0579(.A0(ori_ori_n571_), .A1(ori_ori_n607_), .B0(ori_ori_n568_), .B1(ori_ori_n606_), .Y(ori_ori_n608_));
  NA3        o0580(.A(ori_ori_n463_), .B(ori_ori_n94_), .C(ori_ori_n93_), .Y(ori_ori_n609_));
  AN2        o0581(.A(h), .B(f), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n610_), .B(ori_ori_n36_), .Y(ori_ori_n611_));
  NO2        o0583(.A(ori_ori_n611_), .B(ori_ori_n413_), .Y(ori_ori_n612_));
  AOI210     o0584(.A0(ori_ori_n505_), .A1(ori_ori_n378_), .B0(ori_ori_n46_), .Y(ori_ori_n613_));
  INV        o0585(.A(ori_ori_n612_), .Y(ori_ori_n614_));
  NA4        o0586(.A(ori_ori_n614_), .B(ori_ori_n609_), .C(ori_ori_n608_), .D(ori_ori_n605_), .Y(ori_ori_n615_));
  NA2        o0587(.A(ori_ori_n124_), .B(ori_ori_n46_), .Y(ori_ori_n616_));
  AOI220     o0588(.A0(ori_ori_n616_), .A1(ori_ori_n469_), .B0(ori_ori_n320_), .B1(ori_ori_n108_), .Y(ori_ori_n617_));
  OA220      o0589(.A0(ori_ori_n617_), .A1(ori_ori_n489_), .B0(ori_ori_n318_), .B1(ori_ori_n106_), .Y(ori_ori_n618_));
  INV        o0590(.A(ori_ori_n618_), .Y(ori_ori_n619_));
  NO3        o0591(.A(ori_ori_n361_), .B(ori_ori_n179_), .C(ori_ori_n178_), .Y(ori_ori_n620_));
  NA2        o0592(.A(ori_ori_n620_), .B(ori_ori_n217_), .Y(ori_ori_n621_));
  NA3        o0593(.A(ori_ori_n621_), .B(ori_ori_n238_), .C(j), .Y(ori_ori_n622_));
  NO3        o0594(.A(ori_ori_n409_), .B(ori_ori_n165_), .C(i), .Y(ori_ori_n623_));
  NA2        o0595(.A(ori_ori_n412_), .B(ori_ori_n78_), .Y(ori_ori_n624_));
  NA3        o0596(.A(ori_ori_n622_), .B(ori_ori_n453_), .C(ori_ori_n359_), .Y(ori_ori_n625_));
  NO4        o0597(.A(ori_ori_n625_), .B(ori_ori_n619_), .C(ori_ori_n615_), .D(ori_ori_n602_), .Y(ori_ori_n626_));
  NA4        o0598(.A(ori_ori_n626_), .B(ori_ori_n594_), .C(ori_ori_n551_), .D(ori_ori_n519_), .Y(ori08));
  NO2        o0599(.A(k), .B(h), .Y(ori_ori_n628_));
  AO210      o0600(.A0(ori_ori_n236_), .A1(ori_ori_n399_), .B0(ori_ori_n628_), .Y(ori_ori_n629_));
  NO2        o0601(.A(ori_ori_n629_), .B(ori_ori_n268_), .Y(ori_ori_n630_));
  NA2        o0602(.A(ori_ori_n559_), .B(ori_ori_n78_), .Y(ori_ori_n631_));
  NA2        o0603(.A(ori_ori_n631_), .B(ori_ori_n409_), .Y(ori_ori_n632_));
  NA2        o0604(.A(ori_ori_n632_), .B(ori_ori_n630_), .Y(ori_ori_n633_));
  NA2        o0605(.A(ori_ori_n78_), .B(ori_ori_n105_), .Y(ori_ori_n634_));
  NO2        o0606(.A(ori_ori_n634_), .B(ori_ori_n54_), .Y(ori_ori_n635_));
  NO4        o0607(.A(ori_ori_n336_), .B(ori_ori_n107_), .C(j), .D(ori_ori_n200_), .Y(ori_ori_n636_));
  NA2        o0608(.A(ori_ori_n636_), .B(ori_ori_n635_), .Y(ori_ori_n637_));
  AOI210     o0609(.A0(ori_ori_n515_), .A1(ori_ori_n148_), .B0(ori_ori_n78_), .Y(ori_ori_n638_));
  NA4        o0610(.A(ori_ori_n202_), .B(ori_ori_n131_), .C(ori_ori_n42_), .D(h), .Y(ori_ori_n639_));
  AN2        o0611(.A(l), .B(k), .Y(ori_ori_n640_));
  NA4        o0612(.A(ori_ori_n640_), .B(ori_ori_n103_), .C(ori_ori_n67_), .D(ori_ori_n200_), .Y(ori_ori_n641_));
  OAI210     o0613(.A0(ori_ori_n639_), .A1(g), .B0(ori_ori_n641_), .Y(ori_ori_n642_));
  NA2        o0614(.A(ori_ori_n642_), .B(ori_ori_n638_), .Y(ori_ori_n643_));
  NA4        o0615(.A(ori_ori_n643_), .B(ori_ori_n637_), .C(ori_ori_n633_), .D(ori_ori_n307_), .Y(ori_ori_n644_));
  NO2        o0616(.A(ori_ori_n37_), .B(ori_ori_n199_), .Y(ori_ori_n645_));
  AOI220     o0617(.A0(ori_ori_n561_), .A1(ori_ori_n306_), .B0(ori_ori_n645_), .B1(ori_ori_n502_), .Y(ori_ori_n646_));
  INV        o0618(.A(ori_ori_n646_), .Y(ori_ori_n647_));
  NO2        o0619(.A(ori_ori_n476_), .B(ori_ori_n34_), .Y(ori_ori_n648_));
  OAI210     o0620(.A0(ori_ori_n492_), .A1(ori_ori_n44_), .B0(ori_ori_n590_), .Y(ori_ori_n649_));
  NO2        o0621(.A(ori_ori_n427_), .B(ori_ori_n124_), .Y(ori_ori_n650_));
  AOI210     o0622(.A0(ori_ori_n650_), .A1(ori_ori_n649_), .B0(ori_ori_n648_), .Y(ori_ori_n651_));
  NO3        o0623(.A(ori_ori_n283_), .B(ori_ori_n123_), .C(ori_ori_n40_), .Y(ori_ori_n652_));
  NAi21      o0624(.An(ori_ori_n652_), .B(ori_ori_n641_), .Y(ori_ori_n653_));
  NA2        o0625(.A(ori_ori_n629_), .B(ori_ori_n126_), .Y(ori_ori_n654_));
  AOI220     o0626(.A0(ori_ori_n654_), .A1(ori_ori_n360_), .B0(ori_ori_n653_), .B1(ori_ori_n70_), .Y(ori_ori_n655_));
  OAI210     o0627(.A0(ori_ori_n651_), .A1(ori_ori_n81_), .B0(ori_ori_n655_), .Y(ori_ori_n656_));
  NA3        o0628(.A(ori_ori_n621_), .B(ori_ori_n296_), .C(ori_ori_n341_), .Y(ori_ori_n657_));
  NA3        o0629(.A(m), .B(l), .C(k), .Y(ori_ori_n658_));
  AOI210     o0630(.A0(ori_ori_n599_), .A1(ori_ori_n597_), .B0(ori_ori_n658_), .Y(ori_ori_n659_));
  INV        o0631(.A(ori_ori_n659_), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n660_), .B(ori_ori_n657_), .Y(ori_ori_n661_));
  NO4        o0633(.A(ori_ori_n661_), .B(ori_ori_n656_), .C(ori_ori_n647_), .D(ori_ori_n644_), .Y(ori_ori_n662_));
  NOi31      o0634(.An(g), .B(h), .C(f), .Y(ori_ori_n663_));
  NA2        o0635(.A(ori_ori_n574_), .B(ori_ori_n663_), .Y(ori_ori_n664_));
  AO210      o0636(.A0(ori_ori_n664_), .A1(ori_ori_n529_), .B0(ori_ori_n478_), .Y(ori_ori_n665_));
  NO3        o0637(.A(ori_ori_n354_), .B(ori_ori_n464_), .C(h), .Y(ori_ori_n666_));
  AOI210     o0638(.A0(ori_ori_n666_), .A1(ori_ori_n108_), .B0(ori_ori_n441_), .Y(ori_ori_n667_));
  NA3        o0639(.A(ori_ori_n667_), .B(ori_ori_n665_), .C(ori_ori_n235_), .Y(ori_ori_n668_));
  NA2        o0640(.A(ori_ori_n640_), .B(ori_ori_n67_), .Y(ori_ori_n669_));
  NO4        o0641(.A(ori_ori_n620_), .B(ori_ori_n165_), .C(n), .D(i), .Y(ori_ori_n670_));
  NOi21      o0642(.An(h), .B(j), .Y(ori_ori_n671_));
  NA2        o0643(.A(ori_ori_n671_), .B(f), .Y(ori_ori_n672_));
  NO2        o0644(.A(ori_ori_n672_), .B(ori_ori_n229_), .Y(ori_ori_n673_));
  NO3        o0645(.A(ori_ori_n673_), .B(ori_ori_n670_), .C(ori_ori_n623_), .Y(ori_ori_n674_));
  OAI220     o0646(.A0(ori_ori_n674_), .A1(ori_ori_n669_), .B0(ori_ori_n531_), .B1(ori_ori_n59_), .Y(ori_ori_n675_));
  AOI210     o0647(.A0(ori_ori_n668_), .A1(l), .B0(ori_ori_n675_), .Y(ori_ori_n676_));
  NO2        o0648(.A(j), .B(i), .Y(ori_ori_n677_));
  NA3        o0649(.A(ori_ori_n677_), .B(ori_ori_n74_), .C(l), .Y(ori_ori_n678_));
  NA2        o0650(.A(ori_ori_n677_), .B(ori_ori_n32_), .Y(ori_ori_n679_));
  OR2        o0651(.A(ori_ori_n678_), .B(ori_ori_n527_), .Y(ori_ori_n680_));
  NO3        o0652(.A(ori_ori_n143_), .B(ori_ori_n46_), .C(ori_ori_n105_), .Y(ori_ori_n681_));
  NO3        o0653(.A(ori_ori_n482_), .B(ori_ori_n141_), .C(ori_ori_n67_), .Y(ori_ori_n682_));
  NO2        o0654(.A(ori_ori_n664_), .B(ori_ori_n59_), .Y(ori_ori_n683_));
  INV        o0655(.A(j), .Y(ori_ori_n684_));
  NO3        o0656(.A(ori_ori_n268_), .B(ori_ori_n684_), .C(ori_ori_n39_), .Y(ori_ori_n685_));
  AOI210     o0657(.A0(ori_ori_n469_), .A1(n), .B0(ori_ori_n491_), .Y(ori_ori_n686_));
  NA2        o0658(.A(ori_ori_n686_), .B(ori_ori_n494_), .Y(ori_ori_n687_));
  AN3        o0659(.A(ori_ori_n687_), .B(ori_ori_n685_), .C(ori_ori_n93_), .Y(ori_ori_n688_));
  NO3        o0660(.A(ori_ori_n165_), .B(ori_ori_n349_), .C(ori_ori_n107_), .Y(ori_ori_n689_));
  AOI220     o0661(.A0(ori_ori_n689_), .A1(ori_ori_n230_), .B0(ori_ori_n554_), .B1(ori_ori_n276_), .Y(ori_ori_n690_));
  NAi31      o0662(.An(ori_ori_n547_), .B(ori_ori_n87_), .C(ori_ori_n78_), .Y(ori_ori_n691_));
  NA2        o0663(.A(ori_ori_n691_), .B(ori_ori_n690_), .Y(ori_ori_n692_));
  OR3        o0664(.A(ori_ori_n692_), .B(ori_ori_n688_), .C(ori_ori_n683_), .Y(ori_ori_n693_));
  NA3        o0665(.A(ori_ori_n686_), .B(ori_ori_n494_), .C(ori_ori_n493_), .Y(ori_ori_n694_));
  NA4        o0666(.A(ori_ori_n694_), .B(ori_ori_n202_), .C(ori_ori_n399_), .D(ori_ori_n33_), .Y(ori_ori_n695_));
  NO4        o0667(.A(ori_ori_n427_), .B(ori_ori_n383_), .C(j), .D(f), .Y(ori_ori_n696_));
  NO2        o0668(.A(ori_ori_n639_), .B(ori_ori_n631_), .Y(ori_ori_n697_));
  AOI210     o0669(.A0(ori_ori_n696_), .A1(ori_ori_n242_), .B0(ori_ori_n697_), .Y(ori_ori_n698_));
  NA3        o0670(.A(ori_ori_n485_), .B(ori_ori_n266_), .C(h), .Y(ori_ori_n699_));
  OAI220     o0671(.A0(ori_ori_n699_), .A1(ori_ori_n543_), .B0(ori_ori_n678_), .B1(ori_ori_n606_), .Y(ori_ori_n700_));
  INV        o0672(.A(ori_ori_n700_), .Y(ori_ori_n701_));
  NA3        o0673(.A(ori_ori_n701_), .B(ori_ori_n698_), .C(ori_ori_n695_), .Y(ori_ori_n702_));
  NO2        o0674(.A(ori_ori_n598_), .B(ori_ori_n67_), .Y(ori_ori_n703_));
  AOI210     o0675(.A0(ori_ori_n696_), .A1(ori_ori_n703_), .B0(ori_ori_n298_), .Y(ori_ori_n704_));
  OAI210     o0676(.A0(ori_ori_n658_), .A1(ori_ori_n596_), .B0(ori_ori_n459_), .Y(ori_ori_n705_));
  NA3        o0677(.A(ori_ori_n233_), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n706_));
  AOI220     o0678(.A0(ori_ori_n542_), .A1(ori_ori_n29_), .B0(ori_ori_n412_), .B1(ori_ori_n78_), .Y(ori_ori_n707_));
  NA2        o0679(.A(ori_ori_n707_), .B(ori_ori_n706_), .Y(ori_ori_n708_));
  NA2        o0680(.A(ori_ori_n708_), .B(ori_ori_n705_), .Y(ori_ori_n709_));
  NA2        o0681(.A(ori_ori_n709_), .B(ori_ori_n704_), .Y(ori_ori_n710_));
  NOi41      o0682(.An(ori_ori_n680_), .B(ori_ori_n710_), .C(ori_ori_n702_), .D(ori_ori_n693_), .Y(ori_ori_n711_));
  NO3        o0683(.A(ori_ori_n303_), .B(ori_ori_n269_), .C(ori_ori_n107_), .Y(ori_ori_n712_));
  NA2        o0684(.A(ori_ori_n712_), .B(ori_ori_n687_), .Y(ori_ori_n713_));
  NO3        o0685(.A(ori_ori_n464_), .B(ori_ori_n88_), .C(h), .Y(ori_ori_n714_));
  NA2        o0686(.A(ori_ori_n714_), .B(ori_ori_n635_), .Y(ori_ori_n715_));
  NA3        o0687(.A(ori_ori_n715_), .B(ori_ori_n713_), .C(ori_ori_n362_), .Y(ori_ori_n716_));
  OR2        o0688(.A(ori_ori_n596_), .B(ori_ori_n86_), .Y(ori_ori_n717_));
  NOi31      o0689(.An(b), .B(d), .C(a), .Y(ori_ori_n718_));
  NO2        o0690(.A(ori_ori_n718_), .B(ori_ori_n540_), .Y(ori_ori_n719_));
  NO2        o0691(.A(ori_ori_n719_), .B(n), .Y(ori_ori_n720_));
  BUFFER     o0692(.A(ori_ori_n707_), .Y(ori_ori_n721_));
  OAI220     o0693(.A0(ori_ori_n721_), .A1(ori_ori_n717_), .B0(ori_ori_n699_), .B1(ori_ori_n541_), .Y(ori_ori_n722_));
  NO2        o0694(.A(ori_ori_n492_), .B(ori_ori_n78_), .Y(ori_ori_n723_));
  NO3        o0695(.A(ori_ori_n560_), .B(ori_ori_n292_), .C(ori_ori_n111_), .Y(ori_ori_n724_));
  NOi21      o0696(.An(ori_ori_n724_), .B(ori_ori_n153_), .Y(ori_ori_n725_));
  AOI210     o0697(.A0(ori_ori_n712_), .A1(ori_ori_n723_), .B0(ori_ori_n725_), .Y(ori_ori_n726_));
  INV        o0698(.A(ori_ori_n726_), .Y(ori_ori_n727_));
  NO2        o0699(.A(ori_ori_n620_), .B(n), .Y(ori_ori_n728_));
  NA2        o0700(.A(ori_ori_n728_), .B(ori_ori_n630_), .Y(ori_ori_n729_));
  NO2        o0701(.A(ori_ori_n289_), .B(ori_ori_n223_), .Y(ori_ori_n730_));
  OAI210     o0702(.A0(ori_ori_n90_), .A1(ori_ori_n87_), .B0(ori_ori_n730_), .Y(ori_ori_n731_));
  NA2        o0703(.A(ori_ori_n114_), .B(ori_ori_n78_), .Y(ori_ori_n732_));
  INV        o0704(.A(ori_ori_n731_), .Y(ori_ori_n733_));
  OAI210     o0705(.A0(ori_ori_n534_), .A1(ori_ori_n533_), .B0(ori_ori_n321_), .Y(ori_ori_n734_));
  NAi31      o0706(.An(ori_ori_n733_), .B(ori_ori_n734_), .C(ori_ori_n729_), .Y(ori_ori_n735_));
  NO4        o0707(.A(ori_ori_n735_), .B(ori_ori_n727_), .C(ori_ori_n722_), .D(ori_ori_n716_), .Y(ori_ori_n736_));
  NA4        o0708(.A(ori_ori_n736_), .B(ori_ori_n711_), .C(ori_ori_n676_), .D(ori_ori_n662_), .Y(ori09));
  INV        o0709(.A(ori_ori_n115_), .Y(ori_ori_n738_));
  NA2        o0710(.A(f), .B(e), .Y(ori_ori_n739_));
  NO2        o0711(.A(ori_ori_n212_), .B(ori_ori_n107_), .Y(ori_ori_n740_));
  NA3        o0712(.A(ori_ori_n278_), .B(ori_ori_n1225_), .C(ori_ori_n244_), .Y(ori_ori_n741_));
  AOI210     o0713(.A0(ori_ori_n741_), .A1(g), .B0(ori_ori_n416_), .Y(ori_ori_n742_));
  NO2        o0714(.A(ori_ori_n742_), .B(ori_ori_n739_), .Y(ori_ori_n743_));
  NA2        o0715(.A(ori_ori_n393_), .B(e), .Y(ori_ori_n744_));
  NO2        o0716(.A(ori_ori_n744_), .B(ori_ori_n450_), .Y(ori_ori_n745_));
  AOI210     o0717(.A0(ori_ori_n743_), .A1(ori_ori_n738_), .B0(ori_ori_n745_), .Y(ori_ori_n746_));
  NO2        o0718(.A(ori_ori_n191_), .B(ori_ori_n199_), .Y(ori_ori_n747_));
  NA3        o0719(.A(m), .B(l), .C(i), .Y(ori_ori_n748_));
  OAI220     o0720(.A0(ori_ori_n528_), .A1(ori_ori_n748_), .B0(ori_ori_n311_), .B1(ori_ori_n465_), .Y(ori_ori_n749_));
  NAi21      o0721(.An(ori_ori_n749_), .B(ori_ori_n388_), .Y(ori_ori_n750_));
  OR2        o0722(.A(ori_ori_n750_), .B(ori_ori_n747_), .Y(ori_ori_n751_));
  NA2        o0723(.A(ori_ori_n717_), .B(ori_ori_n504_), .Y(ori_ori_n752_));
  OA210      o0724(.A0(ori_ori_n752_), .A1(ori_ori_n751_), .B0(ori_ori_n720_), .Y(ori_ori_n753_));
  INV        o0725(.A(ori_ori_n301_), .Y(ori_ori_n754_));
  NO2        o0726(.A(ori_ori_n120_), .B(ori_ori_n118_), .Y(ori_ori_n755_));
  NOi31      o0727(.An(k), .B(m), .C(l), .Y(ori_ori_n756_));
  NO2        o0728(.A(ori_ori_n302_), .B(ori_ori_n756_), .Y(ori_ori_n757_));
  AOI210     o0729(.A0(ori_ori_n757_), .A1(ori_ori_n755_), .B0(ori_ori_n537_), .Y(ori_ori_n758_));
  NA2        o0730(.A(ori_ori_n706_), .B(ori_ori_n295_), .Y(ori_ori_n759_));
  NA2        o0731(.A(ori_ori_n304_), .B(ori_ori_n305_), .Y(ori_ori_n760_));
  OAI210     o0732(.A0(ori_ori_n191_), .A1(ori_ori_n199_), .B0(ori_ori_n760_), .Y(ori_ori_n761_));
  AOI220     o0733(.A0(ori_ori_n761_), .A1(ori_ori_n759_), .B0(ori_ori_n758_), .B1(ori_ori_n754_), .Y(ori_ori_n762_));
  NA3        o0734(.A(ori_ori_n762_), .B(ori_ori_n562_), .C(ori_ori_n76_), .Y(ori_ori_n763_));
  NOi21      o0735(.An(f), .B(d), .Y(ori_ori_n764_));
  NA2        o0736(.A(ori_ori_n764_), .B(m), .Y(ori_ori_n765_));
  NO2        o0737(.A(ori_ori_n765_), .B(ori_ori_n49_), .Y(ori_ori_n766_));
  NOi32      o0738(.An(g), .Bn(f), .C(d), .Y(ori_ori_n767_));
  NA4        o0739(.A(ori_ori_n767_), .B(ori_ori_n542_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n768_));
  NOi21      o0740(.An(ori_ori_n279_), .B(ori_ori_n768_), .Y(ori_ori_n769_));
  AOI210     o0741(.A0(ori_ori_n766_), .A1(ori_ori_n483_), .B0(ori_ori_n769_), .Y(ori_ori_n770_));
  NA2        o0742(.A(ori_ori_n278_), .B(ori_ori_n244_), .Y(ori_ori_n771_));
  AN2        o0743(.A(f), .B(d), .Y(ori_ori_n772_));
  NA3        o0744(.A(ori_ori_n421_), .B(ori_ori_n772_), .C(ori_ori_n78_), .Y(ori_ori_n773_));
  NO3        o0745(.A(ori_ori_n773_), .B(ori_ori_n67_), .C(ori_ori_n200_), .Y(ori_ori_n774_));
  NA2        o0746(.A(ori_ori_n771_), .B(ori_ori_n774_), .Y(ori_ori_n775_));
  NAi31      o0747(.An(ori_ori_n432_), .B(ori_ori_n775_), .C(ori_ori_n770_), .Y(ori_ori_n776_));
  NO4        o0748(.A(ori_ori_n560_), .B(ori_ori_n124_), .C(ori_ori_n292_), .D(ori_ori_n144_), .Y(ori_ori_n777_));
  INV        o0749(.A(ori_ori_n777_), .Y(ori_ori_n778_));
  NA2        o0750(.A(ori_ori_n540_), .B(ori_ori_n78_), .Y(ori_ori_n779_));
  NO2        o0751(.A(ori_ori_n760_), .B(ori_ori_n779_), .Y(ori_ori_n780_));
  NA3        o0752(.A(ori_ori_n152_), .B(ori_ori_n103_), .C(ori_ori_n102_), .Y(ori_ori_n781_));
  OAI220     o0753(.A0(ori_ori_n773_), .A1(ori_ori_n380_), .B0(ori_ori_n301_), .B1(ori_ori_n781_), .Y(ori_ori_n782_));
  NOi41      o0754(.An(ori_ori_n210_), .B(ori_ori_n782_), .C(ori_ori_n780_), .D(ori_ori_n274_), .Y(ori_ori_n783_));
  NA2        o0755(.A(c), .B(ori_ori_n110_), .Y(ori_ori_n784_));
  NO2        o0756(.A(ori_ori_n784_), .B(ori_ori_n366_), .Y(ori_ori_n785_));
  NA3        o0757(.A(ori_ori_n785_), .B(ori_ori_n448_), .C(f), .Y(ori_ori_n786_));
  OR2        o0758(.A(ori_ori_n596_), .B(ori_ori_n479_), .Y(ori_ori_n787_));
  INV        o0759(.A(ori_ori_n787_), .Y(ori_ori_n788_));
  NA2        o0760(.A(ori_ori_n719_), .B(ori_ori_n106_), .Y(ori_ori_n789_));
  NA2        o0761(.A(ori_ori_n789_), .B(ori_ori_n788_), .Y(ori_ori_n790_));
  NA4        o0762(.A(ori_ori_n790_), .B(ori_ori_n786_), .C(ori_ori_n783_), .D(ori_ori_n778_), .Y(ori_ori_n791_));
  NO4        o0763(.A(ori_ori_n791_), .B(ori_ori_n776_), .C(ori_ori_n763_), .D(ori_ori_n753_), .Y(ori_ori_n792_));
  NA2        o0764(.A(ori_ori_n107_), .B(j), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n217_), .B(ori_ori_n211_), .Y(ori_ori_n794_));
  NA2        o0766(.A(ori_ori_n794_), .B(ori_ori_n214_), .Y(ori_ori_n795_));
  INV        o0767(.A(ori_ori_n795_), .Y(ori_ori_n796_));
  NA2        o0768(.A(e), .B(d), .Y(ori_ori_n797_));
  OAI220     o0769(.A0(ori_ori_n797_), .A1(c), .B0(ori_ori_n289_), .B1(d), .Y(ori_ori_n798_));
  NA3        o0770(.A(ori_ori_n798_), .B(ori_ori_n402_), .C(ori_ori_n446_), .Y(ori_ori_n799_));
  AOI210     o0771(.A0(ori_ori_n454_), .A1(ori_ori_n172_), .B0(ori_ori_n217_), .Y(ori_ori_n800_));
  AOI210     o0772(.A0(ori_ori_n561_), .A1(ori_ori_n306_), .B0(ori_ori_n800_), .Y(ori_ori_n801_));
  NA2        o0773(.A(ori_ori_n774_), .B(j), .Y(ori_ori_n802_));
  NA3        o0774(.A(ori_ori_n802_), .B(ori_ori_n801_), .C(ori_ori_n799_), .Y(ori_ori_n803_));
  NO2        o0775(.A(ori_ori_n803_), .B(ori_ori_n796_), .Y(ori_ori_n804_));
  OR2        o0776(.A(ori_ori_n631_), .B(ori_ori_n203_), .Y(ori_ori_n805_));
  NA2        o0777(.A(ori_ori_n552_), .B(ori_ori_n559_), .Y(ori_ori_n806_));
  OAI210     o0778(.A0(ori_ori_n744_), .A1(ori_ori_n162_), .B0(ori_ori_n806_), .Y(ori_ori_n807_));
  OAI210     o0779(.A0(ori_ori_n740_), .A1(j), .B0(ori_ori_n767_), .Y(ori_ori_n808_));
  NO2        o0780(.A(ori_ori_n808_), .B(ori_ori_n543_), .Y(ori_ori_n809_));
  NA2        o0781(.A(ori_ori_n112_), .B(ori_ori_n111_), .Y(ori_ori_n810_));
  NO2        o0782(.A(ori_ori_n810_), .B(ori_ori_n768_), .Y(ori_ori_n811_));
  AO210      o0783(.A0(ori_ori_n759_), .A1(ori_ori_n749_), .B0(ori_ori_n811_), .Y(ori_ori_n812_));
  NO3        o0784(.A(ori_ori_n812_), .B(ori_ori_n809_), .C(ori_ori_n807_), .Y(ori_ori_n813_));
  AO220      o0785(.A0(ori_ori_n402_), .A1(ori_ori_n671_), .B0(ori_ori_n167_), .B1(f), .Y(ori_ori_n814_));
  OAI210     o0786(.A0(ori_ori_n814_), .A1(ori_ori_n405_), .B0(ori_ori_n798_), .Y(ori_ori_n815_));
  NO2        o0787(.A(ori_ori_n387_), .B(ori_ori_n64_), .Y(ori_ori_n816_));
  OAI210     o0788(.A0(ori_ori_n752_), .A1(ori_ori_n816_), .B0(ori_ori_n635_), .Y(ori_ori_n817_));
  AN4        o0789(.A(ori_ori_n817_), .B(ori_ori_n815_), .C(ori_ori_n813_), .D(ori_ori_n805_), .Y(ori_ori_n818_));
  NA4        o0790(.A(ori_ori_n818_), .B(ori_ori_n804_), .C(ori_ori_n792_), .D(ori_ori_n746_), .Y(ori12));
  NO2        o0791(.A(ori_ori_n400_), .B(c), .Y(ori_ori_n820_));
  NO4        o0792(.A(ori_ori_n392_), .B(ori_ori_n236_), .C(ori_ori_n520_), .D(ori_ori_n200_), .Y(ori_ori_n821_));
  NA2        o0793(.A(ori_ori_n821_), .B(ori_ori_n820_), .Y(ori_ori_n822_));
  NA2        o0794(.A(ori_ori_n483_), .B(ori_ori_n816_), .Y(ori_ori_n823_));
  NO2        o0795(.A(ori_ori_n400_), .B(ori_ori_n110_), .Y(ori_ori_n824_));
  NO2        o0796(.A(ori_ori_n755_), .B(ori_ori_n311_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n596_), .B(ori_ori_n336_), .Y(ori_ori_n826_));
  AOI220     o0798(.A0(ori_ori_n826_), .A1(ori_ori_n481_), .B0(ori_ori_n825_), .B1(ori_ori_n824_), .Y(ori_ori_n827_));
  NA4        o0799(.A(ori_ori_n827_), .B(ori_ori_n823_), .C(ori_ori_n822_), .D(ori_ori_n391_), .Y(ori_ori_n828_));
  AOI210     o0800(.A0(ori_ori_n220_), .A1(ori_ori_n300_), .B0(ori_ori_n188_), .Y(ori_ori_n829_));
  OR2        o0801(.A(ori_ori_n829_), .B(ori_ori_n821_), .Y(ori_ori_n830_));
  AOI210     o0802(.A0(ori_ori_n297_), .A1(ori_ori_n347_), .B0(ori_ori_n200_), .Y(ori_ori_n831_));
  OAI210     o0803(.A0(ori_ori_n831_), .A1(ori_ori_n830_), .B0(ori_ori_n361_), .Y(ori_ori_n832_));
  NO2        o0804(.A(ori_ori_n576_), .B(ori_ori_n245_), .Y(ori_ori_n833_));
  NO2        o0805(.A(ori_ori_n528_), .B(ori_ori_n748_), .Y(ori_ori_n834_));
  AOI220     o0806(.A0(ori_ori_n834_), .A1(ori_ori_n502_), .B0(ori_ori_n730_), .B1(ori_ori_n833_), .Y(ori_ori_n835_));
  NO2        o0807(.A(ori_ori_n143_), .B(ori_ori_n223_), .Y(ori_ori_n836_));
  NA3        o0808(.A(ori_ori_n836_), .B(ori_ori_n226_), .C(i), .Y(ori_ori_n837_));
  NA3        o0809(.A(ori_ori_n837_), .B(ori_ori_n835_), .C(ori_ori_n832_), .Y(ori_ori_n838_));
  OR2        o0810(.A(ori_ori_n290_), .B(ori_ori_n824_), .Y(ori_ori_n839_));
  NA2        o0811(.A(ori_ori_n839_), .B(ori_ori_n312_), .Y(ori_ori_n840_));
  NO3        o0812(.A(ori_ori_n124_), .B(ori_ori_n144_), .C(ori_ori_n200_), .Y(ori_ori_n841_));
  NA2        o0813(.A(ori_ori_n841_), .B(ori_ori_n469_), .Y(ori_ori_n842_));
  NA4        o0814(.A(ori_ori_n393_), .B(ori_ori_n385_), .C(ori_ori_n173_), .D(g), .Y(ori_ori_n843_));
  NA3        o0815(.A(ori_ori_n843_), .B(ori_ori_n842_), .C(ori_ori_n840_), .Y(ori_ori_n844_));
  NO3        o0816(.A(ori_ori_n601_), .B(ori_ori_n86_), .C(ori_ori_n42_), .Y(ori_ori_n845_));
  NO4        o0817(.A(ori_ori_n845_), .B(ori_ori_n844_), .C(ori_ori_n838_), .D(ori_ori_n828_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n492_), .B(ori_ori_n136_), .Y(ori_ori_n847_));
  NOi21      o0819(.An(ori_ori_n33_), .B(ori_ori_n589_), .Y(ori_ori_n848_));
  NA2        o0820(.A(ori_ori_n848_), .B(ori_ori_n847_), .Y(ori_ori_n849_));
  OAI210     o0821(.A0(ori_ori_n234_), .A1(ori_ori_n42_), .B0(ori_ori_n849_), .Y(ori_ori_n850_));
  INV        o0822(.A(ori_ori_n287_), .Y(ori_ori_n851_));
  NO2        o0823(.A(ori_ori_n46_), .B(ori_ori_n42_), .Y(ori_ori_n852_));
  NO2        o0824(.A(ori_ori_n444_), .B(ori_ori_n269_), .Y(ori_ori_n853_));
  INV        o0825(.A(ori_ori_n853_), .Y(ori_ori_n854_));
  NO2        o0826(.A(ori_ori_n854_), .B(ori_ori_n136_), .Y(ori_ori_n855_));
  INV        o0827(.A(ori_ori_n325_), .Y(ori_ori_n856_));
  NO4        o0828(.A(ori_ori_n856_), .B(ori_ori_n855_), .C(ori_ori_n851_), .D(ori_ori_n850_), .Y(ori_ori_n857_));
  NA2        o0829(.A(ori_ori_n306_), .B(g), .Y(ori_ori_n858_));
  NA2        o0830(.A(ori_ori_n155_), .B(i), .Y(ori_ori_n859_));
  NA2        o0831(.A(ori_ori_n43_), .B(i), .Y(ori_ori_n860_));
  NO2        o0832(.A(ori_ori_n136_), .B(ori_ori_n78_), .Y(ori_ori_n861_));
  OR2        o0833(.A(ori_ori_n861_), .B(ori_ori_n491_), .Y(ori_ori_n862_));
  NA2        o0834(.A(ori_ori_n492_), .B(ori_ori_n339_), .Y(ori_ori_n863_));
  AOI210     o0835(.A0(ori_ori_n863_), .A1(n), .B0(ori_ori_n862_), .Y(ori_ori_n864_));
  NO2        o0836(.A(ori_ori_n864_), .B(ori_ori_n858_), .Y(ori_ori_n865_));
  NA3        o0837(.A(ori_ori_n304_), .B(ori_ori_n565_), .C(i), .Y(ori_ori_n866_));
  OAI210     o0838(.A0(ori_ori_n387_), .A1(ori_ori_n278_), .B0(ori_ori_n866_), .Y(ori_ori_n867_));
  OAI210     o0839(.A0(ori_ori_n613_), .A1(ori_ori_n682_), .B0(ori_ori_n867_), .Y(ori_ori_n868_));
  NA2        o0840(.A(ori_ori_n546_), .B(ori_ori_n108_), .Y(ori_ori_n869_));
  NA3        o0841(.A(ori_ori_n565_), .B(ori_ori_n74_), .C(i), .Y(ori_ori_n870_));
  OR2        o0842(.A(ori_ori_n870_), .B(ori_ori_n869_), .Y(ori_ori_n871_));
  NA3        o0843(.A(ori_ori_n291_), .B(ori_ori_n112_), .C(g), .Y(ori_ori_n872_));
  AOI210     o0844(.A0(ori_ori_n611_), .A1(ori_ori_n872_), .B0(m), .Y(ori_ori_n873_));
  OAI210     o0845(.A0(ori_ori_n873_), .A1(ori_ori_n825_), .B0(ori_ori_n290_), .Y(ori_ori_n874_));
  NA2        o0846(.A(ori_ori_n624_), .B(ori_ori_n779_), .Y(ori_ori_n875_));
  INV        o0847(.A(ori_ori_n388_), .Y(ori_ori_n876_));
  INV        o0848(.A(ori_ori_n870_), .Y(ori_ori_n877_));
  AOI220     o0849(.A0(ori_ori_n877_), .A1(ori_ori_n242_), .B0(ori_ori_n876_), .B1(ori_ori_n875_), .Y(ori_ori_n878_));
  NA4        o0850(.A(ori_ori_n878_), .B(ori_ori_n874_), .C(ori_ori_n871_), .D(ori_ori_n868_), .Y(ori_ori_n879_));
  NO2        o0851(.A(ori_ori_n336_), .B(ori_ori_n85_), .Y(ori_ori_n880_));
  OAI210     o0852(.A0(ori_ori_n880_), .A1(ori_ori_n833_), .B0(ori_ori_n224_), .Y(ori_ori_n881_));
  NA2        o0853(.A(ori_ori_n600_), .B(ori_ori_n82_), .Y(ori_ori_n882_));
  NO2        o0854(.A(ori_ori_n408_), .B(ori_ori_n200_), .Y(ori_ori_n883_));
  AOI220     o0855(.A0(ori_ori_n883_), .A1(ori_ori_n340_), .B0(ori_ori_n839_), .B1(ori_ori_n204_), .Y(ori_ori_n884_));
  AOI220     o0856(.A0(ori_ori_n826_), .A1(ori_ori_n836_), .B0(ori_ori_n526_), .B1(ori_ori_n84_), .Y(ori_ori_n885_));
  NA4        o0857(.A(ori_ori_n885_), .B(ori_ori_n884_), .C(ori_ori_n882_), .D(ori_ori_n881_), .Y(ori_ori_n886_));
  NA2        o0858(.A(ori_ori_n876_), .B(ori_ori_n481_), .Y(ori_ori_n887_));
  AOI210     o0859(.A0(ori_ori_n375_), .A1(ori_ori_n368_), .B0(ori_ori_n732_), .Y(ori_ori_n888_));
  OAI210     o0860(.A0(ori_ori_n327_), .A1(ori_ori_n326_), .B0(ori_ori_n104_), .Y(ori_ori_n889_));
  AOI210     o0861(.A0(ori_ori_n889_), .A1(ori_ori_n473_), .B0(ori_ori_n888_), .Y(ori_ori_n890_));
  NA2        o0862(.A(ori_ori_n873_), .B(ori_ori_n824_), .Y(ori_ori_n891_));
  NO3        o0863(.A(ori_ori_n793_), .B(ori_ori_n46_), .C(ori_ori_n42_), .Y(ori_ori_n892_));
  AOI220     o0864(.A0(ori_ori_n892_), .A1(ori_ori_n564_), .B0(ori_ori_n581_), .B1(ori_ori_n469_), .Y(ori_ori_n893_));
  NA4        o0865(.A(ori_ori_n893_), .B(ori_ori_n891_), .C(ori_ori_n890_), .D(ori_ori_n887_), .Y(ori_ori_n894_));
  NO4        o0866(.A(ori_ori_n894_), .B(ori_ori_n886_), .C(ori_ori_n879_), .D(ori_ori_n865_), .Y(ori_ori_n895_));
  NAi31      o0867(.An(ori_ori_n132_), .B(ori_ori_n376_), .C(n), .Y(ori_ori_n896_));
  NO3        o0868(.A(ori_ori_n118_), .B(ori_ori_n302_), .C(ori_ori_n756_), .Y(ori_ori_n897_));
  NO2        o0869(.A(ori_ori_n897_), .B(ori_ori_n896_), .Y(ori_ori_n898_));
  NA2        o0870(.A(ori_ori_n217_), .B(ori_ori_n163_), .Y(ori_ori_n899_));
  NO3        o0871(.A(ori_ori_n276_), .B(ori_ori_n393_), .C(ori_ori_n167_), .Y(ori_ori_n900_));
  NOi31      o0872(.An(ori_ori_n899_), .B(ori_ori_n900_), .C(ori_ori_n200_), .Y(ori_ori_n901_));
  NAi21      o0873(.An(ori_ori_n492_), .B(ori_ori_n883_), .Y(ori_ori_n902_));
  INV        o0874(.A(ori_ori_n902_), .Y(ori_ori_n903_));
  OAI220     o0875(.A0(ori_ori_n896_), .A1(ori_ori_n220_), .B0(ori_ori_n866_), .B1(ori_ori_n541_), .Y(ori_ori_n904_));
  NO2        o0876(.A(ori_ori_n597_), .B(ori_ori_n336_), .Y(ori_ori_n905_));
  NA2        o0877(.A(ori_ori_n829_), .B(ori_ori_n820_), .Y(ori_ori_n906_));
  OAI220     o0878(.A0(ori_ori_n826_), .A1(ori_ori_n834_), .B0(ori_ori_n483_), .B1(ori_ori_n379_), .Y(ori_ori_n907_));
  NA3        o0879(.A(ori_ori_n907_), .B(ori_ori_n906_), .C(ori_ori_n558_), .Y(ori_ori_n908_));
  OAI210     o0880(.A0(ori_ori_n829_), .A1(ori_ori_n821_), .B0(ori_ori_n899_), .Y(ori_ori_n909_));
  NA3        o0881(.A(ori_ori_n863_), .B(ori_ori_n429_), .C(ori_ori_n43_), .Y(ori_ori_n910_));
  INV        o0882(.A(ori_ori_n294_), .Y(ori_ori_n911_));
  NA4        o0883(.A(ori_ori_n911_), .B(ori_ori_n910_), .C(ori_ori_n909_), .D(ori_ori_n250_), .Y(ori_ori_n912_));
  OR4        o0884(.A(ori_ori_n912_), .B(ori_ori_n908_), .C(ori_ori_n905_), .D(ori_ori_n904_), .Y(ori_ori_n913_));
  NO4        o0885(.A(ori_ori_n913_), .B(ori_ori_n903_), .C(ori_ori_n901_), .D(ori_ori_n898_), .Y(ori_ori_n914_));
  NA4        o0886(.A(ori_ori_n914_), .B(ori_ori_n895_), .C(ori_ori_n857_), .D(ori_ori_n846_), .Y(ori13));
  AN2        o0887(.A(d), .B(c), .Y(ori_ori_n916_));
  NA2        o0888(.A(ori_ori_n916_), .B(ori_ori_n110_), .Y(ori_ori_n917_));
  NAi32      o0889(.An(f), .Bn(e), .C(c), .Y(ori_ori_n918_));
  NO3        o0890(.A(m), .B(i), .C(h), .Y(ori_ori_n919_));
  OR2        o0891(.A(d), .B(c), .Y(ori_ori_n920_));
  NA3        o0892(.A(k), .B(j), .C(i), .Y(ori_ori_n921_));
  NO3        o0893(.A(ori_ori_n921_), .B(ori_ori_n275_), .C(ori_ori_n85_), .Y(ori_ori_n922_));
  NOi21      o0894(.An(ori_ori_n922_), .B(ori_ori_n920_), .Y(ori_ori_n923_));
  NA2        o0895(.A(ori_ori_n414_), .B(ori_ori_n296_), .Y(ori_ori_n924_));
  NO4        o0896(.A(ori_ori_n924_), .B(ori_ori_n524_), .C(ori_ori_n399_), .D(ori_ori_n42_), .Y(ori05));
  OR2        o0897(.A(ori05), .B(ori_ori_n923_), .Y(ori02));
  OR2        o0898(.A(l), .B(k), .Y(ori_ori_n927_));
  OR3        o0899(.A(h), .B(g), .C(f), .Y(ori_ori_n928_));
  OR3        o0900(.A(n), .B(m), .C(i), .Y(ori_ori_n929_));
  NO4        o0901(.A(ori_ori_n929_), .B(ori_ori_n928_), .C(ori_ori_n927_), .D(ori_ori_n920_), .Y(ori03));
  AN3        o0902(.A(g), .B(f), .C(c), .Y(ori_ori_n931_));
  NA3        o0903(.A(l), .B(k), .C(j), .Y(ori_ori_n932_));
  NA2        o0904(.A(i), .B(h), .Y(ori_ori_n933_));
  NO3        o0905(.A(ori_ori_n933_), .B(ori_ori_n932_), .C(ori_ori_n124_), .Y(ori_ori_n934_));
  NO3        o0906(.A(ori_ori_n133_), .B(ori_ori_n258_), .C(ori_ori_n200_), .Y(ori_ori_n935_));
  NA3        o0907(.A(c), .B(b), .C(a), .Y(ori_ori_n936_));
  NO2        o0908(.A(ori_ori_n465_), .B(ori_ori_n537_), .Y(ori_ori_n937_));
  NA4        o0909(.A(ori_ori_n82_), .B(ori_ori_n81_), .C(g), .D(ori_ori_n199_), .Y(ori_ori_n938_));
  NA4        o0910(.A(ori_ori_n512_), .B(m), .C(ori_ori_n107_), .D(ori_ori_n199_), .Y(ori_ori_n939_));
  NA3        o0911(.A(ori_ori_n939_), .B(ori_ori_n328_), .C(ori_ori_n938_), .Y(ori_ori_n940_));
  NO3        o0912(.A(ori_ori_n940_), .B(ori_ori_n937_), .C(ori_ori_n889_), .Y(ori_ori_n941_));
  NOi41      o0913(.An(ori_ori_n717_), .B(ori_ori_n761_), .C(ori_ori_n750_), .D(ori_ori_n645_), .Y(ori_ori_n942_));
  OAI220     o0914(.A0(ori_ori_n942_), .A1(ori_ori_n624_), .B0(ori_ori_n941_), .B1(ori_ori_n525_), .Y(ori_ori_n943_));
  NOi31      o0915(.An(m), .B(n), .C(f), .Y(ori_ori_n944_));
  NA2        o0916(.A(ori_ori_n944_), .B(ori_ori_n48_), .Y(ori_ori_n945_));
  NA2        o0917(.A(ori_ori_n446_), .B(l), .Y(ori_ori_n946_));
  NO2        o0918(.A(ori_ori_n81_), .B(g), .Y(ori_ori_n947_));
  NO4        o0919(.A(ori_ori_n888_), .B(ori_ori_n943_), .C(ori_ori_n733_), .D(ori_ori_n501_), .Y(ori_ori_n948_));
  NA2        o0920(.A(c), .B(b), .Y(ori_ori_n949_));
  NO2        o0921(.A(ori_ori_n634_), .B(ori_ori_n949_), .Y(ori_ori_n950_));
  OAI210     o0922(.A0(ori_ori_n765_), .A1(ori_ori_n742_), .B0(ori_ori_n371_), .Y(ori_ori_n951_));
  OAI210     o0923(.A0(ori_ori_n951_), .A1(ori_ori_n766_), .B0(ori_ori_n950_), .Y(ori_ori_n952_));
  NAi21      o0924(.An(ori_ori_n375_), .B(ori_ori_n950_), .Y(ori_ori_n953_));
  NA3        o0925(.A(ori_ori_n379_), .B(ori_ori_n497_), .C(f), .Y(ori_ori_n954_));
  NA2        o0926(.A(ori_ori_n954_), .B(ori_ori_n953_), .Y(ori_ori_n955_));
  INV        o0927(.A(ori_ori_n244_), .Y(ori_ori_n956_));
  OAI210     o0928(.A0(ori_ori_n956_), .A1(ori_ori_n262_), .B0(g), .Y(ori_ori_n957_));
  NAi21      o0929(.An(f), .B(d), .Y(ori_ori_n958_));
  NO2        o0930(.A(ori_ori_n958_), .B(ori_ori_n936_), .Y(ori_ori_n959_));
  INV        o0931(.A(ori_ori_n959_), .Y(ori_ori_n960_));
  NO2        o0932(.A(ori_ori_n957_), .B(ori_ori_n960_), .Y(ori_ori_n961_));
  AOI210     o0933(.A0(ori_ori_n961_), .A1(ori_ori_n108_), .B0(ori_ori_n955_), .Y(ori_ori_n962_));
  NO2        o0934(.A(ori_ori_n174_), .B(ori_ori_n223_), .Y(ori_ori_n963_));
  NA2        o0935(.A(ori_ori_n963_), .B(m), .Y(ori_ori_n964_));
  NA3        o0936(.A(ori_ori_n810_), .B(ori_ori_n946_), .C(ori_ori_n1225_), .Y(ori_ori_n965_));
  INV        o0937(.A(ori_ori_n417_), .Y(ori_ori_n966_));
  NO2        o0938(.A(ori_ori_n966_), .B(ori_ori_n964_), .Y(ori_ori_n967_));
  NA2        o0939(.A(ori_ori_n396_), .B(ori_ori_n959_), .Y(ori_ori_n968_));
  NO2        o0940(.A(ori_ori_n330_), .B(ori_ori_n329_), .Y(ori_ori_n969_));
  NA2        o0941(.A(ori_ori_n963_), .B(ori_ori_n381_), .Y(ori_ori_n970_));
  NAi31      o0942(.An(ori_ori_n969_), .B(ori_ori_n970_), .C(ori_ori_n968_), .Y(ori_ori_n971_));
  NO2        o0943(.A(ori_ori_n971_), .B(ori_ori_n967_), .Y(ori_ori_n972_));
  NA4        o0944(.A(ori_ori_n972_), .B(ori_ori_n962_), .C(ori_ori_n952_), .D(ori_ori_n948_), .Y(ori00));
  INV        o0945(.A(ori_ori_n890_), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n448_), .B(f), .Y(ori_ori_n975_));
  OAI210     o0947(.A0(ori_ori_n897_), .A1(ori_ori_n39_), .B0(ori_ori_n583_), .Y(ori_ori_n976_));
  NA3        o0948(.A(ori_ori_n976_), .B(ori_ori_n241_), .C(n), .Y(ori_ori_n977_));
  AOI210     o0949(.A0(ori_ori_n977_), .A1(ori_ori_n975_), .B0(ori_ori_n917_), .Y(ori_ori_n978_));
  NO3        o0950(.A(ori_ori_n978_), .B(ori_ori_n974_), .C(ori_ori_n923_), .Y(ori_ori_n979_));
  NA3        o0951(.A(d), .B(ori_ori_n53_), .C(b), .Y(ori_ori_n980_));
  INV        o0952(.A(ori_ori_n514_), .Y(ori_ori_n981_));
  NO2        o0953(.A(ori_ori_n981_), .B(ori_ori_n969_), .Y(ori_ori_n982_));
  NO4        o0954(.A(ori_ori_n430_), .B(ori_ori_n314_), .C(ori_ori_n949_), .D(ori_ori_n56_), .Y(ori_ori_n983_));
  NA3        o0955(.A(ori_ori_n341_), .B(ori_ori_n207_), .C(g), .Y(ori_ori_n984_));
  OA220      o0956(.A0(ori_ori_n984_), .A1(ori_ori_n980_), .B0(ori_ori_n342_), .B1(ori_ori_n125_), .Y(ori_ori_n985_));
  NO2        o0957(.A(h), .B(g), .Y(ori_ori_n986_));
  OAI220     o0958(.A0(ori_ori_n465_), .A1(ori_ori_n537_), .B0(ori_ori_n86_), .B1(ori_ori_n85_), .Y(ori_ori_n987_));
  AOI220     o0959(.A0(ori_ori_n987_), .A1(ori_ori_n473_), .B0(ori_ori_n841_), .B1(ori_ori_n513_), .Y(ori_ori_n988_));
  AOI220     o0960(.A0(ori_ori_n284_), .A1(ori_ori_n230_), .B0(ori_ori_n169_), .B1(ori_ori_n140_), .Y(ori_ori_n989_));
  NA3        o0961(.A(ori_ori_n989_), .B(ori_ori_n988_), .C(ori_ori_n985_), .Y(ori_ori_n990_));
  NO2        o0962(.A(ori_ori_n990_), .B(ori_ori_n983_), .Y(ori_ori_n991_));
  INV        o0963(.A(ori_ori_n288_), .Y(ori_ori_n992_));
  NA2        o0964(.A(ori_ori_n230_), .B(ori_ori_n306_), .Y(ori_ori_n993_));
  NA3        o0965(.A(ori_ori_n993_), .B(ori_ori_n992_), .C(ori_ori_n146_), .Y(ori_ori_n994_));
  NO3        o0966(.A(ori03), .B(ori_ori_n994_), .C(ori_ori_n458_), .Y(ori_ori_n995_));
  AN3        o0967(.A(ori_ori_n995_), .B(ori_ori_n991_), .C(ori_ori_n982_), .Y(ori_ori_n996_));
  NA2        o0968(.A(ori_ori_n473_), .B(ori_ori_n96_), .Y(ori_ori_n997_));
  NA2        o0969(.A(ori_ori_n997_), .B(ori_ori_n227_), .Y(ori_ori_n998_));
  NA2        o0970(.A(ori_ori_n940_), .B(ori_ori_n473_), .Y(ori_ori_n999_));
  NA4        o0971(.A(ori_ori_n586_), .B(ori_ori_n192_), .C(ori_ori_n207_), .D(ori_ori_n155_), .Y(ori_ori_n1000_));
  NA2        o0972(.A(ori_ori_n1000_), .B(ori_ori_n999_), .Y(ori_ori_n1001_));
  OAI210     o0973(.A0(ori_ori_n413_), .A1(ori_ori_n113_), .B0(ori_ori_n768_), .Y(ori_ori_n1002_));
  NA2        o0974(.A(ori_ori_n1002_), .B(ori_ori_n965_), .Y(ori_ori_n1003_));
  NA2        o0975(.A(n), .B(e), .Y(ori_ori_n1004_));
  NO2        o0976(.A(ori_ori_n1004_), .B(ori_ori_n138_), .Y(ori_ori_n1005_));
  NA2        o0977(.A(ori_ori_n1005_), .B(ori_ori_n251_), .Y(ori_ori_n1006_));
  OAI210     o0978(.A0(ori_ori_n315_), .A1(ori_ori_n280_), .B0(ori_ori_n398_), .Y(ori_ori_n1007_));
  NA3        o0979(.A(ori_ori_n1007_), .B(ori_ori_n1006_), .C(ori_ori_n1003_), .Y(ori_ori_n1008_));
  NA2        o0980(.A(ori_ori_n1005_), .B(ori_ori_n758_), .Y(ori_ori_n1009_));
  NA2        o0981(.A(ori_ori_n1009_), .B(ori_ori_n770_), .Y(ori_ori_n1010_));
  NO4        o0982(.A(ori_ori_n1010_), .B(ori_ori_n1008_), .C(ori_ori_n1001_), .D(ori_ori_n998_), .Y(ori_ori_n1011_));
  NA2        o0983(.A(ori_ori_n743_), .B(ori_ori_n681_), .Y(ori_ori_n1012_));
  NA4        o0984(.A(ori_ori_n1012_), .B(ori_ori_n1011_), .C(ori_ori_n996_), .D(ori_ori_n979_), .Y(ori01));
  INV        o0985(.A(ori_ori_n256_), .Y(ori_ori_n1014_));
  NA2        o0986(.A(ori_ori_n352_), .B(i), .Y(ori_ori_n1015_));
  NA3        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1014_), .C(ori_ori_n906_), .Y(ori_ori_n1016_));
  NA2        o0988(.A(ori_ori_n526_), .B(ori_ori_n84_), .Y(ori_ori_n1017_));
  NA2        o0989(.A(ori_ori_n492_), .B(ori_ori_n248_), .Y(ori_ori_n1018_));
  NA2        o0990(.A(ori_ori_n853_), .B(ori_ori_n1018_), .Y(ori_ori_n1019_));
  NA3        o0991(.A(ori_ori_n1019_), .B(ori_ori_n1017_), .C(ori_ori_n806_), .Y(ori_ori_n1020_));
  NA2        o0992(.A(ori_ori_n42_), .B(f), .Y(ori_ori_n1021_));
  NA2        o0993(.A(ori_ori_n640_), .B(ori_ori_n91_), .Y(ori_ori_n1022_));
  NO2        o0994(.A(ori_ori_n1022_), .B(ori_ori_n1021_), .Y(ori_ori_n1023_));
  OAI210     o0995(.A0(ori_ori_n699_), .A1(ori_ori_n541_), .B0(ori_ori_n1000_), .Y(ori_ori_n1024_));
  INV        o0996(.A(ori_ori_n1024_), .Y(ori_ori_n1025_));
  INV        o0997(.A(ori_ori_n112_), .Y(ori_ori_n1026_));
  OA220      o0998(.A0(ori_ori_n1026_), .A1(ori_ori_n523_), .B0(ori_ori_n598_), .B1(ori_ori_n328_), .Y(ori_ori_n1027_));
  NAi41      o0999(.An(ori_ori_n154_), .B(ori_ori_n1027_), .C(ori_ori_n1025_), .D(ori_ori_n795_), .Y(ori_ori_n1028_));
  NO2        o1000(.A(ori_ori_n612_), .B(ori_ori_n451_), .Y(ori_ori_n1029_));
  NA4        o1001(.A(ori_ori_n640_), .B(ori_ori_n91_), .C(ori_ori_n42_), .D(ori_ori_n199_), .Y(ori_ori_n1030_));
  OR2        o1002(.A(ori_ori_n182_), .B(ori_ori_n180_), .Y(ori_ori_n1031_));
  NA3        o1003(.A(ori_ori_n1031_), .B(ori_ori_n1029_), .C(ori_ori_n128_), .Y(ori_ori_n1032_));
  NO4        o1004(.A(ori_ori_n1032_), .B(ori_ori_n1028_), .C(ori_ori_n1020_), .D(ori_ori_n1016_), .Y(ori_ori_n1033_));
  INV        o1005(.A(ori_ori_n984_), .Y(ori_ori_n1034_));
  OAI210     o1006(.A0(ori_ori_n1034_), .A1(ori_ori_n271_), .B0(ori_ori_n469_), .Y(ori_ori_n1035_));
  NA2        o1007(.A(ori_ori_n476_), .B(ori_ori_n354_), .Y(ori_ori_n1036_));
  NOi21      o1008(.An(ori_ori_n498_), .B(ori_ori_n520_), .Y(ori_ori_n1037_));
  NA2        o1009(.A(ori_ori_n1037_), .B(ori_ori_n1036_), .Y(ori_ori_n1038_));
  AOI210     o1010(.A0(ori_ori_n191_), .A1(ori_ori_n83_), .B0(ori_ori_n199_), .Y(ori_ori_n1039_));
  OAI210     o1011(.A0(ori_ori_n720_), .A1(ori_ori_n379_), .B0(ori_ori_n1039_), .Y(ori_ori_n1040_));
  AN3        o1012(.A(m), .B(l), .C(k), .Y(ori_ori_n1041_));
  OAI210     o1013(.A0(ori_ori_n317_), .A1(ori_ori_n33_), .B0(ori_ori_n1041_), .Y(ori_ori_n1042_));
  NA2        o1014(.A(ori_ori_n190_), .B(ori_ori_n33_), .Y(ori_ori_n1043_));
  AO210      o1015(.A0(ori_ori_n1043_), .A1(ori_ori_n1042_), .B0(ori_ori_n295_), .Y(ori_ori_n1044_));
  NA4        o1016(.A(ori_ori_n1044_), .B(ori_ori_n1040_), .C(ori_ori_n1038_), .D(ori_ori_n1035_), .Y(ori_ori_n1045_));
  AOI210     o1017(.A0(ori_ori_n535_), .A1(ori_ori_n112_), .B0(ori_ori_n539_), .Y(ori_ori_n1046_));
  OAI210     o1018(.A0(ori_ori_n1026_), .A1(ori_ori_n532_), .B0(ori_ori_n1046_), .Y(ori_ori_n1047_));
  NA2        o1019(.A(ori_ori_n255_), .B(ori_ori_n182_), .Y(ori_ori_n1048_));
  NA2        o1020(.A(ori_ori_n1048_), .B(ori_ori_n603_), .Y(ori_ori_n1049_));
  NA2        o1021(.A(ori_ori_n1023_), .B(ori_ori_n613_), .Y(ori_ori_n1050_));
  NA3        o1022(.A(ori_ori_n1050_), .B(ori_ori_n1049_), .C(ori_ori_n701_), .Y(ori_ori_n1051_));
  NO3        o1023(.A(ori_ori_n1051_), .B(ori_ori_n1047_), .C(ori_ori_n1045_), .Y(ori_ori_n1052_));
  NA3        o1024(.A(ori_ori_n542_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1053_));
  NO2        o1025(.A(ori_ori_n1053_), .B(ori_ori_n191_), .Y(ori_ori_n1054_));
  AOI210     o1026(.A0(ori_ori_n445_), .A1(ori_ori_n55_), .B0(ori_ori_n1054_), .Y(ori_ori_n1055_));
  OR3        o1027(.A(ori_ori_n1022_), .B(ori_ori_n543_), .C(ori_ori_n1021_), .Y(ori_ori_n1056_));
  NO2        o1028(.A(ori_ori_n1030_), .B(ori_ori_n869_), .Y(ori_ori_n1057_));
  NO2        o1029(.A(ori_ori_n193_), .B(ori_ori_n106_), .Y(ori_ori_n1058_));
  NO2        o1030(.A(ori_ori_n1058_), .B(ori_ori_n1057_), .Y(ori_ori_n1059_));
  NA4        o1031(.A(ori_ori_n1059_), .B(ori_ori_n1056_), .C(ori_ori_n1055_), .D(ori_ori_n680_), .Y(ori_ori_n1060_));
  NO2        o1032(.A(ori_ori_n859_), .B(ori_ori_n219_), .Y(ori_ori_n1061_));
  NO2        o1033(.A(ori_ori_n860_), .B(ori_ori_n494_), .Y(ori_ori_n1062_));
  OAI210     o1034(.A0(ori_ori_n1062_), .A1(ori_ori_n1061_), .B0(ori_ori_n302_), .Y(ori_ori_n1063_));
  NA2        o1035(.A(ori_ori_n508_), .B(ori_ori_n506_), .Y(ori_ori_n1064_));
  NO3        o1036(.A(ori_ori_n73_), .B(ori_ori_n269_), .C(ori_ori_n42_), .Y(ori_ori_n1065_));
  NA2        o1037(.A(ori_ori_n1065_), .B(ori_ori_n491_), .Y(ori_ori_n1066_));
  NA3        o1038(.A(ori_ori_n1066_), .B(ori_ori_n1064_), .C(ori_ori_n608_), .Y(ori_ori_n1067_));
  OR2        o1039(.A(ori_ori_n984_), .B(ori_ori_n980_), .Y(ori_ori_n1068_));
  NO2        o1040(.A(ori_ori_n328_), .B(ori_ori_n66_), .Y(ori_ori_n1069_));
  INV        o1041(.A(ori_ori_n1069_), .Y(ori_ori_n1070_));
  NA2        o1042(.A(ori_ori_n1065_), .B(ori_ori_n723_), .Y(ori_ori_n1071_));
  NA4        o1043(.A(ori_ori_n1071_), .B(ori_ori_n1070_), .C(ori_ori_n1068_), .D(ori_ori_n344_), .Y(ori_ori_n1072_));
  NOi41      o1044(.An(ori_ori_n1063_), .B(ori_ori_n1072_), .C(ori_ori_n1067_), .D(ori_ori_n1060_), .Y(ori_ori_n1073_));
  INV        o1045(.A(ori_ori_n125_), .Y(ori_ori_n1074_));
  NO3        o1046(.A(ori_ori_n933_), .B(ori_ori_n168_), .C(ori_ori_n81_), .Y(ori_ori_n1075_));
  AOI220     o1047(.A0(ori_ori_n1075_), .A1(ori_ori_n1074_), .B0(ori_ori_n1065_), .B1(ori_ori_n861_), .Y(ori_ori_n1076_));
  INV        o1048(.A(ori_ori_n1076_), .Y(ori_ori_n1077_));
  NO2        o1049(.A(ori_ori_n554_), .B(ori_ori_n553_), .Y(ori_ori_n1078_));
  NO4        o1050(.A(ori_ori_n933_), .B(ori_ori_n1078_), .C(ori_ori_n166_), .D(ori_ori_n81_), .Y(ori_ori_n1079_));
  NO3        o1051(.A(ori_ori_n1079_), .B(ori_ori_n1077_), .C(ori_ori_n575_), .Y(ori_ori_n1080_));
  NA4        o1052(.A(ori_ori_n1080_), .B(ori_ori_n1073_), .C(ori_ori_n1052_), .D(ori_ori_n1033_), .Y(ori06));
  NO2        o1053(.A(ori_ori_n211_), .B(ori_ori_n97_), .Y(ori_ori_n1082_));
  OAI210     o1054(.A0(ori_ori_n1082_), .A1(ori_ori_n1075_), .B0(ori_ori_n340_), .Y(ori_ori_n1083_));
  NO3        o1055(.A(ori_ori_n538_), .B(ori_ori_n718_), .C(ori_ori_n540_), .Y(ori_ori_n1084_));
  OR2        o1056(.A(ori_ori_n1084_), .B(ori_ori_n787_), .Y(ori_ori_n1085_));
  NA3        o1057(.A(ori_ori_n1085_), .B(ori_ori_n1083_), .C(ori_ori_n1063_), .Y(ori_ori_n1086_));
  NO3        o1058(.A(ori_ori_n1086_), .B(ori_ori_n1067_), .C(ori_ori_n240_), .Y(ori_ori_n1087_));
  NO2        o1059(.A(ori_ori_n269_), .B(ori_ori_n42_), .Y(ori_ori_n1088_));
  AOI210     o1060(.A0(ori_ori_n1088_), .A1(ori_ori_n862_), .B0(ori_ori_n1061_), .Y(ori_ori_n1089_));
  NA2        o1061(.A(ori_ori_n1088_), .B(ori_ori_n495_), .Y(ori_ori_n1090_));
  AOI210     o1062(.A0(ori_ori_n1090_), .A1(ori_ori_n1089_), .B0(ori_ori_n300_), .Y(ori_ori_n1091_));
  NO2        o1063(.A(ori_ori_n83_), .B(ori_ori_n39_), .Y(ori_ori_n1092_));
  NA2        o1064(.A(ori_ori_n1092_), .B(ori_ori_n579_), .Y(ori_ori_n1093_));
  NOi21      o1065(.An(ori_ori_n127_), .B(ori_ori_n42_), .Y(ori_ori_n1094_));
  NO2        o1066(.A(ori_ori_n547_), .B(ori_ori_n945_), .Y(ori_ori_n1095_));
  NO2        o1067(.A(ori_ori_n409_), .B(ori_ori_n231_), .Y(ori_ori_n1096_));
  NO3        o1068(.A(ori_ori_n1096_), .B(ori_ori_n1095_), .C(ori_ori_n1094_), .Y(ori_ori_n1097_));
  INV        o1069(.A(ori_ori_n539_), .Y(ori_ori_n1098_));
  NA3        o1070(.A(ori_ori_n1098_), .B(ori_ori_n1097_), .C(ori_ori_n1093_), .Y(ori_ori_n1099_));
  AN2        o1071(.A(ori_ori_n848_), .B(ori_ori_n582_), .Y(ori_ori_n1100_));
  NO3        o1072(.A(ori_ori_n1100_), .B(ori_ori_n1099_), .C(ori_ori_n1091_), .Y(ori_ori_n1101_));
  NO3        o1073(.A(h), .B(ori_ori_n97_), .C(ori_ori_n258_), .Y(ori_ori_n1102_));
  OAI220     o1074(.A0(ori_ori_n631_), .A1(ori_ori_n231_), .B0(ori_ori_n450_), .B1(ori_ori_n454_), .Y(ori_ori_n1103_));
  INV        o1075(.A(k), .Y(ori_ori_n1104_));
  NO3        o1076(.A(ori_ori_n1104_), .B(ori_ori_n537_), .C(j), .Y(ori_ori_n1105_));
  NOi21      o1077(.An(ori_ori_n1105_), .B(ori_ori_n606_), .Y(ori_ori_n1106_));
  NO3        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1103_), .C(ori_ori_n1102_), .Y(ori_ori_n1107_));
  NA4        o1079(.A(ori_ori_n707_), .B(ori_ori_n706_), .C(ori_ori_n386_), .D(ori_ori_n779_), .Y(ori_ori_n1108_));
  NAi31      o1080(.An(ori_ori_n672_), .B(ori_ori_n1108_), .C(ori_ori_n190_), .Y(ori_ori_n1109_));
  NA2        o1081(.A(ori_ori_n1109_), .B(ori_ori_n1107_), .Y(ori_ori_n1110_));
  OR3        o1082(.A(ori_ori_n1084_), .B(ori_ori_n699_), .C(ori_ori_n479_), .Y(ori_ori_n1111_));
  AOI210     o1083(.A0(ori_ori_n508_), .A1(ori_ori_n398_), .B0(ori_ori_n331_), .Y(ori_ori_n1112_));
  NA2        o1084(.A(ori_ori_n1105_), .B(ori_ori_n703_), .Y(ori_ori_n1113_));
  NA3        o1085(.A(ori_ori_n1113_), .B(ori_ori_n1112_), .C(ori_ori_n1111_), .Y(ori_ori_n1114_));
  AN2        o1086(.A(ori_ori_n821_), .B(ori_ori_n820_), .Y(ori_ori_n1115_));
  NO2        o1087(.A(ori_ori_n1115_), .B(ori_ori_n441_), .Y(ori_ori_n1116_));
  NA2        o1088(.A(ori_ori_n1116_), .B(ori_ori_n1071_), .Y(ori_ori_n1117_));
  NAi21      o1089(.An(j), .B(i), .Y(ori_ori_n1118_));
  NO4        o1090(.A(ori_ori_n1078_), .B(ori_ori_n1118_), .C(ori_ori_n392_), .D(ori_ori_n221_), .Y(ori_ori_n1119_));
  NO4        o1091(.A(ori_ori_n1119_), .B(ori_ori_n1117_), .C(ori_ori_n1114_), .D(ori_ori_n1110_), .Y(ori_ori_n1120_));
  NA4        o1092(.A(ori_ori_n1120_), .B(ori_ori_n1101_), .C(ori_ori_n1087_), .D(ori_ori_n1080_), .Y(ori07));
  NOi21      o1093(.An(j), .B(k), .Y(ori_ori_n1122_));
  NA4        o1094(.A(ori_ori_n171_), .B(ori_ori_n103_), .C(ori_ori_n1122_), .D(f), .Y(ori_ori_n1123_));
  NAi32      o1095(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1124_));
  NO3        o1096(.A(ori_ori_n1124_), .B(g), .C(f), .Y(ori_ori_n1125_));
  INV        o1097(.A(ori_ori_n1125_), .Y(ori_ori_n1126_));
  OR2        o1098(.A(e), .B(d), .Y(ori_ori_n1127_));
  NOi31      o1099(.An(n), .B(m), .C(b), .Y(ori_ori_n1128_));
  NO3        o1100(.A(ori_ori_n124_), .B(ori_ori_n399_), .C(h), .Y(ori_ori_n1129_));
  NA2        o1101(.A(ori_ori_n1126_), .B(ori_ori_n1123_), .Y(ori_ori_n1130_));
  NOi41      o1102(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1131_));
  NO2        o1103(.A(ori_ori_n918_), .B(ori_ori_n392_), .Y(ori_ori_n1132_));
  INV        o1104(.A(ori_ori_n1132_), .Y(ori_ori_n1133_));
  NO2        o1105(.A(ori_ori_n921_), .B(ori_ori_n275_), .Y(ori_ori_n1134_));
  NA2        o1106(.A(ori_ori_n480_), .B(ori_ori_n74_), .Y(ori_ori_n1135_));
  NA2        o1107(.A(ori_ori_n1135_), .B(ori_ori_n1133_), .Y(ori_ori_n1136_));
  NO2        o1108(.A(ori_ori_n1136_), .B(ori_ori_n1130_), .Y(ori_ori_n1137_));
  NO3        o1109(.A(e), .B(d), .C(c), .Y(ori_ori_n1138_));
  NO2        o1110(.A(ori_ori_n124_), .B(ori_ori_n200_), .Y(ori_ori_n1139_));
  NA2        o1111(.A(ori_ori_n1139_), .B(ori_ori_n1138_), .Y(ori_ori_n1140_));
  INV        o1112(.A(ori_ori_n1140_), .Y(ori_ori_n1141_));
  NA3        o1113(.A(ori_ori_n628_), .B(ori_ori_n616_), .C(ori_ori_n107_), .Y(ori_ori_n1142_));
  NO2        o1114(.A(ori_ori_n1142_), .B(ori_ori_n42_), .Y(ori_ori_n1143_));
  NO2        o1115(.A(l), .B(k), .Y(ori_ori_n1144_));
  NO2        o1116(.A(ori_ori_n1143_), .B(ori_ori_n1141_), .Y(ori_ori_n1145_));
  NO2        o1117(.A(g), .B(c), .Y(ori_ori_n1146_));
  NO2        o1118(.A(ori_ori_n400_), .B(a), .Y(ori_ori_n1147_));
  NA2        o1119(.A(ori_ori_n1147_), .B(ori_ori_n108_), .Y(ori_ori_n1148_));
  NO2        o1120(.A(ori_ori_n679_), .B(ori_ori_n177_), .Y(ori_ori_n1149_));
  NOi31      o1121(.An(m), .B(n), .C(b), .Y(ori_ori_n1150_));
  NOi31      o1122(.An(f), .B(d), .C(c), .Y(ori_ori_n1151_));
  NA2        o1123(.A(ori_ori_n1151_), .B(ori_ori_n1150_), .Y(ori_ori_n1152_));
  INV        o1124(.A(ori_ori_n1152_), .Y(ori_ori_n1153_));
  NO2        o1125(.A(ori_ori_n1153_), .B(ori_ori_n1149_), .Y(ori_ori_n1154_));
  NA2        o1126(.A(ori_ori_n931_), .B(ori_ori_n414_), .Y(ori_ori_n1155_));
  NO2        o1127(.A(ori_ori_n1155_), .B(ori_ori_n392_), .Y(ori_ori_n1156_));
  NO2        o1128(.A(ori_ori_n919_), .B(ori_ori_n1156_), .Y(ori_ori_n1157_));
  AN3        o1129(.A(ori_ori_n1157_), .B(ori_ori_n1154_), .C(ori_ori_n1148_), .Y(ori_ori_n1158_));
  NA2        o1130(.A(ori_ori_n1128_), .B(ori_ori_n337_), .Y(ori_ori_n1159_));
  INV        o1131(.A(ori_ori_n1159_), .Y(ori_ori_n1160_));
  INV        o1132(.A(ori_ori_n934_), .Y(ori_ori_n1161_));
  NAi21      o1133(.An(ori_ori_n1160_), .B(ori_ori_n1161_), .Y(ori_ori_n1162_));
  NO4        o1134(.A(ori_ori_n124_), .B(g), .C(f), .D(e), .Y(ori_ori_n1163_));
  NA2        o1135(.A(ori_ori_n1131_), .B(ori_ori_n1144_), .Y(ori_ori_n1164_));
  INV        o1136(.A(ori_ori_n1164_), .Y(ori_ori_n1165_));
  OR3        o1137(.A(ori_ori_n479_), .B(ori_ori_n478_), .C(ori_ori_n107_), .Y(ori_ori_n1166_));
  NA2        o1138(.A(ori_ori_n944_), .B(ori_ori_n366_), .Y(ori_ori_n1167_));
  NO2        o1139(.A(ori_ori_n1167_), .B(ori_ori_n385_), .Y(ori_ori_n1168_));
  AO210      o1140(.A0(ori_ori_n1168_), .A1(ori_ori_n110_), .B0(ori_ori_n1165_), .Y(ori_ori_n1169_));
  NO2        o1141(.A(ori_ori_n1169_), .B(ori_ori_n1162_), .Y(ori_ori_n1170_));
  NA4        o1142(.A(ori_ori_n1170_), .B(ori_ori_n1158_), .C(ori_ori_n1145_), .D(ori_ori_n1137_), .Y(ori_ori_n1171_));
  NO2        o1143(.A(ori_ori_n949_), .B(ori_ori_n105_), .Y(ori_ori_n1172_));
  NO2        o1144(.A(ori_ori_n349_), .B(j), .Y(ori_ori_n1173_));
  NA2        o1145(.A(ori_ori_n1173_), .B(ori_ori_n151_), .Y(ori_ori_n1174_));
  INV        o1146(.A(ori_ori_n46_), .Y(ori_ori_n1175_));
  NA2        o1147(.A(ori_ori_n1175_), .B(ori_ori_n986_), .Y(ori_ori_n1176_));
  INV        o1148(.A(ori_ori_n1176_), .Y(ori_ori_n1177_));
  NO2        o1149(.A(ori_ori_n211_), .B(ori_ori_n168_), .Y(ori_ori_n1178_));
  NO2        o1150(.A(ori_ori_n1166_), .B(ori_ori_n311_), .Y(ori_ori_n1179_));
  NO3        o1151(.A(ori_ori_n1179_), .B(ori_ori_n1178_), .C(ori_ori_n1177_), .Y(ori_ori_n1180_));
  NO3        o1152(.A(ori_ori_n936_), .B(ori_ori_n1127_), .C(ori_ori_n46_), .Y(ori_ori_n1181_));
  NA3        o1153(.A(ori_ori_n1172_), .B(ori_ori_n414_), .C(f), .Y(ori_ori_n1182_));
  NO2        o1154(.A(ori_ori_n1220_), .B(ori_ori_n1182_), .Y(ori_ori_n1183_));
  NO2        o1155(.A(ori_ori_n1118_), .B(ori_ori_n166_), .Y(ori_ori_n1184_));
  NOi21      o1156(.An(d), .B(f), .Y(ori_ori_n1185_));
  NA2        o1157(.A(h), .B(ori_ori_n1184_), .Y(ori_ori_n1186_));
  INV        o1158(.A(ori_ori_n1186_), .Y(ori_ori_n1187_));
  NO2        o1159(.A(ori_ori_n1187_), .B(ori_ori_n1183_), .Y(ori_ori_n1188_));
  NA3        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1180_), .C(ori_ori_n1174_), .Y(ori_ori_n1189_));
  NA2        o1161(.A(h), .B(ori_ori_n1134_), .Y(ori_ori_n1190_));
  OAI210     o1162(.A0(ori_ori_n1163_), .A1(ori_ori_n1128_), .B0(ori_ori_n784_), .Y(ori_ori_n1191_));
  NA2        o1163(.A(ori_ori_n1191_), .B(ori_ori_n1190_), .Y(ori_ori_n1192_));
  NA2        o1164(.A(ori_ori_n1146_), .B(ori_ori_n1185_), .Y(ori_ori_n1193_));
  NO2        o1165(.A(ori_ori_n1193_), .B(m), .Y(ori_ori_n1194_));
  NA2        o1166(.A(ori_ori_n935_), .B(ori_ori_n207_), .Y(ori_ori_n1195_));
  NO2        o1167(.A(ori_ori_n143_), .B(ori_ori_n173_), .Y(ori_ori_n1196_));
  OAI210     o1168(.A0(ori_ori_n1196_), .A1(ori_ori_n105_), .B0(ori_ori_n1150_), .Y(ori_ori_n1197_));
  NA2        o1169(.A(ori_ori_n1197_), .B(ori_ori_n1195_), .Y(ori_ori_n1198_));
  NO3        o1170(.A(ori_ori_n1198_), .B(ori_ori_n1194_), .C(ori_ori_n1192_), .Y(ori_ori_n1199_));
  NO2        o1171(.A(ori_ori_n173_), .B(c), .Y(ori_ori_n1200_));
  NA2        o1172(.A(ori_ori_n1200_), .B(ori_ori_n171_), .Y(ori_ori_n1201_));
  AOI210     o1173(.A0(ori_ori_n470_), .A1(ori_ori_n326_), .B0(ori_ori_n1201_), .Y(ori_ori_n1202_));
  INV        o1174(.A(ori_ori_n1181_), .Y(ori_ori_n1203_));
  INV        o1175(.A(ori_ori_n947_), .Y(ori_ori_n1204_));
  OAI210     o1176(.A0(ori_ori_n1204_), .A1(ori_ori_n63_), .B0(ori_ori_n1203_), .Y(ori_ori_n1205_));
  NO2        o1177(.A(ori_ori_n46_), .B(l), .Y(ori_ori_n1206_));
  INV        o1178(.A(ori_ori_n426_), .Y(ori_ori_n1207_));
  NA2        o1179(.A(ori_ori_n1207_), .B(ori_ori_n1206_), .Y(ori_ori_n1208_));
  INV        o1180(.A(ori_ori_n1208_), .Y(ori_ori_n1209_));
  NO3        o1181(.A(ori_ori_n1209_), .B(ori_ori_n1205_), .C(ori_ori_n1202_), .Y(ori_ori_n1210_));
  NA2        o1182(.A(ori_ori_n1210_), .B(ori_ori_n1199_), .Y(ori_ori_n1211_));
  NA3        o1183(.A(ori_ori_n852_), .B(ori_ori_n129_), .C(ori_ori_n43_), .Y(ori_ori_n1212_));
  NOi31      o1184(.An(ori_ori_n30_), .B(m), .C(n), .Y(ori_ori_n1213_));
  INV        o1185(.A(ori_ori_n1213_), .Y(ori_ori_n1214_));
  NO2        o1186(.A(ori_ori_n1167_), .B(d), .Y(ori_ori_n1215_));
  NA4        o1187(.A(ori_ori_n1221_), .B(ori_ori_n1214_), .C(ori_ori_n1222_), .D(ori_ori_n1212_), .Y(ori_ori_n1216_));
  OR4        o1188(.A(ori_ori_n1216_), .B(ori_ori_n1211_), .C(ori_ori_n1189_), .D(ori_ori_n1171_), .Y(ori04));
  INV        o1189(.A(ori_ori_n108_), .Y(ori_ori_n1220_));
  INV        o1190(.A(ori_ori_n1215_), .Y(ori_ori_n1221_));
  INV        o1191(.A(ori_ori_n1129_), .Y(ori_ori_n1222_));
  INV        o1192(.A(ori_ori_n277_), .Y(ori_ori_n1223_));
  INV        o1193(.A(ori_ori_n87_), .Y(ori_ori_n1224_));
  INV        o1194(.A(j), .Y(ori_ori_n1225_));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  INV        m0023(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  INV        m0025(.A(mai_mai_n43_), .Y(mai_mai_n54_));
  NO2        m0026(.A(mai_mai_n54_), .B(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA2        m0031(.A(g), .B(mai_mai_n59_), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi41      m0043(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n72_));
  NA2        m0044(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n73_));
  INV        m0045(.A(m), .Y(mai_mai_n74_));
  NOi21      m0046(.An(k), .B(l), .Y(mai_mai_n75_));
  NA2        m0047(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  AN4        m0048(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n77_));
  NOi31      m0049(.An(h), .B(g), .C(f), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n77_), .Y(mai_mai_n79_));
  NAi32      m0051(.An(m), .Bn(k), .C(j), .Y(mai_mai_n80_));
  NOi32      m0052(.An(h), .Bn(g), .C(f), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n77_), .Y(mai_mai_n82_));
  OA220      m0054(.A0(mai_mai_n82_), .A1(mai_mai_n80_), .B0(mai_mai_n79_), .B1(mai_mai_n76_), .Y(mai_mai_n83_));
  NA3        m0055(.A(mai_mai_n83_), .B(mai_mai_n73_), .C(mai_mai_n64_), .Y(mai_mai_n84_));
  INV        m0056(.A(n), .Y(mai_mai_n85_));
  NOi32      m0057(.An(e), .Bn(b), .C(d), .Y(mai_mai_n86_));
  NA2        m0058(.A(mai_mai_n86_), .B(mai_mai_n85_), .Y(mai_mai_n87_));
  INV        m0059(.A(j), .Y(mai_mai_n88_));
  AN3        m0060(.A(m), .B(k), .C(i), .Y(mai_mai_n89_));
  NA3        m0061(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(g), .Y(mai_mai_n90_));
  NAi32      m0062(.An(g), .Bn(f), .C(h), .Y(mai_mai_n91_));
  NAi31      m0063(.An(j), .B(m), .C(l), .Y(mai_mai_n92_));
  NO2        m0064(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n93_));
  NA2        m0065(.A(m), .B(l), .Y(mai_mai_n94_));
  NAi31      m0066(.An(k), .B(j), .C(g), .Y(mai_mai_n95_));
  NO3        m0067(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(f), .Y(mai_mai_n96_));
  AN2        m0068(.A(j), .B(g), .Y(mai_mai_n97_));
  NOi32      m0069(.An(m), .Bn(l), .C(i), .Y(mai_mai_n98_));
  NOi32      m0070(.An(m), .Bn(j), .C(k), .Y(mai_mai_n99_));
  NO2        m0071(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n100_));
  NAi41      m0072(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n101_));
  AN2        m0073(.A(e), .B(b), .Y(mai_mai_n102_));
  NOi31      m0074(.An(c), .B(h), .C(f), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NO2        m0076(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n105_));
  NOi21      m0077(.An(g), .B(f), .Y(mai_mai_n106_));
  NOi21      m0078(.An(i), .B(h), .Y(mai_mai_n107_));
  NA3        m0079(.A(mai_mai_n107_), .B(mai_mai_n106_), .C(mai_mai_n36_), .Y(mai_mai_n108_));
  INV        m0080(.A(a), .Y(mai_mai_n109_));
  NA2        m0081(.A(mai_mai_n102_), .B(mai_mai_n109_), .Y(mai_mai_n110_));
  INV        m0082(.A(l), .Y(mai_mai_n111_));
  NOi21      m0083(.An(m), .B(n), .Y(mai_mai_n112_));
  AN2        m0084(.A(k), .B(h), .Y(mai_mai_n113_));
  NO2        m0085(.A(mai_mai_n108_), .B(mai_mai_n87_), .Y(mai_mai_n114_));
  INV        m0086(.A(b), .Y(mai_mai_n115_));
  NA2        m0087(.A(l), .B(j), .Y(mai_mai_n116_));
  AN2        m0088(.A(k), .B(i), .Y(mai_mai_n117_));
  NA2        m0089(.A(mai_mai_n117_), .B(mai_mai_n116_), .Y(mai_mai_n118_));
  NA2        m0090(.A(g), .B(e), .Y(mai_mai_n119_));
  NOi32      m0091(.An(c), .Bn(a), .C(d), .Y(mai_mai_n120_));
  NA2        m0092(.A(mai_mai_n120_), .B(mai_mai_n112_), .Y(mai_mai_n121_));
  NO4        m0093(.A(mai_mai_n121_), .B(mai_mai_n119_), .C(mai_mai_n118_), .D(mai_mai_n115_), .Y(mai_mai_n122_));
  NO3        m0094(.A(mai_mai_n122_), .B(mai_mai_n114_), .C(mai_mai_n105_), .Y(mai_mai_n123_));
  OAI210     m0095(.A0(mai_mai_n100_), .A1(mai_mai_n87_), .B0(mai_mai_n123_), .Y(mai_mai_n124_));
  NOi31      m0096(.An(k), .B(m), .C(j), .Y(mai_mai_n125_));
  NOi31      m0097(.An(k), .B(m), .C(i), .Y(mai_mai_n126_));
  NOi32      m0098(.An(f), .Bn(b), .C(e), .Y(mai_mai_n127_));
  NAi21      m0099(.An(g), .B(h), .Y(mai_mai_n128_));
  NAi21      m0100(.An(m), .B(n), .Y(mai_mai_n129_));
  NAi21      m0101(.An(j), .B(k), .Y(mai_mai_n130_));
  NO3        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(mai_mai_n128_), .Y(mai_mai_n131_));
  NAi41      m0103(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n132_));
  NAi31      m0104(.An(j), .B(k), .C(h), .Y(mai_mai_n133_));
  NA2        m0105(.A(mai_mai_n131_), .B(mai_mai_n127_), .Y(mai_mai_n134_));
  NO2        m0106(.A(k), .B(j), .Y(mai_mai_n135_));
  NO2        m0107(.A(mai_mai_n135_), .B(mai_mai_n129_), .Y(mai_mai_n136_));
  AN2        m0108(.A(k), .B(j), .Y(mai_mai_n137_));
  NAi21      m0109(.An(c), .B(b), .Y(mai_mai_n138_));
  NA2        m0110(.A(f), .B(d), .Y(mai_mai_n139_));
  NO4        m0111(.A(mai_mai_n139_), .B(mai_mai_n138_), .C(mai_mai_n137_), .D(mai_mai_n128_), .Y(mai_mai_n140_));
  NA2        m0112(.A(h), .B(c), .Y(mai_mai_n141_));
  NAi31      m0113(.An(f), .B(e), .C(b), .Y(mai_mai_n142_));
  NA2        m0114(.A(mai_mai_n140_), .B(mai_mai_n136_), .Y(mai_mai_n143_));
  NA2        m0115(.A(d), .B(b), .Y(mai_mai_n144_));
  NAi21      m0116(.An(e), .B(f), .Y(mai_mai_n145_));
  NO2        m0117(.A(mai_mai_n145_), .B(mai_mai_n144_), .Y(mai_mai_n146_));
  NA2        m0118(.A(b), .B(a), .Y(mai_mai_n147_));
  NAi21      m0119(.An(e), .B(g), .Y(mai_mai_n148_));
  NAi21      m0120(.An(c), .B(d), .Y(mai_mai_n149_));
  NAi31      m0121(.An(l), .B(k), .C(h), .Y(mai_mai_n150_));
  NA2        m0122(.A(mai_mai_n143_), .B(mai_mai_n134_), .Y(mai_mai_n151_));
  NAi31      m0123(.An(e), .B(f), .C(b), .Y(mai_mai_n152_));
  NOi21      m0124(.An(g), .B(d), .Y(mai_mai_n153_));
  NO2        m0125(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m0126(.An(h), .B(i), .Y(mai_mai_n155_));
  NOi21      m0127(.An(k), .B(m), .Y(mai_mai_n156_));
  NA3        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .C(n), .Y(mai_mai_n157_));
  NOi21      m0129(.An(mai_mai_n154_), .B(mai_mai_n157_), .Y(mai_mai_n158_));
  NOi21      m0130(.An(h), .B(g), .Y(mai_mai_n159_));
  NO2        m0131(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n160_));
  NA2        m0132(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  NOi32      m0133(.An(n), .Bn(k), .C(m), .Y(mai_mai_n162_));
  NA2        m0134(.A(l), .B(i), .Y(mai_mai_n163_));
  INV        m0135(.A(mai_mai_n162_), .Y(mai_mai_n164_));
  NO2        m0136(.A(mai_mai_n164_), .B(mai_mai_n161_), .Y(mai_mai_n165_));
  NAi31      m0137(.An(d), .B(f), .C(c), .Y(mai_mai_n166_));
  NAi31      m0138(.An(e), .B(f), .C(c), .Y(mai_mai_n167_));
  NA2        m0139(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  NA2        m0140(.A(j), .B(h), .Y(mai_mai_n169_));
  OR3        m0141(.A(n), .B(m), .C(k), .Y(mai_mai_n170_));
  NO2        m0142(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  NAi32      m0143(.An(m), .Bn(k), .C(n), .Y(mai_mai_n172_));
  NO2        m0144(.A(mai_mai_n172_), .B(mai_mai_n169_), .Y(mai_mai_n173_));
  AOI220     m0145(.A0(mai_mai_n173_), .A1(mai_mai_n154_), .B0(mai_mai_n171_), .B1(mai_mai_n168_), .Y(mai_mai_n174_));
  NO2        m0146(.A(n), .B(m), .Y(mai_mai_n175_));
  NA2        m0147(.A(mai_mai_n175_), .B(mai_mai_n50_), .Y(mai_mai_n176_));
  NAi21      m0148(.An(f), .B(e), .Y(mai_mai_n177_));
  NA2        m0149(.A(d), .B(c), .Y(mai_mai_n178_));
  NAi31      m0150(.An(m), .B(n), .C(b), .Y(mai_mai_n179_));
  NA2        m0151(.A(k), .B(i), .Y(mai_mai_n180_));
  NAi21      m0152(.An(h), .B(f), .Y(mai_mai_n181_));
  NO2        m0153(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NO2        m0154(.A(mai_mai_n179_), .B(mai_mai_n149_), .Y(mai_mai_n183_));
  NA2        m0155(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  NOi32      m0156(.An(f), .Bn(c), .C(d), .Y(mai_mai_n185_));
  NOi32      m0157(.An(f), .Bn(c), .C(e), .Y(mai_mai_n186_));
  NO2        m0158(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NO3        m0159(.A(n), .B(m), .C(j), .Y(mai_mai_n188_));
  NA2        m0160(.A(mai_mai_n188_), .B(mai_mai_n113_), .Y(mai_mai_n189_));
  AO210      m0161(.A0(mai_mai_n189_), .A1(mai_mai_n176_), .B0(mai_mai_n187_), .Y(mai_mai_n190_));
  NA3        m0162(.A(mai_mai_n190_), .B(mai_mai_n184_), .C(mai_mai_n174_), .Y(mai_mai_n191_));
  OR4        m0163(.A(mai_mai_n191_), .B(mai_mai_n165_), .C(mai_mai_n158_), .D(mai_mai_n151_), .Y(mai_mai_n192_));
  NO4        m0164(.A(mai_mai_n192_), .B(mai_mai_n124_), .C(mai_mai_n84_), .D(mai_mai_n55_), .Y(mai_mai_n193_));
  NA3        m0165(.A(m), .B(mai_mai_n111_), .C(j), .Y(mai_mai_n194_));
  NAi31      m0166(.An(n), .B(h), .C(g), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NOi32      m0168(.An(m), .Bn(k), .C(l), .Y(mai_mai_n197_));
  NA3        m0169(.A(mai_mai_n197_), .B(mai_mai_n88_), .C(g), .Y(mai_mai_n198_));
  NO2        m0170(.A(mai_mai_n198_), .B(n), .Y(mai_mai_n199_));
  NOi21      m0171(.An(k), .B(j), .Y(mai_mai_n200_));
  NA4        m0172(.A(mai_mai_n200_), .B(mai_mai_n112_), .C(i), .D(g), .Y(mai_mai_n201_));
  AN2        m0173(.A(i), .B(g), .Y(mai_mai_n202_));
  INV        m0174(.A(mai_mai_n201_), .Y(mai_mai_n203_));
  NAi41      m0175(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n204_));
  INV        m0176(.A(f), .Y(mai_mai_n205_));
  INV        m0177(.A(g), .Y(mai_mai_n206_));
  NOi31      m0178(.An(i), .B(j), .C(h), .Y(mai_mai_n207_));
  NOi21      m0179(.An(l), .B(m), .Y(mai_mai_n208_));
  NA2        m0180(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n209_));
  NO3        m0181(.A(mai_mai_n209_), .B(mai_mai_n206_), .C(mai_mai_n205_), .Y(mai_mai_n210_));
  NO2        m0182(.A(mai_mai_n201_), .B(mai_mai_n32_), .Y(mai_mai_n211_));
  NOi21      m0183(.An(n), .B(m), .Y(mai_mai_n212_));
  NOi32      m0184(.An(l), .Bn(i), .C(j), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n213_), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  OA220      m0186(.A0(mai_mai_n214_), .A1(mai_mai_n104_), .B0(mai_mai_n80_), .B1(mai_mai_n79_), .Y(mai_mai_n215_));
  NAi21      m0187(.An(j), .B(h), .Y(mai_mai_n216_));
  XN2        m0188(.A(i), .B(h), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  NOi31      m0190(.An(k), .B(n), .C(m), .Y(mai_mai_n219_));
  NOi31      m0191(.An(mai_mai_n219_), .B(mai_mai_n178_), .C(mai_mai_n177_), .Y(mai_mai_n220_));
  NA2        m0192(.A(mai_mai_n220_), .B(mai_mai_n218_), .Y(mai_mai_n221_));
  NAi31      m0193(.An(f), .B(e), .C(c), .Y(mai_mai_n222_));
  NO4        m0194(.A(mai_mai_n222_), .B(mai_mai_n170_), .C(mai_mai_n169_), .D(mai_mai_n59_), .Y(mai_mai_n223_));
  NA4        m0195(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n224_));
  NAi32      m0196(.An(m), .Bn(i), .C(k), .Y(mai_mai_n225_));
  NO3        m0197(.A(mai_mai_n225_), .B(mai_mai_n91_), .C(mai_mai_n224_), .Y(mai_mai_n226_));
  INV        m0198(.A(k), .Y(mai_mai_n227_));
  NO2        m0199(.A(mai_mai_n226_), .B(mai_mai_n223_), .Y(mai_mai_n228_));
  NAi21      m0200(.An(n), .B(a), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n229_), .B(mai_mai_n144_), .Y(mai_mai_n230_));
  NAi41      m0202(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n231_));
  NO3        m0203(.A(mai_mai_n145_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n232_));
  NA2        m0204(.A(mai_mai_n232_), .B(mai_mai_n230_), .Y(mai_mai_n233_));
  AN4        m0205(.A(mai_mai_n233_), .B(mai_mai_n228_), .C(mai_mai_n221_), .D(mai_mai_n215_), .Y(mai_mai_n234_));
  OR2        m0206(.A(h), .B(g), .Y(mai_mai_n235_));
  NO2        m0207(.A(mai_mai_n235_), .B(mai_mai_n101_), .Y(mai_mai_n236_));
  NA2        m0208(.A(mai_mai_n236_), .B(mai_mai_n127_), .Y(mai_mai_n237_));
  NAi41      m0209(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n238_));
  NO2        m0210(.A(mai_mai_n238_), .B(mai_mai_n205_), .Y(mai_mai_n239_));
  NA2        m0211(.A(mai_mai_n156_), .B(mai_mai_n107_), .Y(mai_mai_n240_));
  NAi21      m0212(.An(mai_mai_n240_), .B(mai_mai_n239_), .Y(mai_mai_n241_));
  NO2        m0213(.A(n), .B(a), .Y(mai_mai_n242_));
  NAi31      m0214(.An(mai_mai_n231_), .B(mai_mai_n242_), .C(mai_mai_n102_), .Y(mai_mai_n243_));
  AN2        m0215(.A(mai_mai_n243_), .B(mai_mai_n241_), .Y(mai_mai_n244_));
  NAi21      m0216(.An(h), .B(i), .Y(mai_mai_n245_));
  NA2        m0217(.A(mai_mai_n175_), .B(k), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n246_), .B(mai_mai_n245_), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n247_), .B(mai_mai_n185_), .Y(mai_mai_n248_));
  NA3        m0220(.A(mai_mai_n248_), .B(mai_mai_n244_), .C(mai_mai_n237_), .Y(mai_mai_n249_));
  NOi21      m0221(.An(g), .B(e), .Y(mai_mai_n250_));
  NO2        m0222(.A(mai_mai_n72_), .B(mai_mai_n74_), .Y(mai_mai_n251_));
  NOi32      m0223(.An(l), .Bn(j), .C(i), .Y(mai_mai_n252_));
  AOI210     m0224(.A0(mai_mai_n75_), .A1(mai_mai_n88_), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  NAi21      m0225(.An(f), .B(g), .Y(mai_mai_n254_));
  NO2        m0226(.A(mai_mai_n254_), .B(mai_mai_n65_), .Y(mai_mai_n255_));
  NO2        m0227(.A(mai_mai_n69_), .B(mai_mai_n116_), .Y(mai_mai_n256_));
  NA2        m0228(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n257_));
  INV        m0229(.A(mai_mai_n257_), .Y(mai_mai_n258_));
  NO3        m0230(.A(mai_mai_n130_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n259_));
  NOi41      m0231(.An(mai_mai_n234_), .B(mai_mai_n258_), .C(mai_mai_n249_), .D(mai_mai_n211_), .Y(mai_mai_n260_));
  NO4        m0232(.A(mai_mai_n196_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n261_), .B(mai_mai_n110_), .Y(mai_mai_n262_));
  NA3        m0234(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n263_));
  NAi21      m0235(.An(h), .B(g), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n240_), .B(mai_mai_n254_), .Y(mai_mai_n265_));
  NAi31      m0237(.An(g), .B(k), .C(h), .Y(mai_mai_n266_));
  NO3        m0238(.A(mai_mai_n129_), .B(mai_mai_n266_), .C(l), .Y(mai_mai_n267_));
  NAi31      m0239(.An(e), .B(d), .C(a), .Y(mai_mai_n268_));
  NA2        m0240(.A(mai_mai_n267_), .B(mai_mai_n127_), .Y(mai_mai_n269_));
  INV        m0241(.A(mai_mai_n269_), .Y(mai_mai_n270_));
  NA4        m0242(.A(mai_mai_n156_), .B(mai_mai_n81_), .C(mai_mai_n77_), .D(mai_mai_n116_), .Y(mai_mai_n271_));
  NA3        m0243(.A(mai_mai_n156_), .B(mai_mai_n155_), .C(mai_mai_n85_), .Y(mai_mai_n272_));
  NO2        m0244(.A(mai_mai_n272_), .B(mai_mai_n187_), .Y(mai_mai_n273_));
  NOi21      m0245(.An(mai_mai_n271_), .B(mai_mai_n273_), .Y(mai_mai_n274_));
  NA3        m0246(.A(e), .B(c), .C(b), .Y(mai_mai_n275_));
  NAi21      m0247(.An(l), .B(k), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n276_), .B(mai_mai_n49_), .Y(mai_mai_n277_));
  NOi21      m0249(.An(l), .B(j), .Y(mai_mai_n278_));
  NA2        m0250(.A(mai_mai_n159_), .B(mai_mai_n278_), .Y(mai_mai_n279_));
  NA3        m0251(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(g), .Y(mai_mai_n280_));
  OR3        m0252(.A(mai_mai_n72_), .B(mai_mai_n74_), .C(e), .Y(mai_mai_n281_));
  AOI210     m0253(.A0(mai_mai_n280_), .A1(mai_mai_n279_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  INV        m0254(.A(mai_mai_n282_), .Y(mai_mai_n283_));
  NAi32      m0255(.An(j), .Bn(h), .C(i), .Y(mai_mai_n284_));
  NAi21      m0256(.An(m), .B(l), .Y(mai_mai_n285_));
  NO3        m0257(.A(mai_mai_n285_), .B(mai_mai_n284_), .C(mai_mai_n85_), .Y(mai_mai_n286_));
  NA2        m0258(.A(h), .B(g), .Y(mai_mai_n287_));
  NA2        m0259(.A(mai_mai_n286_), .B(mai_mai_n160_), .Y(mai_mai_n288_));
  NA3        m0260(.A(mai_mai_n288_), .B(mai_mai_n283_), .C(mai_mai_n274_), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n142_), .B(d), .Y(mai_mai_n290_));
  NA2        m0262(.A(mai_mai_n290_), .B(mai_mai_n53_), .Y(mai_mai_n291_));
  NO2        m0263(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n292_));
  NAi32      m0264(.An(n), .Bn(m), .C(l), .Y(mai_mai_n293_));
  NO2        m0265(.A(mai_mai_n293_), .B(mai_mai_n284_), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n121_), .B(mai_mai_n115_), .Y(mai_mai_n295_));
  NAi31      m0267(.An(k), .B(l), .C(j), .Y(mai_mai_n296_));
  OAI210     m0268(.A0(mai_mai_n276_), .A1(j), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  NOi21      m0269(.An(mai_mai_n297_), .B(mai_mai_n119_), .Y(mai_mai_n298_));
  NA2        m0270(.A(mai_mai_n298_), .B(mai_mai_n295_), .Y(mai_mai_n299_));
  NA2        m0271(.A(mai_mai_n299_), .B(mai_mai_n291_), .Y(mai_mai_n300_));
  NO4        m0272(.A(mai_mai_n300_), .B(mai_mai_n289_), .C(mai_mai_n270_), .D(mai_mai_n262_), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n247_), .B(mai_mai_n186_), .Y(mai_mai_n302_));
  NAi21      m0274(.An(m), .B(k), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n217_), .B(mai_mai_n303_), .Y(mai_mai_n304_));
  NAi41      m0276(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n305_), .B(mai_mai_n148_), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n306_), .B(mai_mai_n304_), .Y(mai_mai_n307_));
  NAi31      m0279(.An(i), .B(l), .C(h), .Y(mai_mai_n308_));
  NO4        m0280(.A(mai_mai_n308_), .B(mai_mai_n148_), .C(mai_mai_n72_), .D(mai_mai_n74_), .Y(mai_mai_n309_));
  NA2        m0281(.A(e), .B(c), .Y(mai_mai_n310_));
  NO3        m0282(.A(mai_mai_n310_), .B(n), .C(d), .Y(mai_mai_n311_));
  NOi21      m0283(.An(f), .B(h), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n312_), .B(mai_mai_n117_), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n313_), .B(mai_mai_n206_), .Y(mai_mai_n314_));
  NAi31      m0286(.An(d), .B(e), .C(b), .Y(mai_mai_n315_));
  NO2        m0287(.A(mai_mai_n129_), .B(mai_mai_n315_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n316_), .B(mai_mai_n314_), .Y(mai_mai_n317_));
  NAi41      m0289(.An(mai_mai_n309_), .B(mai_mai_n317_), .C(mai_mai_n307_), .D(mai_mai_n302_), .Y(mai_mai_n318_));
  NA2        m0290(.A(mai_mai_n242_), .B(mai_mai_n102_), .Y(mai_mai_n319_));
  OR2        m0291(.A(mai_mai_n319_), .B(mai_mai_n198_), .Y(mai_mai_n320_));
  NOi31      m0292(.An(l), .B(n), .C(m), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n321_), .B(mai_mai_n207_), .Y(mai_mai_n322_));
  NO2        m0294(.A(mai_mai_n322_), .B(mai_mai_n187_), .Y(mai_mai_n323_));
  NAi21      m0295(.An(mai_mai_n323_), .B(mai_mai_n320_), .Y(mai_mai_n324_));
  NAi32      m0296(.An(m), .Bn(j), .C(k), .Y(mai_mai_n325_));
  NAi41      m0297(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n204_), .B(mai_mai_n326_), .Y(mai_mai_n327_));
  NOi31      m0299(.An(j), .B(m), .C(k), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n125_), .B(mai_mai_n328_), .Y(mai_mai_n329_));
  AN3        m0301(.A(h), .B(g), .C(f), .Y(mai_mai_n330_));
  NAi31      m0302(.An(mai_mai_n329_), .B(mai_mai_n330_), .C(mai_mai_n327_), .Y(mai_mai_n331_));
  NOi32      m0303(.An(m), .Bn(j), .C(l), .Y(mai_mai_n332_));
  NO2        m0304(.A(mai_mai_n332_), .B(mai_mai_n98_), .Y(mai_mai_n333_));
  NAi32      m0305(.An(mai_mai_n333_), .Bn(mai_mai_n195_), .C(mai_mai_n290_), .Y(mai_mai_n334_));
  NO2        m0306(.A(mai_mai_n285_), .B(mai_mai_n284_), .Y(mai_mai_n335_));
  NO2        m0307(.A(mai_mai_n209_), .B(g), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n152_), .B(mai_mai_n85_), .Y(mai_mai_n337_));
  AOI220     m0309(.A0(mai_mai_n337_), .A1(mai_mai_n336_), .B0(mai_mai_n239_), .B1(mai_mai_n335_), .Y(mai_mai_n338_));
  NA3        m0310(.A(mai_mai_n338_), .B(mai_mai_n334_), .C(mai_mai_n331_), .Y(mai_mai_n339_));
  NA3        m0311(.A(h), .B(g), .C(f), .Y(mai_mai_n340_));
  NO2        m0312(.A(mai_mai_n340_), .B(mai_mai_n76_), .Y(mai_mai_n341_));
  NA2        m0313(.A(mai_mai_n326_), .B(mai_mai_n204_), .Y(mai_mai_n342_));
  NA2        m0314(.A(mai_mai_n159_), .B(e), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n343_), .B(mai_mai_n41_), .Y(mai_mai_n344_));
  AOI220     m0316(.A0(mai_mai_n344_), .A1(mai_mai_n295_), .B0(mai_mai_n342_), .B1(mai_mai_n341_), .Y(mai_mai_n345_));
  NOi32      m0317(.An(e), .Bn(b), .C(a), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n201_), .B(mai_mai_n35_), .Y(mai_mai_n347_));
  NA2        m0319(.A(mai_mai_n347_), .B(mai_mai_n346_), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n315_), .B(n), .Y(mai_mai_n349_));
  NA2        m0321(.A(mai_mai_n202_), .B(k), .Y(mai_mai_n350_));
  NA3        m0322(.A(m), .B(mai_mai_n111_), .C(mai_mai_n205_), .Y(mai_mai_n351_));
  NA4        m0323(.A(mai_mai_n197_), .B(mai_mai_n88_), .C(g), .D(mai_mai_n205_), .Y(mai_mai_n352_));
  INV        m0324(.A(mai_mai_n352_), .Y(mai_mai_n353_));
  NAi41      m0325(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n51_), .B(mai_mai_n112_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n353_), .B(mai_mai_n349_), .Y(mai_mai_n356_));
  NA3        m0328(.A(mai_mai_n356_), .B(mai_mai_n348_), .C(mai_mai_n345_), .Y(mai_mai_n357_));
  NO4        m0329(.A(mai_mai_n357_), .B(mai_mai_n339_), .C(mai_mai_n324_), .D(mai_mai_n318_), .Y(mai_mai_n358_));
  NA4        m0330(.A(mai_mai_n358_), .B(mai_mai_n301_), .C(mai_mai_n260_), .D(mai_mai_n193_), .Y(mai10));
  NA3        m0331(.A(m), .B(k), .C(i), .Y(mai_mai_n360_));
  NO3        m0332(.A(mai_mai_n360_), .B(j), .C(mai_mai_n206_), .Y(mai_mai_n361_));
  NOi21      m0333(.An(e), .B(f), .Y(mai_mai_n362_));
  NO4        m0334(.A(mai_mai_n149_), .B(mai_mai_n362_), .C(n), .D(mai_mai_n109_), .Y(mai_mai_n363_));
  NAi31      m0335(.An(b), .B(f), .C(c), .Y(mai_mai_n364_));
  INV        m0336(.A(mai_mai_n364_), .Y(mai_mai_n365_));
  NOi32      m0337(.An(k), .Bn(h), .C(j), .Y(mai_mai_n366_));
  NA2        m0338(.A(mai_mai_n366_), .B(mai_mai_n212_), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n157_), .B(mai_mai_n367_), .Y(mai_mai_n368_));
  AOI220     m0340(.A0(mai_mai_n368_), .A1(mai_mai_n365_), .B0(mai_mai_n363_), .B1(mai_mai_n361_), .Y(mai_mai_n369_));
  AN2        m0341(.A(j), .B(h), .Y(mai_mai_n370_));
  NO3        m0342(.A(n), .B(m), .C(k), .Y(mai_mai_n371_));
  NA2        m0343(.A(mai_mai_n371_), .B(mai_mai_n370_), .Y(mai_mai_n372_));
  NO3        m0344(.A(mai_mai_n372_), .B(mai_mai_n149_), .C(mai_mai_n205_), .Y(mai_mai_n373_));
  OR2        m0345(.A(m), .B(k), .Y(mai_mai_n374_));
  NO2        m0346(.A(mai_mai_n169_), .B(mai_mai_n374_), .Y(mai_mai_n375_));
  NA4        m0347(.A(n), .B(f), .C(c), .D(mai_mai_n115_), .Y(mai_mai_n376_));
  NOi21      m0348(.An(mai_mai_n375_), .B(mai_mai_n376_), .Y(mai_mai_n377_));
  NOi32      m0349(.An(d), .Bn(a), .C(c), .Y(mai_mai_n378_));
  NA2        m0350(.A(mai_mai_n378_), .B(mai_mai_n177_), .Y(mai_mai_n379_));
  NAi21      m0351(.An(i), .B(g), .Y(mai_mai_n380_));
  NAi31      m0352(.An(k), .B(m), .C(j), .Y(mai_mai_n381_));
  NO3        m0353(.A(mai_mai_n381_), .B(mai_mai_n380_), .C(n), .Y(mai_mai_n382_));
  NOi21      m0354(.An(mai_mai_n382_), .B(mai_mai_n379_), .Y(mai_mai_n383_));
  NO3        m0355(.A(mai_mai_n383_), .B(mai_mai_n377_), .C(mai_mai_n373_), .Y(mai_mai_n384_));
  NO2        m0356(.A(mai_mai_n376_), .B(mai_mai_n285_), .Y(mai_mai_n385_));
  NOi32      m0357(.An(f), .Bn(d), .C(c), .Y(mai_mai_n386_));
  AOI220     m0358(.A0(mai_mai_n386_), .A1(mai_mai_n294_), .B0(mai_mai_n385_), .B1(mai_mai_n207_), .Y(mai_mai_n387_));
  NA3        m0359(.A(mai_mai_n387_), .B(mai_mai_n384_), .C(mai_mai_n369_), .Y(mai_mai_n388_));
  NO2        m0360(.A(mai_mai_n59_), .B(mai_mai_n115_), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n242_), .B(mai_mai_n389_), .Y(mai_mai_n390_));
  INV        m0362(.A(e), .Y(mai_mai_n391_));
  NA2        m0363(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n392_));
  OAI220     m0364(.A0(mai_mai_n392_), .A1(mai_mai_n194_), .B0(mai_mai_n198_), .B1(mai_mai_n391_), .Y(mai_mai_n393_));
  AN2        m0365(.A(g), .B(e), .Y(mai_mai_n394_));
  NO2        m0366(.A(mai_mai_n90_), .B(mai_mai_n391_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n395_), .B(mai_mai_n393_), .Y(mai_mai_n396_));
  NOi32      m0368(.An(h), .Bn(e), .C(g), .Y(mai_mai_n397_));
  NA3        m0369(.A(mai_mai_n397_), .B(mai_mai_n278_), .C(m), .Y(mai_mai_n398_));
  NOi21      m0370(.An(g), .B(h), .Y(mai_mai_n399_));
  AN3        m0371(.A(m), .B(l), .C(i), .Y(mai_mai_n400_));
  AN3        m0372(.A(h), .B(g), .C(e), .Y(mai_mai_n401_));
  NA2        m0373(.A(mai_mai_n401_), .B(mai_mai_n98_), .Y(mai_mai_n402_));
  AN2        m0374(.A(mai_mai_n402_), .B(mai_mai_n398_), .Y(mai_mai_n403_));
  AOI210     m0375(.A0(mai_mai_n403_), .A1(mai_mai_n396_), .B0(mai_mai_n390_), .Y(mai_mai_n404_));
  NA3        m0376(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n405_));
  NO2        m0377(.A(mai_mai_n405_), .B(mai_mai_n390_), .Y(mai_mai_n406_));
  NA3        m0378(.A(mai_mai_n378_), .B(mai_mai_n177_), .C(mai_mai_n85_), .Y(mai_mai_n407_));
  NAi31      m0379(.An(b), .B(c), .C(a), .Y(mai_mai_n408_));
  NO2        m0380(.A(mai_mai_n408_), .B(n), .Y(mai_mai_n409_));
  NA2        m0381(.A(mai_mai_n51_), .B(m), .Y(mai_mai_n410_));
  NO2        m0382(.A(mai_mai_n410_), .B(mai_mai_n145_), .Y(mai_mai_n411_));
  NA2        m0383(.A(mai_mai_n411_), .B(mai_mai_n409_), .Y(mai_mai_n412_));
  INV        m0384(.A(mai_mai_n412_), .Y(mai_mai_n413_));
  NO4        m0385(.A(mai_mai_n413_), .B(mai_mai_n406_), .C(mai_mai_n404_), .D(mai_mai_n388_), .Y(mai_mai_n414_));
  NA2        m0386(.A(i), .B(g), .Y(mai_mai_n415_));
  NO3        m0387(.A(mai_mai_n268_), .B(mai_mai_n415_), .C(c), .Y(mai_mai_n416_));
  NOi21      m0388(.An(a), .B(n), .Y(mai_mai_n417_));
  NOi21      m0389(.An(d), .B(c), .Y(mai_mai_n418_));
  NA2        m0390(.A(mai_mai_n418_), .B(mai_mai_n417_), .Y(mai_mai_n419_));
  NA3        m0391(.A(i), .B(g), .C(f), .Y(mai_mai_n420_));
  OR2        m0392(.A(mai_mai_n420_), .B(mai_mai_n71_), .Y(mai_mai_n421_));
  NA3        m0393(.A(mai_mai_n400_), .B(mai_mai_n399_), .C(mai_mai_n177_), .Y(mai_mai_n422_));
  AOI210     m0394(.A0(mai_mai_n422_), .A1(mai_mai_n421_), .B0(mai_mai_n419_), .Y(mai_mai_n423_));
  AOI210     m0395(.A0(mai_mai_n416_), .A1(mai_mai_n277_), .B0(mai_mai_n423_), .Y(mai_mai_n424_));
  OR2        m0396(.A(n), .B(m), .Y(mai_mai_n425_));
  NO2        m0397(.A(mai_mai_n425_), .B(mai_mai_n150_), .Y(mai_mai_n426_));
  NO2        m0398(.A(mai_mai_n178_), .B(mai_mai_n145_), .Y(mai_mai_n427_));
  OAI210     m0399(.A0(mai_mai_n426_), .A1(mai_mai_n171_), .B0(mai_mai_n427_), .Y(mai_mai_n428_));
  INV        m0400(.A(mai_mai_n355_), .Y(mai_mai_n429_));
  NA3        m0401(.A(mai_mai_n429_), .B(mai_mai_n346_), .C(d), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n408_), .B(mai_mai_n49_), .Y(mai_mai_n431_));
  NO3        m0403(.A(mai_mai_n66_), .B(mai_mai_n111_), .C(e), .Y(mai_mai_n432_));
  NAi21      m0404(.An(k), .B(j), .Y(mai_mai_n433_));
  NA2        m0405(.A(mai_mai_n245_), .B(mai_mai_n433_), .Y(mai_mai_n434_));
  NA3        m0406(.A(mai_mai_n434_), .B(mai_mai_n432_), .C(mai_mai_n431_), .Y(mai_mai_n435_));
  NAi21      m0407(.An(e), .B(d), .Y(mai_mai_n436_));
  INV        m0408(.A(mai_mai_n436_), .Y(mai_mai_n437_));
  NO2        m0409(.A(mai_mai_n246_), .B(mai_mai_n205_), .Y(mai_mai_n438_));
  NA3        m0410(.A(mai_mai_n438_), .B(mai_mai_n437_), .C(mai_mai_n218_), .Y(mai_mai_n439_));
  NA4        m0411(.A(mai_mai_n439_), .B(mai_mai_n435_), .C(mai_mai_n430_), .D(mai_mai_n428_), .Y(mai_mai_n440_));
  NO2        m0412(.A(mai_mai_n322_), .B(mai_mai_n205_), .Y(mai_mai_n441_));
  NA2        m0413(.A(mai_mai_n441_), .B(mai_mai_n437_), .Y(mai_mai_n442_));
  NOi31      m0414(.An(n), .B(m), .C(k), .Y(mai_mai_n443_));
  AOI220     m0415(.A0(mai_mai_n443_), .A1(mai_mai_n370_), .B0(mai_mai_n212_), .B1(mai_mai_n50_), .Y(mai_mai_n444_));
  NAi31      m0416(.An(g), .B(f), .C(c), .Y(mai_mai_n445_));
  OR3        m0417(.A(mai_mai_n445_), .B(mai_mai_n444_), .C(e), .Y(mai_mai_n446_));
  NA2        m0418(.A(mai_mai_n446_), .B(mai_mai_n442_), .Y(mai_mai_n447_));
  NOi41      m0419(.An(mai_mai_n424_), .B(mai_mai_n447_), .C(mai_mai_n440_), .D(mai_mai_n258_), .Y(mai_mai_n448_));
  NOi32      m0420(.An(c), .Bn(a), .C(b), .Y(mai_mai_n449_));
  NA2        m0421(.A(mai_mai_n449_), .B(mai_mai_n112_), .Y(mai_mai_n450_));
  INV        m0422(.A(mai_mai_n266_), .Y(mai_mai_n451_));
  AN2        m0423(.A(e), .B(d), .Y(mai_mai_n452_));
  NA2        m0424(.A(mai_mai_n452_), .B(mai_mai_n451_), .Y(mai_mai_n453_));
  INV        m0425(.A(mai_mai_n145_), .Y(mai_mai_n454_));
  NO2        m0426(.A(mai_mai_n128_), .B(mai_mai_n41_), .Y(mai_mai_n455_));
  NO2        m0427(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n456_));
  NA3        m0428(.A(mai_mai_n308_), .B(mai_mai_n253_), .C(mai_mai_n118_), .Y(mai_mai_n457_));
  AOI220     m0429(.A0(mai_mai_n457_), .A1(mai_mai_n456_), .B0(mai_mai_n455_), .B1(mai_mai_n454_), .Y(mai_mai_n458_));
  AOI210     m0430(.A0(mai_mai_n458_), .A1(mai_mai_n453_), .B0(mai_mai_n450_), .Y(mai_mai_n459_));
  NO2        m0431(.A(mai_mai_n203_), .B(mai_mai_n199_), .Y(mai_mai_n460_));
  NOi21      m0432(.An(a), .B(b), .Y(mai_mai_n461_));
  NA3        m0433(.A(e), .B(d), .C(c), .Y(mai_mai_n462_));
  NAi21      m0434(.An(mai_mai_n462_), .B(mai_mai_n461_), .Y(mai_mai_n463_));
  NO2        m0435(.A(mai_mai_n407_), .B(mai_mai_n198_), .Y(mai_mai_n464_));
  NOi21      m0436(.An(mai_mai_n463_), .B(mai_mai_n464_), .Y(mai_mai_n465_));
  AOI210     m0437(.A0(mai_mai_n261_), .A1(mai_mai_n460_), .B0(mai_mai_n465_), .Y(mai_mai_n466_));
  NO4        m0438(.A(mai_mai_n181_), .B(mai_mai_n101_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n467_));
  OR2        m0439(.A(k), .B(j), .Y(mai_mai_n468_));
  NA2        m0440(.A(l), .B(k), .Y(mai_mai_n469_));
  NA3        m0441(.A(mai_mai_n469_), .B(mai_mai_n468_), .C(mai_mai_n212_), .Y(mai_mai_n470_));
  AOI210     m0442(.A0(mai_mai_n225_), .A1(mai_mai_n325_), .B0(mai_mai_n85_), .Y(mai_mai_n471_));
  NOi21      m0443(.An(mai_mai_n470_), .B(mai_mai_n471_), .Y(mai_mai_n472_));
  OR3        m0444(.A(mai_mai_n472_), .B(mai_mai_n141_), .C(mai_mai_n132_), .Y(mai_mai_n473_));
  INV        m0445(.A(mai_mai_n271_), .Y(mai_mai_n474_));
  NA2        m0446(.A(mai_mai_n378_), .B(mai_mai_n112_), .Y(mai_mai_n475_));
  NO4        m0447(.A(mai_mai_n475_), .B(mai_mai_n95_), .C(mai_mai_n111_), .D(e), .Y(mai_mai_n476_));
  NO3        m0448(.A(mai_mai_n407_), .B(mai_mai_n92_), .C(mai_mai_n128_), .Y(mai_mai_n477_));
  NO4        m0449(.A(mai_mai_n477_), .B(mai_mai_n476_), .C(mai_mai_n474_), .D(mai_mai_n309_), .Y(mai_mai_n478_));
  NA2        m0450(.A(mai_mai_n478_), .B(mai_mai_n473_), .Y(mai_mai_n479_));
  NO4        m0451(.A(mai_mai_n479_), .B(mai_mai_n467_), .C(mai_mai_n466_), .D(mai_mai_n459_), .Y(mai_mai_n480_));
  NA2        m0452(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n481_));
  NOi21      m0453(.An(d), .B(e), .Y(mai_mai_n482_));
  NO2        m0454(.A(mai_mai_n181_), .B(mai_mai_n56_), .Y(mai_mai_n483_));
  NAi31      m0455(.An(j), .B(l), .C(i), .Y(mai_mai_n484_));
  OAI210     m0456(.A0(mai_mai_n484_), .A1(mai_mai_n129_), .B0(mai_mai_n101_), .Y(mai_mai_n485_));
  NA3        m0457(.A(mai_mai_n485_), .B(mai_mai_n483_), .C(mai_mai_n482_), .Y(mai_mai_n486_));
  NO3        m0458(.A(mai_mai_n379_), .B(mai_mai_n333_), .C(mai_mai_n195_), .Y(mai_mai_n487_));
  NO2        m0459(.A(mai_mai_n379_), .B(mai_mai_n355_), .Y(mai_mai_n488_));
  NO3        m0460(.A(mai_mai_n488_), .B(mai_mai_n487_), .C(mai_mai_n292_), .Y(mai_mai_n489_));
  NA4        m0461(.A(mai_mai_n489_), .B(mai_mai_n486_), .C(mai_mai_n481_), .D(mai_mai_n234_), .Y(mai_mai_n490_));
  OAI210     m0462(.A0(mai_mai_n126_), .A1(mai_mai_n125_), .B0(n), .Y(mai_mai_n491_));
  NO2        m0463(.A(mai_mai_n491_), .B(mai_mai_n128_), .Y(mai_mai_n492_));
  BUFFER     m0464(.A(mai_mai_n236_), .Y(mai_mai_n493_));
  OA210      m0465(.A0(mai_mai_n493_), .A1(mai_mai_n492_), .B0(mai_mai_n186_), .Y(mai_mai_n494_));
  XO2        m0466(.A(i), .B(h), .Y(mai_mai_n495_));
  NA3        m0467(.A(mai_mai_n495_), .B(mai_mai_n156_), .C(n), .Y(mai_mai_n496_));
  NAi41      m0468(.An(mai_mai_n286_), .B(mai_mai_n496_), .C(mai_mai_n444_), .D(mai_mai_n367_), .Y(mai_mai_n497_));
  NAi31      m0469(.An(c), .B(f), .C(d), .Y(mai_mai_n498_));
  AOI210     m0470(.A0(mai_mai_n272_), .A1(mai_mai_n189_), .B0(mai_mai_n498_), .Y(mai_mai_n499_));
  NOi21      m0471(.An(mai_mai_n83_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NA3        m0472(.A(mai_mai_n363_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n501_));
  NA2        m0473(.A(mai_mai_n219_), .B(mai_mai_n107_), .Y(mai_mai_n502_));
  AOI210     m0474(.A0(mai_mai_n502_), .A1(mai_mai_n176_), .B0(mai_mai_n498_), .Y(mai_mai_n503_));
  NOi21      m0475(.An(mai_mai_n501_), .B(mai_mai_n503_), .Y(mai_mai_n504_));
  NA3        m0476(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n505_));
  NO2        m0477(.A(mai_mai_n505_), .B(mai_mai_n419_), .Y(mai_mai_n506_));
  NO2        m0478(.A(mai_mai_n506_), .B(mai_mai_n282_), .Y(mai_mai_n507_));
  NA3        m0479(.A(mai_mai_n507_), .B(mai_mai_n504_), .C(mai_mai_n500_), .Y(mai_mai_n508_));
  NO3        m0480(.A(mai_mai_n508_), .B(mai_mai_n494_), .C(mai_mai_n490_), .Y(mai_mai_n509_));
  NA4        m0481(.A(mai_mai_n509_), .B(mai_mai_n480_), .C(mai_mai_n448_), .D(mai_mai_n414_), .Y(mai11));
  NO2        m0482(.A(mai_mai_n72_), .B(f), .Y(mai_mai_n511_));
  NA2        m0483(.A(j), .B(g), .Y(mai_mai_n512_));
  NAi31      m0484(.An(i), .B(m), .C(l), .Y(mai_mai_n513_));
  NA3        m0485(.A(m), .B(k), .C(j), .Y(mai_mai_n514_));
  NOi32      m0486(.An(e), .Bn(b), .C(f), .Y(mai_mai_n515_));
  NA2        m0487(.A(mai_mai_n252_), .B(mai_mai_n112_), .Y(mai_mai_n516_));
  NA2        m0488(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n517_));
  NAi31      m0489(.An(d), .B(e), .C(a), .Y(mai_mai_n518_));
  NO2        m0490(.A(mai_mai_n518_), .B(n), .Y(mai_mai_n519_));
  NAi41      m0491(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n520_));
  AN2        m0492(.A(mai_mai_n520_), .B(mai_mai_n354_), .Y(mai_mai_n521_));
  AOI210     m0493(.A0(mai_mai_n521_), .A1(mai_mai_n379_), .B0(mai_mai_n264_), .Y(mai_mai_n522_));
  NA2        m0494(.A(j), .B(i), .Y(mai_mai_n523_));
  NAi31      m0495(.An(n), .B(m), .C(k), .Y(mai_mai_n524_));
  NO3        m0496(.A(mai_mai_n524_), .B(mai_mai_n523_), .C(mai_mai_n111_), .Y(mai_mai_n525_));
  NO4        m0497(.A(n), .B(d), .C(mai_mai_n115_), .D(a), .Y(mai_mai_n526_));
  OR2        m0498(.A(n), .B(c), .Y(mai_mai_n527_));
  NO2        m0499(.A(mai_mai_n527_), .B(mai_mai_n147_), .Y(mai_mai_n528_));
  NOi32      m0500(.An(g), .Bn(f), .C(i), .Y(mai_mai_n529_));
  NO2        m0501(.A(mai_mai_n266_), .B(mai_mai_n49_), .Y(mai_mai_n530_));
  NA2        m0502(.A(mai_mai_n525_), .B(mai_mai_n522_), .Y(mai_mai_n531_));
  NA2        m0503(.A(mai_mai_n137_), .B(mai_mai_n34_), .Y(mai_mai_n532_));
  OAI220     m0504(.A0(mai_mai_n532_), .A1(m), .B0(mai_mai_n517_), .B1(mai_mai_n225_), .Y(mai_mai_n533_));
  NOi41      m0505(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n534_));
  NAi32      m0506(.An(e), .Bn(b), .C(c), .Y(mai_mai_n535_));
  OR2        m0507(.A(mai_mai_n535_), .B(mai_mai_n85_), .Y(mai_mai_n536_));
  AN2        m0508(.A(mai_mai_n326_), .B(mai_mai_n305_), .Y(mai_mai_n537_));
  NA2        m0509(.A(mai_mai_n537_), .B(mai_mai_n536_), .Y(mai_mai_n538_));
  AN2        m0510(.A(mai_mai_n538_), .B(mai_mai_n533_), .Y(mai_mai_n539_));
  OAI220     m0511(.A0(mai_mai_n381_), .A1(mai_mai_n380_), .B0(mai_mai_n513_), .B1(mai_mai_n512_), .Y(mai_mai_n540_));
  NAi31      m0512(.An(d), .B(c), .C(a), .Y(mai_mai_n541_));
  NO2        m0513(.A(mai_mai_n541_), .B(n), .Y(mai_mai_n542_));
  NA3        m0514(.A(mai_mai_n542_), .B(mai_mai_n540_), .C(e), .Y(mai_mai_n543_));
  NO3        m0515(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n206_), .Y(mai_mai_n544_));
  NO2        m0516(.A(mai_mai_n222_), .B(mai_mai_n109_), .Y(mai_mai_n545_));
  OAI210     m0517(.A0(mai_mai_n544_), .A1(mai_mai_n382_), .B0(mai_mai_n545_), .Y(mai_mai_n546_));
  NA2        m0518(.A(mai_mai_n546_), .B(mai_mai_n543_), .Y(mai_mai_n547_));
  NO2        m0519(.A(mai_mai_n268_), .B(n), .Y(mai_mai_n548_));
  NAi32      m0520(.An(d), .Bn(a), .C(b), .Y(mai_mai_n549_));
  NA2        m0521(.A(h), .B(f), .Y(mai_mai_n550_));
  NO2        m0522(.A(mai_mai_n550_), .B(mai_mai_n95_), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n144_), .B(c), .Y(mai_mai_n552_));
  NA3        m0524(.A(f), .B(d), .C(b), .Y(mai_mai_n553_));
  NO4        m0525(.A(mai_mai_n553_), .B(mai_mai_n172_), .C(mai_mai_n169_), .D(g), .Y(mai_mai_n554_));
  NO3        m0526(.A(mai_mai_n554_), .B(mai_mai_n547_), .C(mai_mai_n539_), .Y(mai_mai_n555_));
  AN2        m0527(.A(mai_mai_n555_), .B(mai_mai_n531_), .Y(mai_mai_n556_));
  INV        m0528(.A(k), .Y(mai_mai_n557_));
  NA3        m0529(.A(l), .B(mai_mai_n557_), .C(i), .Y(mai_mai_n558_));
  INV        m0530(.A(mai_mai_n558_), .Y(mai_mai_n559_));
  NA3        m0531(.A(mai_mai_n378_), .B(mai_mai_n399_), .C(mai_mai_n112_), .Y(mai_mai_n560_));
  NAi32      m0532(.An(h), .Bn(f), .C(g), .Y(mai_mai_n561_));
  NAi41      m0533(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n562_));
  OAI210     m0534(.A0(mai_mai_n518_), .A1(n), .B0(mai_mai_n562_), .Y(mai_mai_n563_));
  NA2        m0535(.A(mai_mai_n563_), .B(m), .Y(mai_mai_n564_));
  NAi31      m0536(.An(h), .B(g), .C(f), .Y(mai_mai_n565_));
  NAi31      m0537(.An(f), .B(h), .C(g), .Y(mai_mai_n566_));
  NO4        m0538(.A(mai_mai_n296_), .B(mai_mai_n566_), .C(mai_mai_n72_), .D(mai_mai_n74_), .Y(mai_mai_n567_));
  NOi32      m0539(.An(d), .Bn(a), .C(e), .Y(mai_mai_n568_));
  NO2        m0540(.A(n), .B(c), .Y(mai_mai_n569_));
  NOi32      m0541(.An(e), .Bn(a), .C(d), .Y(mai_mai_n570_));
  AOI210     m0542(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n570_), .Y(mai_mai_n571_));
  OAI210     m0543(.A0(mai_mai_n241_), .A1(mai_mai_n88_), .B0(mai_mai_n1430_), .Y(mai_mai_n572_));
  AOI210     m0544(.A0(mai_mai_n1433_), .A1(mai_mai_n559_), .B0(mai_mai_n572_), .Y(mai_mai_n573_));
  NO3        m0545(.A(mai_mai_n303_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n574_));
  NA3        m0546(.A(mai_mai_n498_), .B(mai_mai_n167_), .C(mai_mai_n166_), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n445_), .B(mai_mai_n222_), .Y(mai_mai_n576_));
  OR2        m0548(.A(mai_mai_n576_), .B(mai_mai_n575_), .Y(mai_mai_n577_));
  NA2        m0549(.A(mai_mai_n75_), .B(mai_mai_n112_), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n578_), .B(mai_mai_n45_), .Y(mai_mai_n579_));
  AOI220     m0551(.A0(mai_mai_n579_), .A1(mai_mai_n522_), .B0(mai_mai_n577_), .B1(mai_mai_n574_), .Y(mai_mai_n580_));
  NO2        m0552(.A(mai_mai_n580_), .B(mai_mai_n88_), .Y(mai_mai_n581_));
  NA3        m0553(.A(mai_mai_n534_), .B(mai_mai_n328_), .C(mai_mai_n46_), .Y(mai_mai_n582_));
  NOi32      m0554(.An(e), .Bn(c), .C(f), .Y(mai_mai_n583_));
  NOi21      m0555(.An(f), .B(g), .Y(mai_mai_n584_));
  NO2        m0556(.A(mai_mai_n584_), .B(mai_mai_n204_), .Y(mai_mai_n585_));
  AOI220     m0557(.A0(mai_mai_n585_), .A1(mai_mai_n375_), .B0(mai_mai_n583_), .B1(mai_mai_n171_), .Y(mai_mai_n586_));
  NA3        m0558(.A(mai_mai_n586_), .B(mai_mai_n582_), .C(mai_mai_n174_), .Y(mai_mai_n587_));
  AOI210     m0559(.A0(mai_mai_n521_), .A1(mai_mai_n379_), .B0(mai_mai_n287_), .Y(mai_mai_n588_));
  NA2        m0560(.A(mai_mai_n588_), .B(mai_mai_n256_), .Y(mai_mai_n589_));
  NO2        m0561(.A(k), .B(mai_mai_n254_), .Y(mai_mai_n590_));
  NOi31      m0562(.An(m), .B(n), .C(k), .Y(mai_mai_n591_));
  NA2        m0563(.A(j), .B(mai_mai_n591_), .Y(mai_mai_n592_));
  AOI210     m0564(.A0(mai_mai_n379_), .A1(mai_mai_n354_), .B0(mai_mai_n287_), .Y(mai_mai_n593_));
  NAi21      m0565(.An(mai_mai_n592_), .B(mai_mai_n593_), .Y(mai_mai_n594_));
  NO2        m0566(.A(mai_mai_n268_), .B(mai_mai_n49_), .Y(mai_mai_n595_));
  NO2        m0567(.A(mai_mai_n296_), .B(mai_mai_n566_), .Y(mai_mai_n596_));
  NO2        m0568(.A(mai_mai_n518_), .B(mai_mai_n49_), .Y(mai_mai_n597_));
  AOI220     m0569(.A0(mai_mai_n597_), .A1(mai_mai_n596_), .B0(mai_mai_n595_), .B1(mai_mai_n551_), .Y(mai_mai_n598_));
  NA3        m0570(.A(mai_mai_n598_), .B(mai_mai_n594_), .C(mai_mai_n589_), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n107_), .B(mai_mai_n36_), .Y(mai_mai_n600_));
  INV        m0572(.A(mai_mai_n346_), .Y(mai_mai_n601_));
  NO2        m0573(.A(mai_mai_n601_), .B(n), .Y(mai_mai_n602_));
  NO2        m0574(.A(mai_mai_n517_), .B(mai_mai_n172_), .Y(mai_mai_n603_));
  NA3        m0575(.A(mai_mai_n535_), .B(mai_mai_n263_), .C(mai_mai_n142_), .Y(mai_mai_n604_));
  NA2        m0576(.A(mai_mai_n495_), .B(mai_mai_n156_), .Y(mai_mai_n605_));
  NO3        m0577(.A(mai_mai_n376_), .B(mai_mai_n605_), .C(mai_mai_n88_), .Y(mai_mai_n606_));
  AOI210     m0578(.A0(mai_mai_n604_), .A1(mai_mai_n603_), .B0(mai_mai_n606_), .Y(mai_mai_n607_));
  AN3        m0579(.A(f), .B(d), .C(b), .Y(mai_mai_n608_));
  OAI210     m0580(.A0(mai_mai_n608_), .A1(mai_mai_n127_), .B0(n), .Y(mai_mai_n609_));
  NA3        m0581(.A(mai_mai_n495_), .B(mai_mai_n156_), .C(mai_mai_n206_), .Y(mai_mai_n610_));
  AOI210     m0582(.A0(mai_mai_n609_), .A1(mai_mai_n224_), .B0(mai_mai_n610_), .Y(mai_mai_n611_));
  NAi31      m0583(.An(m), .B(n), .C(k), .Y(mai_mai_n612_));
  OR2        m0584(.A(mai_mai_n132_), .B(mai_mai_n61_), .Y(mai_mai_n613_));
  OAI210     m0585(.A0(mai_mai_n613_), .A1(mai_mai_n612_), .B0(mai_mai_n243_), .Y(mai_mai_n614_));
  OAI210     m0586(.A0(mai_mai_n614_), .A1(mai_mai_n611_), .B0(j), .Y(mai_mai_n615_));
  NA2        m0587(.A(mai_mai_n615_), .B(mai_mai_n607_), .Y(mai_mai_n616_));
  NO4        m0588(.A(mai_mai_n616_), .B(mai_mai_n599_), .C(mai_mai_n587_), .D(mai_mai_n581_), .Y(mai_mai_n617_));
  NA2        m0589(.A(mai_mai_n363_), .B(mai_mai_n159_), .Y(mai_mai_n618_));
  NAi31      m0590(.An(g), .B(h), .C(f), .Y(mai_mai_n619_));
  OA210      m0591(.A0(mai_mai_n518_), .A1(n), .B0(mai_mai_n562_), .Y(mai_mai_n620_));
  NO2        m0592(.A(mai_mai_n620_), .B(mai_mai_n91_), .Y(mai_mai_n621_));
  INV        m0593(.A(mai_mai_n621_), .Y(mai_mai_n622_));
  AOI210     m0594(.A0(mai_mai_n622_), .A1(mai_mai_n618_), .B0(mai_mai_n514_), .Y(mai_mai_n623_));
  NO3        m0595(.A(g), .B(mai_mai_n205_), .C(mai_mai_n56_), .Y(mai_mai_n624_));
  NAi21      m0596(.An(h), .B(j), .Y(mai_mai_n625_));
  NO2        m0597(.A(mai_mai_n502_), .B(mai_mai_n88_), .Y(mai_mai_n626_));
  OAI210     m0598(.A0(mai_mai_n626_), .A1(mai_mai_n375_), .B0(mai_mai_n624_), .Y(mai_mai_n627_));
  OR2        m0599(.A(mai_mai_n72_), .B(mai_mai_n74_), .Y(mai_mai_n628_));
  AN2        m0600(.A(h), .B(f), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n629_), .B(mai_mai_n37_), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n99_), .B(mai_mai_n46_), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n631_), .B(mai_mai_n319_), .Y(mai_mai_n632_));
  AOI210     m0604(.A0(mai_mai_n549_), .A1(mai_mai_n408_), .B0(mai_mai_n49_), .Y(mai_mai_n633_));
  OAI220     m0605(.A0(mai_mai_n565_), .A1(mai_mai_n558_), .B0(mai_mai_n313_), .B1(mai_mai_n512_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(mai_mai_n634_), .A1(mai_mai_n633_), .B0(mai_mai_n632_), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n635_), .B(mai_mai_n627_), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n245_), .B(f), .Y(mai_mai_n637_));
  NO2        m0609(.A(mai_mai_n584_), .B(mai_mai_n61_), .Y(mai_mai_n638_));
  NO3        m0610(.A(mai_mai_n638_), .B(mai_mai_n637_), .C(mai_mai_n34_), .Y(mai_mai_n639_));
  NA2        m0611(.A(mai_mai_n316_), .B(mai_mai_n137_), .Y(mai_mai_n640_));
  NA2        m0612(.A(mai_mai_n129_), .B(mai_mai_n49_), .Y(mai_mai_n641_));
  AOI220     m0613(.A0(mai_mai_n641_), .A1(mai_mai_n515_), .B0(mai_mai_n346_), .B1(mai_mai_n112_), .Y(mai_mai_n642_));
  OR2        m0614(.A(mai_mai_n642_), .B(mai_mai_n532_), .Y(mai_mai_n643_));
  OAI210     m0615(.A0(mai_mai_n640_), .A1(mai_mai_n639_), .B0(mai_mai_n643_), .Y(mai_mai_n644_));
  NO3        m0616(.A(mai_mai_n386_), .B(mai_mai_n186_), .C(mai_mai_n185_), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n645_), .B(mai_mai_n222_), .Y(mai_mai_n646_));
  NA3        m0618(.A(mai_mai_n646_), .B(mai_mai_n247_), .C(j), .Y(mai_mai_n647_));
  NO3        m0619(.A(mai_mai_n445_), .B(mai_mai_n169_), .C(i), .Y(mai_mai_n648_));
  NA2        m0620(.A(mai_mai_n449_), .B(mai_mai_n85_), .Y(mai_mai_n649_));
  NO4        m0621(.A(mai_mai_n514_), .B(mai_mai_n649_), .C(mai_mai_n128_), .D(mai_mai_n205_), .Y(mai_mai_n650_));
  INV        m0622(.A(mai_mai_n650_), .Y(mai_mai_n651_));
  NA4        m0623(.A(mai_mai_n651_), .B(mai_mai_n647_), .C(mai_mai_n501_), .D(mai_mai_n384_), .Y(mai_mai_n652_));
  NO4        m0624(.A(mai_mai_n652_), .B(mai_mai_n644_), .C(mai_mai_n636_), .D(mai_mai_n623_), .Y(mai_mai_n653_));
  NA4        m0625(.A(mai_mai_n653_), .B(mai_mai_n617_), .C(mai_mai_n573_), .D(mai_mai_n556_), .Y(mai08));
  NO2        m0626(.A(k), .B(h), .Y(mai_mai_n655_));
  AO210      m0627(.A0(mai_mai_n245_), .A1(mai_mai_n433_), .B0(mai_mai_n655_), .Y(mai_mai_n656_));
  NO2        m0628(.A(mai_mai_n656_), .B(mai_mai_n285_), .Y(mai_mai_n657_));
  NA2        m0629(.A(mai_mai_n583_), .B(mai_mai_n85_), .Y(mai_mai_n658_));
  NA2        m0630(.A(mai_mai_n658_), .B(mai_mai_n445_), .Y(mai_mai_n659_));
  AOI210     m0631(.A0(mai_mai_n659_), .A1(mai_mai_n657_), .B0(mai_mai_n477_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n85_), .B(mai_mai_n109_), .Y(mai_mai_n661_));
  NO2        m0633(.A(mai_mai_n661_), .B(mai_mai_n57_), .Y(mai_mai_n662_));
  NO3        m0634(.A(mai_mai_n360_), .B(mai_mai_n111_), .C(mai_mai_n206_), .Y(mai_mai_n663_));
  NA2        m0635(.A(mai_mai_n553_), .B(mai_mai_n224_), .Y(mai_mai_n664_));
  AOI220     m0636(.A0(mai_mai_n664_), .A1(mai_mai_n336_), .B0(mai_mai_n663_), .B1(mai_mai_n662_), .Y(mai_mai_n665_));
  AOI210     m0637(.A0(mai_mai_n553_), .A1(mai_mai_n152_), .B0(mai_mai_n85_), .Y(mai_mai_n666_));
  NA4        m0638(.A(mai_mai_n208_), .B(mai_mai_n137_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n667_));
  AN2        m0639(.A(l), .B(k), .Y(mai_mai_n668_));
  NA3        m0640(.A(mai_mai_n665_), .B(mai_mai_n660_), .C(mai_mai_n338_), .Y(mai_mai_n669_));
  AN2        m0641(.A(mai_mai_n519_), .B(mai_mai_n96_), .Y(mai_mai_n670_));
  NO4        m0642(.A(mai_mai_n169_), .B(mai_mai_n374_), .C(mai_mai_n111_), .D(g), .Y(mai_mai_n671_));
  AOI210     m0643(.A0(mai_mai_n671_), .A1(mai_mai_n664_), .B0(mai_mai_n506_), .Y(mai_mai_n672_));
  NO2        m0644(.A(mai_mai_n38_), .B(mai_mai_n205_), .Y(mai_mai_n673_));
  NA2        m0645(.A(mai_mai_n673_), .B(mai_mai_n548_), .Y(mai_mai_n674_));
  NAi31      m0646(.An(mai_mai_n670_), .B(mai_mai_n674_), .C(mai_mai_n672_), .Y(mai_mai_n675_));
  NO2        m0647(.A(mai_mai_n521_), .B(mai_mai_n35_), .Y(mai_mai_n676_));
  OAI210     m0648(.A0(mai_mai_n535_), .A1(mai_mai_n47_), .B0(mai_mai_n613_), .Y(mai_mai_n677_));
  NO2        m0649(.A(mai_mai_n469_), .B(mai_mai_n129_), .Y(mai_mai_n678_));
  AOI210     m0650(.A0(mai_mai_n678_), .A1(mai_mai_n677_), .B0(mai_mai_n676_), .Y(mai_mai_n679_));
  NO3        m0651(.A(mai_mai_n303_), .B(mai_mai_n128_), .C(mai_mai_n41_), .Y(mai_mai_n680_));
  NA2        m0652(.A(mai_mai_n656_), .B(mai_mai_n133_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n681_), .B(mai_mai_n385_), .Y(mai_mai_n682_));
  NA2        m0654(.A(mai_mai_n679_), .B(mai_mai_n682_), .Y(mai_mai_n683_));
  NA2        m0655(.A(mai_mai_n346_), .B(mai_mai_n43_), .Y(mai_mai_n684_));
  NA3        m0656(.A(mai_mai_n646_), .B(mai_mai_n321_), .C(mai_mai_n366_), .Y(mai_mai_n685_));
  NA2        m0657(.A(mai_mai_n668_), .B(mai_mai_n212_), .Y(mai_mai_n686_));
  NO2        m0658(.A(mai_mai_n686_), .B(mai_mai_n315_), .Y(mai_mai_n687_));
  AOI210     m0659(.A0(mai_mai_n687_), .A1(mai_mai_n637_), .B0(mai_mai_n476_), .Y(mai_mai_n688_));
  NA3        m0660(.A(m), .B(l), .C(k), .Y(mai_mai_n689_));
  NO2        m0661(.A(mai_mai_n520_), .B(mai_mai_n264_), .Y(mai_mai_n690_));
  NOi21      m0662(.An(mai_mai_n690_), .B(mai_mai_n516_), .Y(mai_mai_n691_));
  NA4        m0663(.A(mai_mai_n112_), .B(l), .C(k), .D(mai_mai_n88_), .Y(mai_mai_n692_));
  NA3        m0664(.A(mai_mai_n120_), .B(mai_mai_n394_), .C(i), .Y(mai_mai_n693_));
  NO2        m0665(.A(mai_mai_n693_), .B(mai_mai_n692_), .Y(mai_mai_n694_));
  NO2        m0666(.A(mai_mai_n694_), .B(mai_mai_n691_), .Y(mai_mai_n695_));
  NA4        m0667(.A(mai_mai_n695_), .B(mai_mai_n688_), .C(mai_mai_n685_), .D(mai_mai_n684_), .Y(mai_mai_n696_));
  NO4        m0668(.A(mai_mai_n696_), .B(mai_mai_n683_), .C(mai_mai_n675_), .D(mai_mai_n669_), .Y(mai_mai_n697_));
  NA2        m0669(.A(mai_mai_n585_), .B(mai_mai_n375_), .Y(mai_mai_n698_));
  NO3        m0670(.A(mai_mai_n379_), .B(mai_mai_n512_), .C(h), .Y(mai_mai_n699_));
  AOI210     m0671(.A0(mai_mai_n699_), .A1(mai_mai_n112_), .B0(mai_mai_n488_), .Y(mai_mai_n700_));
  NA3        m0672(.A(mai_mai_n700_), .B(mai_mai_n698_), .C(mai_mai_n244_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n668_), .B(mai_mai_n74_), .Y(mai_mai_n702_));
  NO4        m0674(.A(mai_mai_n645_), .B(mai_mai_n169_), .C(n), .D(i), .Y(mai_mai_n703_));
  NOi21      m0675(.An(h), .B(j), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n704_), .B(f), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n705_), .B(mai_mai_n238_), .Y(mai_mai_n706_));
  NO3        m0678(.A(mai_mai_n706_), .B(mai_mai_n703_), .C(mai_mai_n648_), .Y(mai_mai_n707_));
  NO2        m0679(.A(mai_mai_n707_), .B(mai_mai_n702_), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n701_), .A1(l), .B0(mai_mai_n708_), .Y(mai_mai_n709_));
  NO2        m0681(.A(j), .B(i), .Y(mai_mai_n710_));
  NA3        m0682(.A(mai_mai_n710_), .B(mai_mai_n81_), .C(l), .Y(mai_mai_n711_));
  NA2        m0683(.A(mai_mai_n710_), .B(mai_mai_n33_), .Y(mai_mai_n712_));
  NA2        m0684(.A(mai_mai_n401_), .B(mai_mai_n120_), .Y(mai_mai_n713_));
  OA220      m0685(.A0(mai_mai_n713_), .A1(mai_mai_n712_), .B0(mai_mai_n711_), .B1(mai_mai_n564_), .Y(mai_mai_n714_));
  NO3        m0686(.A(mai_mai_n149_), .B(mai_mai_n49_), .C(mai_mai_n109_), .Y(mai_mai_n715_));
  NO3        m0687(.A(mai_mai_n527_), .B(mai_mai_n147_), .C(mai_mai_n74_), .Y(mai_mai_n716_));
  NO3        m0688(.A(mai_mai_n469_), .B(mai_mai_n420_), .C(j), .Y(mai_mai_n717_));
  OAI210     m0689(.A0(mai_mai_n716_), .A1(mai_mai_n715_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  INV        m0690(.A(mai_mai_n718_), .Y(mai_mai_n719_));
  NA2        m0691(.A(k), .B(j), .Y(mai_mai_n720_));
  AOI210     m0692(.A0(mai_mai_n515_), .A1(n), .B0(mai_mai_n534_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n721_), .B(mai_mai_n537_), .Y(mai_mai_n722_));
  NO3        m0694(.A(mai_mai_n169_), .B(mai_mai_n374_), .C(mai_mai_n111_), .Y(mai_mai_n723_));
  NA2        m0695(.A(mai_mai_n723_), .B(mai_mai_n239_), .Y(mai_mai_n724_));
  NAi31      m0696(.An(mai_mai_n571_), .B(mai_mai_n93_), .C(mai_mai_n85_), .Y(mai_mai_n725_));
  NA2        m0697(.A(mai_mai_n725_), .B(mai_mai_n724_), .Y(mai_mai_n726_));
  NO2        m0698(.A(mai_mai_n285_), .B(mai_mai_n133_), .Y(mai_mai_n727_));
  AOI220     m0699(.A0(mai_mai_n727_), .A1(mai_mai_n585_), .B0(mai_mai_n680_), .B1(mai_mai_n666_), .Y(mai_mai_n728_));
  NO2        m0700(.A(mai_mai_n689_), .B(mai_mai_n91_), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n729_), .B(mai_mai_n563_), .Y(mai_mai_n730_));
  NO2        m0702(.A(mai_mai_n565_), .B(mai_mai_n116_), .Y(mai_mai_n731_));
  OAI210     m0703(.A0(mai_mai_n731_), .A1(mai_mai_n717_), .B0(mai_mai_n633_), .Y(mai_mai_n732_));
  NA3        m0704(.A(mai_mai_n732_), .B(mai_mai_n730_), .C(mai_mai_n728_), .Y(mai_mai_n733_));
  OR3        m0705(.A(mai_mai_n733_), .B(mai_mai_n726_), .C(mai_mai_n719_), .Y(mai_mai_n734_));
  NA3        m0706(.A(mai_mai_n721_), .B(mai_mai_n537_), .C(mai_mai_n536_), .Y(mai_mai_n735_));
  NA4        m0707(.A(mai_mai_n735_), .B(mai_mai_n208_), .C(mai_mai_n433_), .D(mai_mai_n34_), .Y(mai_mai_n736_));
  NO4        m0708(.A(mai_mai_n469_), .B(mai_mai_n415_), .C(j), .D(f), .Y(mai_mai_n737_));
  OAI220     m0709(.A0(mai_mai_n667_), .A1(mai_mai_n658_), .B0(mai_mai_n319_), .B1(mai_mai_n38_), .Y(mai_mai_n738_));
  AOI210     m0710(.A0(mai_mai_n737_), .A1(mai_mai_n251_), .B0(mai_mai_n738_), .Y(mai_mai_n739_));
  NA3        m0711(.A(mai_mai_n529_), .B(mai_mai_n278_), .C(h), .Y(mai_mai_n740_));
  NOi21      m0712(.An(mai_mai_n633_), .B(mai_mai_n740_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n92_), .B(mai_mai_n47_), .Y(mai_mai_n742_));
  NO2        m0714(.A(mai_mai_n711_), .B(mai_mai_n628_), .Y(mai_mai_n743_));
  AOI210     m0715(.A0(mai_mai_n742_), .A1(mai_mai_n602_), .B0(mai_mai_n743_), .Y(mai_mai_n744_));
  NAi41      m0716(.An(mai_mai_n741_), .B(mai_mai_n744_), .C(mai_mai_n739_), .D(mai_mai_n736_), .Y(mai_mai_n745_));
  OR2        m0717(.A(mai_mai_n729_), .B(mai_mai_n96_), .Y(mai_mai_n746_));
  AOI220     m0718(.A0(mai_mai_n746_), .A1(mai_mai_n230_), .B0(mai_mai_n717_), .B1(mai_mai_n595_), .Y(mai_mai_n747_));
  NO2        m0719(.A(mai_mai_n620_), .B(mai_mai_n74_), .Y(mai_mai_n748_));
  AOI210     m0720(.A0(mai_mai_n737_), .A1(mai_mai_n748_), .B0(mai_mai_n323_), .Y(mai_mai_n749_));
  AOI220     m0721(.A0(mai_mai_n569_), .A1(mai_mai_n29_), .B0(mai_mai_n449_), .B1(mai_mai_n85_), .Y(mai_mai_n750_));
  NO2        m0722(.A(mai_mai_n740_), .B(mai_mai_n475_), .Y(mai_mai_n751_));
  INV        m0723(.A(mai_mai_n751_), .Y(mai_mai_n752_));
  NA3        m0724(.A(mai_mai_n752_), .B(mai_mai_n749_), .C(mai_mai_n747_), .Y(mai_mai_n753_));
  NOi41      m0725(.An(mai_mai_n714_), .B(mai_mai_n753_), .C(mai_mai_n745_), .D(mai_mai_n734_), .Y(mai_mai_n754_));
  OR2        m0726(.A(mai_mai_n667_), .B(mai_mai_n224_), .Y(mai_mai_n755_));
  NO3        m0727(.A(mai_mai_n329_), .B(mai_mai_n287_), .C(mai_mai_n111_), .Y(mai_mai_n756_));
  NA2        m0728(.A(mai_mai_n756_), .B(mai_mai_n722_), .Y(mai_mai_n757_));
  NA2        m0729(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n758_));
  NO3        m0730(.A(mai_mai_n758_), .B(mai_mai_n712_), .C(mai_mai_n268_), .Y(mai_mai_n759_));
  INV        m0731(.A(mai_mai_n759_), .Y(mai_mai_n760_));
  NA4        m0732(.A(mai_mai_n760_), .B(mai_mai_n757_), .C(mai_mai_n755_), .D(mai_mai_n387_), .Y(mai_mai_n761_));
  OR2        m0733(.A(mai_mai_n619_), .B(mai_mai_n92_), .Y(mai_mai_n762_));
  NOi31      m0734(.An(b), .B(d), .C(a), .Y(mai_mai_n763_));
  NO2        m0735(.A(mai_mai_n763_), .B(mai_mai_n568_), .Y(mai_mai_n764_));
  NO2        m0736(.A(mai_mai_n764_), .B(n), .Y(mai_mai_n765_));
  NOi21      m0737(.An(mai_mai_n750_), .B(mai_mai_n765_), .Y(mai_mai_n766_));
  NO2        m0738(.A(mai_mai_n766_), .B(mai_mai_n762_), .Y(mai_mai_n767_));
  NO2        m0739(.A(mai_mai_n535_), .B(mai_mai_n85_), .Y(mai_mai_n768_));
  NA2        m0740(.A(mai_mai_n756_), .B(mai_mai_n768_), .Y(mai_mai_n769_));
  OAI210     m0741(.A0(mai_mai_n667_), .A1(mai_mai_n376_), .B0(mai_mai_n769_), .Y(mai_mai_n770_));
  NO2        m0742(.A(mai_mai_n645_), .B(n), .Y(mai_mai_n771_));
  BUFFER     m0743(.A(mai_mai_n727_), .Y(mai_mai_n772_));
  AOI220     m0744(.A0(mai_mai_n772_), .A1(mai_mai_n624_), .B0(mai_mai_n771_), .B1(mai_mai_n657_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n310_), .B(mai_mai_n229_), .Y(mai_mai_n774_));
  OAI210     m0746(.A0(mai_mai_n96_), .A1(mai_mai_n93_), .B0(mai_mai_n774_), .Y(mai_mai_n775_));
  NA2        m0747(.A(mai_mai_n120_), .B(mai_mai_n85_), .Y(mai_mai_n776_));
  AOI210     m0748(.A0(mai_mai_n405_), .A1(mai_mai_n398_), .B0(mai_mai_n776_), .Y(mai_mai_n777_));
  NAi21      m0749(.An(mai_mai_n777_), .B(mai_mai_n775_), .Y(mai_mai_n778_));
  NA2        m0750(.A(mai_mai_n687_), .B(mai_mai_n34_), .Y(mai_mai_n779_));
  NAi21      m0751(.An(mai_mai_n692_), .B(mai_mai_n416_), .Y(mai_mai_n780_));
  NO2        m0752(.A(mai_mai_n264_), .B(i), .Y(mai_mai_n781_));
  NA2        m0753(.A(mai_mai_n671_), .B(mai_mai_n337_), .Y(mai_mai_n782_));
  AN2        m0754(.A(mai_mai_n782_), .B(mai_mai_n780_), .Y(mai_mai_n783_));
  NAi41      m0755(.An(mai_mai_n778_), .B(mai_mai_n783_), .C(mai_mai_n779_), .D(mai_mai_n773_), .Y(mai_mai_n784_));
  NO4        m0756(.A(mai_mai_n784_), .B(mai_mai_n770_), .C(mai_mai_n767_), .D(mai_mai_n761_), .Y(mai_mai_n785_));
  NA4        m0757(.A(mai_mai_n785_), .B(mai_mai_n754_), .C(mai_mai_n709_), .D(mai_mai_n697_), .Y(mai09));
  INV        m0758(.A(mai_mai_n121_), .Y(mai_mai_n787_));
  NA2        m0759(.A(f), .B(e), .Y(mai_mai_n788_));
  NO2        m0760(.A(mai_mai_n217_), .B(mai_mai_n111_), .Y(mai_mai_n789_));
  NA2        m0761(.A(mai_mai_n789_), .B(g), .Y(mai_mai_n790_));
  NA3        m0762(.A(mai_mai_n296_), .B(mai_mai_n253_), .C(mai_mai_n118_), .Y(mai_mai_n791_));
  AOI210     m0763(.A0(mai_mai_n791_), .A1(g), .B0(mai_mai_n455_), .Y(mai_mai_n792_));
  AOI210     m0764(.A0(mai_mai_n792_), .A1(mai_mai_n790_), .B0(mai_mai_n788_), .Y(mai_mai_n793_));
  NA2        m0765(.A(mai_mai_n426_), .B(e), .Y(mai_mai_n794_));
  NO2        m0766(.A(mai_mai_n794_), .B(mai_mai_n498_), .Y(mai_mai_n795_));
  AOI210     m0767(.A0(mai_mai_n793_), .A1(mai_mai_n787_), .B0(mai_mai_n795_), .Y(mai_mai_n796_));
  NA3        m0768(.A(m), .B(l), .C(i), .Y(mai_mai_n797_));
  OAI220     m0769(.A0(mai_mai_n565_), .A1(mai_mai_n797_), .B0(mai_mai_n340_), .B1(mai_mai_n513_), .Y(mai_mai_n798_));
  NA4        m0770(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(g), .D(f), .Y(mai_mai_n799_));
  NAi31      m0771(.An(mai_mai_n798_), .B(mai_mai_n799_), .C(mai_mai_n421_), .Y(mai_mai_n800_));
  NA2        m0772(.A(mai_mai_n762_), .B(mai_mai_n505_), .Y(mai_mai_n801_));
  OA210      m0773(.A0(mai_mai_n801_), .A1(mai_mai_n800_), .B0(mai_mai_n765_), .Y(mai_mai_n802_));
  INV        m0774(.A(mai_mai_n326_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n126_), .B(mai_mai_n125_), .Y(mai_mai_n804_));
  NOi31      m0776(.An(k), .B(m), .C(l), .Y(mai_mai_n805_));
  NO2        m0777(.A(mai_mai_n328_), .B(mai_mai_n805_), .Y(mai_mai_n806_));
  AOI210     m0778(.A0(mai_mai_n806_), .A1(mai_mai_n804_), .B0(mai_mai_n566_), .Y(mai_mai_n807_));
  INV        m0779(.A(mai_mai_n319_), .Y(mai_mai_n808_));
  NA2        m0780(.A(mai_mai_n807_), .B(mai_mai_n803_), .Y(mai_mai_n809_));
  NA2        m0781(.A(mai_mai_n163_), .B(mai_mai_n113_), .Y(mai_mai_n810_));
  NA3        m0782(.A(mai_mai_n810_), .B(mai_mai_n656_), .C(mai_mai_n133_), .Y(mai_mai_n811_));
  NA3        m0783(.A(mai_mai_n811_), .B(mai_mai_n183_), .C(mai_mai_n31_), .Y(mai_mai_n812_));
  NA4        m0784(.A(mai_mai_n812_), .B(mai_mai_n809_), .C(mai_mai_n586_), .D(mai_mai_n83_), .Y(mai_mai_n813_));
  NO2        m0785(.A(mai_mai_n561_), .B(mai_mai_n484_), .Y(mai_mai_n814_));
  NA2        m0786(.A(mai_mai_n814_), .B(mai_mai_n183_), .Y(mai_mai_n815_));
  NOi21      m0787(.An(f), .B(d), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n816_), .B(m), .Y(mai_mai_n817_));
  NA3        m0789(.A(mai_mai_n296_), .B(mai_mai_n253_), .C(mai_mai_n118_), .Y(mai_mai_n818_));
  AN2        m0790(.A(f), .B(d), .Y(mai_mai_n819_));
  NA3        m0791(.A(mai_mai_n461_), .B(mai_mai_n819_), .C(mai_mai_n85_), .Y(mai_mai_n820_));
  NO3        m0792(.A(mai_mai_n820_), .B(mai_mai_n74_), .C(mai_mai_n206_), .Y(mai_mai_n821_));
  NO2        m0793(.A(k), .B(mai_mai_n56_), .Y(mai_mai_n822_));
  NA2        m0794(.A(mai_mai_n818_), .B(mai_mai_n821_), .Y(mai_mai_n823_));
  NAi31      m0795(.An(mai_mai_n474_), .B(mai_mai_n823_), .C(mai_mai_n815_), .Y(mai_mai_n824_));
  NO4        m0796(.A(mai_mai_n584_), .B(mai_mai_n129_), .C(mai_mai_n315_), .D(mai_mai_n150_), .Y(mai_mai_n825_));
  NO2        m0797(.A(mai_mai_n612_), .B(mai_mai_n315_), .Y(mai_mai_n826_));
  AN2        m0798(.A(mai_mai_n826_), .B(mai_mai_n637_), .Y(mai_mai_n827_));
  NO3        m0799(.A(mai_mai_n827_), .B(mai_mai_n825_), .C(mai_mai_n226_), .Y(mai_mai_n828_));
  NA2        m0800(.A(mai_mai_n568_), .B(mai_mai_n85_), .Y(mai_mai_n829_));
  NA3        m0801(.A(mai_mai_n156_), .B(mai_mai_n107_), .C(mai_mai_n106_), .Y(mai_mai_n830_));
  OAI220     m0802(.A0(mai_mai_n820_), .A1(mai_mai_n410_), .B0(mai_mai_n326_), .B1(mai_mai_n830_), .Y(mai_mai_n831_));
  NOi31      m0803(.An(mai_mai_n215_), .B(mai_mai_n831_), .C(mai_mai_n292_), .Y(mai_mai_n832_));
  NA2        m0804(.A(c), .B(mai_mai_n115_), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n833_), .B(mai_mai_n391_), .Y(mai_mai_n834_));
  NA3        m0806(.A(mai_mai_n834_), .B(mai_mai_n497_), .C(f), .Y(mai_mai_n835_));
  OR2        m0807(.A(mai_mai_n619_), .B(mai_mai_n524_), .Y(mai_mai_n836_));
  INV        m0808(.A(mai_mai_n836_), .Y(mai_mai_n837_));
  NA2        m0809(.A(mai_mai_n764_), .B(mai_mai_n110_), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n838_), .B(mai_mai_n837_), .Y(mai_mai_n839_));
  NA4        m0811(.A(mai_mai_n839_), .B(mai_mai_n835_), .C(mai_mai_n832_), .D(mai_mai_n828_), .Y(mai_mai_n840_));
  NO4        m0812(.A(mai_mai_n840_), .B(mai_mai_n824_), .C(mai_mai_n813_), .D(mai_mai_n802_), .Y(mai_mai_n841_));
  OR2        m0813(.A(mai_mai_n820_), .B(mai_mai_n74_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n111_), .B(j), .Y(mai_mai_n843_));
  NA2        m0815(.A(mai_mai_n789_), .B(g), .Y(mai_mai_n844_));
  AOI210     m0816(.A0(mai_mai_n844_), .A1(mai_mai_n279_), .B0(mai_mai_n842_), .Y(mai_mai_n845_));
  NO2        m0817(.A(mai_mai_n319_), .B(mai_mai_n799_), .Y(mai_mai_n846_));
  NO2        m0818(.A(mai_mai_n133_), .B(mai_mai_n129_), .Y(mai_mai_n847_));
  NO2        m0819(.A(mai_mai_n222_), .B(mai_mai_n216_), .Y(mai_mai_n848_));
  AOI220     m0820(.A0(mai_mai_n848_), .A1(mai_mai_n219_), .B0(mai_mai_n290_), .B1(mai_mai_n847_), .Y(mai_mai_n849_));
  NO2        m0821(.A(mai_mai_n410_), .B(mai_mai_n788_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n850_), .B(mai_mai_n542_), .Y(mai_mai_n851_));
  NA2        m0823(.A(mai_mai_n851_), .B(mai_mai_n849_), .Y(mai_mai_n852_));
  NA2        m0824(.A(e), .B(d), .Y(mai_mai_n853_));
  OAI220     m0825(.A0(mai_mai_n853_), .A1(c), .B0(mai_mai_n310_), .B1(d), .Y(mai_mai_n854_));
  NA3        m0826(.A(mai_mai_n854_), .B(mai_mai_n438_), .C(mai_mai_n495_), .Y(mai_mai_n855_));
  AOI210     m0827(.A0(mai_mai_n502_), .A1(mai_mai_n176_), .B0(mai_mai_n222_), .Y(mai_mai_n856_));
  INV        m0828(.A(mai_mai_n856_), .Y(mai_mai_n857_));
  NA3        m0829(.A(mai_mai_n162_), .B(mai_mai_n86_), .C(mai_mai_n34_), .Y(mai_mai_n858_));
  NA3        m0830(.A(mai_mai_n858_), .B(mai_mai_n857_), .C(mai_mai_n855_), .Y(mai_mai_n859_));
  NO4        m0831(.A(mai_mai_n859_), .B(mai_mai_n852_), .C(mai_mai_n846_), .D(mai_mai_n845_), .Y(mai_mai_n860_));
  NA2        m0832(.A(mai_mai_n803_), .B(mai_mai_n31_), .Y(mai_mai_n861_));
  OR2        m0833(.A(mai_mai_n861_), .B(mai_mai_n209_), .Y(mai_mai_n862_));
  OAI220     m0834(.A0(mai_mai_n584_), .A1(mai_mai_n61_), .B0(mai_mai_n287_), .B1(j), .Y(mai_mai_n863_));
  AOI220     m0835(.A0(mai_mai_n863_), .A1(mai_mai_n826_), .B0(mai_mai_n574_), .B1(mai_mai_n583_), .Y(mai_mai_n864_));
  OAI210     m0836(.A0(mai_mai_n794_), .A1(mai_mai_n166_), .B0(mai_mai_n864_), .Y(mai_mai_n865_));
  AN2        m0837(.A(mai_mai_n808_), .B(mai_mai_n798_), .Y(mai_mai_n866_));
  NOi31      m0838(.An(mai_mai_n528_), .B(mai_mai_n817_), .C(mai_mai_n279_), .Y(mai_mai_n867_));
  NO3        m0839(.A(mai_mai_n867_), .B(mai_mai_n866_), .C(mai_mai_n865_), .Y(mai_mai_n868_));
  AO220      m0840(.A0(mai_mai_n438_), .A1(mai_mai_n704_), .B0(mai_mai_n171_), .B1(f), .Y(mai_mai_n869_));
  OAI210     m0841(.A0(mai_mai_n869_), .A1(mai_mai_n441_), .B0(mai_mai_n854_), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n420_), .B(mai_mai_n71_), .Y(mai_mai_n871_));
  OAI210     m0843(.A0(mai_mai_n801_), .A1(mai_mai_n871_), .B0(mai_mai_n662_), .Y(mai_mai_n872_));
  AN4        m0844(.A(mai_mai_n872_), .B(mai_mai_n870_), .C(mai_mai_n868_), .D(mai_mai_n862_), .Y(mai_mai_n873_));
  NA4        m0845(.A(mai_mai_n873_), .B(mai_mai_n860_), .C(mai_mai_n841_), .D(mai_mai_n796_), .Y(mai12));
  NO4        m0846(.A(mai_mai_n425_), .B(mai_mai_n245_), .C(mai_mai_n557_), .D(mai_mai_n206_), .Y(mai_mai_n875_));
  NA2        m0847(.A(mai_mai_n528_), .B(mai_mai_n871_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n436_), .B(mai_mai_n115_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n804_), .B(mai_mai_n340_), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n619_), .B(mai_mai_n360_), .Y(mai_mai_n879_));
  NA2        m0851(.A(mai_mai_n876_), .B(mai_mai_n424_), .Y(mai_mai_n880_));
  AOI210     m0852(.A0(mai_mai_n225_), .A1(mai_mai_n325_), .B0(mai_mai_n195_), .Y(mai_mai_n881_));
  OR2        m0853(.A(mai_mai_n881_), .B(mai_mai_n875_), .Y(mai_mai_n882_));
  AOI210     m0854(.A0(mai_mai_n322_), .A1(mai_mai_n372_), .B0(mai_mai_n206_), .Y(mai_mai_n883_));
  OAI210     m0855(.A0(mai_mai_n883_), .A1(mai_mai_n882_), .B0(mai_mai_n386_), .Y(mai_mai_n884_));
  NO2        m0856(.A(mai_mai_n600_), .B(mai_mai_n254_), .Y(mai_mai_n885_));
  NO2        m0857(.A(mai_mai_n565_), .B(mai_mai_n797_), .Y(mai_mai_n886_));
  NA2        m0858(.A(mai_mai_n774_), .B(mai_mai_n885_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n149_), .B(mai_mai_n229_), .Y(mai_mai_n888_));
  NA2        m0860(.A(mai_mai_n887_), .B(mai_mai_n884_), .Y(mai_mai_n889_));
  OR2        m0861(.A(mai_mai_n311_), .B(mai_mai_n877_), .Y(mai_mai_n890_));
  NA2        m0862(.A(mai_mai_n890_), .B(mai_mai_n341_), .Y(mai_mai_n891_));
  NO3        m0863(.A(mai_mai_n129_), .B(mai_mai_n150_), .C(mai_mai_n206_), .Y(mai_mai_n892_));
  NA2        m0864(.A(mai_mai_n892_), .B(mai_mai_n515_), .Y(mai_mai_n893_));
  NA4        m0865(.A(mai_mai_n426_), .B(mai_mai_n418_), .C(mai_mai_n177_), .D(g), .Y(mai_mai_n894_));
  NA3        m0866(.A(mai_mai_n894_), .B(mai_mai_n893_), .C(mai_mai_n891_), .Y(mai_mai_n895_));
  NO3        m0867(.A(mai_mai_n895_), .B(mai_mai_n889_), .C(mai_mai_n880_), .Y(mai_mai_n896_));
  NO2        m0868(.A(mai_mai_n351_), .B(mai_mai_n350_), .Y(mai_mai_n897_));
  NA2        m0869(.A(mai_mai_n562_), .B(mai_mai_n72_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n535_), .B(mai_mai_n142_), .Y(mai_mai_n899_));
  NOi21      m0871(.An(mai_mai_n34_), .B(mai_mai_n612_), .Y(mai_mai_n900_));
  AOI220     m0872(.A0(mai_mai_n900_), .A1(mai_mai_n899_), .B0(mai_mai_n898_), .B1(mai_mai_n897_), .Y(mai_mai_n901_));
  OAI210     m0873(.A0(mai_mai_n243_), .A1(mai_mai_n45_), .B0(mai_mai_n901_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n416_), .B(mai_mai_n256_), .Y(mai_mai_n903_));
  NO3        m0875(.A(mai_mai_n776_), .B(mai_mai_n90_), .C(mai_mai_n391_), .Y(mai_mai_n904_));
  NAi31      m0876(.An(mai_mai_n904_), .B(mai_mai_n903_), .C(mai_mai_n307_), .Y(mai_mai_n905_));
  NO2        m0877(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n906_));
  NO2        m0878(.A(mai_mai_n491_), .B(mai_mai_n287_), .Y(mai_mai_n907_));
  INV        m0879(.A(mai_mai_n907_), .Y(mai_mai_n908_));
  NO2        m0880(.A(mai_mai_n908_), .B(mai_mai_n142_), .Y(mai_mai_n909_));
  NA2        m0881(.A(mai_mai_n591_), .B(j), .Y(mai_mai_n910_));
  OAI210     m0882(.A0(mai_mai_n693_), .A1(mai_mai_n910_), .B0(mai_mai_n348_), .Y(mai_mai_n911_));
  NO4        m0883(.A(mai_mai_n911_), .B(mai_mai_n909_), .C(mai_mai_n905_), .D(mai_mai_n902_), .Y(mai_mai_n912_));
  NA2        m0884(.A(mai_mai_n335_), .B(g), .Y(mai_mai_n913_));
  NA2        m0885(.A(mai_mai_n159_), .B(i), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n915_));
  OAI220     m0887(.A0(mai_mai_n915_), .A1(mai_mai_n194_), .B0(mai_mai_n914_), .B1(mai_mai_n92_), .Y(mai_mai_n916_));
  AOI210     m0888(.A0(mai_mai_n400_), .A1(mai_mai_n37_), .B0(mai_mai_n916_), .Y(mai_mai_n917_));
  NO2        m0889(.A(mai_mai_n142_), .B(mai_mai_n85_), .Y(mai_mai_n918_));
  OR2        m0890(.A(mai_mai_n918_), .B(mai_mai_n534_), .Y(mai_mai_n919_));
  NA2        m0891(.A(mai_mai_n535_), .B(mai_mai_n364_), .Y(mai_mai_n920_));
  AOI210     m0892(.A0(mai_mai_n920_), .A1(n), .B0(mai_mai_n919_), .Y(mai_mai_n921_));
  OAI220     m0893(.A0(mai_mai_n921_), .A1(mai_mai_n913_), .B0(mai_mai_n917_), .B1(mai_mai_n319_), .Y(mai_mai_n922_));
  NO2        m0894(.A(mai_mai_n619_), .B(mai_mai_n484_), .Y(mai_mai_n923_));
  OAI210     m0895(.A0(mai_mai_n633_), .A1(mai_mai_n716_), .B0(mai_mai_n923_), .Y(mai_mai_n924_));
  OR3        m0896(.A(mai_mai_n296_), .B(mai_mai_n415_), .C(f), .Y(mai_mai_n925_));
  OR2        m0897(.A(mai_mai_n925_), .B(mai_mai_n564_), .Y(mai_mai_n926_));
  NA3        m0898(.A(mai_mai_n312_), .B(mai_mai_n117_), .C(g), .Y(mai_mai_n927_));
  AOI210     m0899(.A0(mai_mai_n630_), .A1(mai_mai_n927_), .B0(m), .Y(mai_mai_n928_));
  OAI210     m0900(.A0(mai_mai_n928_), .A1(mai_mai_n878_), .B0(mai_mai_n311_), .Y(mai_mai_n929_));
  NA2        m0901(.A(mai_mai_n649_), .B(mai_mai_n829_), .Y(mai_mai_n930_));
  NA2        m0902(.A(mai_mai_n799_), .B(mai_mai_n421_), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n213_), .B(mai_mai_n78_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n932_), .B(mai_mai_n925_), .Y(mai_mai_n933_));
  AOI220     m0905(.A0(mai_mai_n933_), .A1(mai_mai_n251_), .B0(mai_mai_n931_), .B1(mai_mai_n930_), .Y(mai_mai_n934_));
  NA4        m0906(.A(mai_mai_n934_), .B(mai_mai_n929_), .C(mai_mai_n926_), .D(mai_mai_n924_), .Y(mai_mai_n935_));
  NA2        m0907(.A(mai_mai_n621_), .B(mai_mai_n89_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n444_), .B(mai_mai_n206_), .Y(mai_mai_n937_));
  AOI220     m0909(.A0(mai_mai_n937_), .A1(mai_mai_n365_), .B0(mai_mai_n890_), .B1(mai_mai_n210_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n879_), .B(mai_mai_n888_), .Y(mai_mai_n939_));
  NA3        m0911(.A(mai_mai_n939_), .B(mai_mai_n938_), .C(mai_mai_n936_), .Y(mai_mai_n940_));
  OAI210     m0912(.A0(mai_mai_n931_), .A1(mai_mai_n886_), .B0(mai_mai_n526_), .Y(mai_mai_n941_));
  OAI210     m0913(.A0(mai_mai_n351_), .A1(mai_mai_n350_), .B0(mai_mai_n108_), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n942_), .B(mai_mai_n519_), .Y(mai_mai_n943_));
  NA2        m0915(.A(mai_mai_n928_), .B(mai_mai_n877_), .Y(mai_mai_n944_));
  NO3        m0916(.A(mai_mai_n843_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n945_));
  AOI220     m0917(.A0(mai_mai_n945_), .A1(mai_mai_n588_), .B0(mai_mai_n603_), .B1(mai_mai_n515_), .Y(mai_mai_n946_));
  NA4        m0918(.A(mai_mai_n946_), .B(mai_mai_n944_), .C(mai_mai_n943_), .D(mai_mai_n941_), .Y(mai_mai_n947_));
  NO4        m0919(.A(mai_mai_n947_), .B(mai_mai_n940_), .C(mai_mai_n935_), .D(mai_mai_n922_), .Y(mai_mai_n948_));
  NAi31      m0920(.An(mai_mai_n138_), .B(mai_mai_n401_), .C(n), .Y(mai_mai_n949_));
  NO3        m0921(.A(mai_mai_n125_), .B(mai_mai_n328_), .C(mai_mai_n805_), .Y(mai_mai_n950_));
  NO2        m0922(.A(mai_mai_n950_), .B(mai_mai_n949_), .Y(mai_mai_n951_));
  NO3        m0923(.A(mai_mai_n264_), .B(mai_mai_n138_), .C(mai_mai_n391_), .Y(mai_mai_n952_));
  AOI210     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n485_), .B0(mai_mai_n951_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n477_), .B(i), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n954_), .B(mai_mai_n953_), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n222_), .B(mai_mai_n167_), .Y(mai_mai_n956_));
  NO3        m0928(.A(mai_mai_n294_), .B(mai_mai_n426_), .C(mai_mai_n171_), .Y(mai_mai_n957_));
  NOi31      m0929(.An(mai_mai_n956_), .B(mai_mai_n957_), .C(mai_mai_n206_), .Y(mai_mai_n958_));
  NAi21      m0930(.An(mai_mai_n535_), .B(mai_mai_n937_), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n419_), .B(mai_mai_n829_), .Y(mai_mai_n960_));
  NO3        m0932(.A(mai_mai_n420_), .B(mai_mai_n296_), .C(mai_mai_n74_), .Y(mai_mai_n961_));
  AOI220     m0933(.A0(mai_mai_n961_), .A1(mai_mai_n960_), .B0(mai_mai_n467_), .B1(g), .Y(mai_mai_n962_));
  NA2        m0934(.A(mai_mai_n962_), .B(mai_mai_n959_), .Y(mai_mai_n963_));
  NO3        m0935(.A(mai_mai_n527_), .B(mai_mai_n147_), .C(mai_mai_n205_), .Y(mai_mai_n964_));
  OAI210     m0936(.A0(mai_mai_n964_), .A1(mai_mai_n511_), .B0(mai_mai_n361_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n965_), .B(mai_mai_n582_), .Y(mai_mai_n966_));
  OAI210     m0938(.A0(mai_mai_n881_), .A1(mai_mai_n875_), .B0(mai_mai_n956_), .Y(mai_mai_n967_));
  NA3        m0939(.A(mai_mai_n920_), .B(mai_mai_n471_), .C(mai_mai_n46_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n363_), .B(mai_mai_n361_), .Y(mai_mai_n969_));
  NA3        m0941(.A(mai_mai_n969_), .B(mai_mai_n968_), .C(mai_mai_n967_), .Y(mai_mai_n970_));
  OR2        m0942(.A(mai_mai_n970_), .B(mai_mai_n966_), .Y(mai_mai_n971_));
  NO4        m0943(.A(mai_mai_n971_), .B(mai_mai_n963_), .C(mai_mai_n958_), .D(mai_mai_n955_), .Y(mai_mai_n972_));
  NA4        m0944(.A(mai_mai_n972_), .B(mai_mai_n948_), .C(mai_mai_n912_), .D(mai_mai_n896_), .Y(mai13));
  INV        m0945(.A(mai_mai_n46_), .Y(mai_mai_n974_));
  AN2        m0946(.A(c), .B(b), .Y(mai_mai_n975_));
  NA3        m0947(.A(mai_mai_n242_), .B(mai_mai_n975_), .C(m), .Y(mai_mai_n976_));
  NA2        m0948(.A(mai_mai_n482_), .B(f), .Y(mai_mai_n977_));
  NO4        m0949(.A(mai_mai_n977_), .B(mai_mai_n976_), .C(mai_mai_n974_), .D(mai_mai_n558_), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n256_), .B(mai_mai_n975_), .Y(mai_mai_n979_));
  NO3        m0951(.A(mai_mai_n979_), .B(mai_mai_n977_), .C(mai_mai_n914_), .Y(mai_mai_n980_));
  NAi32      m0952(.An(d), .Bn(c), .C(e), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n137_), .B(mai_mai_n45_), .Y(mai_mai_n982_));
  NO4        m0954(.A(mai_mai_n982_), .B(mai_mai_n981_), .C(mai_mai_n565_), .D(mai_mai_n293_), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n625_), .B(mai_mai_n216_), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n394_), .B(mai_mai_n205_), .Y(mai_mai_n985_));
  AN2        m0957(.A(d), .B(c), .Y(mai_mai_n986_));
  NA2        m0958(.A(mai_mai_n986_), .B(mai_mai_n115_), .Y(mai_mai_n987_));
  NO4        m0959(.A(mai_mai_n987_), .B(mai_mai_n985_), .C(mai_mai_n172_), .D(mai_mai_n163_), .Y(mai_mai_n988_));
  NA2        m0960(.A(mai_mai_n482_), .B(c), .Y(mai_mai_n989_));
  NO4        m0961(.A(mai_mai_n982_), .B(mai_mai_n561_), .C(mai_mai_n989_), .D(mai_mai_n293_), .Y(mai_mai_n990_));
  AO210      m0962(.A0(mai_mai_n988_), .A1(mai_mai_n984_), .B0(mai_mai_n990_), .Y(mai_mai_n991_));
  OR4        m0963(.A(mai_mai_n991_), .B(mai_mai_n983_), .C(mai_mai_n980_), .D(mai_mai_n978_), .Y(mai_mai_n992_));
  NAi32      m0964(.An(f), .Bn(e), .C(c), .Y(mai_mai_n993_));
  NO2        m0965(.A(mai_mai_n993_), .B(mai_mai_n144_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n994_), .B(g), .Y(mai_mai_n995_));
  OR3        m0967(.A(mai_mai_n216_), .B(mai_mai_n172_), .C(mai_mai_n163_), .Y(mai_mai_n996_));
  NO2        m0968(.A(mai_mai_n996_), .B(mai_mai_n995_), .Y(mai_mai_n997_));
  NO2        m0969(.A(mai_mai_n989_), .B(mai_mai_n293_), .Y(mai_mai_n998_));
  NO2        m0970(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n590_), .B(mai_mai_n999_), .Y(mai_mai_n1000_));
  NOi21      m0972(.An(mai_mai_n998_), .B(mai_mai_n1000_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(mai_mai_n720_), .B(mai_mai_n111_), .Y(mai_mai_n1002_));
  NOi41      m0974(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1003_));
  NA2        m0975(.A(mai_mai_n1003_), .B(mai_mai_n1002_), .Y(mai_mai_n1004_));
  NO2        m0976(.A(mai_mai_n1004_), .B(mai_mai_n995_), .Y(mai_mai_n1005_));
  NA3        m0977(.A(k), .B(j), .C(i), .Y(mai_mai_n1006_));
  NO3        m0978(.A(mai_mai_n1006_), .B(mai_mai_n293_), .C(mai_mai_n91_), .Y(mai_mai_n1007_));
  OR3        m0979(.A(mai_mai_n1005_), .B(mai_mai_n1001_), .C(mai_mai_n997_), .Y(mai_mai_n1008_));
  NA3        m0980(.A(mai_mai_n452_), .B(mai_mai_n321_), .C(mai_mai_n56_), .Y(mai_mai_n1009_));
  NO2        m0981(.A(mai_mai_n1009_), .B(mai_mai_n1000_), .Y(mai_mai_n1010_));
  NO3        m0982(.A(mai_mai_n1009_), .B(mai_mai_n561_), .C(mai_mai_n433_), .Y(mai_mai_n1011_));
  NO2        m0983(.A(f), .B(c), .Y(mai_mai_n1012_));
  NOi21      m0984(.An(mai_mai_n1012_), .B(mai_mai_n425_), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n1013_), .B(mai_mai_n59_), .Y(mai_mai_n1014_));
  OR2        m0986(.A(k), .B(i), .Y(mai_mai_n1015_));
  NO3        m0987(.A(mai_mai_n1015_), .B(mai_mai_n235_), .C(l), .Y(mai_mai_n1016_));
  NOi31      m0988(.An(mai_mai_n1016_), .B(mai_mai_n1014_), .C(j), .Y(mai_mai_n1017_));
  OR3        m0989(.A(mai_mai_n1017_), .B(mai_mai_n1011_), .C(mai_mai_n1010_), .Y(mai_mai_n1018_));
  OR3        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1008_), .C(mai_mai_n992_), .Y(mai02));
  OR3        m0991(.A(n), .B(m), .C(i), .Y(mai_mai_n1020_));
  NOi31      m0992(.An(e), .B(d), .C(c), .Y(mai_mai_n1021_));
  AOI210     m0993(.A0(mai_mai_n1007_), .A1(mai_mai_n1021_), .B0(mai_mai_n983_), .Y(mai_mai_n1022_));
  AN3        m0994(.A(g), .B(f), .C(c), .Y(mai_mai_n1023_));
  NA2        m0995(.A(mai_mai_n1023_), .B(mai_mai_n452_), .Y(mai_mai_n1024_));
  OR2        m0996(.A(mai_mai_n1006_), .B(mai_mai_n293_), .Y(mai_mai_n1025_));
  OR2        m0997(.A(mai_mai_n1025_), .B(mai_mai_n1024_), .Y(mai_mai_n1026_));
  NO3        m0998(.A(mai_mai_n1009_), .B(mai_mai_n982_), .C(mai_mai_n561_), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n1027_), .B(mai_mai_n997_), .Y(mai_mai_n1028_));
  NA3        m1000(.A(l), .B(k), .C(j), .Y(mai_mai_n1029_));
  NA2        m1001(.A(i), .B(h), .Y(mai_mai_n1030_));
  NO3        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1029_), .C(mai_mai_n129_), .Y(mai_mai_n1031_));
  NO3        m1003(.A(mai_mai_n139_), .B(mai_mai_n275_), .C(mai_mai_n206_), .Y(mai_mai_n1032_));
  AOI210     m1004(.A0(mai_mai_n1032_), .A1(mai_mai_n1031_), .B0(mai_mai_n1001_), .Y(mai_mai_n1033_));
  NA3        m1005(.A(c), .B(b), .C(a), .Y(mai_mai_n1034_));
  NO3        m1006(.A(mai_mai_n1034_), .B(mai_mai_n853_), .C(mai_mai_n205_), .Y(mai_mai_n1035_));
  NO3        m1007(.A(mai_mai_n1006_), .B(mai_mai_n287_), .C(mai_mai_n49_), .Y(mai_mai_n1036_));
  AOI210     m1008(.A0(mai_mai_n1036_), .A1(mai_mai_n1035_), .B0(mai_mai_n1010_), .Y(mai_mai_n1037_));
  AN4        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1033_), .C(mai_mai_n1028_), .D(mai_mai_n1026_), .Y(mai_mai_n1038_));
  NO2        m1010(.A(mai_mai_n987_), .B(mai_mai_n985_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n1004_), .B(mai_mai_n996_), .Y(mai_mai_n1040_));
  AOI210     m1012(.A0(mai_mai_n1040_), .A1(mai_mai_n1039_), .B0(mai_mai_n978_), .Y(mai_mai_n1041_));
  NA3        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1038_), .C(mai_mai_n1022_), .Y(mai03));
  NO2        m1014(.A(mai_mai_n513_), .B(mai_mai_n566_), .Y(mai_mai_n1043_));
  INV        m1015(.A(mai_mai_n352_), .Y(mai_mai_n1044_));
  NO3        m1016(.A(mai_mai_n1044_), .B(mai_mai_n1043_), .C(mai_mai_n942_), .Y(mai_mai_n1045_));
  NOi31      m1017(.An(mai_mai_n762_), .B(mai_mai_n800_), .C(mai_mai_n673_), .Y(mai_mai_n1046_));
  OAI220     m1018(.A0(mai_mai_n1046_), .A1(mai_mai_n649_), .B0(mai_mai_n1045_), .B1(mai_mai_n562_), .Y(mai_mai_n1047_));
  NA4        m1019(.A(i), .B(mai_mai_n1021_), .C(mai_mai_n330_), .D(mai_mai_n321_), .Y(mai_mai_n1048_));
  OAI210     m1020(.A0(mai_mai_n776_), .A1(mai_mai_n402_), .B0(mai_mai_n1048_), .Y(mai_mai_n1049_));
  NOi31      m1021(.An(m), .B(n), .C(f), .Y(mai_mai_n1050_));
  NA2        m1022(.A(mai_mai_n1050_), .B(mai_mai_n51_), .Y(mai_mai_n1051_));
  AN2        m1023(.A(e), .B(c), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n1052_), .B(a), .Y(mai_mai_n1053_));
  OAI220     m1025(.A0(mai_mai_n1053_), .A1(mai_mai_n1051_), .B0(mai_mai_n836_), .B1(mai_mai_n408_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n495_), .B(l), .Y(mai_mai_n1055_));
  NOi31      m1027(.An(g), .B(mai_mai_n976_), .C(mai_mai_n1055_), .Y(mai_mai_n1056_));
  NO3        m1028(.A(mai_mai_n1056_), .B(mai_mai_n1054_), .C(mai_mai_n1049_), .Y(mai_mai_n1057_));
  NO2        m1029(.A(mai_mai_n275_), .B(a), .Y(mai_mai_n1058_));
  INV        m1030(.A(mai_mai_n983_), .Y(mai_mai_n1059_));
  NO2        m1031(.A(mai_mai_n1030_), .B(mai_mai_n469_), .Y(mai_mai_n1060_));
  NO2        m1032(.A(mai_mai_n88_), .B(g), .Y(mai_mai_n1061_));
  AOI210     m1033(.A0(mai_mai_n1061_), .A1(mai_mai_n1060_), .B0(mai_mai_n1016_), .Y(mai_mai_n1062_));
  OR2        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1014_), .Y(mai_mai_n1063_));
  NA3        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1059_), .C(mai_mai_n1057_), .Y(mai_mai_n1064_));
  NO4        m1036(.A(mai_mai_n1064_), .B(mai_mai_n1047_), .C(mai_mai_n778_), .D(mai_mai_n547_), .Y(mai_mai_n1065_));
  NA2        m1037(.A(c), .B(b), .Y(mai_mai_n1066_));
  NO2        m1038(.A(mai_mai_n661_), .B(mai_mai_n1066_), .Y(mai_mai_n1067_));
  OAI210     m1039(.A0(mai_mai_n817_), .A1(mai_mai_n792_), .B0(mai_mai_n396_), .Y(mai_mai_n1068_));
  NA2        m1040(.A(mai_mai_n1068_), .B(mai_mai_n1067_), .Y(mai_mai_n1069_));
  NAi21      m1041(.An(mai_mai_n403_), .B(mai_mai_n1067_), .Y(mai_mai_n1070_));
  OAI210     m1042(.A0(mai_mai_n530_), .A1(mai_mai_n39_), .B0(mai_mai_n1058_), .Y(mai_mai_n1071_));
  NA2        m1043(.A(mai_mai_n1071_), .B(mai_mai_n1070_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n253_), .B(mai_mai_n118_), .Y(mai_mai_n1073_));
  NA2        m1045(.A(mai_mai_n1073_), .B(g), .Y(mai_mai_n1074_));
  NAi21      m1046(.An(f), .B(d), .Y(mai_mai_n1075_));
  NO2        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1034_), .Y(mai_mai_n1076_));
  INV        m1048(.A(mai_mai_n1076_), .Y(mai_mai_n1077_));
  AOI210     m1049(.A0(mai_mai_n1074_), .A1(mai_mai_n279_), .B0(mai_mai_n1077_), .Y(mai_mai_n1078_));
  AOI210     m1050(.A0(mai_mai_n1078_), .A1(mai_mai_n112_), .B0(mai_mai_n1072_), .Y(mai_mai_n1079_));
  NA2        m1051(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n1080_));
  NO2        m1052(.A(mai_mai_n178_), .B(mai_mai_n229_), .Y(mai_mai_n1081_));
  NA2        m1053(.A(mai_mai_n1081_), .B(m), .Y(mai_mai_n1082_));
  NO2        m1054(.A(mai_mai_n1080_), .B(mai_mai_n1082_), .Y(mai_mai_n1083_));
  NA2        m1055(.A(mai_mai_n542_), .B(mai_mai_n393_), .Y(mai_mai_n1084_));
  NA2        m1056(.A(mai_mai_n155_), .B(mai_mai_n33_), .Y(mai_mai_n1085_));
  AOI210     m1057(.A0(mai_mai_n910_), .A1(mai_mai_n1085_), .B0(mai_mai_n206_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n1076_), .Y(mai_mai_n1087_));
  INV        m1059(.A(mai_mai_n904_), .Y(mai_mai_n1088_));
  NA3        m1060(.A(mai_mai_n1088_), .B(mai_mai_n1087_), .C(mai_mai_n1084_), .Y(mai_mai_n1089_));
  NO2        m1061(.A(mai_mai_n1089_), .B(mai_mai_n1083_), .Y(mai_mai_n1090_));
  NA4        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1079_), .C(mai_mai_n1069_), .D(mai_mai_n1065_), .Y(mai00));
  AOI210     m1063(.A0(mai_mai_n286_), .A1(mai_mai_n206_), .B0(mai_mai_n267_), .Y(mai_mai_n1092_));
  NO2        m1064(.A(mai_mai_n1092_), .B(mai_mai_n553_), .Y(mai_mai_n1093_));
  AOI210     m1065(.A0(mai_mai_n850_), .A1(mai_mai_n888_), .B0(mai_mai_n1049_), .Y(mai_mai_n1094_));
  NO3        m1066(.A(mai_mai_n1027_), .B(mai_mai_n904_), .C(mai_mai_n670_), .Y(mai_mai_n1095_));
  NA3        m1067(.A(mai_mai_n1095_), .B(mai_mai_n1094_), .C(mai_mai_n943_), .Y(mai_mai_n1096_));
  NA2        m1068(.A(mai_mai_n497_), .B(f), .Y(mai_mai_n1097_));
  OAI210     m1069(.A0(mai_mai_n950_), .A1(mai_mai_n40_), .B0(mai_mai_n605_), .Y(mai_mai_n1098_));
  NA3        m1070(.A(mai_mai_n1098_), .B(mai_mai_n250_), .C(n), .Y(mai_mai_n1099_));
  AOI210     m1071(.A0(mai_mai_n1099_), .A1(mai_mai_n1097_), .B0(mai_mai_n987_), .Y(mai_mai_n1100_));
  NO4        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1096_), .C(mai_mai_n1093_), .D(mai_mai_n1008_), .Y(mai_mai_n1101_));
  NA3        m1073(.A(mai_mai_n162_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1102_));
  NA3        m1074(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1103_));
  NOi31      m1075(.An(n), .B(m), .C(i), .Y(mai_mai_n1104_));
  NA3        m1076(.A(mai_mai_n1104_), .B(mai_mai_n608_), .C(mai_mai_n51_), .Y(mai_mai_n1105_));
  OAI210     m1077(.A0(mai_mai_n1103_), .A1(mai_mai_n1102_), .B0(mai_mai_n1105_), .Y(mai_mai_n1106_));
  NO2        m1078(.A(mai_mai_n1106_), .B(mai_mai_n867_), .Y(mai_mai_n1107_));
  NO4        m1079(.A(mai_mai_n472_), .B(mai_mai_n343_), .C(mai_mai_n1066_), .D(mai_mai_n59_), .Y(mai_mai_n1108_));
  NA3        m1080(.A(mai_mai_n366_), .B(mai_mai_n212_), .C(g), .Y(mai_mai_n1109_));
  OR2        m1081(.A(mai_mai_n1109_), .B(mai_mai_n1103_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(h), .B(g), .Y(mai_mai_n1111_));
  NA4        m1083(.A(mai_mai_n485_), .B(mai_mai_n452_), .C(mai_mai_n1111_), .D(mai_mai_n975_), .Y(mai_mai_n1112_));
  OAI220     m1084(.A0(mai_mai_n513_), .A1(mai_mai_n566_), .B0(mai_mai_n92_), .B1(mai_mai_n91_), .Y(mai_mai_n1113_));
  AOI220     m1085(.A0(mai_mai_n1113_), .A1(mai_mai_n519_), .B0(mai_mai_n892_), .B1(mai_mai_n552_), .Y(mai_mai_n1114_));
  AOI220     m1086(.A0(mai_mai_n304_), .A1(mai_mai_n239_), .B0(mai_mai_n173_), .B1(mai_mai_n146_), .Y(mai_mai_n1115_));
  NA4        m1087(.A(mai_mai_n1115_), .B(mai_mai_n1114_), .C(mai_mai_n1112_), .D(mai_mai_n1110_), .Y(mai_mai_n1116_));
  NO3        m1088(.A(mai_mai_n1116_), .B(mai_mai_n1108_), .C(mai_mai_n258_), .Y(mai_mai_n1117_));
  INV        m1089(.A(mai_mai_n309_), .Y(mai_mai_n1118_));
  AOI210     m1090(.A0(mai_mai_n239_), .A1(mai_mai_n335_), .B0(mai_mai_n554_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n1119_), .B(mai_mai_n1118_), .Y(mai_mai_n1120_));
  NO2        m1092(.A(mai_mai_n231_), .B(mai_mai_n177_), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n1121_), .B(mai_mai_n409_), .Y(mai_mai_n1122_));
  NA3        m1094(.A(mai_mai_n175_), .B(mai_mai_n111_), .C(g), .Y(mai_mai_n1123_));
  NA3        m1095(.A(mai_mai_n452_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1124_));
  NOi31      m1096(.An(mai_mai_n822_), .B(mai_mai_n1124_), .C(mai_mai_n1123_), .Y(mai_mai_n1125_));
  NAi31      m1097(.An(mai_mai_n179_), .B(mai_mai_n814_), .C(mai_mai_n452_), .Y(mai_mai_n1126_));
  NAi31      m1098(.An(mai_mai_n1125_), .B(mai_mai_n1126_), .C(mai_mai_n1122_), .Y(mai_mai_n1127_));
  NO2        m1099(.A(mai_mai_n266_), .B(mai_mai_n74_), .Y(mai_mai_n1128_));
  NO3        m1100(.A(mai_mai_n408_), .B(mai_mai_n788_), .C(n), .Y(mai_mai_n1129_));
  NA2        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1128_), .Y(mai_mai_n1130_));
  NAi31      m1102(.An(mai_mai_n990_), .B(mai_mai_n1130_), .C(mai_mai_n73_), .Y(mai_mai_n1131_));
  NO3        m1103(.A(mai_mai_n1131_), .B(mai_mai_n1127_), .C(mai_mai_n1120_), .Y(mai_mai_n1132_));
  AN3        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1117_), .C(mai_mai_n1107_), .Y(mai_mai_n1133_));
  NA3        m1105(.A(mai_mai_n1050_), .B(mai_mai_n570_), .C(mai_mai_n451_), .Y(mai_mai_n1134_));
  NA3        m1106(.A(mai_mai_n1134_), .B(mai_mai_n543_), .C(mai_mai_n233_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n1044_), .B(mai_mai_n519_), .Y(mai_mai_n1136_));
  NA4        m1108(.A(mai_mai_n608_), .B(mai_mai_n200_), .C(mai_mai_n212_), .D(mai_mai_n159_), .Y(mai_mai_n1137_));
  NA3        m1109(.A(mai_mai_n1137_), .B(mai_mai_n1136_), .C(mai_mai_n283_), .Y(mai_mai_n1138_));
  NA2        m1110(.A(mai_mai_n542_), .B(mai_mai_n393_), .Y(mai_mai_n1139_));
  OR4        m1111(.A(mai_mai_n987_), .B(mai_mai_n264_), .C(mai_mai_n214_), .D(e), .Y(mai_mai_n1140_));
  NO2        m1112(.A(mai_mai_n209_), .B(mai_mai_n206_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(n), .B(e), .Y(mai_mai_n1142_));
  NO2        m1114(.A(mai_mai_n1142_), .B(mai_mai_n144_), .Y(mai_mai_n1143_));
  AOI220     m1115(.A0(mai_mai_n1143_), .A1(mai_mai_n265_), .B0(mai_mai_n803_), .B1(mai_mai_n1141_), .Y(mai_mai_n1144_));
  OAI210     m1116(.A0(mai_mai_n344_), .A1(mai_mai_n298_), .B0(mai_mai_n431_), .Y(mai_mai_n1145_));
  NA4        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1144_), .C(mai_mai_n1140_), .D(mai_mai_n1139_), .Y(mai_mai_n1146_));
  AOI210     m1118(.A0(mai_mai_n1143_), .A1(mai_mai_n807_), .B0(mai_mai_n777_), .Y(mai_mai_n1147_));
  AOI220     m1119(.A0(mai_mai_n900_), .A1(mai_mai_n552_), .B0(mai_mai_n608_), .B1(mai_mai_n236_), .Y(mai_mai_n1148_));
  NO2        m1120(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1149_));
  NO3        m1121(.A(mai_mai_n987_), .B(mai_mai_n985_), .C(mai_mai_n686_), .Y(mai_mai_n1150_));
  INV        m1122(.A(mai_mai_n129_), .Y(mai_mai_n1151_));
  AN2        m1123(.A(mai_mai_n1151_), .B(mai_mai_n1032_), .Y(mai_mai_n1152_));
  OAI210     m1124(.A0(mai_mai_n1152_), .A1(mai_mai_n1150_), .B0(mai_mai_n1149_), .Y(mai_mai_n1153_));
  NA3        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1148_), .C(mai_mai_n1147_), .Y(mai_mai_n1154_));
  NO4        m1126(.A(mai_mai_n1154_), .B(mai_mai_n1146_), .C(mai_mai_n1138_), .D(mai_mai_n1135_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n793_), .B(mai_mai_n715_), .Y(mai_mai_n1156_));
  NA4        m1128(.A(mai_mai_n1156_), .B(mai_mai_n1155_), .C(mai_mai_n1133_), .D(mai_mai_n1101_), .Y(mai01));
  NO4        m1129(.A(mai_mai_n759_), .B(mai_mai_n751_), .C(mai_mai_n464_), .D(mai_mai_n273_), .Y(mai_mai_n1158_));
  NA2        m1130(.A(mai_mai_n377_), .B(i), .Y(mai_mai_n1159_));
  NA3        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1158_), .C(mai_mai_n965_), .Y(mai_mai_n1160_));
  NA2        m1132(.A(mai_mai_n535_), .B(mai_mai_n263_), .Y(mai_mai_n1161_));
  NA2        m1133(.A(mai_mai_n907_), .B(mai_mai_n1161_), .Y(mai_mai_n1162_));
  NA3        m1134(.A(mai_mai_n1162_), .B(mai_mai_n864_), .C(mai_mai_n320_), .Y(mai_mai_n1163_));
  OR2        m1135(.A(mai_mai_n620_), .B(mai_mai_n352_), .Y(mai_mai_n1164_));
  NAi41      m1136(.An(mai_mai_n158_), .B(mai_mai_n1164_), .C(mai_mai_n1137_), .D(mai_mai_n849_), .Y(mai_mai_n1165_));
  NO3        m1137(.A(mai_mai_n741_), .B(mai_mai_n632_), .C(mai_mai_n499_), .Y(mai_mai_n1166_));
  NA3        m1138(.A(mai_mai_n668_), .B(mai_mai_n97_), .C(mai_mai_n45_), .Y(mai_mai_n1167_));
  OA220      m1139(.A0(mai_mai_n1167_), .A1(mai_mai_n628_), .B0(mai_mai_n189_), .B1(mai_mai_n187_), .Y(mai_mai_n1168_));
  NA3        m1140(.A(mai_mai_n1168_), .B(mai_mai_n1166_), .C(mai_mai_n134_), .Y(mai_mai_n1169_));
  NO4        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1165_), .C(mai_mai_n1163_), .D(mai_mai_n1160_), .Y(mai_mai_n1170_));
  INV        m1142(.A(mai_mai_n1109_), .Y(mai_mai_n1171_));
  NA2        m1143(.A(mai_mai_n1171_), .B(mai_mai_n515_), .Y(mai_mai_n1172_));
  NA2        m1144(.A(mai_mai_n521_), .B(mai_mai_n379_), .Y(mai_mai_n1173_));
  NOi21      m1145(.An(mai_mai_n544_), .B(mai_mai_n557_), .Y(mai_mai_n1174_));
  NA2        m1146(.A(mai_mai_n1174_), .B(mai_mai_n1173_), .Y(mai_mai_n1175_));
  NA2        m1147(.A(mai_mai_n1175_), .B(mai_mai_n1172_), .Y(mai_mai_n1176_));
  NA2        m1148(.A(mai_mai_n272_), .B(mai_mai_n189_), .Y(mai_mai_n1177_));
  NA2        m1149(.A(mai_mai_n1177_), .B(mai_mai_n624_), .Y(mai_mai_n1178_));
  NO3        m1150(.A(mai_mai_n776_), .B(mai_mai_n198_), .C(mai_mai_n391_), .Y(mai_mai_n1179_));
  NO2        m1151(.A(mai_mai_n1179_), .B(mai_mai_n904_), .Y(mai_mai_n1180_));
  NA2        m1152(.A(mai_mai_n314_), .B(mai_mai_n633_), .Y(mai_mai_n1181_));
  NA4        m1153(.A(mai_mai_n1181_), .B(mai_mai_n1180_), .C(mai_mai_n1178_), .D(mai_mai_n744_), .Y(mai_mai_n1182_));
  NO3        m1154(.A(mai_mai_n1182_), .B(mai_mai_n567_), .C(mai_mai_n1176_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n492_), .B(mai_mai_n58_), .Y(mai_mai_n1184_));
  NO2        m1156(.A(mai_mai_n201_), .B(mai_mai_n110_), .Y(mai_mai_n1185_));
  NO2        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1106_), .Y(mai_mai_n1186_));
  NA3        m1158(.A(mai_mai_n1186_), .B(mai_mai_n1184_), .C(mai_mai_n714_), .Y(mai_mai_n1187_));
  NO3        m1159(.A(mai_mai_n80_), .B(mai_mai_n287_), .C(mai_mai_n45_), .Y(mai_mai_n1188_));
  NA2        m1160(.A(mai_mai_n1188_), .B(mai_mai_n534_), .Y(mai_mai_n1189_));
  INV        m1161(.A(mai_mai_n1189_), .Y(mai_mai_n1190_));
  OR2        m1162(.A(mai_mai_n1109_), .B(mai_mai_n1103_), .Y(mai_mai_n1191_));
  NO2        m1163(.A(mai_mai_n352_), .B(mai_mai_n72_), .Y(mai_mai_n1192_));
  INV        m1164(.A(mai_mai_n1192_), .Y(mai_mai_n1193_));
  NA2        m1165(.A(mai_mai_n1188_), .B(mai_mai_n768_), .Y(mai_mai_n1194_));
  NA4        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1193_), .C(mai_mai_n1191_), .D(mai_mai_n369_), .Y(mai_mai_n1195_));
  NO3        m1167(.A(mai_mai_n1195_), .B(mai_mai_n1190_), .C(mai_mai_n1187_), .Y(mai_mai_n1196_));
  NO2        m1168(.A(mai_mai_n128_), .B(mai_mai_n45_), .Y(mai_mai_n1197_));
  NO2        m1169(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1198_));
  AO220      m1170(.A0(mai_mai_n1198_), .A1(mai_mai_n585_), .B0(mai_mai_n1197_), .B1(mai_mai_n666_), .Y(mai_mai_n1199_));
  NA2        m1171(.A(mai_mai_n1199_), .B(mai_mai_n328_), .Y(mai_mai_n1200_));
  INV        m1172(.A(mai_mai_n132_), .Y(mai_mai_n1201_));
  NO3        m1173(.A(mai_mai_n1030_), .B(mai_mai_n172_), .C(mai_mai_n88_), .Y(mai_mai_n1202_));
  AOI220     m1174(.A0(mai_mai_n1202_), .A1(mai_mai_n1201_), .B0(mai_mai_n1188_), .B1(mai_mai_n918_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n1203_), .B(mai_mai_n1200_), .Y(mai_mai_n1204_));
  NO2        m1176(.A(mai_mai_n576_), .B(mai_mai_n575_), .Y(mai_mai_n1205_));
  NO4        m1177(.A(mai_mai_n1030_), .B(mai_mai_n1205_), .C(mai_mai_n170_), .D(mai_mai_n88_), .Y(mai_mai_n1206_));
  NO3        m1178(.A(mai_mai_n1206_), .B(mai_mai_n1204_), .C(mai_mai_n599_), .Y(mai_mai_n1207_));
  NA4        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1196_), .C(mai_mai_n1183_), .D(mai_mai_n1170_), .Y(mai06));
  NO2        m1180(.A(mai_mai_n392_), .B(mai_mai_n541_), .Y(mai_mai_n1209_));
  INV        m1181(.A(mai_mai_n692_), .Y(mai_mai_n1210_));
  OAI210     m1182(.A0(mai_mai_n1210_), .A1(mai_mai_n259_), .B0(mai_mai_n1209_), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n216_), .B(mai_mai_n101_), .Y(mai_mai_n1212_));
  OAI210     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n1202_), .B0(mai_mai_n365_), .Y(mai_mai_n1213_));
  NA2        m1185(.A(mai_mai_n1213_), .B(mai_mai_n1211_), .Y(mai_mai_n1214_));
  NO3        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1190_), .C(mai_mai_n249_), .Y(mai_mai_n1215_));
  NO2        m1187(.A(mai_mai_n287_), .B(mai_mai_n45_), .Y(mai_mai_n1216_));
  NA2        m1188(.A(mai_mai_n1216_), .B(mai_mai_n919_), .Y(mai_mai_n1217_));
  AOI210     m1189(.A0(mai_mai_n1216_), .A1(mai_mai_n538_), .B0(mai_mai_n1199_), .Y(mai_mai_n1218_));
  AOI210     m1190(.A0(mai_mai_n1218_), .A1(mai_mai_n1217_), .B0(mai_mai_n325_), .Y(mai_mai_n1219_));
  OAI210     m1191(.A0(mai_mai_n90_), .A1(mai_mai_n40_), .B0(mai_mai_n631_), .Y(mai_mai_n1220_));
  NA2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n602_), .Y(mai_mai_n1221_));
  NO2        m1193(.A(mai_mai_n502_), .B(mai_mai_n167_), .Y(mai_mai_n1222_));
  NO2        m1194(.A(mai_mai_n571_), .B(mai_mai_n1051_), .Y(mai_mai_n1223_));
  OAI210     m1195(.A0(mai_mai_n445_), .A1(mai_mai_n240_), .B0(mai_mai_n858_), .Y(mai_mai_n1224_));
  NO3        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1223_), .C(mai_mai_n1222_), .Y(mai_mai_n1225_));
  INV        m1197(.A(mai_mai_n567_), .Y(mai_mai_n1226_));
  NA3        m1198(.A(mai_mai_n1226_), .B(mai_mai_n1225_), .C(mai_mai_n1221_), .Y(mai_mai_n1227_));
  NO2        m1199(.A(mai_mai_n705_), .B(mai_mai_n350_), .Y(mai_mai_n1228_));
  NO3        m1200(.A(mai_mai_n633_), .B(mai_mai_n716_), .C(mai_mai_n595_), .Y(mai_mai_n1229_));
  NOi21      m1201(.An(mai_mai_n1228_), .B(mai_mai_n1229_), .Y(mai_mai_n1230_));
  AN2        m1202(.A(mai_mai_n900_), .B(mai_mai_n604_), .Y(mai_mai_n1231_));
  NO4        m1203(.A(mai_mai_n1231_), .B(mai_mai_n1230_), .C(mai_mai_n1227_), .D(mai_mai_n1219_), .Y(mai_mai_n1232_));
  NO2        m1204(.A(mai_mai_n758_), .B(mai_mai_n268_), .Y(mai_mai_n1233_));
  OAI220     m1205(.A0(mai_mai_n692_), .A1(mai_mai_n47_), .B0(mai_mai_n216_), .B1(mai_mai_n578_), .Y(mai_mai_n1234_));
  OAI210     m1206(.A0(mai_mai_n268_), .A1(c), .B0(mai_mai_n601_), .Y(mai_mai_n1235_));
  AOI220     m1207(.A0(mai_mai_n1235_), .A1(mai_mai_n1234_), .B0(mai_mai_n1233_), .B1(mai_mai_n259_), .Y(mai_mai_n1236_));
  OAI220     m1208(.A0(mai_mai_n658_), .A1(mai_mai_n240_), .B0(mai_mai_n498_), .B1(mai_mai_n502_), .Y(mai_mai_n1237_));
  INV        m1209(.A(k), .Y(mai_mai_n1238_));
  NO3        m1210(.A(mai_mai_n1238_), .B(mai_mai_n566_), .C(j), .Y(mai_mai_n1239_));
  NOi21      m1211(.An(mai_mai_n1239_), .B(mai_mai_n628_), .Y(mai_mai_n1240_));
  NO3        m1212(.A(mai_mai_n1240_), .B(mai_mai_n1237_), .C(mai_mai_n1054_), .Y(mai_mai_n1241_));
  NA3        m1213(.A(mai_mai_n1241_), .B(mai_mai_n1236_), .C(mai_mai_n1148_), .Y(mai_mai_n1242_));
  NO2        m1214(.A(mai_mai_n449_), .B(mai_mai_n378_), .Y(mai_mai_n1243_));
  OR3        m1215(.A(mai_mai_n1243_), .B(mai_mai_n740_), .C(mai_mai_n524_), .Y(mai_mai_n1244_));
  OR3        m1216(.A(mai_mai_n354_), .B(mai_mai_n216_), .C(mai_mai_n578_), .Y(mai_mai_n1245_));
  NA2        m1217(.A(mai_mai_n1239_), .B(mai_mai_n748_), .Y(mai_mai_n1246_));
  NA3        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1245_), .C(mai_mai_n1244_), .Y(mai_mai_n1247_));
  NA2        m1219(.A(mai_mai_n1228_), .B(mai_mai_n715_), .Y(mai_mai_n1248_));
  NO3        m1220(.A(mai_mai_n827_), .B(mai_mai_n488_), .C(mai_mai_n467_), .Y(mai_mai_n1249_));
  NA3        m1221(.A(mai_mai_n1249_), .B(mai_mai_n1248_), .C(mai_mai_n1194_), .Y(mai_mai_n1250_));
  NAi21      m1222(.An(j), .B(i), .Y(mai_mai_n1251_));
  NO4        m1223(.A(mai_mai_n1205_), .B(mai_mai_n1251_), .C(mai_mai_n425_), .D(mai_mai_n227_), .Y(mai_mai_n1252_));
  NO4        m1224(.A(mai_mai_n1252_), .B(mai_mai_n1250_), .C(mai_mai_n1247_), .D(mai_mai_n1242_), .Y(mai_mai_n1253_));
  NA4        m1225(.A(mai_mai_n1253_), .B(mai_mai_n1232_), .C(mai_mai_n1215_), .D(mai_mai_n1207_), .Y(mai07));
  NOi21      m1226(.An(j), .B(k), .Y(mai_mai_n1255_));
  NA4        m1227(.A(mai_mai_n175_), .B(mai_mai_n107_), .C(mai_mai_n1255_), .D(f), .Y(mai_mai_n1256_));
  NAi32      m1228(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1257_));
  NO3        m1229(.A(mai_mai_n1257_), .B(g), .C(f), .Y(mai_mai_n1258_));
  OAI210     m1230(.A0(mai_mai_n308_), .A1(mai_mai_n468_), .B0(mai_mai_n1258_), .Y(mai_mai_n1259_));
  NAi21      m1231(.An(f), .B(c), .Y(mai_mai_n1260_));
  OR2        m1232(.A(e), .B(d), .Y(mai_mai_n1261_));
  OAI220     m1233(.A0(mai_mai_n1261_), .A1(mai_mai_n1260_), .B0(k), .B1(mai_mai_n310_), .Y(mai_mai_n1262_));
  NA3        m1234(.A(mai_mai_n1262_), .B(mai_mai_n999_), .C(mai_mai_n175_), .Y(mai_mai_n1263_));
  NOi31      m1235(.An(n), .B(m), .C(b), .Y(mai_mai_n1264_));
  NO3        m1236(.A(mai_mai_n129_), .B(mai_mai_n433_), .C(h), .Y(mai_mai_n1265_));
  NA3        m1237(.A(mai_mai_n1263_), .B(mai_mai_n1259_), .C(mai_mai_n1256_), .Y(mai_mai_n1266_));
  NO2        m1238(.A(k), .B(i), .Y(mai_mai_n1267_));
  NA3        m1239(.A(mai_mai_n1267_), .B(mai_mai_n848_), .C(mai_mai_n175_), .Y(mai_mai_n1268_));
  NA2        m1240(.A(mai_mai_n88_), .B(mai_mai_n45_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n993_), .B(mai_mai_n425_), .Y(mai_mai_n1270_));
  NA3        m1242(.A(mai_mai_n1270_), .B(mai_mai_n1269_), .C(mai_mai_n206_), .Y(mai_mai_n1271_));
  NO2        m1243(.A(mai_mai_n1006_), .B(mai_mai_n293_), .Y(mai_mai_n1272_));
  NA2        m1244(.A(mai_mai_n525_), .B(mai_mai_n81_), .Y(mai_mai_n1273_));
  NA2        m1245(.A(mai_mai_n1149_), .B(mai_mai_n277_), .Y(mai_mai_n1274_));
  NA4        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1273_), .C(mai_mai_n1271_), .D(mai_mai_n1268_), .Y(mai_mai_n1275_));
  NO2        m1247(.A(mai_mai_n1275_), .B(mai_mai_n1266_), .Y(mai_mai_n1276_));
  NO3        m1248(.A(e), .B(d), .C(c), .Y(mai_mai_n1277_));
  NO2        m1249(.A(mai_mai_n129_), .B(mai_mai_n206_), .Y(mai_mai_n1278_));
  NA2        m1250(.A(mai_mai_n1278_), .B(mai_mai_n1277_), .Y(mai_mai_n1279_));
  INV        m1251(.A(mai_mai_n1279_), .Y(mai_mai_n1280_));
  NA3        m1252(.A(mai_mai_n655_), .B(mai_mai_n641_), .C(mai_mai_n111_), .Y(mai_mai_n1281_));
  NO2        m1253(.A(mai_mai_n1281_), .B(mai_mai_n45_), .Y(mai_mai_n1282_));
  NO2        m1254(.A(l), .B(k), .Y(mai_mai_n1283_));
  NOi41      m1255(.An(mai_mai_n529_), .B(mai_mai_n1283_), .C(mai_mai_n462_), .D(mai_mai_n425_), .Y(mai_mai_n1284_));
  NO3        m1256(.A(mai_mai_n425_), .B(d), .C(c), .Y(mai_mai_n1285_));
  NO3        m1257(.A(mai_mai_n1284_), .B(mai_mai_n1282_), .C(mai_mai_n1280_), .Y(mai_mai_n1286_));
  NO2        m1258(.A(mai_mai_n145_), .B(h), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n1015_), .B(l), .Y(mai_mai_n1288_));
  NO2        m1260(.A(g), .B(c), .Y(mai_mai_n1289_));
  NA3        m1261(.A(mai_mai_n1289_), .B(mai_mai_n139_), .C(mai_mai_n180_), .Y(mai_mai_n1290_));
  NO2        m1262(.A(mai_mai_n1290_), .B(mai_mai_n1288_), .Y(mai_mai_n1291_));
  NA2        m1263(.A(mai_mai_n1291_), .B(mai_mai_n175_), .Y(mai_mai_n1292_));
  NO2        m1264(.A(mai_mai_n436_), .B(a), .Y(mai_mai_n1293_));
  NA3        m1265(.A(mai_mai_n1293_), .B(mai_mai_n1432_), .C(mai_mai_n112_), .Y(mai_mai_n1294_));
  NO2        m1266(.A(i), .B(h), .Y(mai_mai_n1295_));
  NA2        m1267(.A(mai_mai_n1075_), .B(h), .Y(mai_mai_n1296_));
  NA2        m1268(.A(mai_mai_n135_), .B(mai_mai_n212_), .Y(mai_mai_n1297_));
  NO2        m1269(.A(mai_mai_n1297_), .B(mai_mai_n1296_), .Y(mai_mai_n1298_));
  NO2        m1270(.A(mai_mai_n712_), .B(mai_mai_n181_), .Y(mai_mai_n1299_));
  NOi31      m1271(.An(m), .B(n), .C(b), .Y(mai_mai_n1300_));
  NOi31      m1272(.An(f), .B(d), .C(c), .Y(mai_mai_n1301_));
  NA2        m1273(.A(mai_mai_n1301_), .B(mai_mai_n1300_), .Y(mai_mai_n1302_));
  INV        m1274(.A(mai_mai_n1302_), .Y(mai_mai_n1303_));
  NO3        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1299_), .C(mai_mai_n1298_), .Y(mai_mai_n1304_));
  NA2        m1276(.A(mai_mai_n1023_), .B(mai_mai_n452_), .Y(mai_mai_n1305_));
  NO4        m1277(.A(mai_mai_n1305_), .B(mai_mai_n1002_), .C(mai_mai_n425_), .D(mai_mai_n45_), .Y(mai_mai_n1306_));
  OAI210     m1278(.A0(mai_mai_n178_), .A1(mai_mai_n512_), .B0(mai_mai_n1003_), .Y(mai_mai_n1307_));
  NO3        m1279(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1308_));
  INV        m1280(.A(mai_mai_n1307_), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n1309_), .B(mai_mai_n1306_), .Y(mai_mai_n1310_));
  AN4        m1282(.A(mai_mai_n1310_), .B(mai_mai_n1304_), .C(mai_mai_n1294_), .D(mai_mai_n1292_), .Y(mai_mai_n1311_));
  NA2        m1283(.A(mai_mai_n1264_), .B(mai_mai_n362_), .Y(mai_mai_n1312_));
  NO2        m1284(.A(mai_mai_n1312_), .B(mai_mai_n984_), .Y(mai_mai_n1313_));
  NA2        m1285(.A(mai_mai_n1285_), .B(mai_mai_n207_), .Y(mai_mai_n1314_));
  NO2        m1286(.A(mai_mai_n181_), .B(b), .Y(mai_mai_n1315_));
  AOI220     m1287(.A0(mai_mai_n1104_), .A1(mai_mai_n1315_), .B0(mai_mai_n1031_), .B1(mai_mai_n1305_), .Y(mai_mai_n1316_));
  NAi31      m1288(.An(mai_mai_n1313_), .B(mai_mai_n1316_), .C(mai_mai_n1314_), .Y(mai_mai_n1317_));
  NO4        m1289(.A(mai_mai_n129_), .B(g), .C(f), .D(e), .Y(mai_mai_n1318_));
  NA3        m1290(.A(mai_mai_n1267_), .B(mai_mai_n278_), .C(h), .Y(mai_mai_n1319_));
  OR2        m1291(.A(e), .B(a), .Y(mai_mai_n1320_));
  NO2        m1292(.A(mai_mai_n1261_), .B(mai_mai_n1260_), .Y(mai_mai_n1321_));
  AOI210     m1293(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1321_), .Y(mai_mai_n1322_));
  NO2        m1294(.A(mai_mai_n1322_), .B(mai_mai_n1020_), .Y(mai_mai_n1323_));
  OR3        m1295(.A(mai_mai_n524_), .B(mai_mai_n523_), .C(mai_mai_n111_), .Y(mai_mai_n1324_));
  NA2        m1296(.A(mai_mai_n1050_), .B(mai_mai_n391_), .Y(mai_mai_n1325_));
  NO2        m1297(.A(mai_mai_n1325_), .B(mai_mai_n418_), .Y(mai_mai_n1326_));
  AN2        m1298(.A(mai_mai_n1326_), .B(mai_mai_n115_), .Y(mai_mai_n1327_));
  NO3        m1299(.A(mai_mai_n1327_), .B(mai_mai_n1323_), .C(mai_mai_n1317_), .Y(mai_mai_n1328_));
  NA4        m1300(.A(mai_mai_n1328_), .B(mai_mai_n1311_), .C(mai_mai_n1286_), .D(mai_mai_n1276_), .Y(mai_mai_n1329_));
  NO2        m1301(.A(mai_mai_n1066_), .B(mai_mai_n109_), .Y(mai_mai_n1330_));
  NA2        m1302(.A(mai_mai_n362_), .B(mai_mai_n56_), .Y(mai_mai_n1331_));
  NA2        m1303(.A(mai_mai_n207_), .B(mai_mai_n175_), .Y(mai_mai_n1332_));
  AOI210     m1304(.A0(mai_mai_n1332_), .A1(mai_mai_n1123_), .B0(mai_mai_n1331_), .Y(mai_mai_n1333_));
  NO2        m1305(.A(mai_mai_n374_), .B(j), .Y(mai_mai_n1334_));
  NA3        m1306(.A(mai_mai_n1308_), .B(mai_mai_n1261_), .C(mai_mai_n1050_), .Y(mai_mai_n1335_));
  NAi41      m1307(.An(mai_mai_n1295_), .B(mai_mai_n1013_), .C(mai_mai_n163_), .D(mai_mai_n148_), .Y(mai_mai_n1336_));
  NA2        m1308(.A(mai_mai_n1336_), .B(mai_mai_n1335_), .Y(mai_mai_n1337_));
  NA3        m1309(.A(g), .B(mai_mai_n1334_), .C(mai_mai_n155_), .Y(mai_mai_n1338_));
  INV        m1310(.A(mai_mai_n1338_), .Y(mai_mai_n1339_));
  NO3        m1311(.A(mai_mai_n705_), .B(mai_mai_n170_), .C(mai_mai_n394_), .Y(mai_mai_n1340_));
  NO3        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1339_), .C(mai_mai_n1337_), .Y(mai_mai_n1341_));
  OR2        m1313(.A(n), .B(i), .Y(mai_mai_n1342_));
  OAI210     m1314(.A0(mai_mai_n1342_), .A1(mai_mai_n1012_), .B0(mai_mai_n49_), .Y(mai_mai_n1343_));
  AOI220     m1315(.A0(mai_mai_n1343_), .A1(mai_mai_n1111_), .B0(mai_mai_n781_), .B1(mai_mai_n188_), .Y(mai_mai_n1344_));
  INV        m1316(.A(mai_mai_n1344_), .Y(mai_mai_n1345_));
  OAI220     m1317(.A0(mai_mai_n625_), .A1(g), .B0(mai_mai_n216_), .B1(c), .Y(mai_mai_n1346_));
  AOI210     m1318(.A0(mai_mai_n1315_), .A1(mai_mai_n41_), .B0(mai_mai_n1346_), .Y(mai_mai_n1347_));
  NO2        m1319(.A(mai_mai_n129_), .B(l), .Y(mai_mai_n1348_));
  NO2        m1320(.A(mai_mai_n216_), .B(k), .Y(mai_mai_n1349_));
  OAI210     m1321(.A0(mai_mai_n1349_), .A1(mai_mai_n1295_), .B0(mai_mai_n1348_), .Y(mai_mai_n1350_));
  OAI220     m1322(.A0(mai_mai_n1350_), .A1(mai_mai_n31_), .B0(mai_mai_n1347_), .B1(mai_mai_n172_), .Y(mai_mai_n1351_));
  NO3        m1323(.A(mai_mai_n1324_), .B(mai_mai_n452_), .C(mai_mai_n340_), .Y(mai_mai_n1352_));
  NO3        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1351_), .C(mai_mai_n1345_), .Y(mai_mai_n1353_));
  NO3        m1325(.A(mai_mai_n1034_), .B(mai_mai_n1261_), .C(mai_mai_n49_), .Y(mai_mai_n1354_));
  NA3        m1326(.A(mai_mai_n1330_), .B(mai_mai_n452_), .C(f), .Y(mai_mai_n1355_));
  NA2        m1327(.A(mai_mai_n175_), .B(mai_mai_n111_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n1255_), .B(mai_mai_n42_), .Y(mai_mai_n1357_));
  AOI210     m1329(.A0(mai_mai_n112_), .A1(mai_mai_n40_), .B0(mai_mai_n1357_), .Y(mai_mai_n1358_));
  NO2        m1330(.A(mai_mai_n1358_), .B(mai_mai_n1355_), .Y(mai_mai_n1359_));
  NOi21      m1331(.An(d), .B(f), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n1293_), .B(mai_mai_n1357_), .Y(mai_mai_n1361_));
  INV        m1333(.A(mai_mai_n1361_), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1362_), .B(mai_mai_n1359_), .Y(mai_mai_n1363_));
  NA4        m1335(.A(mai_mai_n1363_), .B(mai_mai_n1353_), .C(mai_mai_n1341_), .D(mai_mai_n1431_), .Y(mai_mai_n1364_));
  NO3        m1336(.A(mai_mai_n1023_), .B(mai_mai_n1012_), .C(mai_mai_n40_), .Y(mai_mai_n1365_));
  NO2        m1337(.A(mai_mai_n452_), .B(mai_mai_n287_), .Y(mai_mai_n1366_));
  OAI210     m1338(.A0(mai_mai_n1366_), .A1(mai_mai_n1365_), .B0(mai_mai_n1272_), .Y(mai_mai_n1367_));
  OAI210     m1339(.A0(mai_mai_n1318_), .A1(mai_mai_n1264_), .B0(mai_mai_n833_), .Y(mai_mai_n1368_));
  NO2        m1340(.A(mai_mai_n981_), .B(mai_mai_n129_), .Y(mai_mai_n1369_));
  NA2        m1341(.A(mai_mai_n1369_), .B(mai_mai_n584_), .Y(mai_mai_n1370_));
  NA3        m1342(.A(mai_mai_n1370_), .B(mai_mai_n1368_), .C(mai_mai_n1367_), .Y(mai_mai_n1371_));
  NA2        m1343(.A(mai_mai_n1289_), .B(mai_mai_n1360_), .Y(mai_mai_n1372_));
  NO2        m1344(.A(mai_mai_n1372_), .B(m), .Y(mai_mai_n1373_));
  NO2        m1345(.A(mai_mai_n149_), .B(mai_mai_n177_), .Y(mai_mai_n1374_));
  OAI210     m1346(.A0(mai_mai_n1374_), .A1(mai_mai_n109_), .B0(mai_mai_n1300_), .Y(mai_mai_n1375_));
  INV        m1347(.A(mai_mai_n1375_), .Y(mai_mai_n1376_));
  NO3        m1348(.A(mai_mai_n1376_), .B(mai_mai_n1373_), .C(mai_mai_n1371_), .Y(mai_mai_n1377_));
  NO2        m1349(.A(mai_mai_n1260_), .B(e), .Y(mai_mai_n1378_));
  NA2        m1350(.A(mai_mai_n1378_), .B(mai_mai_n389_), .Y(mai_mai_n1379_));
  NA2        m1351(.A(mai_mai_n1061_), .B(mai_mai_n591_), .Y(mai_mai_n1380_));
  OR3        m1352(.A(mai_mai_n1349_), .B(mai_mai_n1149_), .C(mai_mai_n129_), .Y(mai_mai_n1381_));
  OAI220     m1353(.A0(mai_mai_n1381_), .A1(mai_mai_n1379_), .B0(mai_mai_n1380_), .B1(mai_mai_n427_), .Y(mai_mai_n1382_));
  INV        m1354(.A(mai_mai_n1382_), .Y(mai_mai_n1383_));
  NO2        m1355(.A(mai_mai_n177_), .B(c), .Y(mai_mai_n1384_));
  OAI210     m1356(.A0(mai_mai_n1384_), .A1(mai_mai_n1378_), .B0(mai_mai_n175_), .Y(mai_mai_n1385_));
  AOI220     m1357(.A0(mai_mai_n1385_), .A1(mai_mai_n1014_), .B0(mai_mai_n517_), .B1(mai_mai_n350_), .Y(mai_mai_n1386_));
  NA2        m1358(.A(mai_mai_n523_), .B(g), .Y(mai_mai_n1387_));
  AOI210     m1359(.A0(mai_mai_n1387_), .A1(mai_mai_n1285_), .B0(mai_mai_n1354_), .Y(mai_mai_n1388_));
  NO2        m1360(.A(mai_mai_n1320_), .B(f), .Y(mai_mai_n1389_));
  AOI210     m1361(.A0(mai_mai_n1061_), .A1(a), .B0(mai_mai_n1389_), .Y(mai_mai_n1390_));
  OAI220     m1362(.A0(mai_mai_n1390_), .A1(mai_mai_n69_), .B0(mai_mai_n1388_), .B1(mai_mai_n205_), .Y(mai_mai_n1391_));
  AOI210     m1363(.A0(mai_mai_n853_), .A1(mai_mai_n399_), .B0(mai_mai_n103_), .Y(mai_mai_n1392_));
  NA2        m1364(.A(mai_mai_n1389_), .B(mai_mai_n1269_), .Y(mai_mai_n1393_));
  OAI220     m1365(.A0(mai_mai_n1393_), .A1(mai_mai_n49_), .B0(mai_mai_n1392_), .B1(mai_mai_n170_), .Y(mai_mai_n1394_));
  NA4        m1366(.A(mai_mai_n1032_), .B(mai_mai_n1029_), .C(mai_mai_n212_), .D(mai_mai_n68_), .Y(mai_mai_n1395_));
  NA2        m1367(.A(mai_mai_n1265_), .B(mai_mai_n178_), .Y(mai_mai_n1396_));
  NO2        m1368(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1397_));
  OAI210     m1369(.A0(mai_mai_n1320_), .A1(mai_mai_n816_), .B0(mai_mai_n468_), .Y(mai_mai_n1398_));
  OAI210     m1370(.A0(mai_mai_n1398_), .A1(mai_mai_n1035_), .B0(mai_mai_n1397_), .Y(mai_mai_n1399_));
  NO2        m1371(.A(m), .B(i), .Y(mai_mai_n1400_));
  BUFFER     m1372(.A(mai_mai_n1400_), .Y(mai_mai_n1401_));
  NA2        m1373(.A(mai_mai_n1401_), .B(mai_mai_n1287_), .Y(mai_mai_n1402_));
  NA4        m1374(.A(mai_mai_n1402_), .B(mai_mai_n1399_), .C(mai_mai_n1396_), .D(mai_mai_n1395_), .Y(mai_mai_n1403_));
  NO4        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1394_), .C(mai_mai_n1391_), .D(mai_mai_n1386_), .Y(mai_mai_n1404_));
  NA3        m1376(.A(mai_mai_n1404_), .B(mai_mai_n1383_), .C(mai_mai_n1377_), .Y(mai_mai_n1405_));
  NA3        m1377(.A(mai_mai_n906_), .B(mai_mai_n135_), .C(mai_mai_n46_), .Y(mai_mai_n1406_));
  AOI210     m1378(.A0(mai_mai_n146_), .A1(c), .B0(mai_mai_n1406_), .Y(mai_mai_n1407_));
  INV        m1379(.A(mai_mai_n1407_), .Y(mai_mai_n1408_));
  AOI210     m1380(.A0(mai_mai_n153_), .A1(mai_mai_n56_), .B0(mai_mai_n1378_), .Y(mai_mai_n1409_));
  NO2        m1381(.A(mai_mai_n1409_), .B(mai_mai_n1356_), .Y(mai_mai_n1410_));
  INV        m1382(.A(mai_mai_n1410_), .Y(mai_mai_n1411_));
  NO2        m1383(.A(mai_mai_n1355_), .B(mai_mai_n69_), .Y(mai_mai_n1412_));
  NA2        m1384(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1413_));
  NO2        m1385(.A(mai_mai_n1267_), .B(mai_mai_n117_), .Y(mai_mai_n1414_));
  OAI220     m1386(.A0(mai_mai_n1414_), .A1(mai_mai_n1312_), .B0(mai_mai_n1325_), .B1(mai_mai_n1413_), .Y(mai_mai_n1415_));
  NO2        m1387(.A(mai_mai_n1415_), .B(mai_mai_n1412_), .Y(mai_mai_n1416_));
  NA3        m1388(.A(mai_mai_n1416_), .B(mai_mai_n1411_), .C(mai_mai_n1408_), .Y(mai_mai_n1417_));
  OR4        m1389(.A(mai_mai_n1417_), .B(mai_mai_n1405_), .C(mai_mai_n1364_), .D(mai_mai_n1329_), .Y(mai04));
  NOi31      m1390(.An(mai_mai_n1318_), .B(mai_mai_n1319_), .C(mai_mai_n987_), .Y(mai_mai_n1419_));
  INV        m1391(.A(mai_mai_n781_), .Y(mai_mai_n1420_));
  NO3        m1392(.A(mai_mai_n1420_), .B(mai_mai_n976_), .C(mai_mai_n469_), .Y(mai_mai_n1421_));
  OR3        m1393(.A(mai_mai_n1421_), .B(mai_mai_n1419_), .C(mai_mai_n1005_), .Y(mai_mai_n1422_));
  NO2        m1394(.A(mai_mai_n1269_), .B(mai_mai_n91_), .Y(mai_mai_n1423_));
  AOI210     m1395(.A0(mai_mai_n1423_), .A1(mai_mai_n998_), .B0(mai_mai_n1125_), .Y(mai_mai_n1424_));
  NA2        m1396(.A(mai_mai_n1424_), .B(mai_mai_n1153_), .Y(mai_mai_n1425_));
  NO4        m1397(.A(mai_mai_n1425_), .B(mai_mai_n1422_), .C(mai_mai_n1011_), .D(mai_mai_n992_), .Y(mai_mai_n1426_));
  NA4        m1398(.A(mai_mai_n1426_), .B(mai_mai_n1063_), .C(mai_mai_n1048_), .D(mai_mai_n1038_), .Y(mai05));
  INV        m1399(.A(mai_mai_n567_), .Y(mai_mai_n1430_));
  INV        m1400(.A(mai_mai_n1333_), .Y(mai_mai_n1431_));
  INV        m1401(.A(i), .Y(mai_mai_n1432_));
  INV        m1402(.A(mai_mai_n560_), .Y(mai_mai_n1433_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA2        u0031(.A(g), .B(men_men_n59_), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NA2        u0033(.A(l), .B(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi21      u0042(.An(e), .B(h), .Y(men_men_n71_));
  NAi41      u0043(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n73_));
  INV        u0045(.A(m), .Y(men_men_n74_));
  NOi21      u0046(.An(k), .B(l), .Y(men_men_n75_));
  AN4        u0047(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n76_));
  NOi31      u0048(.An(h), .B(g), .C(f), .Y(men_men_n77_));
  NOi32      u0049(.An(h), .Bn(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n73_), .B(men_men_n64_), .Y(men_men_n79_));
  INV        u0051(.A(n), .Y(men_men_n80_));
  NOi32      u0052(.An(e), .Bn(b), .C(d), .Y(men_men_n81_));
  NA2        u0053(.A(men_men_n81_), .B(men_men_n80_), .Y(men_men_n82_));
  INV        u0054(.A(j), .Y(men_men_n83_));
  AN3        u0055(.A(m), .B(k), .C(i), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n83_), .C(g), .Y(men_men_n85_));
  NO2        u0057(.A(men_men_n85_), .B(f), .Y(men_men_n86_));
  NAi32      u0058(.An(g), .Bn(f), .C(h), .Y(men_men_n87_));
  NAi31      u0059(.An(j), .B(m), .C(l), .Y(men_men_n88_));
  NA2        u0060(.A(m), .B(l), .Y(men_men_n89_));
  NAi31      u0061(.An(k), .B(j), .C(g), .Y(men_men_n90_));
  NO3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(f), .Y(men_men_n91_));
  AN2        u0063(.A(j), .B(g), .Y(men_men_n92_));
  NOi32      u0064(.An(m), .Bn(l), .C(i), .Y(men_men_n93_));
  NOi21      u0065(.An(g), .B(i), .Y(men_men_n94_));
  NOi32      u0066(.An(m), .Bn(j), .C(k), .Y(men_men_n95_));
  AOI220     u0067(.A0(men_men_n95_), .A1(men_men_n94_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n96_));
  NO2        u0068(.A(men_men_n96_), .B(f), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n91_), .C(men_men_n86_), .Y(men_men_n98_));
  NAi41      u0070(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n99_));
  AN2        u0071(.A(e), .B(b), .Y(men_men_n100_));
  NOi21      u0072(.An(i), .B(h), .Y(men_men_n101_));
  INV        u0073(.A(a), .Y(men_men_n102_));
  NA2        u0074(.A(men_men_n100_), .B(men_men_n102_), .Y(men_men_n103_));
  INV        u0075(.A(l), .Y(men_men_n104_));
  NOi21      u0076(.An(m), .B(n), .Y(men_men_n105_));
  AN2        u0077(.A(k), .B(h), .Y(men_men_n106_));
  INV        u0078(.A(b), .Y(men_men_n107_));
  NA2        u0079(.A(l), .B(j), .Y(men_men_n108_));
  AN2        u0080(.A(k), .B(i), .Y(men_men_n109_));
  NA2        u0081(.A(men_men_n109_), .B(men_men_n108_), .Y(men_men_n110_));
  NA2        u0082(.A(g), .B(e), .Y(men_men_n111_));
  NOi32      u0083(.An(c), .Bn(a), .C(d), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n112_), .B(men_men_n105_), .Y(men_men_n113_));
  NO4        u0085(.A(men_men_n113_), .B(men_men_n111_), .C(men_men_n110_), .D(men_men_n107_), .Y(men_men_n114_));
  INV        u0086(.A(men_men_n114_), .Y(men_men_n115_));
  OAI210     u0087(.A0(men_men_n98_), .A1(men_men_n82_), .B0(men_men_n115_), .Y(men_men_n116_));
  NOi31      u0088(.An(k), .B(m), .C(j), .Y(men_men_n117_));
  NA3        u0089(.A(men_men_n117_), .B(men_men_n77_), .C(men_men_n76_), .Y(men_men_n118_));
  NOi31      u0090(.An(k), .B(m), .C(i), .Y(men_men_n119_));
  NA3        u0091(.A(men_men_n119_), .B(men_men_n78_), .C(men_men_n76_), .Y(men_men_n120_));
  NA2        u0092(.A(men_men_n120_), .B(men_men_n118_), .Y(men_men_n121_));
  NOi32      u0093(.An(f), .Bn(b), .C(e), .Y(men_men_n122_));
  NAi21      u0094(.An(g), .B(h), .Y(men_men_n123_));
  NAi21      u0095(.An(m), .B(n), .Y(men_men_n124_));
  NAi21      u0096(.An(j), .B(k), .Y(men_men_n125_));
  NO3        u0097(.A(men_men_n125_), .B(men_men_n124_), .C(men_men_n123_), .Y(men_men_n126_));
  NAi41      u0098(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n127_));
  NAi31      u0099(.An(j), .B(k), .C(h), .Y(men_men_n128_));
  NO3        u0100(.A(men_men_n128_), .B(men_men_n127_), .C(men_men_n124_), .Y(men_men_n129_));
  AOI210     u0101(.A0(men_men_n126_), .A1(men_men_n122_), .B0(men_men_n129_), .Y(men_men_n130_));
  NO2        u0102(.A(k), .B(j), .Y(men_men_n131_));
  AN2        u0103(.A(k), .B(j), .Y(men_men_n132_));
  NAi21      u0104(.An(c), .B(b), .Y(men_men_n133_));
  NA2        u0105(.A(f), .B(d), .Y(men_men_n134_));
  NAi31      u0106(.An(f), .B(e), .C(b), .Y(men_men_n135_));
  NA2        u0107(.A(d), .B(b), .Y(men_men_n136_));
  NAi21      u0108(.An(e), .B(f), .Y(men_men_n137_));
  NO2        u0109(.A(men_men_n137_), .B(men_men_n136_), .Y(men_men_n138_));
  NA2        u0110(.A(b), .B(a), .Y(men_men_n139_));
  NAi21      u0111(.An(c), .B(d), .Y(men_men_n140_));
  NAi31      u0112(.An(l), .B(k), .C(h), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n124_), .B(men_men_n141_), .Y(men_men_n142_));
  NA2        u0114(.A(men_men_n142_), .B(men_men_n138_), .Y(men_men_n143_));
  NAi31      u0115(.An(men_men_n121_), .B(men_men_n143_), .C(men_men_n130_), .Y(men_men_n144_));
  NAi31      u0116(.An(e), .B(f), .C(b), .Y(men_men_n145_));
  NOi21      u0117(.An(g), .B(d), .Y(men_men_n146_));
  NO2        u0118(.A(men_men_n146_), .B(men_men_n145_), .Y(men_men_n147_));
  NOi21      u0119(.An(h), .B(i), .Y(men_men_n148_));
  NOi21      u0120(.An(k), .B(m), .Y(men_men_n149_));
  NA3        u0121(.A(men_men_n149_), .B(men_men_n148_), .C(n), .Y(men_men_n150_));
  NOi21      u0122(.An(h), .B(g), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n152_));
  NA2        u0124(.A(men_men_n152_), .B(men_men_n151_), .Y(men_men_n153_));
  NAi31      u0125(.An(l), .B(j), .C(h), .Y(men_men_n154_));
  NO2        u0126(.A(men_men_n154_), .B(men_men_n49_), .Y(men_men_n155_));
  NA2        u0127(.A(men_men_n155_), .B(men_men_n67_), .Y(men_men_n156_));
  NOi32      u0128(.An(n), .Bn(k), .C(m), .Y(men_men_n157_));
  NA2        u0129(.A(l), .B(i), .Y(men_men_n158_));
  NA2        u0130(.A(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  OAI210     u0131(.A0(men_men_n159_), .A1(men_men_n153_), .B0(men_men_n156_), .Y(men_men_n160_));
  NAi31      u0132(.An(d), .B(f), .C(c), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(c), .Y(men_men_n162_));
  NA2        u0134(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  NA2        u0135(.A(j), .B(h), .Y(men_men_n164_));
  OR3        u0136(.A(n), .B(m), .C(k), .Y(men_men_n165_));
  NO2        u0137(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  NAi32      u0138(.An(m), .Bn(k), .C(n), .Y(men_men_n167_));
  NO2        u0139(.A(men_men_n167_), .B(men_men_n164_), .Y(men_men_n168_));
  AOI220     u0140(.A0(men_men_n168_), .A1(men_men_n147_), .B0(men_men_n166_), .B1(men_men_n163_), .Y(men_men_n169_));
  NO2        u0141(.A(n), .B(m), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n50_), .Y(men_men_n171_));
  NAi21      u0143(.An(f), .B(e), .Y(men_men_n172_));
  NA2        u0144(.A(d), .B(c), .Y(men_men_n173_));
  NO2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NOi21      u0146(.An(men_men_n174_), .B(men_men_n171_), .Y(men_men_n175_));
  NAi21      u0147(.An(d), .B(c), .Y(men_men_n176_));
  NAi31      u0148(.An(m), .B(n), .C(b), .Y(men_men_n177_));
  NA2        u0149(.A(k), .B(i), .Y(men_men_n178_));
  NAi21      u0150(.An(h), .B(f), .Y(men_men_n179_));
  NO2        u0151(.A(men_men_n179_), .B(men_men_n178_), .Y(men_men_n180_));
  NO2        u0152(.A(men_men_n177_), .B(men_men_n140_), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  NOi32      u0154(.An(f), .Bn(c), .C(d), .Y(men_men_n183_));
  NOi32      u0155(.An(f), .Bn(c), .C(e), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NO3        u0157(.A(n), .B(m), .C(j), .Y(men_men_n186_));
  NA2        u0158(.A(men_men_n186_), .B(men_men_n106_), .Y(men_men_n187_));
  AO210      u0159(.A0(men_men_n187_), .A1(men_men_n171_), .B0(men_men_n185_), .Y(men_men_n188_));
  NAi41      u0160(.An(men_men_n175_), .B(men_men_n188_), .C(men_men_n182_), .D(men_men_n169_), .Y(men_men_n189_));
  OR3        u0161(.A(men_men_n189_), .B(men_men_n160_), .C(men_men_n144_), .Y(men_men_n190_));
  NO4        u0162(.A(men_men_n190_), .B(men_men_n116_), .C(men_men_n79_), .D(men_men_n55_), .Y(men_men_n191_));
  NA3        u0163(.A(m), .B(men_men_n104_), .C(j), .Y(men_men_n192_));
  NAi31      u0164(.An(n), .B(h), .C(g), .Y(men_men_n193_));
  NO2        u0165(.A(men_men_n193_), .B(men_men_n192_), .Y(men_men_n194_));
  NOi32      u0166(.An(m), .Bn(k), .C(l), .Y(men_men_n195_));
  NA3        u0167(.A(men_men_n195_), .B(men_men_n83_), .C(g), .Y(men_men_n196_));
  NO2        u0168(.A(men_men_n196_), .B(n), .Y(men_men_n197_));
  AN2        u0169(.A(i), .B(g), .Y(men_men_n198_));
  NA3        u0170(.A(men_men_n75_), .B(men_men_n198_), .C(men_men_n105_), .Y(men_men_n199_));
  INV        u0171(.A(men_men_n199_), .Y(men_men_n200_));
  NO3        u0172(.A(men_men_n200_), .B(men_men_n197_), .C(men_men_n194_), .Y(men_men_n201_));
  NAi41      u0173(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n202_));
  INV        u0174(.A(men_men_n202_), .Y(men_men_n203_));
  INV        u0175(.A(f), .Y(men_men_n204_));
  INV        u0176(.A(g), .Y(men_men_n205_));
  NOi31      u0177(.An(i), .B(j), .C(h), .Y(men_men_n206_));
  NOi21      u0178(.An(l), .B(m), .Y(men_men_n207_));
  NA2        u0179(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NO3        u0180(.A(men_men_n208_), .B(men_men_n205_), .C(men_men_n204_), .Y(men_men_n209_));
  NA2        u0181(.A(men_men_n209_), .B(men_men_n203_), .Y(men_men_n210_));
  OAI210     u0182(.A0(men_men_n201_), .A1(men_men_n32_), .B0(men_men_n210_), .Y(men_men_n211_));
  NOi21      u0183(.An(n), .B(m), .Y(men_men_n212_));
  NOi32      u0184(.An(l), .Bn(i), .C(j), .Y(men_men_n213_));
  NA2        u0185(.A(men_men_n213_), .B(men_men_n212_), .Y(men_men_n214_));
  NAi21      u0186(.An(j), .B(h), .Y(men_men_n215_));
  XN2        u0187(.A(i), .B(h), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NOi31      u0189(.An(k), .B(n), .C(m), .Y(men_men_n218_));
  NOi31      u0190(.An(men_men_n218_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n217_), .Y(men_men_n220_));
  NAi31      u0192(.An(f), .B(e), .C(c), .Y(men_men_n221_));
  NO4        u0193(.A(men_men_n221_), .B(men_men_n165_), .C(men_men_n164_), .D(men_men_n59_), .Y(men_men_n222_));
  NA4        u0194(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n223_));
  NAi32      u0195(.An(m), .Bn(i), .C(k), .Y(men_men_n224_));
  NO3        u0196(.A(men_men_n224_), .B(men_men_n87_), .C(men_men_n223_), .Y(men_men_n225_));
  INV        u0197(.A(k), .Y(men_men_n226_));
  NO2        u0198(.A(men_men_n225_), .B(men_men_n222_), .Y(men_men_n227_));
  NAi21      u0199(.An(n), .B(a), .Y(men_men_n228_));
  NO2        u0200(.A(men_men_n228_), .B(men_men_n136_), .Y(men_men_n229_));
  NAi41      u0201(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n230_));
  NO2        u0202(.A(men_men_n230_), .B(e), .Y(men_men_n231_));
  NO3        u0203(.A(men_men_n137_), .B(men_men_n90_), .C(men_men_n89_), .Y(men_men_n232_));
  OAI210     u0204(.A0(men_men_n232_), .A1(men_men_n231_), .B0(men_men_n229_), .Y(men_men_n233_));
  AN3        u0205(.A(men_men_n233_), .B(men_men_n227_), .C(men_men_n220_), .Y(men_men_n234_));
  OR2        u0206(.A(h), .B(g), .Y(men_men_n235_));
  NO2        u0207(.A(men_men_n235_), .B(men_men_n99_), .Y(men_men_n236_));
  NA2        u0208(.A(men_men_n236_), .B(men_men_n122_), .Y(men_men_n237_));
  NA2        u0209(.A(men_men_n149_), .B(men_men_n101_), .Y(men_men_n238_));
  NO2        u0210(.A(n), .B(a), .Y(men_men_n239_));
  NAi31      u0211(.An(men_men_n230_), .B(men_men_n239_), .C(men_men_n100_), .Y(men_men_n240_));
  NAi21      u0212(.An(h), .B(i), .Y(men_men_n241_));
  NA2        u0213(.A(men_men_n170_), .B(k), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n242_), .B(men_men_n241_), .Y(men_men_n243_));
  NA2        u0215(.A(men_men_n243_), .B(men_men_n183_), .Y(men_men_n244_));
  NA3        u0216(.A(men_men_n244_), .B(men_men_n240_), .C(men_men_n237_), .Y(men_men_n245_));
  NOi21      u0217(.An(g), .B(e), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n247_));
  NA2        u0219(.A(men_men_n247_), .B(men_men_n246_), .Y(men_men_n248_));
  NOi32      u0220(.An(l), .Bn(j), .C(i), .Y(men_men_n249_));
  AOI210     u0221(.A0(men_men_n75_), .A1(men_men_n83_), .B0(men_men_n249_), .Y(men_men_n250_));
  NO2        u0222(.A(men_men_n241_), .B(men_men_n44_), .Y(men_men_n251_));
  NAi21      u0223(.An(f), .B(g), .Y(men_men_n252_));
  NO2        u0224(.A(men_men_n252_), .B(men_men_n65_), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n69_), .B(men_men_n108_), .Y(men_men_n254_));
  AOI220     u0226(.A0(men_men_n254_), .A1(men_men_n253_), .B0(men_men_n251_), .B1(men_men_n67_), .Y(men_men_n255_));
  OAI210     u0227(.A0(men_men_n250_), .A1(men_men_n248_), .B0(men_men_n255_), .Y(men_men_n256_));
  NO3        u0228(.A(men_men_n125_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n257_));
  NOi41      u0229(.An(men_men_n234_), .B(men_men_n256_), .C(men_men_n245_), .D(men_men_n211_), .Y(men_men_n258_));
  NO4        u0230(.A(men_men_n194_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n103_), .Y(men_men_n260_));
  NAi21      u0232(.An(h), .B(g), .Y(men_men_n261_));
  OR4        u0233(.A(men_men_n261_), .B(men_men_n1468_), .C(men_men_n214_), .D(e), .Y(men_men_n262_));
  NAi31      u0234(.An(g), .B(k), .C(h), .Y(men_men_n263_));
  NO3        u0235(.A(men_men_n124_), .B(men_men_n263_), .C(l), .Y(men_men_n264_));
  NAi31      u0236(.An(e), .B(d), .C(a), .Y(men_men_n265_));
  NA2        u0237(.A(men_men_n264_), .B(men_men_n122_), .Y(men_men_n266_));
  NA2        u0238(.A(men_men_n266_), .B(men_men_n262_), .Y(men_men_n267_));
  NA3        u0239(.A(men_men_n149_), .B(men_men_n148_), .C(men_men_n80_), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n268_), .B(men_men_n185_), .Y(men_men_n269_));
  INV        u0241(.A(men_men_n269_), .Y(men_men_n270_));
  NA3        u0242(.A(e), .B(c), .C(b), .Y(men_men_n271_));
  NO2        u0243(.A(men_men_n60_), .B(men_men_n271_), .Y(men_men_n272_));
  NAi32      u0244(.An(k), .Bn(i), .C(j), .Y(men_men_n273_));
  NAi31      u0245(.An(h), .B(l), .C(i), .Y(men_men_n274_));
  NA3        u0246(.A(men_men_n274_), .B(men_men_n273_), .C(men_men_n154_), .Y(men_men_n275_));
  NOi21      u0247(.An(men_men_n275_), .B(men_men_n49_), .Y(men_men_n276_));
  OAI210     u0248(.A0(men_men_n253_), .A1(men_men_n272_), .B0(men_men_n276_), .Y(men_men_n277_));
  NAi21      u0249(.An(l), .B(k), .Y(men_men_n278_));
  NO2        u0250(.A(men_men_n278_), .B(men_men_n49_), .Y(men_men_n279_));
  NOi21      u0251(.An(l), .B(j), .Y(men_men_n280_));
  NA2        u0252(.A(men_men_n151_), .B(men_men_n280_), .Y(men_men_n281_));
  NA3        u0253(.A(men_men_n109_), .B(men_men_n108_), .C(g), .Y(men_men_n282_));
  OR3        u0254(.A(men_men_n72_), .B(men_men_n74_), .C(e), .Y(men_men_n283_));
  AOI210     u0255(.A0(men_men_n282_), .A1(men_men_n281_), .B0(men_men_n283_), .Y(men_men_n284_));
  INV        u0256(.A(men_men_n284_), .Y(men_men_n285_));
  NAi32      u0257(.An(j), .Bn(h), .C(i), .Y(men_men_n286_));
  NAi21      u0258(.An(m), .B(l), .Y(men_men_n287_));
  NO3        u0259(.A(men_men_n287_), .B(men_men_n286_), .C(men_men_n80_), .Y(men_men_n288_));
  NA2        u0260(.A(h), .B(g), .Y(men_men_n289_));
  NA2        u0261(.A(men_men_n157_), .B(men_men_n45_), .Y(men_men_n290_));
  NO2        u0262(.A(men_men_n290_), .B(men_men_n289_), .Y(men_men_n291_));
  OAI210     u0263(.A0(men_men_n291_), .A1(men_men_n288_), .B0(men_men_n152_), .Y(men_men_n292_));
  NA4        u0264(.A(men_men_n292_), .B(men_men_n285_), .C(men_men_n277_), .D(men_men_n270_), .Y(men_men_n293_));
  NO2        u0265(.A(men_men_n135_), .B(d), .Y(men_men_n294_));
  NA2        u0266(.A(men_men_n294_), .B(men_men_n53_), .Y(men_men_n295_));
  NAi32      u0267(.An(n), .Bn(m), .C(l), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n296_), .B(men_men_n286_), .Y(men_men_n297_));
  NA2        u0269(.A(men_men_n297_), .B(men_men_n174_), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n113_), .B(men_men_n107_), .Y(men_men_n299_));
  NAi31      u0271(.An(k), .B(l), .C(j), .Y(men_men_n300_));
  OAI210     u0272(.A0(men_men_n278_), .A1(j), .B0(men_men_n300_), .Y(men_men_n301_));
  NOi21      u0273(.An(men_men_n301_), .B(men_men_n111_), .Y(men_men_n302_));
  NA2        u0274(.A(men_men_n302_), .B(men_men_n299_), .Y(men_men_n303_));
  NA3        u0275(.A(men_men_n303_), .B(men_men_n298_), .C(men_men_n295_), .Y(men_men_n304_));
  NO4        u0276(.A(men_men_n304_), .B(men_men_n293_), .C(men_men_n267_), .D(men_men_n260_), .Y(men_men_n305_));
  NA2        u0277(.A(men_men_n243_), .B(men_men_n184_), .Y(men_men_n306_));
  NAi21      u0278(.An(m), .B(k), .Y(men_men_n307_));
  NAi41      u0279(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n308_));
  NAi31      u0280(.An(i), .B(l), .C(h), .Y(men_men_n309_));
  NA2        u0281(.A(e), .B(c), .Y(men_men_n310_));
  NO3        u0282(.A(men_men_n310_), .B(n), .C(d), .Y(men_men_n311_));
  NOi21      u0283(.An(f), .B(h), .Y(men_men_n312_));
  NA2        u0284(.A(men_men_n312_), .B(men_men_n109_), .Y(men_men_n313_));
  NO2        u0285(.A(men_men_n313_), .B(men_men_n205_), .Y(men_men_n314_));
  NAi31      u0286(.An(d), .B(e), .C(b), .Y(men_men_n315_));
  NO2        u0287(.A(men_men_n124_), .B(men_men_n315_), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n316_), .B(men_men_n314_), .Y(men_men_n317_));
  NA2        u0289(.A(men_men_n317_), .B(men_men_n306_), .Y(men_men_n318_));
  NO4        u0290(.A(men_men_n308_), .B(m), .C(men_men_n71_), .D(men_men_n205_), .Y(men_men_n319_));
  NA2        u0291(.A(men_men_n239_), .B(men_men_n100_), .Y(men_men_n320_));
  OR2        u0292(.A(men_men_n320_), .B(men_men_n196_), .Y(men_men_n321_));
  NOi31      u0293(.An(l), .B(n), .C(m), .Y(men_men_n322_));
  NAi21      u0294(.An(men_men_n319_), .B(men_men_n321_), .Y(men_men_n323_));
  NAi32      u0295(.An(m), .Bn(j), .C(k), .Y(men_men_n324_));
  NAi41      u0296(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n325_));
  NA2        u0297(.A(men_men_n202_), .B(men_men_n325_), .Y(men_men_n326_));
  NOi31      u0298(.An(j), .B(m), .C(k), .Y(men_men_n327_));
  NO2        u0299(.A(men_men_n117_), .B(men_men_n327_), .Y(men_men_n328_));
  AN3        u0300(.A(h), .B(g), .C(f), .Y(men_men_n329_));
  NAi31      u0301(.An(men_men_n328_), .B(men_men_n329_), .C(men_men_n326_), .Y(men_men_n330_));
  NOi32      u0302(.An(m), .Bn(j), .C(l), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n331_), .B(men_men_n93_), .Y(men_men_n332_));
  NO2        u0304(.A(men_men_n287_), .B(men_men_n286_), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n208_), .B(g), .Y(men_men_n334_));
  NO2        u0306(.A(men_men_n145_), .B(men_men_n80_), .Y(men_men_n335_));
  NA2        u0307(.A(men_men_n335_), .B(men_men_n334_), .Y(men_men_n336_));
  INV        u0308(.A(men_men_n224_), .Y(men_men_n337_));
  NA3        u0309(.A(men_men_n337_), .B(men_men_n329_), .C(men_men_n203_), .Y(men_men_n338_));
  NA3        u0310(.A(men_men_n338_), .B(men_men_n336_), .C(men_men_n330_), .Y(men_men_n339_));
  NA3        u0311(.A(h), .B(g), .C(f), .Y(men_men_n340_));
  NA2        u0312(.A(men_men_n151_), .B(e), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n341_), .B(men_men_n41_), .Y(men_men_n342_));
  NA2        u0314(.A(men_men_n342_), .B(men_men_n299_), .Y(men_men_n343_));
  NOi32      u0315(.An(j), .Bn(g), .C(i), .Y(men_men_n344_));
  NA3        u0316(.A(men_men_n344_), .B(men_men_n278_), .C(men_men_n105_), .Y(men_men_n345_));
  AO210      u0317(.A0(men_men_n103_), .A1(men_men_n32_), .B0(men_men_n345_), .Y(men_men_n346_));
  NOi32      u0318(.An(e), .Bn(b), .C(a), .Y(men_men_n347_));
  AN2        u0319(.A(l), .B(j), .Y(men_men_n348_));
  NA2        u0320(.A(men_men_n199_), .B(men_men_n35_), .Y(men_men_n349_));
  NA2        u0321(.A(men_men_n349_), .B(men_men_n347_), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n315_), .B(n), .Y(men_men_n351_));
  NA2        u0323(.A(men_men_n198_), .B(k), .Y(men_men_n352_));
  NA3        u0324(.A(m), .B(men_men_n104_), .C(men_men_n204_), .Y(men_men_n353_));
  NO2        u0325(.A(men_men_n353_), .B(men_men_n352_), .Y(men_men_n354_));
  NAi41      u0326(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n355_));
  NA2        u0327(.A(men_men_n51_), .B(men_men_n105_), .Y(men_men_n356_));
  NO2        u0328(.A(men_men_n356_), .B(men_men_n355_), .Y(men_men_n357_));
  AOI220     u0329(.A0(men_men_n357_), .A1(b), .B0(men_men_n354_), .B1(men_men_n351_), .Y(men_men_n358_));
  NA4        u0330(.A(men_men_n358_), .B(men_men_n350_), .C(men_men_n346_), .D(men_men_n343_), .Y(men_men_n359_));
  NO4        u0331(.A(men_men_n359_), .B(men_men_n339_), .C(men_men_n323_), .D(men_men_n318_), .Y(men_men_n360_));
  NA4        u0332(.A(men_men_n360_), .B(men_men_n305_), .C(men_men_n258_), .D(men_men_n191_), .Y(men10));
  NA3        u0333(.A(m), .B(k), .C(i), .Y(men_men_n362_));
  NO3        u0334(.A(men_men_n362_), .B(j), .C(men_men_n205_), .Y(men_men_n363_));
  NOi21      u0335(.An(e), .B(f), .Y(men_men_n364_));
  NO4        u0336(.A(men_men_n140_), .B(men_men_n364_), .C(n), .D(men_men_n102_), .Y(men_men_n365_));
  NAi31      u0337(.An(b), .B(f), .C(c), .Y(men_men_n366_));
  INV        u0338(.A(men_men_n366_), .Y(men_men_n367_));
  NOi32      u0339(.An(k), .Bn(h), .C(j), .Y(men_men_n368_));
  NA2        u0340(.A(men_men_n368_), .B(men_men_n212_), .Y(men_men_n369_));
  NA2        u0341(.A(men_men_n150_), .B(men_men_n369_), .Y(men_men_n370_));
  AOI220     u0342(.A0(men_men_n370_), .A1(men_men_n367_), .B0(men_men_n365_), .B1(men_men_n363_), .Y(men_men_n371_));
  AN2        u0343(.A(j), .B(h), .Y(men_men_n372_));
  NO3        u0344(.A(n), .B(m), .C(k), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n373_), .B(men_men_n372_), .Y(men_men_n374_));
  NO3        u0346(.A(men_men_n374_), .B(men_men_n140_), .C(men_men_n204_), .Y(men_men_n375_));
  OR2        u0347(.A(m), .B(k), .Y(men_men_n376_));
  NO2        u0348(.A(men_men_n164_), .B(men_men_n376_), .Y(men_men_n377_));
  NA4        u0349(.A(n), .B(f), .C(c), .D(men_men_n107_), .Y(men_men_n378_));
  NOi21      u0350(.An(men_men_n377_), .B(men_men_n378_), .Y(men_men_n379_));
  NOi32      u0351(.An(d), .Bn(a), .C(c), .Y(men_men_n380_));
  NA2        u0352(.A(men_men_n380_), .B(men_men_n172_), .Y(men_men_n381_));
  NAi21      u0353(.An(i), .B(g), .Y(men_men_n382_));
  NAi31      u0354(.An(k), .B(m), .C(j), .Y(men_men_n383_));
  NO2        u0355(.A(men_men_n379_), .B(men_men_n375_), .Y(men_men_n384_));
  NO2        u0356(.A(men_men_n378_), .B(men_men_n287_), .Y(men_men_n385_));
  NOi32      u0357(.An(f), .Bn(d), .C(c), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n384_), .B(men_men_n371_), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n59_), .B(men_men_n107_), .Y(men_men_n388_));
  NA2        u0360(.A(men_men_n239_), .B(men_men_n388_), .Y(men_men_n389_));
  INV        u0361(.A(e), .Y(men_men_n390_));
  NA2        u0362(.A(men_men_n46_), .B(e), .Y(men_men_n391_));
  OAI220     u0363(.A0(men_men_n391_), .A1(men_men_n192_), .B0(men_men_n196_), .B1(men_men_n390_), .Y(men_men_n392_));
  AN2        u0364(.A(g), .B(e), .Y(men_men_n393_));
  NA3        u0365(.A(men_men_n393_), .B(men_men_n195_), .C(i), .Y(men_men_n394_));
  INV        u0366(.A(men_men_n394_), .Y(men_men_n395_));
  NO2        u0367(.A(men_men_n96_), .B(men_men_n390_), .Y(men_men_n396_));
  NO3        u0368(.A(men_men_n396_), .B(men_men_n395_), .C(men_men_n392_), .Y(men_men_n397_));
  NOi32      u0369(.An(h), .Bn(e), .C(g), .Y(men_men_n398_));
  NA3        u0370(.A(men_men_n398_), .B(men_men_n280_), .C(m), .Y(men_men_n399_));
  NOi21      u0371(.An(g), .B(h), .Y(men_men_n400_));
  AN3        u0372(.A(m), .B(l), .C(i), .Y(men_men_n401_));
  NA3        u0373(.A(men_men_n401_), .B(men_men_n400_), .C(e), .Y(men_men_n402_));
  AN3        u0374(.A(h), .B(g), .C(e), .Y(men_men_n403_));
  NA2        u0375(.A(men_men_n403_), .B(men_men_n93_), .Y(men_men_n404_));
  AN3        u0376(.A(men_men_n404_), .B(men_men_n402_), .C(men_men_n399_), .Y(men_men_n405_));
  AOI210     u0377(.A0(men_men_n405_), .A1(men_men_n397_), .B0(men_men_n389_), .Y(men_men_n406_));
  NA3        u0378(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n407_));
  NO2        u0379(.A(men_men_n407_), .B(men_men_n389_), .Y(men_men_n408_));
  NA3        u0380(.A(men_men_n380_), .B(men_men_n172_), .C(men_men_n80_), .Y(men_men_n409_));
  NAi31      u0381(.An(b), .B(c), .C(a), .Y(men_men_n410_));
  NO2        u0382(.A(men_men_n410_), .B(n), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n51_), .B(m), .Y(men_men_n412_));
  NO2        u0384(.A(men_men_n412_), .B(men_men_n137_), .Y(men_men_n413_));
  NA2        u0385(.A(men_men_n413_), .B(men_men_n411_), .Y(men_men_n414_));
  INV        u0386(.A(men_men_n414_), .Y(men_men_n415_));
  NO4        u0387(.A(men_men_n415_), .B(men_men_n408_), .C(men_men_n406_), .D(men_men_n387_), .Y(men_men_n416_));
  NA2        u0388(.A(i), .B(g), .Y(men_men_n417_));
  NO3        u0389(.A(men_men_n265_), .B(men_men_n417_), .C(c), .Y(men_men_n418_));
  NOi21      u0390(.An(a), .B(n), .Y(men_men_n419_));
  NOi21      u0391(.An(d), .B(c), .Y(men_men_n420_));
  NA2        u0392(.A(men_men_n420_), .B(men_men_n419_), .Y(men_men_n421_));
  NA3        u0393(.A(i), .B(g), .C(f), .Y(men_men_n422_));
  NA2        u0394(.A(men_men_n418_), .B(men_men_n279_), .Y(men_men_n423_));
  OR2        u0395(.A(n), .B(m), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n424_), .B(men_men_n141_), .Y(men_men_n425_));
  NO2        u0397(.A(men_men_n173_), .B(men_men_n137_), .Y(men_men_n426_));
  OAI210     u0398(.A0(men_men_n425_), .A1(men_men_n166_), .B0(men_men_n426_), .Y(men_men_n427_));
  INV        u0399(.A(men_men_n356_), .Y(men_men_n428_));
  NA3        u0400(.A(men_men_n428_), .B(men_men_n347_), .C(d), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n410_), .B(men_men_n49_), .Y(men_men_n430_));
  NAi21      u0402(.An(k), .B(j), .Y(men_men_n431_));
  NAi21      u0403(.An(e), .B(d), .Y(men_men_n432_));
  INV        u0404(.A(men_men_n432_), .Y(men_men_n433_));
  NO2        u0405(.A(men_men_n242_), .B(men_men_n204_), .Y(men_men_n434_));
  NA3        u0406(.A(men_men_n434_), .B(men_men_n433_), .C(men_men_n217_), .Y(men_men_n435_));
  NA3        u0407(.A(men_men_n435_), .B(men_men_n429_), .C(men_men_n427_), .Y(men_men_n436_));
  NOi31      u0408(.An(n), .B(m), .C(k), .Y(men_men_n437_));
  AOI220     u0409(.A0(men_men_n437_), .A1(men_men_n372_), .B0(men_men_n212_), .B1(men_men_n50_), .Y(men_men_n438_));
  NAi31      u0410(.An(g), .B(f), .C(c), .Y(men_men_n439_));
  OR3        u0411(.A(men_men_n439_), .B(men_men_n438_), .C(e), .Y(men_men_n440_));
  NA2        u0412(.A(men_men_n440_), .B(men_men_n298_), .Y(men_men_n441_));
  NOi41      u0413(.An(men_men_n423_), .B(men_men_n441_), .C(men_men_n436_), .D(men_men_n256_), .Y(men_men_n442_));
  NOi32      u0414(.An(c), .Bn(a), .C(b), .Y(men_men_n443_));
  NA2        u0415(.A(men_men_n443_), .B(men_men_n105_), .Y(men_men_n444_));
  INV        u0416(.A(men_men_n263_), .Y(men_men_n445_));
  AN2        u0417(.A(e), .B(d), .Y(men_men_n446_));
  NA2        u0418(.A(men_men_n446_), .B(men_men_n445_), .Y(men_men_n447_));
  NO2        u0419(.A(men_men_n123_), .B(men_men_n41_), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n66_), .B(e), .Y(men_men_n449_));
  NOi31      u0421(.An(j), .B(k), .C(i), .Y(men_men_n450_));
  NOi21      u0422(.An(men_men_n154_), .B(men_men_n450_), .Y(men_men_n451_));
  NA4        u0423(.A(men_men_n309_), .B(men_men_n451_), .C(men_men_n250_), .D(men_men_n110_), .Y(men_men_n452_));
  NA2        u0424(.A(men_men_n452_), .B(men_men_n449_), .Y(men_men_n453_));
  AOI210     u0425(.A0(men_men_n453_), .A1(men_men_n447_), .B0(men_men_n444_), .Y(men_men_n454_));
  NO2        u0426(.A(men_men_n200_), .B(men_men_n197_), .Y(men_men_n455_));
  NOi21      u0427(.An(a), .B(b), .Y(men_men_n456_));
  NA3        u0428(.A(e), .B(d), .C(c), .Y(men_men_n457_));
  NAi21      u0429(.An(men_men_n457_), .B(men_men_n456_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n409_), .B(men_men_n196_), .Y(men_men_n459_));
  NOi21      u0431(.An(men_men_n458_), .B(men_men_n459_), .Y(men_men_n460_));
  AOI210     u0432(.A0(men_men_n259_), .A1(men_men_n455_), .B0(men_men_n460_), .Y(men_men_n461_));
  NO4        u0433(.A(men_men_n179_), .B(men_men_n99_), .C(men_men_n56_), .D(b), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n367_), .B(men_men_n142_), .Y(men_men_n463_));
  OR2        u0435(.A(k), .B(j), .Y(men_men_n464_));
  NA2        u0436(.A(l), .B(k), .Y(men_men_n465_));
  NA2        u0437(.A(men_men_n120_), .B(men_men_n118_), .Y(men_men_n466_));
  NA2        u0438(.A(men_men_n380_), .B(men_men_n105_), .Y(men_men_n467_));
  NO4        u0439(.A(men_men_n467_), .B(men_men_n90_), .C(men_men_n104_), .D(e), .Y(men_men_n468_));
  NO3        u0440(.A(men_men_n409_), .B(men_men_n88_), .C(men_men_n123_), .Y(men_men_n469_));
  NO3        u0441(.A(men_men_n469_), .B(men_men_n468_), .C(men_men_n466_), .Y(men_men_n470_));
  NA2        u0442(.A(men_men_n470_), .B(men_men_n463_), .Y(men_men_n471_));
  NO4        u0443(.A(men_men_n471_), .B(men_men_n462_), .C(men_men_n461_), .D(men_men_n454_), .Y(men_men_n472_));
  NA2        u0444(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n473_));
  NAi31      u0445(.An(j), .B(l), .C(i), .Y(men_men_n474_));
  OAI210     u0446(.A0(men_men_n474_), .A1(men_men_n124_), .B0(men_men_n99_), .Y(men_men_n475_));
  NO3        u0447(.A(men_men_n381_), .B(men_men_n332_), .C(men_men_n193_), .Y(men_men_n476_));
  NO2        u0448(.A(men_men_n381_), .B(men_men_n356_), .Y(men_men_n477_));
  NO3        u0449(.A(men_men_n477_), .B(men_men_n476_), .C(men_men_n175_), .Y(men_men_n478_));
  NA3        u0450(.A(men_men_n478_), .B(men_men_n473_), .C(men_men_n234_), .Y(men_men_n479_));
  OAI210     u0451(.A0(men_men_n119_), .A1(men_men_n117_), .B0(n), .Y(men_men_n480_));
  NO2        u0452(.A(men_men_n480_), .B(men_men_n123_), .Y(men_men_n481_));
  OR2        u0453(.A(men_men_n288_), .B(men_men_n236_), .Y(men_men_n482_));
  OA210      u0454(.A0(men_men_n482_), .A1(men_men_n481_), .B0(men_men_n184_), .Y(men_men_n483_));
  XO2        u0455(.A(i), .B(h), .Y(men_men_n484_));
  NA3        u0456(.A(men_men_n484_), .B(men_men_n149_), .C(n), .Y(men_men_n485_));
  NAi41      u0457(.An(men_men_n288_), .B(men_men_n485_), .C(men_men_n438_), .D(men_men_n369_), .Y(men_men_n486_));
  NOi32      u0458(.An(men_men_n486_), .Bn(men_men_n449_), .C(men_men_n1468_), .Y(men_men_n487_));
  NAi31      u0459(.An(c), .B(f), .C(d), .Y(men_men_n488_));
  AOI210     u0460(.A0(men_men_n268_), .A1(men_men_n187_), .B0(men_men_n488_), .Y(men_men_n489_));
  INV        u0461(.A(men_men_n489_), .Y(men_men_n490_));
  NA2        u0462(.A(men_men_n218_), .B(men_men_n101_), .Y(men_men_n491_));
  AOI210     u0463(.A0(men_men_n491_), .A1(men_men_n171_), .B0(men_men_n488_), .Y(men_men_n492_));
  AOI210     u0464(.A0(men_men_n345_), .A1(men_men_n35_), .B0(men_men_n458_), .Y(men_men_n493_));
  NO2        u0465(.A(men_men_n493_), .B(men_men_n492_), .Y(men_men_n494_));
  AO220      u0466(.A0(men_men_n276_), .A1(men_men_n253_), .B0(men_men_n155_), .B1(men_men_n67_), .Y(men_men_n495_));
  NA3        u0467(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n496_));
  NO2        u0468(.A(men_men_n496_), .B(men_men_n421_), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n497_), .B(men_men_n284_), .Y(men_men_n498_));
  NAi41      u0470(.An(men_men_n495_), .B(men_men_n498_), .C(men_men_n494_), .D(men_men_n490_), .Y(men_men_n499_));
  NO4        u0471(.A(men_men_n499_), .B(men_men_n487_), .C(men_men_n483_), .D(men_men_n479_), .Y(men_men_n500_));
  NA4        u0472(.A(men_men_n500_), .B(men_men_n472_), .C(men_men_n442_), .D(men_men_n416_), .Y(men11));
  NO2        u0473(.A(men_men_n72_), .B(f), .Y(men_men_n502_));
  NA2        u0474(.A(j), .B(g), .Y(men_men_n503_));
  NAi31      u0475(.An(i), .B(m), .C(l), .Y(men_men_n504_));
  NA3        u0476(.A(m), .B(k), .C(j), .Y(men_men_n505_));
  OAI220     u0477(.A0(men_men_n505_), .A1(men_men_n123_), .B0(men_men_n504_), .B1(men_men_n503_), .Y(men_men_n506_));
  NA2        u0478(.A(men_men_n506_), .B(men_men_n502_), .Y(men_men_n507_));
  NOi32      u0479(.An(e), .Bn(b), .C(f), .Y(men_men_n508_));
  NA2        u0480(.A(men_men_n249_), .B(men_men_n105_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n46_), .B(j), .Y(men_men_n510_));
  NO2        u0482(.A(men_men_n510_), .B(men_men_n290_), .Y(men_men_n511_));
  NAi31      u0483(.An(d), .B(e), .C(a), .Y(men_men_n512_));
  NO2        u0484(.A(men_men_n512_), .B(n), .Y(men_men_n513_));
  AOI220     u0485(.A0(men_men_n513_), .A1(men_men_n97_), .B0(men_men_n511_), .B1(men_men_n508_), .Y(men_men_n514_));
  NAi41      u0486(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n515_));
  AN2        u0487(.A(men_men_n515_), .B(men_men_n355_), .Y(men_men_n516_));
  AOI210     u0488(.A0(men_men_n516_), .A1(men_men_n381_), .B0(men_men_n261_), .Y(men_men_n517_));
  NA2        u0489(.A(j), .B(i), .Y(men_men_n518_));
  NAi31      u0490(.An(n), .B(m), .C(k), .Y(men_men_n519_));
  NO3        u0491(.A(men_men_n519_), .B(men_men_n518_), .C(men_men_n104_), .Y(men_men_n520_));
  NO4        u0492(.A(n), .B(d), .C(men_men_n107_), .D(a), .Y(men_men_n521_));
  OR2        u0493(.A(n), .B(c), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n522_), .B(men_men_n139_), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n523_), .B(men_men_n521_), .Y(men_men_n524_));
  NOi32      u0496(.An(g), .Bn(f), .C(i), .Y(men_men_n525_));
  AOI220     u0497(.A0(men_men_n525_), .A1(men_men_n95_), .B0(men_men_n506_), .B1(f), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n263_), .B(men_men_n49_), .Y(men_men_n527_));
  NO2        u0499(.A(men_men_n526_), .B(men_men_n524_), .Y(men_men_n528_));
  INV        u0500(.A(men_men_n528_), .Y(men_men_n529_));
  NA2        u0501(.A(men_men_n132_), .B(men_men_n34_), .Y(men_men_n530_));
  OAI220     u0502(.A0(men_men_n530_), .A1(m), .B0(men_men_n510_), .B1(men_men_n224_), .Y(men_men_n531_));
  NOi41      u0503(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n532_));
  AN2        u0504(.A(men_men_n325_), .B(men_men_n308_), .Y(men_men_n533_));
  INV        u0505(.A(men_men_n533_), .Y(men_men_n534_));
  OA210      u0506(.A0(men_men_n534_), .A1(men_men_n532_), .B0(men_men_n531_), .Y(men_men_n535_));
  OAI220     u0507(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n504_), .B1(men_men_n503_), .Y(men_men_n536_));
  NAi31      u0508(.An(d), .B(c), .C(a), .Y(men_men_n537_));
  NO2        u0509(.A(men_men_n537_), .B(n), .Y(men_men_n538_));
  NA3        u0510(.A(men_men_n538_), .B(men_men_n536_), .C(e), .Y(men_men_n539_));
  INV        u0511(.A(men_men_n539_), .Y(men_men_n540_));
  NO2        u0512(.A(men_men_n265_), .B(n), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n411_), .B(men_men_n541_), .Y(men_men_n542_));
  NA2        u0514(.A(men_men_n536_), .B(f), .Y(men_men_n543_));
  NAi32      u0515(.An(d), .Bn(a), .C(b), .Y(men_men_n544_));
  NO2        u0516(.A(men_men_n544_), .B(men_men_n49_), .Y(men_men_n545_));
  NA2        u0517(.A(h), .B(f), .Y(men_men_n546_));
  NO2        u0518(.A(men_men_n546_), .B(men_men_n90_), .Y(men_men_n547_));
  NO3        u0519(.A(men_men_n167_), .B(men_men_n164_), .C(g), .Y(men_men_n548_));
  AOI220     u0520(.A0(men_men_n548_), .A1(men_men_n58_), .B0(men_men_n547_), .B1(men_men_n545_), .Y(men_men_n549_));
  OAI210     u0521(.A0(men_men_n543_), .A1(men_men_n542_), .B0(men_men_n549_), .Y(men_men_n550_));
  AN3        u0522(.A(j), .B(h), .C(g), .Y(men_men_n551_));
  NO2        u0523(.A(men_men_n136_), .B(c), .Y(men_men_n552_));
  NA3        u0524(.A(men_men_n552_), .B(men_men_n551_), .C(men_men_n437_), .Y(men_men_n553_));
  NA3        u0525(.A(f), .B(d), .C(b), .Y(men_men_n554_));
  NO4        u0526(.A(men_men_n554_), .B(men_men_n167_), .C(men_men_n164_), .D(g), .Y(men_men_n555_));
  INV        u0527(.A(men_men_n553_), .Y(men_men_n556_));
  NO4        u0528(.A(men_men_n556_), .B(men_men_n550_), .C(men_men_n540_), .D(men_men_n535_), .Y(men_men_n557_));
  AN4        u0529(.A(men_men_n557_), .B(men_men_n529_), .C(men_men_n514_), .D(men_men_n507_), .Y(men_men_n558_));
  INV        u0530(.A(k), .Y(men_men_n559_));
  NA3        u0531(.A(l), .B(men_men_n559_), .C(i), .Y(men_men_n560_));
  INV        u0532(.A(men_men_n560_), .Y(men_men_n561_));
  NA4        u0533(.A(men_men_n380_), .B(men_men_n400_), .C(men_men_n172_), .D(men_men_n105_), .Y(men_men_n562_));
  NAi32      u0534(.An(h), .Bn(f), .C(g), .Y(men_men_n563_));
  NAi41      u0535(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n564_));
  OAI210     u0536(.A0(men_men_n512_), .A1(n), .B0(men_men_n564_), .Y(men_men_n565_));
  NA2        u0537(.A(men_men_n565_), .B(m), .Y(men_men_n566_));
  NAi31      u0538(.An(h), .B(g), .C(f), .Y(men_men_n567_));
  OR3        u0539(.A(men_men_n567_), .B(men_men_n265_), .C(men_men_n49_), .Y(men_men_n568_));
  NA4        u0540(.A(men_men_n400_), .B(men_men_n112_), .C(men_men_n105_), .D(e), .Y(men_men_n569_));
  AN2        u0541(.A(men_men_n569_), .B(men_men_n568_), .Y(men_men_n570_));
  OA210      u0542(.A0(men_men_n566_), .A1(men_men_n563_), .B0(men_men_n570_), .Y(men_men_n571_));
  NO3        u0543(.A(men_men_n563_), .B(men_men_n72_), .C(men_men_n74_), .Y(men_men_n572_));
  NO4        u0544(.A(men_men_n567_), .B(men_men_n522_), .C(men_men_n139_), .D(men_men_n74_), .Y(men_men_n573_));
  OR2        u0545(.A(men_men_n573_), .B(men_men_n572_), .Y(men_men_n574_));
  NAi21      u0546(.An(men_men_n574_), .B(men_men_n571_), .Y(men_men_n575_));
  NAi31      u0547(.An(f), .B(h), .C(g), .Y(men_men_n576_));
  NO4        u0548(.A(men_men_n300_), .B(men_men_n576_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n577_));
  NOi32      u0549(.An(b), .Bn(a), .C(c), .Y(men_men_n578_));
  NOi41      u0550(.An(men_men_n578_), .B(men_men_n340_), .C(men_men_n69_), .D(men_men_n108_), .Y(men_men_n579_));
  OR2        u0551(.A(men_men_n579_), .B(men_men_n577_), .Y(men_men_n580_));
  NOi32      u0552(.An(d), .Bn(a), .C(e), .Y(men_men_n581_));
  NA2        u0553(.A(men_men_n581_), .B(men_men_n105_), .Y(men_men_n582_));
  NO2        u0554(.A(n), .B(c), .Y(men_men_n583_));
  NA3        u0555(.A(men_men_n583_), .B(men_men_n29_), .C(m), .Y(men_men_n584_));
  NAi32      u0556(.An(n), .Bn(f), .C(m), .Y(men_men_n585_));
  NA3        u0557(.A(men_men_n585_), .B(men_men_n584_), .C(men_men_n582_), .Y(men_men_n586_));
  NOi32      u0558(.An(e), .Bn(a), .C(d), .Y(men_men_n587_));
  AOI210     u0559(.A0(men_men_n29_), .A1(d), .B0(men_men_n587_), .Y(men_men_n588_));
  AOI210     u0560(.A0(men_men_n588_), .A1(men_men_n204_), .B0(men_men_n530_), .Y(men_men_n589_));
  AOI210     u0561(.A0(men_men_n589_), .A1(men_men_n586_), .B0(men_men_n580_), .Y(men_men_n590_));
  INV        u0562(.A(men_men_n590_), .Y(men_men_n591_));
  AOI210     u0563(.A0(men_men_n575_), .A1(men_men_n561_), .B0(men_men_n591_), .Y(men_men_n592_));
  NO3        u0564(.A(men_men_n307_), .B(men_men_n61_), .C(n), .Y(men_men_n593_));
  NA3        u0565(.A(men_men_n488_), .B(men_men_n162_), .C(men_men_n161_), .Y(men_men_n594_));
  NA2        u0566(.A(men_men_n439_), .B(men_men_n221_), .Y(men_men_n595_));
  OR2        u0567(.A(men_men_n595_), .B(men_men_n594_), .Y(men_men_n596_));
  NA2        u0568(.A(men_men_n75_), .B(men_men_n105_), .Y(men_men_n597_));
  NO2        u0569(.A(men_men_n597_), .B(men_men_n45_), .Y(men_men_n598_));
  AOI220     u0570(.A0(men_men_n598_), .A1(men_men_n517_), .B0(men_men_n596_), .B1(men_men_n593_), .Y(men_men_n599_));
  NO2        u0571(.A(men_men_n599_), .B(men_men_n83_), .Y(men_men_n600_));
  NOi32      u0572(.An(e), .Bn(c), .C(f), .Y(men_men_n601_));
  NOi21      u0573(.An(f), .B(g), .Y(men_men_n602_));
  NO2        u0574(.A(men_men_n602_), .B(men_men_n202_), .Y(men_men_n603_));
  AOI220     u0575(.A0(men_men_n603_), .A1(men_men_n377_), .B0(men_men_n601_), .B1(men_men_n166_), .Y(men_men_n604_));
  NA2        u0576(.A(men_men_n604_), .B(men_men_n169_), .Y(men_men_n605_));
  AOI210     u0577(.A0(men_men_n516_), .A1(men_men_n381_), .B0(men_men_n289_), .Y(men_men_n606_));
  NA2        u0578(.A(men_men_n606_), .B(men_men_n254_), .Y(men_men_n607_));
  NOi21      u0579(.An(j), .B(l), .Y(men_men_n608_));
  NAi21      u0580(.An(k), .B(h), .Y(men_men_n609_));
  NO2        u0581(.A(men_men_n609_), .B(men_men_n252_), .Y(men_men_n610_));
  NA2        u0582(.A(men_men_n610_), .B(men_men_n608_), .Y(men_men_n611_));
  OR2        u0583(.A(men_men_n611_), .B(men_men_n566_), .Y(men_men_n612_));
  NOi31      u0584(.An(m), .B(n), .C(k), .Y(men_men_n613_));
  NA2        u0585(.A(men_men_n608_), .B(men_men_n613_), .Y(men_men_n614_));
  NO2        u0586(.A(men_men_n265_), .B(men_men_n49_), .Y(men_men_n615_));
  NO2        u0587(.A(men_men_n300_), .B(men_men_n576_), .Y(men_men_n616_));
  NO2        u0588(.A(men_men_n512_), .B(men_men_n49_), .Y(men_men_n617_));
  AOI220     u0589(.A0(men_men_n617_), .A1(men_men_n616_), .B0(men_men_n615_), .B1(men_men_n547_), .Y(men_men_n618_));
  NA3        u0590(.A(men_men_n618_), .B(men_men_n612_), .C(men_men_n607_), .Y(men_men_n619_));
  NA2        u0591(.A(men_men_n101_), .B(men_men_n36_), .Y(men_men_n620_));
  NO2        u0592(.A(k), .B(men_men_n205_), .Y(men_men_n621_));
  NO2        u0593(.A(men_men_n508_), .B(men_men_n347_), .Y(men_men_n622_));
  NO2        u0594(.A(men_men_n622_), .B(n), .Y(men_men_n623_));
  NAi31      u0595(.An(men_men_n620_), .B(men_men_n623_), .C(men_men_n621_), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n484_), .B(men_men_n149_), .Y(men_men_n625_));
  NO3        u0597(.A(men_men_n378_), .B(men_men_n625_), .C(men_men_n83_), .Y(men_men_n626_));
  INV        u0598(.A(men_men_n626_), .Y(men_men_n627_));
  AN3        u0599(.A(f), .B(d), .C(b), .Y(men_men_n628_));
  OAI210     u0600(.A0(men_men_n628_), .A1(men_men_n122_), .B0(n), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n484_), .B(men_men_n149_), .C(men_men_n205_), .Y(men_men_n630_));
  AOI210     u0602(.A0(men_men_n629_), .A1(men_men_n223_), .B0(men_men_n630_), .Y(men_men_n631_));
  NAi31      u0603(.An(m), .B(n), .C(k), .Y(men_men_n632_));
  INV        u0604(.A(men_men_n240_), .Y(men_men_n633_));
  OAI210     u0605(.A0(men_men_n633_), .A1(men_men_n631_), .B0(j), .Y(men_men_n634_));
  NA3        u0606(.A(men_men_n634_), .B(men_men_n627_), .C(men_men_n624_), .Y(men_men_n635_));
  NO4        u0607(.A(men_men_n635_), .B(men_men_n619_), .C(men_men_n605_), .D(men_men_n600_), .Y(men_men_n636_));
  NAi31      u0608(.An(g), .B(h), .C(f), .Y(men_men_n637_));
  OR3        u0609(.A(men_men_n637_), .B(men_men_n265_), .C(n), .Y(men_men_n638_));
  OA210      u0610(.A0(men_men_n512_), .A1(n), .B0(men_men_n564_), .Y(men_men_n639_));
  NA3        u0611(.A(men_men_n398_), .B(men_men_n112_), .C(men_men_n80_), .Y(men_men_n640_));
  OAI210     u0612(.A0(men_men_n639_), .A1(men_men_n87_), .B0(men_men_n640_), .Y(men_men_n641_));
  NOi21      u0613(.An(men_men_n638_), .B(men_men_n641_), .Y(men_men_n642_));
  NO2        u0614(.A(men_men_n642_), .B(men_men_n505_), .Y(men_men_n643_));
  NO3        u0615(.A(g), .B(men_men_n204_), .C(men_men_n56_), .Y(men_men_n644_));
  NA2        u0616(.A(men_men_n377_), .B(men_men_n644_), .Y(men_men_n645_));
  BUFFER     u0617(.A(men_men_n72_), .Y(men_men_n646_));
  NA2        u0618(.A(men_men_n578_), .B(men_men_n329_), .Y(men_men_n647_));
  OA220      u0619(.A0(men_men_n614_), .A1(men_men_n647_), .B0(men_men_n611_), .B1(men_men_n646_), .Y(men_men_n648_));
  NA3        u0620(.A(men_men_n502_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n649_));
  AN2        u0621(.A(h), .B(f), .Y(men_men_n650_));
  NA2        u0622(.A(men_men_n650_), .B(men_men_n37_), .Y(men_men_n651_));
  NA2        u0623(.A(men_men_n95_), .B(men_men_n46_), .Y(men_men_n652_));
  OAI220     u0624(.A0(men_men_n652_), .A1(men_men_n320_), .B0(men_men_n651_), .B1(men_men_n444_), .Y(men_men_n653_));
  AOI210     u0625(.A0(men_men_n544_), .A1(men_men_n410_), .B0(men_men_n49_), .Y(men_men_n654_));
  OAI220     u0626(.A0(men_men_n567_), .A1(men_men_n560_), .B0(men_men_n313_), .B1(men_men_n503_), .Y(men_men_n655_));
  AOI210     u0627(.A0(men_men_n655_), .A1(men_men_n654_), .B0(men_men_n653_), .Y(men_men_n656_));
  NA4        u0628(.A(men_men_n656_), .B(men_men_n649_), .C(men_men_n648_), .D(men_men_n645_), .Y(men_men_n657_));
  NO2        u0629(.A(men_men_n241_), .B(f), .Y(men_men_n658_));
  INV        u0630(.A(men_men_n61_), .Y(men_men_n659_));
  NO3        u0631(.A(men_men_n659_), .B(men_men_n658_), .C(men_men_n34_), .Y(men_men_n660_));
  NA2        u0632(.A(men_men_n316_), .B(men_men_n132_), .Y(men_men_n661_));
  NA2        u0633(.A(men_men_n124_), .B(men_men_n49_), .Y(men_men_n662_));
  OR2        u0634(.A(men_men_n345_), .B(men_men_n103_), .Y(men_men_n663_));
  OAI210     u0635(.A0(men_men_n661_), .A1(men_men_n660_), .B0(men_men_n663_), .Y(men_men_n664_));
  NO3        u0636(.A(men_men_n386_), .B(men_men_n184_), .C(men_men_n183_), .Y(men_men_n665_));
  NA2        u0637(.A(men_men_n665_), .B(men_men_n221_), .Y(men_men_n666_));
  NA3        u0638(.A(men_men_n666_), .B(men_men_n243_), .C(j), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n443_), .B(men_men_n80_), .Y(men_men_n668_));
  NO4        u0640(.A(men_men_n505_), .B(men_men_n668_), .C(men_men_n123_), .D(men_men_n204_), .Y(men_men_n669_));
  INV        u0641(.A(men_men_n669_), .Y(men_men_n670_));
  NA3        u0642(.A(men_men_n670_), .B(men_men_n667_), .C(men_men_n384_), .Y(men_men_n671_));
  NO4        u0643(.A(men_men_n671_), .B(men_men_n664_), .C(men_men_n657_), .D(men_men_n643_), .Y(men_men_n672_));
  NA4        u0644(.A(men_men_n672_), .B(men_men_n636_), .C(men_men_n592_), .D(men_men_n558_), .Y(men08));
  NO2        u0645(.A(k), .B(h), .Y(men_men_n674_));
  AO210      u0646(.A0(men_men_n241_), .A1(men_men_n431_), .B0(men_men_n674_), .Y(men_men_n675_));
  NO2        u0647(.A(men_men_n675_), .B(men_men_n287_), .Y(men_men_n676_));
  NA2        u0648(.A(men_men_n601_), .B(men_men_n80_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n677_), .B(men_men_n439_), .Y(men_men_n678_));
  AOI210     u0650(.A0(men_men_n678_), .A1(men_men_n676_), .B0(men_men_n469_), .Y(men_men_n679_));
  NA2        u0651(.A(men_men_n80_), .B(men_men_n102_), .Y(men_men_n680_));
  NO2        u0652(.A(men_men_n680_), .B(men_men_n57_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n554_), .B(men_men_n223_), .Y(men_men_n682_));
  NA2        u0654(.A(men_men_n682_), .B(men_men_n334_), .Y(men_men_n683_));
  AOI210     u0655(.A0(men_men_n554_), .A1(men_men_n145_), .B0(men_men_n80_), .Y(men_men_n684_));
  NA4        u0656(.A(men_men_n207_), .B(men_men_n132_), .C(men_men_n45_), .D(h), .Y(men_men_n685_));
  AN2        u0657(.A(l), .B(k), .Y(men_men_n686_));
  NA4        u0658(.A(men_men_n686_), .B(men_men_n101_), .C(men_men_n74_), .D(men_men_n205_), .Y(men_men_n687_));
  OAI210     u0659(.A0(men_men_n685_), .A1(g), .B0(men_men_n687_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n688_), .B(men_men_n684_), .Y(men_men_n689_));
  NA4        u0661(.A(men_men_n689_), .B(men_men_n683_), .C(men_men_n679_), .D(men_men_n336_), .Y(men_men_n690_));
  AN2        u0662(.A(men_men_n513_), .B(men_men_n91_), .Y(men_men_n691_));
  NO4        u0663(.A(men_men_n164_), .B(men_men_n376_), .C(men_men_n104_), .D(g), .Y(men_men_n692_));
  AOI210     u0664(.A0(men_men_n692_), .A1(men_men_n682_), .B0(men_men_n497_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n603_), .B(men_men_n333_), .Y(men_men_n694_));
  NAi31      u0666(.An(men_men_n691_), .B(men_men_n694_), .C(men_men_n693_), .Y(men_men_n695_));
  NO3        u0667(.A(men_men_n307_), .B(men_men_n123_), .C(men_men_n41_), .Y(men_men_n696_));
  NAi21      u0668(.An(men_men_n696_), .B(men_men_n687_), .Y(men_men_n697_));
  NA2        u0669(.A(men_men_n675_), .B(men_men_n128_), .Y(men_men_n698_));
  AOI220     u0670(.A0(men_men_n698_), .A1(men_men_n385_), .B0(men_men_n697_), .B1(men_men_n76_), .Y(men_men_n699_));
  INV        u0671(.A(men_men_n699_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n347_), .B(men_men_n43_), .Y(men_men_n701_));
  NA3        u0673(.A(men_men_n666_), .B(men_men_n322_), .C(men_men_n368_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n686_), .B(men_men_n212_), .Y(men_men_n703_));
  NO2        u0675(.A(men_men_n703_), .B(men_men_n315_), .Y(men_men_n704_));
  AOI210     u0676(.A0(men_men_n704_), .A1(men_men_n658_), .B0(men_men_n468_), .Y(men_men_n705_));
  NA3        u0677(.A(m), .B(l), .C(k), .Y(men_men_n706_));
  AOI210     u0678(.A0(men_men_n640_), .A1(men_men_n638_), .B0(men_men_n706_), .Y(men_men_n707_));
  NO2        u0679(.A(men_men_n515_), .B(men_men_n261_), .Y(men_men_n708_));
  NOi21      u0680(.An(men_men_n708_), .B(men_men_n509_), .Y(men_men_n709_));
  NA4        u0681(.A(men_men_n105_), .B(l), .C(k), .D(men_men_n83_), .Y(men_men_n710_));
  NA3        u0682(.A(men_men_n112_), .B(men_men_n393_), .C(i), .Y(men_men_n711_));
  NO2        u0683(.A(men_men_n711_), .B(men_men_n710_), .Y(men_men_n712_));
  NO3        u0684(.A(men_men_n712_), .B(men_men_n709_), .C(men_men_n707_), .Y(men_men_n713_));
  NA4        u0685(.A(men_men_n713_), .B(men_men_n705_), .C(men_men_n702_), .D(men_men_n701_), .Y(men_men_n714_));
  NO4        u0686(.A(men_men_n714_), .B(men_men_n700_), .C(men_men_n695_), .D(men_men_n690_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n603_), .B(men_men_n377_), .Y(men_men_n716_));
  NOi31      u0688(.An(g), .B(h), .C(f), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n617_), .B(men_men_n717_), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n716_), .B(men_men_n240_), .Y(men_men_n719_));
  NA2        u0691(.A(men_men_n686_), .B(men_men_n74_), .Y(men_men_n720_));
  NO4        u0692(.A(men_men_n665_), .B(men_men_n164_), .C(n), .D(i), .Y(men_men_n721_));
  NOi21      u0693(.An(h), .B(j), .Y(men_men_n722_));
  NA2        u0694(.A(men_men_n722_), .B(f), .Y(men_men_n723_));
  INV        u0695(.A(men_men_n721_), .Y(men_men_n724_));
  OAI220     u0696(.A0(men_men_n724_), .A1(men_men_n720_), .B0(men_men_n570_), .B1(men_men_n62_), .Y(men_men_n725_));
  AOI210     u0697(.A0(men_men_n719_), .A1(l), .B0(men_men_n725_), .Y(men_men_n726_));
  NO2        u0698(.A(j), .B(i), .Y(men_men_n727_));
  NA2        u0699(.A(men_men_n727_), .B(men_men_n33_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n403_), .B(men_men_n112_), .Y(men_men_n729_));
  OR2        u0701(.A(men_men_n729_), .B(men_men_n728_), .Y(men_men_n730_));
  NO3        u0702(.A(men_men_n140_), .B(men_men_n49_), .C(men_men_n102_), .Y(men_men_n731_));
  NO3        u0703(.A(men_men_n522_), .B(men_men_n139_), .C(men_men_n74_), .Y(men_men_n732_));
  NO3        u0704(.A(men_men_n465_), .B(men_men_n422_), .C(j), .Y(men_men_n733_));
  OAI210     u0705(.A0(men_men_n732_), .A1(men_men_n731_), .B0(men_men_n733_), .Y(men_men_n734_));
  OAI210     u0706(.A0(men_men_n718_), .A1(men_men_n62_), .B0(men_men_n734_), .Y(men_men_n735_));
  NA2        u0707(.A(k), .B(j), .Y(men_men_n736_));
  NO3        u0708(.A(men_men_n287_), .B(men_men_n736_), .C(men_men_n40_), .Y(men_men_n737_));
  INV        u0709(.A(men_men_n532_), .Y(men_men_n738_));
  NA2        u0710(.A(men_men_n738_), .B(men_men_n533_), .Y(men_men_n739_));
  AN3        u0711(.A(men_men_n739_), .B(men_men_n737_), .C(men_men_n94_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n595_), .B(men_men_n297_), .Y(men_men_n741_));
  INV        u0713(.A(men_men_n741_), .Y(men_men_n742_));
  NO2        u0714(.A(men_men_n287_), .B(men_men_n128_), .Y(men_men_n743_));
  AOI220     u0715(.A0(men_men_n743_), .A1(men_men_n603_), .B0(men_men_n696_), .B1(men_men_n684_), .Y(men_men_n744_));
  NO2        u0716(.A(men_men_n706_), .B(men_men_n87_), .Y(men_men_n745_));
  NA2        u0717(.A(men_men_n745_), .B(men_men_n565_), .Y(men_men_n746_));
  NO2        u0718(.A(men_men_n567_), .B(men_men_n108_), .Y(men_men_n747_));
  OAI210     u0719(.A0(men_men_n747_), .A1(men_men_n733_), .B0(men_men_n654_), .Y(men_men_n748_));
  NA3        u0720(.A(men_men_n748_), .B(men_men_n746_), .C(men_men_n744_), .Y(men_men_n749_));
  OR4        u0721(.A(men_men_n749_), .B(men_men_n742_), .C(men_men_n740_), .D(men_men_n735_), .Y(men_men_n750_));
  NA2        u0722(.A(men_men_n738_), .B(men_men_n533_), .Y(men_men_n751_));
  NA4        u0723(.A(men_men_n751_), .B(men_men_n207_), .C(men_men_n431_), .D(men_men_n34_), .Y(men_men_n752_));
  OAI220     u0724(.A0(men_men_n685_), .A1(men_men_n677_), .B0(men_men_n320_), .B1(men_men_n38_), .Y(men_men_n753_));
  INV        u0725(.A(men_men_n753_), .Y(men_men_n754_));
  NA3        u0726(.A(men_men_n525_), .B(men_men_n280_), .C(h), .Y(men_men_n755_));
  NOi21      u0727(.An(men_men_n654_), .B(men_men_n755_), .Y(men_men_n756_));
  NO2        u0728(.A(men_men_n88_), .B(men_men_n47_), .Y(men_men_n757_));
  NO2        u0729(.A(men_men_n755_), .B(men_men_n584_), .Y(men_men_n758_));
  AOI210     u0730(.A0(men_men_n757_), .A1(men_men_n623_), .B0(men_men_n758_), .Y(men_men_n759_));
  NAi41      u0731(.An(men_men_n756_), .B(men_men_n759_), .C(men_men_n754_), .D(men_men_n752_), .Y(men_men_n760_));
  OR2        u0732(.A(men_men_n745_), .B(men_men_n91_), .Y(men_men_n761_));
  AOI220     u0733(.A0(men_men_n761_), .A1(men_men_n229_), .B0(men_men_n733_), .B1(men_men_n615_), .Y(men_men_n762_));
  OAI210     u0734(.A0(men_men_n706_), .A1(men_men_n637_), .B0(men_men_n496_), .Y(men_men_n763_));
  NA3        u0735(.A(men_men_n239_), .B(men_men_n59_), .C(b), .Y(men_men_n764_));
  AOI220     u0736(.A0(men_men_n583_), .A1(men_men_n29_), .B0(men_men_n443_), .B1(men_men_n80_), .Y(men_men_n765_));
  NA2        u0737(.A(men_men_n765_), .B(men_men_n764_), .Y(men_men_n766_));
  NO2        u0738(.A(men_men_n755_), .B(men_men_n467_), .Y(men_men_n767_));
  AOI210     u0739(.A0(men_men_n766_), .A1(men_men_n763_), .B0(men_men_n767_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n768_), .B(men_men_n762_), .Y(men_men_n769_));
  NOi41      u0741(.An(men_men_n730_), .B(men_men_n769_), .C(men_men_n760_), .D(men_men_n750_), .Y(men_men_n770_));
  OR3        u0742(.A(men_men_n685_), .B(men_men_n223_), .C(g), .Y(men_men_n771_));
  NO3        u0743(.A(men_men_n328_), .B(men_men_n289_), .C(men_men_n104_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n772_), .B(men_men_n739_), .Y(men_men_n773_));
  NA2        u0745(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n774_));
  NO3        u0746(.A(men_men_n774_), .B(men_men_n728_), .C(men_men_n265_), .Y(men_men_n775_));
  NO3        u0747(.A(men_men_n503_), .B(men_men_n89_), .C(h), .Y(men_men_n776_));
  AOI210     u0748(.A0(men_men_n776_), .A1(men_men_n681_), .B0(men_men_n775_), .Y(men_men_n777_));
  NA3        u0749(.A(men_men_n777_), .B(men_men_n773_), .C(men_men_n771_), .Y(men_men_n778_));
  OR2        u0750(.A(men_men_n637_), .B(men_men_n88_), .Y(men_men_n779_));
  NOi31      u0751(.An(b), .B(d), .C(a), .Y(men_men_n780_));
  NO2        u0752(.A(men_men_n780_), .B(men_men_n581_), .Y(men_men_n781_));
  NO2        u0753(.A(men_men_n781_), .B(n), .Y(men_men_n782_));
  INV        u0754(.A(men_men_n782_), .Y(men_men_n783_));
  OAI220     u0755(.A0(men_men_n783_), .A1(men_men_n779_), .B0(men_men_n755_), .B1(men_men_n582_), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n315_), .B(men_men_n108_), .Y(men_men_n785_));
  NOi21      u0757(.An(men_men_n785_), .B(men_men_n150_), .Y(men_men_n786_));
  INV        u0758(.A(men_men_n786_), .Y(men_men_n787_));
  OAI210     u0759(.A0(men_men_n685_), .A1(men_men_n378_), .B0(men_men_n787_), .Y(men_men_n788_));
  NO2        u0760(.A(men_men_n665_), .B(n), .Y(men_men_n789_));
  AOI220     u0761(.A0(men_men_n743_), .A1(men_men_n644_), .B0(men_men_n789_), .B1(men_men_n676_), .Y(men_men_n790_));
  NA2        u0762(.A(men_men_n112_), .B(men_men_n80_), .Y(men_men_n791_));
  AOI210     u0763(.A0(men_men_n407_), .A1(men_men_n399_), .B0(men_men_n791_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n704_), .B(men_men_n34_), .Y(men_men_n793_));
  NAi21      u0765(.An(men_men_n710_), .B(men_men_n418_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n261_), .B(i), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n692_), .B(men_men_n335_), .Y(men_men_n796_));
  OAI210     u0768(.A0(men_men_n573_), .A1(men_men_n572_), .B0(men_men_n348_), .Y(men_men_n797_));
  AN3        u0769(.A(men_men_n797_), .B(men_men_n796_), .C(men_men_n794_), .Y(men_men_n798_));
  NAi41      u0770(.An(men_men_n792_), .B(men_men_n798_), .C(men_men_n793_), .D(men_men_n790_), .Y(men_men_n799_));
  NO4        u0771(.A(men_men_n799_), .B(men_men_n788_), .C(men_men_n784_), .D(men_men_n778_), .Y(men_men_n800_));
  NA4        u0772(.A(men_men_n800_), .B(men_men_n770_), .C(men_men_n726_), .D(men_men_n715_), .Y(men09));
  INV        u0773(.A(men_men_n113_), .Y(men_men_n802_));
  NA2        u0774(.A(f), .B(e), .Y(men_men_n803_));
  NO2        u0775(.A(men_men_n216_), .B(men_men_n104_), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n804_), .B(g), .Y(men_men_n805_));
  NA4        u0777(.A(men_men_n300_), .B(men_men_n451_), .C(men_men_n250_), .D(men_men_n110_), .Y(men_men_n806_));
  AOI210     u0778(.A0(men_men_n806_), .A1(g), .B0(men_men_n448_), .Y(men_men_n807_));
  AOI210     u0779(.A0(men_men_n807_), .A1(men_men_n805_), .B0(men_men_n803_), .Y(men_men_n808_));
  NA2        u0780(.A(men_men_n808_), .B(men_men_n802_), .Y(men_men_n809_));
  NO2        u0781(.A(men_men_n196_), .B(men_men_n204_), .Y(men_men_n810_));
  NA3        u0782(.A(m), .B(l), .C(i), .Y(men_men_n811_));
  OAI220     u0783(.A0(men_men_n567_), .A1(men_men_n811_), .B0(men_men_n340_), .B1(men_men_n504_), .Y(men_men_n812_));
  NA4        u0784(.A(men_men_n84_), .B(men_men_n83_), .C(g), .D(f), .Y(men_men_n813_));
  NAi21      u0785(.An(men_men_n812_), .B(men_men_n813_), .Y(men_men_n814_));
  OR2        u0786(.A(men_men_n814_), .B(men_men_n810_), .Y(men_men_n815_));
  NA3        u0787(.A(men_men_n779_), .B(men_men_n543_), .C(men_men_n496_), .Y(men_men_n816_));
  OA210      u0788(.A0(men_men_n816_), .A1(men_men_n815_), .B0(men_men_n782_), .Y(men_men_n817_));
  INV        u0789(.A(men_men_n325_), .Y(men_men_n818_));
  NO2        u0790(.A(men_men_n119_), .B(men_men_n117_), .Y(men_men_n819_));
  INV        u0791(.A(men_men_n327_), .Y(men_men_n820_));
  AOI210     u0792(.A0(men_men_n820_), .A1(men_men_n819_), .B0(men_men_n576_), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n764_), .B(men_men_n320_), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n329_), .B(men_men_n331_), .Y(men_men_n823_));
  OAI210     u0795(.A0(men_men_n196_), .A1(men_men_n204_), .B0(men_men_n823_), .Y(men_men_n824_));
  AOI220     u0796(.A0(men_men_n824_), .A1(men_men_n822_), .B0(men_men_n821_), .B1(men_men_n818_), .Y(men_men_n825_));
  NA2        u0797(.A(men_men_n158_), .B(men_men_n106_), .Y(men_men_n826_));
  NA3        u0798(.A(men_men_n826_), .B(men_men_n675_), .C(men_men_n128_), .Y(men_men_n827_));
  NA3        u0799(.A(men_men_n827_), .B(men_men_n181_), .C(men_men_n31_), .Y(men_men_n828_));
  NA3        u0800(.A(men_men_n828_), .B(men_men_n825_), .C(men_men_n604_), .Y(men_men_n829_));
  NO2        u0801(.A(men_men_n563_), .B(men_men_n474_), .Y(men_men_n830_));
  NA2        u0802(.A(men_men_n830_), .B(men_men_n181_), .Y(men_men_n831_));
  NOi21      u0803(.An(f), .B(d), .Y(men_men_n832_));
  NA2        u0804(.A(men_men_n832_), .B(m), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n833_), .B(men_men_n52_), .Y(men_men_n834_));
  NOi32      u0806(.An(g), .Bn(f), .C(d), .Y(men_men_n835_));
  NA4        u0807(.A(men_men_n835_), .B(men_men_n583_), .C(men_men_n29_), .D(m), .Y(men_men_n836_));
  NOi21      u0808(.An(men_men_n301_), .B(men_men_n836_), .Y(men_men_n837_));
  AOI210     u0809(.A0(men_men_n834_), .A1(men_men_n523_), .B0(men_men_n837_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n250_), .B(men_men_n110_), .Y(men_men_n839_));
  AN2        u0811(.A(f), .B(d), .Y(men_men_n840_));
  NA3        u0812(.A(men_men_n456_), .B(men_men_n840_), .C(men_men_n80_), .Y(men_men_n841_));
  NO3        u0813(.A(men_men_n841_), .B(men_men_n74_), .C(men_men_n205_), .Y(men_men_n842_));
  NO2        u0814(.A(men_men_n273_), .B(men_men_n56_), .Y(men_men_n843_));
  NA2        u0815(.A(men_men_n839_), .B(men_men_n842_), .Y(men_men_n844_));
  NAi41      u0816(.An(men_men_n466_), .B(men_men_n844_), .C(men_men_n838_), .D(men_men_n831_), .Y(men_men_n845_));
  NO2        u0817(.A(men_men_n632_), .B(men_men_n315_), .Y(men_men_n846_));
  AN2        u0818(.A(men_men_n846_), .B(men_men_n658_), .Y(men_men_n847_));
  NO2        u0819(.A(men_men_n847_), .B(men_men_n225_), .Y(men_men_n848_));
  NA2        u0820(.A(men_men_n581_), .B(men_men_n80_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n823_), .B(men_men_n849_), .Y(men_men_n850_));
  INV        u0822(.A(men_men_n850_), .Y(men_men_n851_));
  NA2        u0823(.A(c), .B(men_men_n107_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n852_), .B(men_men_n390_), .Y(men_men_n853_));
  NA3        u0825(.A(men_men_n853_), .B(men_men_n486_), .C(f), .Y(men_men_n854_));
  OR2        u0826(.A(men_men_n637_), .B(men_men_n519_), .Y(men_men_n855_));
  INV        u0827(.A(men_men_n855_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n781_), .B(men_men_n103_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n857_), .B(men_men_n856_), .Y(men_men_n858_));
  NA4        u0830(.A(men_men_n858_), .B(men_men_n854_), .C(men_men_n851_), .D(men_men_n848_), .Y(men_men_n859_));
  NO4        u0831(.A(men_men_n859_), .B(men_men_n845_), .C(men_men_n829_), .D(men_men_n817_), .Y(men_men_n860_));
  OR2        u0832(.A(men_men_n841_), .B(men_men_n74_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n804_), .B(g), .Y(men_men_n862_));
  AOI210     u0834(.A0(men_men_n862_), .A1(men_men_n281_), .B0(men_men_n861_), .Y(men_men_n863_));
  NO2        u0835(.A(men_men_n320_), .B(men_men_n813_), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n128_), .B(men_men_n124_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n221_), .B(men_men_n215_), .Y(men_men_n866_));
  AOI220     u0838(.A0(men_men_n866_), .A1(men_men_n218_), .B0(men_men_n294_), .B1(men_men_n865_), .Y(men_men_n867_));
  NO2        u0839(.A(men_men_n412_), .B(men_men_n803_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n868_), .B(men_men_n538_), .Y(men_men_n869_));
  NA2        u0841(.A(men_men_n869_), .B(men_men_n867_), .Y(men_men_n870_));
  NA2        u0842(.A(e), .B(d), .Y(men_men_n871_));
  OAI220     u0843(.A0(men_men_n871_), .A1(c), .B0(men_men_n310_), .B1(d), .Y(men_men_n872_));
  NA3        u0844(.A(men_men_n872_), .B(men_men_n434_), .C(men_men_n484_), .Y(men_men_n873_));
  AOI210     u0845(.A0(men_men_n491_), .A1(men_men_n171_), .B0(men_men_n221_), .Y(men_men_n874_));
  AOI210     u0846(.A0(men_men_n603_), .A1(men_men_n333_), .B0(men_men_n874_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n273_), .B(men_men_n154_), .Y(men_men_n876_));
  NA2        u0848(.A(men_men_n842_), .B(men_men_n876_), .Y(men_men_n877_));
  NA3        u0849(.A(men_men_n157_), .B(men_men_n81_), .C(men_men_n34_), .Y(men_men_n878_));
  NA4        u0850(.A(men_men_n878_), .B(men_men_n877_), .C(men_men_n875_), .D(men_men_n873_), .Y(men_men_n879_));
  NO4        u0851(.A(men_men_n879_), .B(men_men_n870_), .C(men_men_n864_), .D(men_men_n863_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n818_), .B(men_men_n31_), .Y(men_men_n881_));
  AO210      u0853(.A0(men_men_n881_), .A1(men_men_n677_), .B0(men_men_n208_), .Y(men_men_n882_));
  OAI220     u0854(.A0(men_men_n602_), .A1(men_men_n61_), .B0(men_men_n289_), .B1(j), .Y(men_men_n883_));
  AOI220     u0855(.A0(men_men_n883_), .A1(men_men_n846_), .B0(men_men_n593_), .B1(men_men_n601_), .Y(men_men_n884_));
  INV        u0856(.A(men_men_n884_), .Y(men_men_n885_));
  OAI210     u0857(.A0(men_men_n804_), .A1(men_men_n876_), .B0(men_men_n835_), .Y(men_men_n886_));
  NO2        u0858(.A(men_men_n886_), .B(men_men_n584_), .Y(men_men_n887_));
  AOI210     u0859(.A0(men_men_n109_), .A1(men_men_n108_), .B0(men_men_n249_), .Y(men_men_n888_));
  NO2        u0860(.A(men_men_n888_), .B(men_men_n836_), .Y(men_men_n889_));
  BUFFER     u0861(.A(men_men_n889_), .Y(men_men_n890_));
  NOi31      u0862(.An(men_men_n523_), .B(men_men_n833_), .C(men_men_n281_), .Y(men_men_n891_));
  NO4        u0863(.A(men_men_n891_), .B(men_men_n890_), .C(men_men_n887_), .D(men_men_n885_), .Y(men_men_n892_));
  AO220      u0864(.A0(men_men_n434_), .A1(men_men_n722_), .B0(men_men_n166_), .B1(f), .Y(men_men_n893_));
  NA2        u0865(.A(men_men_n893_), .B(men_men_n872_), .Y(men_men_n894_));
  NA2        u0866(.A(men_men_n816_), .B(men_men_n681_), .Y(men_men_n895_));
  AN4        u0867(.A(men_men_n895_), .B(men_men_n894_), .C(men_men_n892_), .D(men_men_n882_), .Y(men_men_n896_));
  NA4        u0868(.A(men_men_n896_), .B(men_men_n880_), .C(men_men_n860_), .D(men_men_n809_), .Y(men12));
  NO2        u0869(.A(men_men_n432_), .B(c), .Y(men_men_n898_));
  NO4        u0870(.A(men_men_n424_), .B(men_men_n241_), .C(men_men_n559_), .D(men_men_n205_), .Y(men_men_n899_));
  NA2        u0871(.A(men_men_n899_), .B(men_men_n898_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n432_), .B(men_men_n107_), .Y(men_men_n901_));
  NO2        u0873(.A(men_men_n819_), .B(men_men_n340_), .Y(men_men_n902_));
  NO2        u0874(.A(men_men_n637_), .B(men_men_n362_), .Y(men_men_n903_));
  AOI220     u0875(.A0(men_men_n903_), .A1(men_men_n521_), .B0(men_men_n902_), .B1(men_men_n901_), .Y(men_men_n904_));
  NA3        u0876(.A(men_men_n904_), .B(men_men_n900_), .C(men_men_n423_), .Y(men_men_n905_));
  AOI210     u0877(.A0(men_men_n224_), .A1(men_men_n324_), .B0(men_men_n193_), .Y(men_men_n906_));
  OR2        u0878(.A(men_men_n906_), .B(men_men_n899_), .Y(men_men_n907_));
  NO2        u0879(.A(men_men_n374_), .B(men_men_n205_), .Y(men_men_n908_));
  OAI210     u0880(.A0(men_men_n908_), .A1(men_men_n907_), .B0(men_men_n386_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n620_), .B(men_men_n252_), .Y(men_men_n910_));
  NO2        u0882(.A(men_men_n567_), .B(men_men_n811_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n911_), .B(men_men_n541_), .Y(men_men_n912_));
  NO2        u0884(.A(men_men_n140_), .B(men_men_n228_), .Y(men_men_n913_));
  NA3        u0885(.A(men_men_n913_), .B(men_men_n231_), .C(i), .Y(men_men_n914_));
  NA3        u0886(.A(men_men_n914_), .B(men_men_n912_), .C(men_men_n909_), .Y(men_men_n915_));
  NO3        u0887(.A(men_men_n642_), .B(men_men_n88_), .C(men_men_n45_), .Y(men_men_n916_));
  NO3        u0888(.A(men_men_n916_), .B(men_men_n915_), .C(men_men_n905_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n353_), .B(men_men_n352_), .Y(men_men_n918_));
  NA2        u0890(.A(men_men_n564_), .B(men_men_n72_), .Y(men_men_n919_));
  NOi21      u0891(.An(men_men_n34_), .B(men_men_n632_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n919_), .B(men_men_n918_), .Y(men_men_n921_));
  OAI210     u0893(.A0(men_men_n240_), .A1(men_men_n45_), .B0(men_men_n921_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n418_), .B(men_men_n254_), .Y(men_men_n923_));
  NO3        u0895(.A(men_men_n791_), .B(men_men_n85_), .C(men_men_n390_), .Y(men_men_n924_));
  NAi21      u0896(.An(men_men_n924_), .B(men_men_n923_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n926_));
  INV        u0898(.A(men_men_n350_), .Y(men_men_n927_));
  NO3        u0899(.A(men_men_n927_), .B(men_men_n925_), .C(men_men_n922_), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n151_), .B(i), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n46_), .B(i), .Y(men_men_n930_));
  OAI220     u0902(.A0(men_men_n930_), .A1(men_men_n192_), .B0(men_men_n929_), .B1(men_men_n88_), .Y(men_men_n931_));
  AOI210     u0903(.A0(men_men_n401_), .A1(men_men_n37_), .B0(men_men_n931_), .Y(men_men_n932_));
  NO2        u0904(.A(men_men_n932_), .B(men_men_n320_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n637_), .B(men_men_n474_), .Y(men_men_n934_));
  NA3        u0906(.A(men_men_n329_), .B(men_men_n608_), .C(i), .Y(men_men_n935_));
  OAI210     u0907(.A0(men_men_n422_), .A1(men_men_n300_), .B0(men_men_n935_), .Y(men_men_n936_));
  OAI220     u0908(.A0(men_men_n936_), .A1(men_men_n934_), .B0(men_men_n654_), .B1(men_men_n732_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n587_), .B(men_men_n105_), .Y(men_men_n938_));
  OR3        u0910(.A(men_men_n300_), .B(men_men_n417_), .C(f), .Y(men_men_n939_));
  NA3        u0911(.A(men_men_n608_), .B(men_men_n78_), .C(i), .Y(men_men_n940_));
  OA220      u0912(.A0(men_men_n940_), .A1(men_men_n938_), .B0(men_men_n939_), .B1(men_men_n566_), .Y(men_men_n941_));
  NA3        u0913(.A(men_men_n312_), .B(men_men_n109_), .C(g), .Y(men_men_n942_));
  AOI210     u0914(.A0(men_men_n651_), .A1(men_men_n942_), .B0(m), .Y(men_men_n943_));
  OAI210     u0915(.A0(men_men_n943_), .A1(men_men_n902_), .B0(men_men_n311_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n668_), .B(men_men_n849_), .Y(men_men_n945_));
  INV        u0917(.A(men_men_n813_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n213_), .B(men_men_n77_), .Y(men_men_n947_));
  NA3        u0919(.A(men_men_n947_), .B(men_men_n940_), .C(men_men_n939_), .Y(men_men_n948_));
  AOI220     u0920(.A0(men_men_n948_), .A1(men_men_n247_), .B0(men_men_n946_), .B1(men_men_n945_), .Y(men_men_n949_));
  NA4        u0921(.A(men_men_n949_), .B(men_men_n944_), .C(men_men_n941_), .D(men_men_n937_), .Y(men_men_n950_));
  NO2        u0922(.A(men_men_n362_), .B(men_men_n87_), .Y(men_men_n951_));
  OAI210     u0923(.A0(men_men_n951_), .A1(men_men_n910_), .B0(men_men_n229_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n641_), .B(men_men_n84_), .Y(men_men_n953_));
  NO2        u0925(.A(men_men_n438_), .B(men_men_n205_), .Y(men_men_n954_));
  NA2        u0926(.A(men_men_n954_), .B(men_men_n367_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n565_), .B(men_men_n86_), .Y(men_men_n956_));
  NA4        u0928(.A(men_men_n956_), .B(men_men_n955_), .C(men_men_n953_), .D(men_men_n952_), .Y(men_men_n957_));
  OAI210     u0929(.A0(men_men_n946_), .A1(men_men_n911_), .B0(men_men_n521_), .Y(men_men_n958_));
  AOI210     u0930(.A0(men_men_n402_), .A1(men_men_n394_), .B0(men_men_n791_), .Y(men_men_n959_));
  INV        u0931(.A(men_men_n959_), .Y(men_men_n960_));
  NA2        u0932(.A(men_men_n943_), .B(men_men_n901_), .Y(men_men_n961_));
  NA3        u0933(.A(men_men_n961_), .B(men_men_n960_), .C(men_men_n958_), .Y(men_men_n962_));
  NO4        u0934(.A(men_men_n962_), .B(men_men_n957_), .C(men_men_n950_), .D(men_men_n933_), .Y(men_men_n963_));
  NAi31      u0935(.An(men_men_n133_), .B(men_men_n403_), .C(n), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n117_), .B(men_men_n327_), .Y(men_men_n965_));
  NO2        u0937(.A(men_men_n965_), .B(men_men_n964_), .Y(men_men_n966_));
  NO3        u0938(.A(men_men_n261_), .B(men_men_n133_), .C(men_men_n390_), .Y(men_men_n967_));
  AOI210     u0939(.A0(men_men_n967_), .A1(men_men_n475_), .B0(men_men_n966_), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n469_), .B(i), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n969_), .B(men_men_n968_), .Y(men_men_n970_));
  NA2        u0942(.A(men_men_n221_), .B(men_men_n162_), .Y(men_men_n971_));
  NO3        u0943(.A(men_men_n297_), .B(men_men_n425_), .C(men_men_n166_), .Y(men_men_n972_));
  NOi31      u0944(.An(men_men_n971_), .B(men_men_n972_), .C(men_men_n205_), .Y(men_men_n973_));
  NO3        u0945(.A(men_men_n422_), .B(men_men_n300_), .C(men_men_n74_), .Y(men_men_n974_));
  AOI220     u0946(.A0(men_men_n974_), .A1(men_men_n419_), .B0(men_men_n462_), .B1(g), .Y(men_men_n975_));
  INV        u0947(.A(men_men_n975_), .Y(men_men_n976_));
  OAI220     u0948(.A0(men_men_n964_), .A1(men_men_n224_), .B0(men_men_n935_), .B1(men_men_n582_), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n638_), .B(men_men_n362_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n906_), .B(men_men_n898_), .Y(men_men_n979_));
  NO3        u0951(.A(men_men_n522_), .B(men_men_n139_), .C(men_men_n204_), .Y(men_men_n980_));
  OAI210     u0952(.A0(men_men_n980_), .A1(men_men_n502_), .B0(men_men_n363_), .Y(men_men_n981_));
  OAI220     u0953(.A0(men_men_n903_), .A1(men_men_n911_), .B0(men_men_n523_), .B1(men_men_n411_), .Y(men_men_n982_));
  NA3        u0954(.A(men_men_n982_), .B(men_men_n981_), .C(men_men_n979_), .Y(men_men_n983_));
  OAI210     u0955(.A0(men_men_n906_), .A1(men_men_n899_), .B0(men_men_n971_), .Y(men_men_n984_));
  AOI210     u0956(.A0(men_men_n365_), .A1(men_men_n363_), .B0(men_men_n319_), .Y(men_men_n985_));
  NA3        u0957(.A(men_men_n985_), .B(men_men_n984_), .C(men_men_n262_), .Y(men_men_n986_));
  OR4        u0958(.A(men_men_n986_), .B(men_men_n983_), .C(men_men_n978_), .D(men_men_n977_), .Y(men_men_n987_));
  NO4        u0959(.A(men_men_n987_), .B(men_men_n976_), .C(men_men_n973_), .D(men_men_n970_), .Y(men_men_n988_));
  NA4        u0960(.A(men_men_n988_), .B(men_men_n963_), .C(men_men_n928_), .D(men_men_n917_), .Y(men13));
  AN2        u0961(.A(c), .B(b), .Y(men_men_n990_));
  NA3        u0962(.A(men_men_n239_), .B(men_men_n990_), .C(m), .Y(men_men_n991_));
  NA2        u0963(.A(d), .B(f), .Y(men_men_n992_));
  NO4        u0964(.A(men_men_n992_), .B(men_men_n991_), .C(j), .D(men_men_n560_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n254_), .B(men_men_n990_), .Y(men_men_n994_));
  NO4        u0966(.A(men_men_n994_), .B(men_men_n992_), .C(men_men_n929_), .D(a), .Y(men_men_n995_));
  NAi32      u0967(.An(d), .Bn(c), .C(e), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n132_), .B(men_men_n45_), .Y(men_men_n997_));
  NO4        u0969(.A(men_men_n997_), .B(men_men_n996_), .C(men_men_n567_), .D(men_men_n296_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n393_), .B(men_men_n204_), .Y(men_men_n999_));
  AN2        u0971(.A(d), .B(c), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n1000_), .B(men_men_n107_), .Y(men_men_n1001_));
  NO4        u0973(.A(men_men_n1001_), .B(men_men_n999_), .C(men_men_n167_), .D(men_men_n158_), .Y(men_men_n1002_));
  NA2        u0974(.A(d), .B(c), .Y(men_men_n1003_));
  NO4        u0975(.A(men_men_n997_), .B(men_men_n563_), .C(men_men_n1003_), .D(men_men_n296_), .Y(men_men_n1004_));
  OR2        u0976(.A(men_men_n1002_), .B(men_men_n1004_), .Y(men_men_n1005_));
  OR4        u0977(.A(men_men_n1005_), .B(men_men_n998_), .C(men_men_n995_), .D(men_men_n993_), .Y(men_men_n1006_));
  NAi32      u0978(.An(f), .Bn(e), .C(c), .Y(men_men_n1007_));
  NO2        u0979(.A(men_men_n1007_), .B(men_men_n136_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n1008_), .B(g), .Y(men_men_n1009_));
  OR3        u0981(.A(men_men_n215_), .B(men_men_n167_), .C(men_men_n158_), .Y(men_men_n1010_));
  NO2        u0982(.A(men_men_n1010_), .B(men_men_n1009_), .Y(men_men_n1011_));
  NO2        u0983(.A(men_men_n1003_), .B(men_men_n296_), .Y(men_men_n1012_));
  NO2        u0984(.A(j), .B(men_men_n45_), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n610_), .B(men_men_n1013_), .Y(men_men_n1014_));
  NOi21      u0986(.An(men_men_n1012_), .B(men_men_n1014_), .Y(men_men_n1015_));
  NO2        u0987(.A(men_men_n736_), .B(men_men_n104_), .Y(men_men_n1016_));
  NOi41      u0988(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n1017_), .B(men_men_n1016_), .Y(men_men_n1018_));
  NO2        u0990(.A(men_men_n1018_), .B(men_men_n1009_), .Y(men_men_n1019_));
  OR3        u0991(.A(e), .B(d), .C(c), .Y(men_men_n1020_));
  NA3        u0992(.A(k), .B(j), .C(i), .Y(men_men_n1021_));
  NO3        u0993(.A(men_men_n1021_), .B(men_men_n296_), .C(men_men_n87_), .Y(men_men_n1022_));
  NOi21      u0994(.An(men_men_n1022_), .B(men_men_n1020_), .Y(men_men_n1023_));
  OR4        u0995(.A(men_men_n1023_), .B(men_men_n1019_), .C(men_men_n1015_), .D(men_men_n1011_), .Y(men_men_n1024_));
  NA3        u0996(.A(men_men_n446_), .B(men_men_n322_), .C(men_men_n56_), .Y(men_men_n1025_));
  NO2        u0997(.A(men_men_n1025_), .B(men_men_n1014_), .Y(men_men_n1026_));
  NO2        u0998(.A(f), .B(c), .Y(men_men_n1027_));
  NOi21      u0999(.An(men_men_n1027_), .B(men_men_n424_), .Y(men_men_n1028_));
  NA2        u1000(.A(men_men_n1028_), .B(men_men_n59_), .Y(men_men_n1029_));
  OR2        u1001(.A(k), .B(i), .Y(men_men_n1030_));
  NO3        u1002(.A(men_men_n1030_), .B(men_men_n235_), .C(l), .Y(men_men_n1031_));
  NOi31      u1003(.An(men_men_n1031_), .B(men_men_n1029_), .C(j), .Y(men_men_n1032_));
  OR2        u1004(.A(men_men_n1032_), .B(men_men_n1026_), .Y(men_men_n1033_));
  OR3        u1005(.A(men_men_n1033_), .B(men_men_n1024_), .C(men_men_n1006_), .Y(men02));
  OR2        u1006(.A(l), .B(k), .Y(men_men_n1035_));
  OR3        u1007(.A(h), .B(g), .C(f), .Y(men_men_n1036_));
  OR3        u1008(.A(n), .B(m), .C(i), .Y(men_men_n1037_));
  NO4        u1009(.A(men_men_n1037_), .B(men_men_n1036_), .C(men_men_n1035_), .D(men_men_n1020_), .Y(men_men_n1038_));
  NOi31      u1010(.An(e), .B(d), .C(c), .Y(men_men_n1039_));
  AOI210     u1011(.A0(men_men_n1022_), .A1(men_men_n1039_), .B0(men_men_n998_), .Y(men_men_n1040_));
  AN3        u1012(.A(g), .B(f), .C(c), .Y(men_men_n1041_));
  NA3        u1013(.A(men_men_n1041_), .B(men_men_n446_), .C(h), .Y(men_men_n1042_));
  OR2        u1014(.A(men_men_n1021_), .B(men_men_n296_), .Y(men_men_n1043_));
  OR2        u1015(.A(men_men_n1043_), .B(men_men_n1042_), .Y(men_men_n1044_));
  NO3        u1016(.A(men_men_n1025_), .B(men_men_n997_), .C(men_men_n563_), .Y(men_men_n1045_));
  NO2        u1017(.A(men_men_n1045_), .B(men_men_n1011_), .Y(men_men_n1046_));
  NA3        u1018(.A(l), .B(k), .C(j), .Y(men_men_n1047_));
  NA2        u1019(.A(i), .B(h), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n1048_), .B(men_men_n1047_), .C(men_men_n124_), .Y(men_men_n1049_));
  NO3        u1021(.A(men_men_n134_), .B(men_men_n271_), .C(men_men_n205_), .Y(men_men_n1050_));
  AOI210     u1022(.A0(men_men_n1050_), .A1(men_men_n1049_), .B0(men_men_n1015_), .Y(men_men_n1051_));
  NA3        u1023(.A(c), .B(b), .C(a), .Y(men_men_n1052_));
  NO3        u1024(.A(men_men_n1052_), .B(men_men_n871_), .C(men_men_n204_), .Y(men_men_n1053_));
  NO3        u1025(.A(men_men_n1021_), .B(men_men_n49_), .C(men_men_n104_), .Y(men_men_n1054_));
  AOI210     u1026(.A0(men_men_n1054_), .A1(men_men_n1053_), .B0(men_men_n1026_), .Y(men_men_n1055_));
  AN4        u1027(.A(men_men_n1055_), .B(men_men_n1051_), .C(men_men_n1046_), .D(men_men_n1044_), .Y(men_men_n1056_));
  NO2        u1028(.A(men_men_n1001_), .B(men_men_n999_), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n1018_), .B(men_men_n1010_), .Y(men_men_n1058_));
  AOI210     u1030(.A0(men_men_n1058_), .A1(men_men_n1057_), .B0(men_men_n993_), .Y(men_men_n1059_));
  NAi41      u1031(.An(men_men_n1038_), .B(men_men_n1059_), .C(men_men_n1056_), .D(men_men_n1040_), .Y(men03));
  NA4        u1032(.A(men_men_n84_), .B(men_men_n83_), .C(g), .D(men_men_n204_), .Y(men_men_n1061_));
  NA4        u1033(.A(men_men_n551_), .B(m), .C(men_men_n104_), .D(men_men_n204_), .Y(men_men_n1062_));
  NA2        u1034(.A(men_men_n1062_), .B(men_men_n1061_), .Y(men_men_n1063_));
  INV        u1035(.A(men_men_n1063_), .Y(men_men_n1064_));
  NO2        u1036(.A(men_men_n824_), .B(men_men_n814_), .Y(men_men_n1065_));
  OAI220     u1037(.A0(men_men_n1065_), .A1(men_men_n668_), .B0(men_men_n1064_), .B1(men_men_n564_), .Y(men_men_n1066_));
  NOi31      u1038(.An(i), .B(k), .C(j), .Y(men_men_n1067_));
  NA4        u1039(.A(men_men_n1067_), .B(men_men_n1039_), .C(men_men_n329_), .D(men_men_n322_), .Y(men_men_n1068_));
  OAI210     u1040(.A0(men_men_n791_), .A1(men_men_n404_), .B0(men_men_n1068_), .Y(men_men_n1069_));
  NOi31      u1041(.An(m), .B(n), .C(f), .Y(men_men_n1070_));
  NA2        u1042(.A(men_men_n1070_), .B(men_men_n51_), .Y(men_men_n1071_));
  AN2        u1043(.A(e), .B(c), .Y(men_men_n1072_));
  NA2        u1044(.A(men_men_n1072_), .B(a), .Y(men_men_n1073_));
  OAI220     u1045(.A0(men_men_n1073_), .A1(men_men_n1071_), .B0(men_men_n855_), .B1(men_men_n410_), .Y(men_men_n1074_));
  NA2        u1046(.A(men_men_n484_), .B(l), .Y(men_men_n1075_));
  NOi31      u1047(.An(men_men_n835_), .B(men_men_n991_), .C(men_men_n1075_), .Y(men_men_n1076_));
  NO4        u1048(.A(men_men_n1076_), .B(men_men_n1074_), .C(men_men_n1069_), .D(men_men_n959_), .Y(men_men_n1077_));
  NO2        u1049(.A(men_men_n271_), .B(a), .Y(men_men_n1078_));
  INV        u1050(.A(men_men_n998_), .Y(men_men_n1079_));
  NO2        u1051(.A(men_men_n1048_), .B(men_men_n465_), .Y(men_men_n1080_));
  NO2        u1052(.A(men_men_n83_), .B(g), .Y(men_men_n1081_));
  AOI210     u1053(.A0(men_men_n1081_), .A1(men_men_n1080_), .B0(men_men_n1031_), .Y(men_men_n1082_));
  OR2        u1054(.A(men_men_n1082_), .B(men_men_n1029_), .Y(men_men_n1083_));
  NA3        u1055(.A(men_men_n1083_), .B(men_men_n1079_), .C(men_men_n1077_), .Y(men_men_n1084_));
  NO4        u1056(.A(men_men_n1084_), .B(men_men_n1066_), .C(men_men_n792_), .D(men_men_n540_), .Y(men_men_n1085_));
  NA2        u1057(.A(c), .B(b), .Y(men_men_n1086_));
  NO2        u1058(.A(men_men_n680_), .B(men_men_n1086_), .Y(men_men_n1087_));
  OAI210     u1059(.A0(men_men_n833_), .A1(men_men_n807_), .B0(men_men_n397_), .Y(men_men_n1088_));
  OAI210     u1060(.A0(men_men_n1088_), .A1(men_men_n834_), .B0(men_men_n1087_), .Y(men_men_n1089_));
  NAi21      u1061(.An(men_men_n405_), .B(men_men_n1087_), .Y(men_men_n1090_));
  NA3        u1062(.A(men_men_n411_), .B(men_men_n536_), .C(f), .Y(men_men_n1091_));
  OAI210     u1063(.A0(men_men_n527_), .A1(men_men_n39_), .B0(men_men_n1078_), .Y(men_men_n1092_));
  NA3        u1064(.A(men_men_n1092_), .B(men_men_n1091_), .C(men_men_n1090_), .Y(men_men_n1093_));
  OAI210     u1065(.A0(men_men_n109_), .A1(men_men_n275_), .B0(g), .Y(men_men_n1094_));
  NAi21      u1066(.An(f), .B(d), .Y(men_men_n1095_));
  NO2        u1067(.A(men_men_n1095_), .B(men_men_n1052_), .Y(men_men_n1096_));
  INV        u1068(.A(men_men_n1096_), .Y(men_men_n1097_));
  AOI210     u1069(.A0(men_men_n1094_), .A1(men_men_n281_), .B0(men_men_n1097_), .Y(men_men_n1098_));
  AOI210     u1070(.A0(men_men_n1098_), .A1(men_men_n105_), .B0(men_men_n1093_), .Y(men_men_n1099_));
  NA2        u1071(.A(men_men_n448_), .B(f), .Y(men_men_n1100_));
  NO2        u1072(.A(men_men_n173_), .B(men_men_n228_), .Y(men_men_n1101_));
  NA2        u1073(.A(men_men_n1101_), .B(m), .Y(men_men_n1102_));
  NA3        u1074(.A(men_men_n888_), .B(men_men_n1075_), .C(men_men_n451_), .Y(men_men_n1103_));
  OAI210     u1075(.A0(men_men_n1103_), .A1(men_men_n301_), .B0(men_men_n449_), .Y(men_men_n1104_));
  AOI210     u1076(.A0(men_men_n1104_), .A1(men_men_n1100_), .B0(men_men_n1102_), .Y(men_men_n1105_));
  NA2        u1077(.A(men_men_n538_), .B(men_men_n392_), .Y(men_men_n1106_));
  OAI210     u1078(.A0(men_men_n33_), .A1(men_men_n428_), .B0(men_men_n1096_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n356_), .B(men_men_n355_), .Y(men_men_n1108_));
  AOI210     u1080(.A0(men_men_n1101_), .A1(men_men_n413_), .B0(men_men_n924_), .Y(men_men_n1109_));
  NAi41      u1081(.An(men_men_n1108_), .B(men_men_n1109_), .C(men_men_n1107_), .D(men_men_n1106_), .Y(men_men_n1110_));
  NO2        u1082(.A(men_men_n1110_), .B(men_men_n1105_), .Y(men_men_n1111_));
  NA4        u1083(.A(men_men_n1111_), .B(men_men_n1099_), .C(men_men_n1089_), .D(men_men_n1085_), .Y(men00));
  AOI210     u1084(.A0(men_men_n288_), .A1(men_men_n205_), .B0(men_men_n264_), .Y(men_men_n1113_));
  NO2        u1085(.A(men_men_n1113_), .B(men_men_n554_), .Y(men_men_n1114_));
  AOI210     u1086(.A0(men_men_n868_), .A1(men_men_n913_), .B0(men_men_n1069_), .Y(men_men_n1115_));
  NO3        u1087(.A(men_men_n1045_), .B(men_men_n924_), .C(men_men_n691_), .Y(men_men_n1116_));
  NA3        u1088(.A(men_men_n1116_), .B(men_men_n1115_), .C(men_men_n960_), .Y(men_men_n1117_));
  NA2        u1089(.A(men_men_n486_), .B(f), .Y(men_men_n1118_));
  NO2        u1090(.A(men_men_n1118_), .B(men_men_n1001_), .Y(men_men_n1119_));
  NO4        u1091(.A(men_men_n1119_), .B(men_men_n1117_), .C(men_men_n1114_), .D(men_men_n1024_), .Y(men_men_n1120_));
  NA3        u1092(.A(men_men_n157_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1121_));
  NA3        u1093(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1122_));
  NOi31      u1094(.An(n), .B(m), .C(i), .Y(men_men_n1123_));
  NA3        u1095(.A(men_men_n1123_), .B(men_men_n628_), .C(men_men_n51_), .Y(men_men_n1124_));
  OAI210     u1096(.A0(men_men_n1122_), .A1(men_men_n1121_), .B0(men_men_n1124_), .Y(men_men_n1125_));
  INV        u1097(.A(men_men_n553_), .Y(men_men_n1126_));
  NO4        u1098(.A(men_men_n1126_), .B(men_men_n1125_), .C(men_men_n1108_), .D(men_men_n891_), .Y(men_men_n1127_));
  OR2        u1099(.A(men_men_n369_), .B(men_men_n127_), .Y(men_men_n1128_));
  NO2        u1100(.A(h), .B(g), .Y(men_men_n1129_));
  NA4        u1101(.A(men_men_n475_), .B(men_men_n446_), .C(men_men_n1129_), .D(men_men_n990_), .Y(men_men_n1130_));
  NA2        u1102(.A(men_men_n1130_), .B(men_men_n1128_), .Y(men_men_n1131_));
  NO2        u1103(.A(men_men_n1131_), .B(men_men_n256_), .Y(men_men_n1132_));
  INV        u1104(.A(men_men_n555_), .Y(men_men_n1133_));
  NA2        u1105(.A(men_men_n1133_), .B(men_men_n143_), .Y(men_men_n1134_));
  NO2        u1106(.A(men_men_n230_), .B(men_men_n172_), .Y(men_men_n1135_));
  NA2        u1107(.A(men_men_n1135_), .B(men_men_n411_), .Y(men_men_n1136_));
  NA3        u1108(.A(men_men_n170_), .B(men_men_n104_), .C(g), .Y(men_men_n1137_));
  NA3        u1109(.A(men_men_n446_), .B(men_men_n40_), .C(f), .Y(men_men_n1138_));
  NOi31      u1110(.An(men_men_n843_), .B(men_men_n1138_), .C(men_men_n1137_), .Y(men_men_n1139_));
  NAi31      u1111(.An(men_men_n177_), .B(men_men_n830_), .C(men_men_n446_), .Y(men_men_n1140_));
  NAi31      u1112(.An(men_men_n1139_), .B(men_men_n1140_), .C(men_men_n1136_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n263_), .B(men_men_n74_), .Y(men_men_n1142_));
  NO3        u1114(.A(men_men_n410_), .B(men_men_n803_), .C(n), .Y(men_men_n1143_));
  AOI210     u1115(.A0(men_men_n1143_), .A1(men_men_n1142_), .B0(men_men_n1038_), .Y(men_men_n1144_));
  NAi31      u1116(.An(men_men_n1004_), .B(men_men_n1144_), .C(men_men_n73_), .Y(men_men_n1145_));
  NO4        u1117(.A(men_men_n1145_), .B(men_men_n1141_), .C(men_men_n1134_), .D(men_men_n495_), .Y(men_men_n1146_));
  AN3        u1118(.A(men_men_n1146_), .B(men_men_n1132_), .C(men_men_n1127_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n513_), .B(men_men_n97_), .Y(men_men_n1148_));
  NA3        u1120(.A(men_men_n1070_), .B(men_men_n587_), .C(men_men_n445_), .Y(men_men_n1149_));
  NA4        u1121(.A(men_men_n1149_), .B(men_men_n539_), .C(men_men_n1148_), .D(men_men_n233_), .Y(men_men_n1150_));
  NA2        u1122(.A(men_men_n1063_), .B(men_men_n513_), .Y(men_men_n1151_));
  NA2        u1123(.A(men_men_n1151_), .B(men_men_n285_), .Y(men_men_n1152_));
  OAI210     u1124(.A0(men_men_n444_), .A1(men_men_n111_), .B0(men_men_n836_), .Y(men_men_n1153_));
  AOI220     u1125(.A0(men_men_n1153_), .A1(men_men_n1103_), .B0(men_men_n538_), .B1(men_men_n392_), .Y(men_men_n1154_));
  OR3        u1126(.A(men_men_n1001_), .B(men_men_n261_), .C(men_men_n214_), .Y(men_men_n1155_));
  NO2        u1127(.A(men_men_n208_), .B(men_men_n205_), .Y(men_men_n1156_));
  NA2        u1128(.A(men_men_n818_), .B(men_men_n1156_), .Y(men_men_n1157_));
  NA3        u1129(.A(men_men_n1157_), .B(men_men_n1155_), .C(men_men_n1154_), .Y(men_men_n1158_));
  INV        u1130(.A(men_men_n792_), .Y(men_men_n1159_));
  AOI220     u1131(.A0(men_men_n920_), .A1(men_men_n552_), .B0(men_men_n628_), .B1(men_men_n236_), .Y(men_men_n1160_));
  NO2        u1132(.A(men_men_n68_), .B(h), .Y(men_men_n1161_));
  NO3        u1133(.A(men_men_n1001_), .B(men_men_n999_), .C(men_men_n703_), .Y(men_men_n1162_));
  NO2        u1134(.A(men_men_n1035_), .B(men_men_n124_), .Y(men_men_n1163_));
  AN2        u1135(.A(men_men_n1163_), .B(men_men_n1050_), .Y(men_men_n1164_));
  OAI210     u1136(.A0(men_men_n1164_), .A1(men_men_n1162_), .B0(men_men_n1161_), .Y(men_men_n1165_));
  NA4        u1137(.A(men_men_n1165_), .B(men_men_n1160_), .C(men_men_n1159_), .D(men_men_n838_), .Y(men_men_n1166_));
  NO4        u1138(.A(men_men_n1166_), .B(men_men_n1158_), .C(men_men_n1152_), .D(men_men_n1150_), .Y(men_men_n1167_));
  NA2        u1139(.A(men_men_n808_), .B(men_men_n731_), .Y(men_men_n1168_));
  NA4        u1140(.A(men_men_n1168_), .B(men_men_n1167_), .C(men_men_n1147_), .D(men_men_n1120_), .Y(men01));
  AN2        u1141(.A(men_men_n981_), .B(men_men_n979_), .Y(men_men_n1170_));
  NO4        u1142(.A(men_men_n775_), .B(men_men_n767_), .C(men_men_n459_), .D(men_men_n269_), .Y(men_men_n1171_));
  NA2        u1143(.A(men_men_n379_), .B(i), .Y(men_men_n1172_));
  NA3        u1144(.A(men_men_n1172_), .B(men_men_n1171_), .C(men_men_n1170_), .Y(men_men_n1173_));
  NA2        u1145(.A(men_men_n565_), .B(men_men_n86_), .Y(men_men_n1174_));
  NA3        u1146(.A(men_men_n1174_), .B(men_men_n884_), .C(men_men_n321_), .Y(men_men_n1175_));
  NA2        u1147(.A(men_men_n45_), .B(f), .Y(men_men_n1176_));
  NA2        u1148(.A(men_men_n686_), .B(men_men_n92_), .Y(men_men_n1177_));
  NO2        u1149(.A(men_men_n1177_), .B(men_men_n1176_), .Y(men_men_n1178_));
  NO2        u1150(.A(men_men_n755_), .B(men_men_n582_), .Y(men_men_n1179_));
  AOI210     u1151(.A0(men_men_n1178_), .A1(men_men_n615_), .B0(men_men_n1179_), .Y(men_men_n1180_));
  INV        u1152(.A(men_men_n109_), .Y(men_men_n1181_));
  OR2        u1153(.A(men_men_n1181_), .B(men_men_n562_), .Y(men_men_n1182_));
  NA3        u1154(.A(men_men_n1182_), .B(men_men_n1180_), .C(men_men_n867_), .Y(men_men_n1183_));
  NO3        u1155(.A(men_men_n756_), .B(men_men_n653_), .C(men_men_n489_), .Y(men_men_n1184_));
  NA4        u1156(.A(men_men_n686_), .B(men_men_n92_), .C(men_men_n45_), .D(men_men_n204_), .Y(men_men_n1185_));
  OA220      u1157(.A0(men_men_n1185_), .A1(men_men_n646_), .B0(men_men_n187_), .B1(men_men_n185_), .Y(men_men_n1186_));
  NA3        u1158(.A(men_men_n1186_), .B(men_men_n1184_), .C(men_men_n130_), .Y(men_men_n1187_));
  NO4        u1159(.A(men_men_n1187_), .B(men_men_n1183_), .C(men_men_n1175_), .D(men_men_n1173_), .Y(men_men_n1188_));
  NA2        u1160(.A(men_men_n291_), .B(men_men_n508_), .Y(men_men_n1189_));
  AOI210     u1161(.A0(men_men_n196_), .A1(men_men_n85_), .B0(men_men_n204_), .Y(men_men_n1190_));
  OAI210     u1162(.A0(men_men_n782_), .A1(men_men_n411_), .B0(men_men_n1190_), .Y(men_men_n1191_));
  AN3        u1163(.A(m), .B(l), .C(k), .Y(men_men_n1192_));
  OAI210     u1164(.A0(men_men_n344_), .A1(men_men_n34_), .B0(men_men_n1192_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n195_), .B(men_men_n34_), .Y(men_men_n1194_));
  AO210      u1166(.A0(men_men_n1194_), .A1(men_men_n1193_), .B0(men_men_n320_), .Y(men_men_n1195_));
  NA3        u1167(.A(men_men_n1195_), .B(men_men_n1191_), .C(men_men_n1189_), .Y(men_men_n1196_));
  AOI210     u1168(.A0(men_men_n574_), .A1(men_men_n109_), .B0(men_men_n580_), .Y(men_men_n1197_));
  OAI210     u1169(.A0(men_men_n1181_), .A1(men_men_n571_), .B0(men_men_n1197_), .Y(men_men_n1198_));
  NO3        u1170(.A(men_men_n791_), .B(men_men_n196_), .C(men_men_n390_), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n1199_), .B(men_men_n924_), .Y(men_men_n1200_));
  OAI210     u1172(.A0(men_men_n1178_), .A1(men_men_n314_), .B0(men_men_n654_), .Y(men_men_n1201_));
  NA3        u1173(.A(men_men_n1201_), .B(men_men_n1200_), .C(men_men_n759_), .Y(men_men_n1202_));
  NO3        u1174(.A(men_men_n1202_), .B(men_men_n1198_), .C(men_men_n1196_), .Y(men_men_n1203_));
  NA3        u1175(.A(men_men_n583_), .B(men_men_n29_), .C(f), .Y(men_men_n1204_));
  NO2        u1176(.A(men_men_n1204_), .B(men_men_n196_), .Y(men_men_n1205_));
  AOI210     u1177(.A0(men_men_n481_), .A1(men_men_n58_), .B0(men_men_n1205_), .Y(men_men_n1206_));
  OR3        u1178(.A(men_men_n1177_), .B(men_men_n584_), .C(men_men_n1176_), .Y(men_men_n1207_));
  NO2        u1179(.A(men_men_n1185_), .B(men_men_n938_), .Y(men_men_n1208_));
  NO2        u1180(.A(men_men_n1208_), .B(men_men_n1125_), .Y(men_men_n1209_));
  NA4        u1181(.A(men_men_n1209_), .B(men_men_n1207_), .C(men_men_n1206_), .D(men_men_n730_), .Y(men_men_n1210_));
  NO2        u1182(.A(men_men_n929_), .B(men_men_n223_), .Y(men_men_n1211_));
  NO2        u1183(.A(men_men_n930_), .B(men_men_n533_), .Y(men_men_n1212_));
  OAI210     u1184(.A0(men_men_n1212_), .A1(men_men_n1211_), .B0(men_men_n327_), .Y(men_men_n1213_));
  NA2        u1185(.A(men_men_n547_), .B(men_men_n545_), .Y(men_men_n1214_));
  NA2        u1186(.A(men_men_n1214_), .B(men_men_n648_), .Y(men_men_n1215_));
  INV        u1187(.A(men_men_n371_), .Y(men_men_n1216_));
  NOi41      u1188(.An(men_men_n1213_), .B(men_men_n1216_), .C(men_men_n1215_), .D(men_men_n1210_), .Y(men_men_n1217_));
  NO2        u1189(.A(men_men_n123_), .B(men_men_n45_), .Y(men_men_n1218_));
  NO2        u1190(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1219_));
  AO220      u1191(.A0(men_men_n1219_), .A1(men_men_n603_), .B0(men_men_n1218_), .B1(men_men_n684_), .Y(men_men_n1220_));
  NA2        u1192(.A(men_men_n1220_), .B(men_men_n327_), .Y(men_men_n1221_));
  NO3        u1193(.A(men_men_n1048_), .B(men_men_n167_), .C(men_men_n83_), .Y(men_men_n1222_));
  INV        u1194(.A(men_men_n1221_), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n595_), .B(men_men_n594_), .Y(men_men_n1224_));
  NO4        u1196(.A(men_men_n1048_), .B(men_men_n1224_), .C(men_men_n165_), .D(men_men_n83_), .Y(men_men_n1225_));
  NO3        u1197(.A(men_men_n1225_), .B(men_men_n1223_), .C(men_men_n619_), .Y(men_men_n1226_));
  NA4        u1198(.A(men_men_n1226_), .B(men_men_n1217_), .C(men_men_n1203_), .D(men_men_n1188_), .Y(men06));
  NO2        u1199(.A(men_men_n391_), .B(men_men_n537_), .Y(men_men_n1228_));
  NA2        u1200(.A(men_men_n257_), .B(men_men_n1228_), .Y(men_men_n1229_));
  NO2        u1201(.A(men_men_n215_), .B(men_men_n99_), .Y(men_men_n1230_));
  OAI210     u1202(.A0(men_men_n1230_), .A1(men_men_n1222_), .B0(men_men_n367_), .Y(men_men_n1231_));
  NO3        u1203(.A(men_men_n578_), .B(men_men_n780_), .C(men_men_n581_), .Y(men_men_n1232_));
  OR2        u1204(.A(men_men_n1232_), .B(men_men_n855_), .Y(men_men_n1233_));
  NA4        u1205(.A(men_men_n1233_), .B(men_men_n1231_), .C(men_men_n1229_), .D(men_men_n1213_), .Y(men_men_n1234_));
  NO3        u1206(.A(men_men_n1234_), .B(men_men_n1215_), .C(men_men_n245_), .Y(men_men_n1235_));
  INV        u1207(.A(men_men_n1211_), .Y(men_men_n1236_));
  INV        u1208(.A(men_men_n1220_), .Y(men_men_n1237_));
  AOI210     u1209(.A0(men_men_n1237_), .A1(men_men_n1236_), .B0(men_men_n324_), .Y(men_men_n1238_));
  INV        u1210(.A(men_men_n652_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n1239_), .B(men_men_n623_), .Y(men_men_n1240_));
  NO2        u1212(.A(men_men_n491_), .B(men_men_n162_), .Y(men_men_n1241_));
  NOi21      u1213(.An(men_men_n129_), .B(men_men_n45_), .Y(men_men_n1242_));
  NO2        u1214(.A(men_men_n588_), .B(men_men_n1071_), .Y(men_men_n1243_));
  INV        u1215(.A(men_men_n878_), .Y(men_men_n1244_));
  NO4        u1216(.A(men_men_n1244_), .B(men_men_n1243_), .C(men_men_n1242_), .D(men_men_n1241_), .Y(men_men_n1245_));
  OR2        u1217(.A(men_men_n579_), .B(men_men_n577_), .Y(men_men_n1246_));
  INV        u1218(.A(men_men_n1246_), .Y(men_men_n1247_));
  NA3        u1219(.A(men_men_n1247_), .B(men_men_n1245_), .C(men_men_n1240_), .Y(men_men_n1248_));
  NO2        u1220(.A(men_men_n723_), .B(men_men_n352_), .Y(men_men_n1249_));
  NO3        u1221(.A(men_men_n654_), .B(men_men_n732_), .C(men_men_n615_), .Y(men_men_n1250_));
  NOi21      u1222(.An(men_men_n1249_), .B(men_men_n1250_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n1251_), .B(men_men_n1248_), .C(men_men_n1238_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n774_), .B(men_men_n265_), .Y(men_men_n1253_));
  OAI220     u1225(.A0(men_men_n710_), .A1(men_men_n47_), .B0(men_men_n215_), .B1(men_men_n597_), .Y(men_men_n1254_));
  OAI210     u1226(.A0(men_men_n265_), .A1(c), .B0(men_men_n622_), .Y(men_men_n1255_));
  AOI220     u1227(.A0(men_men_n1255_), .A1(men_men_n1254_), .B0(men_men_n1253_), .B1(men_men_n257_), .Y(men_men_n1256_));
  NO3        u1228(.A(men_men_n235_), .B(men_men_n99_), .C(men_men_n271_), .Y(men_men_n1257_));
  OAI220     u1229(.A0(men_men_n677_), .A1(men_men_n238_), .B0(men_men_n488_), .B1(men_men_n491_), .Y(men_men_n1258_));
  NO3        u1230(.A(men_men_n1258_), .B(men_men_n1257_), .C(men_men_n1074_), .Y(men_men_n1259_));
  NA4        u1231(.A(men_men_n765_), .B(men_men_n764_), .C(men_men_n421_), .D(men_men_n849_), .Y(men_men_n1260_));
  NAi31      u1232(.An(men_men_n723_), .B(men_men_n1260_), .C(men_men_n195_), .Y(men_men_n1261_));
  NA4        u1233(.A(men_men_n1261_), .B(men_men_n1259_), .C(men_men_n1256_), .D(men_men_n1160_), .Y(men_men_n1262_));
  OR2        u1234(.A(men_men_n755_), .B(men_men_n519_), .Y(men_men_n1263_));
  OR3        u1235(.A(men_men_n355_), .B(men_men_n215_), .C(men_men_n597_), .Y(men_men_n1264_));
  AOI210     u1236(.A0(men_men_n547_), .A1(men_men_n430_), .B0(men_men_n357_), .Y(men_men_n1265_));
  NA3        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .C(men_men_n1263_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n1249_), .B(men_men_n731_), .Y(men_men_n1267_));
  AN2        u1239(.A(men_men_n899_), .B(men_men_n898_), .Y(men_men_n1268_));
  NO4        u1240(.A(men_men_n1268_), .B(men_men_n847_), .C(men_men_n477_), .D(men_men_n462_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n1267_), .Y(men_men_n1270_));
  NAi21      u1242(.An(j), .B(i), .Y(men_men_n1271_));
  NO4        u1243(.A(men_men_n1224_), .B(men_men_n1271_), .C(men_men_n424_), .D(men_men_n226_), .Y(men_men_n1272_));
  NO4        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n1266_), .D(men_men_n1262_), .Y(men_men_n1273_));
  NA4        u1245(.A(men_men_n1273_), .B(men_men_n1252_), .C(men_men_n1235_), .D(men_men_n1226_), .Y(men07));
  NAi32      u1246(.An(m), .Bn(b), .C(n), .Y(men_men_n1275_));
  NO3        u1247(.A(men_men_n1275_), .B(g), .C(f), .Y(men_men_n1276_));
  OAI210     u1248(.A0(men_men_n309_), .A1(men_men_n464_), .B0(men_men_n1276_), .Y(men_men_n1277_));
  NAi21      u1249(.An(f), .B(c), .Y(men_men_n1278_));
  OR2        u1250(.A(e), .B(d), .Y(men_men_n1279_));
  NOi31      u1251(.An(n), .B(m), .C(b), .Y(men_men_n1280_));
  NO3        u1252(.A(men_men_n124_), .B(men_men_n431_), .C(h), .Y(men_men_n1281_));
  INV        u1253(.A(men_men_n1277_), .Y(men_men_n1282_));
  NOi41      u1254(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1283_));
  NA3        u1255(.A(men_men_n1283_), .B(men_men_n840_), .C(men_men_n393_), .Y(men_men_n1284_));
  NO2        u1256(.A(men_men_n1284_), .B(men_men_n56_), .Y(men_men_n1285_));
  NA2        u1257(.A(men_men_n1050_), .B(men_men_n212_), .Y(men_men_n1286_));
  NO2        u1258(.A(men_men_n1286_), .B(men_men_n61_), .Y(men_men_n1287_));
  NA2        u1259(.A(men_men_n83_), .B(men_men_n45_), .Y(men_men_n1288_));
  NO2        u1260(.A(men_men_n1007_), .B(men_men_n424_), .Y(men_men_n1289_));
  NA3        u1261(.A(men_men_n1289_), .B(men_men_n1288_), .C(men_men_n205_), .Y(men_men_n1290_));
  NO2        u1262(.A(men_men_n1021_), .B(men_men_n296_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n1161_), .B(men_men_n279_), .Y(men_men_n1292_));
  NA2        u1264(.A(men_men_n1292_), .B(men_men_n1290_), .Y(men_men_n1293_));
  NO4        u1265(.A(men_men_n1293_), .B(men_men_n1287_), .C(men_men_n1285_), .D(men_men_n1282_), .Y(men_men_n1294_));
  NO3        u1266(.A(e), .B(d), .C(c), .Y(men_men_n1295_));
  OAI210     u1267(.A0(men_men_n124_), .A1(men_men_n205_), .B0(men_men_n585_), .Y(men_men_n1296_));
  NA2        u1268(.A(men_men_n1296_), .B(men_men_n1295_), .Y(men_men_n1297_));
  INV        u1269(.A(men_men_n1297_), .Y(men_men_n1298_));
  OR2        u1270(.A(h), .B(f), .Y(men_men_n1299_));
  NO3        u1271(.A(n), .B(m), .C(i), .Y(men_men_n1300_));
  OAI210     u1272(.A0(men_men_n1072_), .A1(men_men_n146_), .B0(men_men_n1300_), .Y(men_men_n1301_));
  NO2        u1273(.A(i), .B(g), .Y(men_men_n1302_));
  OR3        u1274(.A(men_men_n1302_), .B(men_men_n1275_), .C(men_men_n71_), .Y(men_men_n1303_));
  OAI220     u1275(.A0(men_men_n1303_), .A1(men_men_n464_), .B0(men_men_n1301_), .B1(men_men_n1299_), .Y(men_men_n1304_));
  NA3        u1276(.A(men_men_n674_), .B(men_men_n662_), .C(men_men_n104_), .Y(men_men_n1305_));
  NA3        u1277(.A(men_men_n1280_), .B(men_men_n1016_), .C(men_men_n650_), .Y(men_men_n1306_));
  AOI210     u1278(.A0(men_men_n1306_), .A1(men_men_n1305_), .B0(men_men_n45_), .Y(men_men_n1307_));
  NA2        u1279(.A(men_men_n1300_), .B(men_men_n621_), .Y(men_men_n1308_));
  NO2        u1280(.A(l), .B(k), .Y(men_men_n1309_));
  NO3        u1281(.A(men_men_n424_), .B(d), .C(c), .Y(men_men_n1310_));
  NO3        u1282(.A(men_men_n1307_), .B(men_men_n1304_), .C(men_men_n1298_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n137_), .B(h), .Y(men_men_n1312_));
  NO2        u1284(.A(men_men_n1030_), .B(l), .Y(men_men_n1313_));
  NO2        u1285(.A(g), .B(c), .Y(men_men_n1314_));
  NA3        u1286(.A(men_men_n1314_), .B(men_men_n134_), .C(men_men_n178_), .Y(men_men_n1315_));
  NO2        u1287(.A(men_men_n1315_), .B(men_men_n1313_), .Y(men_men_n1316_));
  NA2        u1288(.A(men_men_n1316_), .B(men_men_n170_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n432_), .B(a), .Y(men_men_n1318_));
  NA3        u1290(.A(men_men_n1318_), .B(k), .C(men_men_n105_), .Y(men_men_n1319_));
  NO2        u1291(.A(i), .B(h), .Y(men_men_n1320_));
  NA2        u1292(.A(men_men_n1320_), .B(men_men_n212_), .Y(men_men_n1321_));
  NA2        u1293(.A(men_men_n1095_), .B(h), .Y(men_men_n1322_));
  NA2        u1294(.A(men_men_n131_), .B(men_men_n212_), .Y(men_men_n1323_));
  AOI210     u1295(.A0(men_men_n246_), .A1(men_men_n107_), .B0(men_men_n508_), .Y(men_men_n1324_));
  OAI220     u1296(.A0(men_men_n1324_), .A1(men_men_n1321_), .B0(men_men_n1323_), .B1(men_men_n1322_), .Y(men_men_n1325_));
  NO2        u1297(.A(men_men_n728_), .B(men_men_n179_), .Y(men_men_n1326_));
  NOi31      u1298(.An(m), .B(n), .C(b), .Y(men_men_n1327_));
  NOi31      u1299(.An(f), .B(d), .C(c), .Y(men_men_n1328_));
  NA2        u1300(.A(men_men_n1328_), .B(men_men_n1327_), .Y(men_men_n1329_));
  INV        u1301(.A(men_men_n1329_), .Y(men_men_n1330_));
  NO3        u1302(.A(men_men_n1330_), .B(men_men_n1326_), .C(men_men_n1325_), .Y(men_men_n1331_));
  NA2        u1303(.A(men_men_n1041_), .B(men_men_n446_), .Y(men_men_n1332_));
  OAI210     u1304(.A0(men_men_n173_), .A1(men_men_n503_), .B0(men_men_n1017_), .Y(men_men_n1333_));
  NO3        u1305(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1334_));
  AN4        u1306(.A(men_men_n1333_), .B(men_men_n1331_), .C(men_men_n1319_), .D(men_men_n1317_), .Y(men_men_n1335_));
  NA2        u1307(.A(men_men_n1280_), .B(men_men_n364_), .Y(men_men_n1336_));
  NA2        u1308(.A(men_men_n1310_), .B(men_men_n206_), .Y(men_men_n1337_));
  NA2        u1309(.A(men_men_n1049_), .B(men_men_n1332_), .Y(men_men_n1338_));
  NO2        u1310(.A(i), .B(men_men_n204_), .Y(men_men_n1339_));
  NA4        u1311(.A(men_men_n1101_), .B(men_men_n1339_), .C(men_men_n100_), .D(m), .Y(men_men_n1340_));
  NA3        u1312(.A(men_men_n1340_), .B(men_men_n1338_), .C(men_men_n1337_), .Y(men_men_n1341_));
  NO4        u1313(.A(men_men_n124_), .B(g), .C(f), .D(e), .Y(men_men_n1342_));
  NA2        u1314(.A(men_men_n280_), .B(h), .Y(men_men_n1343_));
  NA2        u1315(.A(men_men_n186_), .B(men_men_n94_), .Y(men_men_n1344_));
  NA2        u1316(.A(men_men_n30_), .B(h), .Y(men_men_n1345_));
  NO2        u1317(.A(men_men_n1345_), .B(men_men_n1037_), .Y(men_men_n1346_));
  NOi41      u1318(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1347_));
  NA2        u1319(.A(men_men_n1347_), .B(men_men_n105_), .Y(men_men_n1348_));
  NA2        u1320(.A(men_men_n1283_), .B(men_men_n1309_), .Y(men_men_n1349_));
  NA2        u1321(.A(men_men_n1349_), .B(men_men_n1348_), .Y(men_men_n1350_));
  OR3        u1322(.A(men_men_n519_), .B(men_men_n518_), .C(men_men_n104_), .Y(men_men_n1351_));
  NA2        u1323(.A(men_men_n1070_), .B(men_men_n390_), .Y(men_men_n1352_));
  OAI220     u1324(.A0(men_men_n1352_), .A1(men_men_n420_), .B0(men_men_n1351_), .B1(men_men_n289_), .Y(men_men_n1353_));
  AO210      u1325(.A0(men_men_n1353_), .A1(men_men_n107_), .B0(men_men_n1350_), .Y(men_men_n1354_));
  NO3        u1326(.A(men_men_n1354_), .B(men_men_n1346_), .C(men_men_n1341_), .Y(men_men_n1355_));
  NA4        u1327(.A(men_men_n1355_), .B(men_men_n1335_), .C(men_men_n1311_), .D(men_men_n1294_), .Y(men_men_n1356_));
  NA2        u1328(.A(men_men_n364_), .B(men_men_n56_), .Y(men_men_n1357_));
  AOI210     u1329(.A0(men_men_n1357_), .A1(men_men_n1007_), .B0(men_men_n1308_), .Y(men_men_n1358_));
  NA2        u1330(.A(men_men_n206_), .B(men_men_n170_), .Y(men_men_n1359_));
  AOI210     u1331(.A0(men_men_n1359_), .A1(men_men_n1137_), .B0(men_men_n1357_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n1042_), .B(men_men_n1037_), .Y(men_men_n1361_));
  NO3        u1333(.A(men_men_n1361_), .B(men_men_n1360_), .C(men_men_n1358_), .Y(men_men_n1362_));
  NO2        u1334(.A(men_men_n376_), .B(j), .Y(men_men_n1363_));
  NA3        u1335(.A(men_men_n1334_), .B(men_men_n1279_), .C(men_men_n1070_), .Y(men_men_n1364_));
  NAi41      u1336(.An(men_men_n1320_), .B(men_men_n1028_), .C(men_men_n158_), .D(e), .Y(men_men_n1365_));
  NA2        u1337(.A(men_men_n1365_), .B(men_men_n1364_), .Y(men_men_n1366_));
  NA3        u1338(.A(g), .B(men_men_n1363_), .C(men_men_n148_), .Y(men_men_n1367_));
  INV        u1339(.A(men_men_n1367_), .Y(men_men_n1368_));
  NO3        u1340(.A(men_men_n723_), .B(men_men_n165_), .C(men_men_n393_), .Y(men_men_n1369_));
  NO3        u1341(.A(men_men_n1369_), .B(men_men_n1368_), .C(men_men_n1366_), .Y(men_men_n1370_));
  NO3        u1342(.A(men_men_n1037_), .B(men_men_n559_), .C(g), .Y(men_men_n1371_));
  NOi21      u1343(.An(men_men_n1359_), .B(men_men_n1371_), .Y(men_men_n1372_));
  AOI210     u1344(.A0(men_men_n1372_), .A1(men_men_n1344_), .B0(men_men_n1007_), .Y(men_men_n1373_));
  OR2        u1345(.A(n), .B(i), .Y(men_men_n1374_));
  OAI210     u1346(.A0(men_men_n1374_), .A1(men_men_n1027_), .B0(men_men_n49_), .Y(men_men_n1375_));
  AOI220     u1347(.A0(men_men_n1375_), .A1(men_men_n1129_), .B0(men_men_n795_), .B1(men_men_n186_), .Y(men_men_n1376_));
  INV        u1348(.A(men_men_n1376_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n215_), .B(k), .Y(men_men_n1378_));
  NO2        u1350(.A(men_men_n1377_), .B(men_men_n1373_), .Y(men_men_n1379_));
  INV        u1351(.A(men_men_n49_), .Y(men_men_n1380_));
  NO3        u1352(.A(men_men_n1052_), .B(men_men_n1279_), .C(men_men_n49_), .Y(men_men_n1381_));
  NA2        u1353(.A(men_men_n1053_), .B(men_men_n1380_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n1037_), .B(h), .Y(men_men_n1383_));
  NA3        u1355(.A(men_men_n1383_), .B(d), .C(men_men_n999_), .Y(men_men_n1384_));
  OAI220     u1356(.A0(men_men_n1384_), .A1(c), .B0(men_men_n1382_), .B1(j), .Y(men_men_n1385_));
  AOI210     u1357(.A0(men_men_n503_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1386_));
  NA2        u1358(.A(men_men_n1386_), .B(men_men_n1318_), .Y(men_men_n1387_));
  NO2        u1359(.A(men_men_n1271_), .B(men_men_n165_), .Y(men_men_n1388_));
  NOi21      u1360(.An(d), .B(f), .Y(men_men_n1389_));
  NO3        u1361(.A(men_men_n1328_), .B(men_men_n1389_), .C(men_men_n40_), .Y(men_men_n1390_));
  NA2        u1362(.A(men_men_n1390_), .B(men_men_n1388_), .Y(men_men_n1391_));
  NO2        u1363(.A(men_men_n1279_), .B(f), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n289_), .B(c), .Y(men_men_n1393_));
  NA2        u1365(.A(men_men_n1393_), .B(men_men_n520_), .Y(men_men_n1394_));
  NA3        u1366(.A(men_men_n1394_), .B(men_men_n1391_), .C(men_men_n1387_), .Y(men_men_n1395_));
  NO2        u1367(.A(men_men_n1395_), .B(men_men_n1385_), .Y(men_men_n1396_));
  NA4        u1368(.A(men_men_n1396_), .B(men_men_n1379_), .C(men_men_n1370_), .D(men_men_n1362_), .Y(men_men_n1397_));
  NO3        u1369(.A(men_men_n1041_), .B(men_men_n1027_), .C(men_men_n40_), .Y(men_men_n1398_));
  NO2        u1370(.A(men_men_n446_), .B(men_men_n289_), .Y(men_men_n1399_));
  OAI210     u1371(.A0(men_men_n1399_), .A1(men_men_n1398_), .B0(men_men_n1291_), .Y(men_men_n1400_));
  OAI210     u1372(.A0(men_men_n1342_), .A1(men_men_n1280_), .B0(men_men_n852_), .Y(men_men_n1401_));
  NO2        u1373(.A(men_men_n996_), .B(men_men_n124_), .Y(men_men_n1402_));
  NA2        u1374(.A(men_men_n1402_), .B(men_men_n602_), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1403_), .B(men_men_n1401_), .C(men_men_n1400_), .Y(men_men_n1404_));
  NA2        u1376(.A(men_men_n1314_), .B(men_men_n1389_), .Y(men_men_n1405_));
  NO2        u1377(.A(men_men_n1405_), .B(m), .Y(men_men_n1406_));
  NA3        u1378(.A(men_men_n1050_), .B(men_men_n101_), .C(men_men_n212_), .Y(men_men_n1407_));
  NO2        u1379(.A(men_men_n140_), .B(men_men_n172_), .Y(men_men_n1408_));
  OAI210     u1380(.A0(men_men_n1408_), .A1(men_men_n102_), .B0(men_men_n1327_), .Y(men_men_n1409_));
  NA2        u1381(.A(men_men_n1409_), .B(men_men_n1407_), .Y(men_men_n1410_));
  NO3        u1382(.A(men_men_n1410_), .B(men_men_n1406_), .C(men_men_n1404_), .Y(men_men_n1411_));
  NO2        u1383(.A(men_men_n1278_), .B(e), .Y(men_men_n1412_));
  NA2        u1384(.A(men_men_n1412_), .B(men_men_n388_), .Y(men_men_n1413_));
  OAI210     u1385(.A0(men_men_n1392_), .A1(men_men_n1081_), .B0(men_men_n613_), .Y(men_men_n1414_));
  OR3        u1386(.A(men_men_n1378_), .B(men_men_n1161_), .C(men_men_n124_), .Y(men_men_n1415_));
  OAI220     u1387(.A0(men_men_n1415_), .A1(men_men_n1413_), .B0(men_men_n1414_), .B1(men_men_n426_), .Y(men_men_n1416_));
  NO3        u1388(.A(men_men_n1351_), .B(men_men_n340_), .C(a), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n1417_), .B(men_men_n1416_), .Y(men_men_n1418_));
  NO2        u1390(.A(men_men_n172_), .B(c), .Y(men_men_n1419_));
  OAI210     u1391(.A0(men_men_n1419_), .A1(men_men_n1412_), .B0(men_men_n170_), .Y(men_men_n1420_));
  AOI220     u1392(.A0(men_men_n1420_), .A1(men_men_n1029_), .B0(men_men_n510_), .B1(men_men_n352_), .Y(men_men_n1421_));
  NA2        u1393(.A(men_men_n518_), .B(g), .Y(men_men_n1422_));
  AOI210     u1394(.A0(men_men_n1422_), .A1(men_men_n1310_), .B0(men_men_n1381_), .Y(men_men_n1423_));
  NO2        u1395(.A(men_men_n1423_), .B(men_men_n204_), .Y(men_men_n1424_));
  OR2        u1396(.A(h), .B(men_men_n518_), .Y(men_men_n1425_));
  NO2        u1397(.A(men_men_n1425_), .B(men_men_n165_), .Y(men_men_n1426_));
  NA2        u1398(.A(men_men_n1281_), .B(men_men_n173_), .Y(men_men_n1427_));
  NO2        u1399(.A(men_men_n49_), .B(l), .Y(men_men_n1428_));
  INV        u1400(.A(men_men_n464_), .Y(men_men_n1429_));
  OAI210     u1401(.A0(men_men_n1429_), .A1(men_men_n1053_), .B0(men_men_n1428_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n241_), .B(g), .Y(men_men_n1431_));
  NO2        u1403(.A(m), .B(i), .Y(men_men_n1432_));
  BUFFER     u1404(.A(men_men_n1432_), .Y(men_men_n1433_));
  AOI220     u1405(.A0(men_men_n1433_), .A1(men_men_n1312_), .B0(men_men_n1028_), .B1(men_men_n1431_), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1434_), .B(men_men_n1430_), .C(men_men_n1427_), .Y(men_men_n1435_));
  NO4        u1407(.A(men_men_n1435_), .B(men_men_n1426_), .C(men_men_n1424_), .D(men_men_n1421_), .Y(men_men_n1436_));
  NA3        u1408(.A(men_men_n1436_), .B(men_men_n1418_), .C(men_men_n1411_), .Y(men_men_n1437_));
  NA3        u1409(.A(men_men_n926_), .B(men_men_n131_), .C(men_men_n46_), .Y(men_men_n1438_));
  INV        u1410(.A(men_men_n176_), .Y(men_men_n1439_));
  NA2        u1411(.A(men_men_n1439_), .B(men_men_n1383_), .Y(men_men_n1440_));
  AO210      u1412(.A0(men_men_n125_), .A1(l), .B0(men_men_n1336_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n71_), .B(c), .Y(men_men_n1442_));
  NO4        u1414(.A(men_men_n1299_), .B(men_men_n177_), .C(men_men_n431_), .D(men_men_n45_), .Y(men_men_n1443_));
  AOI210     u1415(.A0(men_men_n1388_), .A1(men_men_n1442_), .B0(men_men_n1443_), .Y(men_men_n1444_));
  NA3        u1416(.A(men_men_n1444_), .B(men_men_n1441_), .C(men_men_n1440_), .Y(men_men_n1445_));
  INV        u1417(.A(men_men_n1445_), .Y(men_men_n1446_));
  NO4        u1418(.A(men_men_n215_), .B(men_men_n177_), .C(men_men_n246_), .D(k), .Y(men_men_n1447_));
  NO2        u1419(.A(men_men_n1438_), .B(men_men_n102_), .Y(men_men_n1448_));
  NOi21      u1420(.An(men_men_n1281_), .B(e), .Y(men_men_n1449_));
  NO3        u1421(.A(men_men_n1449_), .B(men_men_n1448_), .C(men_men_n1447_), .Y(men_men_n1450_));
  AN2        u1422(.A(men_men_n1050_), .B(men_men_n1035_), .Y(men_men_n1451_));
  AOI220     u1423(.A0(men_men_n1432_), .A1(men_men_n621_), .B0(men_men_n1013_), .B1(men_men_n149_), .Y(men_men_n1452_));
  NOi31      u1424(.An(men_men_n30_), .B(men_men_n1452_), .C(n), .Y(men_men_n1453_));
  AOI210     u1425(.A0(men_men_n1451_), .A1(men_men_n1123_), .B0(men_men_n1453_), .Y(men_men_n1454_));
  NA3        u1426(.A(men_men_n1454_), .B(men_men_n1450_), .C(men_men_n1446_), .Y(men_men_n1455_));
  OR4        u1427(.A(men_men_n1455_), .B(men_men_n1437_), .C(men_men_n1397_), .D(men_men_n1356_), .Y(men04));
  NOi31      u1428(.An(men_men_n1342_), .B(men_men_n1343_), .C(men_men_n1001_), .Y(men_men_n1457_));
  NA2        u1429(.A(men_men_n1392_), .B(men_men_n795_), .Y(men_men_n1458_));
  NO4        u1430(.A(men_men_n1458_), .B(men_men_n991_), .C(men_men_n465_), .D(j), .Y(men_men_n1459_));
  OR3        u1431(.A(men_men_n1459_), .B(men_men_n1457_), .C(men_men_n1019_), .Y(men_men_n1460_));
  NO3        u1432(.A(men_men_n1288_), .B(men_men_n87_), .C(k), .Y(men_men_n1461_));
  AOI210     u1433(.A0(men_men_n1461_), .A1(men_men_n1012_), .B0(men_men_n1139_), .Y(men_men_n1462_));
  NA2        u1434(.A(men_men_n1462_), .B(men_men_n1165_), .Y(men_men_n1463_));
  NO3        u1435(.A(men_men_n1463_), .B(men_men_n1460_), .C(men_men_n1006_), .Y(men_men_n1464_));
  NA4        u1436(.A(men_men_n1464_), .B(men_men_n1083_), .C(men_men_n1068_), .D(men_men_n1056_), .Y(men05));
  INV        u1437(.A(c), .Y(men_men_n1468_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule