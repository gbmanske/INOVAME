module tb_alu_32bit;

    reg [31:0] A, B;
    reg [2:0] ALUOp;
    wire [31:0] Result;
    wire Overflow, Zero, Negative;

    // Instância da ALU
    ula uut (
        .a(A),
        .b(B),
        .sel(ALUOp),
        .s(Result),
        .fov(Overflow),
        .fz(Zero),
        .fn(Negative)
    );

    initial begin
        // Teste AND
        $display("Teste AND");
        A = 32'hFFFFFFFF; B = 32'h0000FFFF; ALUOp = 3'b000; #10;
        $display("AND: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);
        A = 32'h00000000; B = 32'hFFFFFFFF; ALUOp = 3'b000; #10;
        $display("AND: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Teste OR
        $display("Teste OR");
        A = 32'h0000F0F0; B = 32'h0F0F0000; ALUOp = 3'b001; #10;
        $display("OR: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);
        A = 32'h00000000; B = 32'h00000000; ALUOp = 3'b001; #10;
        $display("OR: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Teste Soma
        $display("Teste Soma");
        A = 32'h7FFFFFFF; B = 32'h00000001; ALUOp = 3'b010; #10;
        $display("ADD: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);
        A = 32'h80000000; B = 32'hFFFFFFFF; ALUOp = 3'b010; #10;
        $display("ADD: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Teste Subtração
        $display("Teste Subtração");
        A = 32'h80000000; B = 32'h00000001; ALUOp = 3'b110; #10;
        $display("SUB: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);
        A = 32'h7FFFFFFF; B = 32'hFFFFFFFF; ALUOp = 3'b110; #10;
        $display("SUB: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Teste A AND !B
        $display("Teste A AND !B");
        A = 32'hFFFF0000; B = 32'h0000FFFF; ALUOp = 3'b100; #10;
        $display("A AND !B: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Teste A OR !B
        $display("Teste A OR !B");
        A = 32'h0F0F0F0F; B = 32'hF0F0F0F0; ALUOp = 3'b101; #10;
        $display("A OR !B: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Teste SLT
        $display("Teste SLT");
        A = 32'h00000001; B = 32'h00000002; ALUOp = 3'b111; #10;
        $display("SLT: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);
        A = 32'hFFFFFFFF; B = 32'h00000000; ALUOp = 3'b111; #10;
        $display("SLT: A=%h, B=%h, Result=%h, Overflow=%b, Zero=%b, Negative=%b", A, B, Result, Overflow, Zero, Negative);

        // Finaliza a simulação
        $stop;
    end

endmodule
