// Benchmark "top" written by ABC on Thu Jun 20 14:00:09 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n781_,
    new_new_n782_, new_new_n783_, new_new_n784_, new_new_n785_,
    new_new_n786_, new_new_n787_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1109_, new_new_n1110_, new_new_n1111_,
    new_new_n1112_, new_new_n1113_, new_new_n1114_, new_new_n1115_,
    new_new_n1116_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  OR4        g0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g0066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  AOI210     g0067(.A0(new_new_n88_), .A1(new_new_n86_), .B0(new_new_n89_), .Y(new_new_n90_));
  OAI210     g0068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g0069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g0070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g0072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g0073(.A(new_new_n95_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g0074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g0075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n98_));
  AN3        g0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g0077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g0078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g0079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  NA2        g0080(.A(new_new_n102_), .B(new_new_n62_), .Y(new_new_n103_));
  INV        g0081(.A(i_7_), .Y(new_new_n104_));
  NA2        g0082(.A(new_new_n46_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g0083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g0084(.A(new_new_n106_), .B(new_new_n86_), .Y(new_new_n107_));
  NA2        g0085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  NAi21      g0086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g0087(.A(new_new_n109_), .B(new_new_n92_), .C(new_new_n53_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  OR2        g0089(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n112_));
  NO2        g0090(.A(i_8_), .B(new_new_n104_), .Y(new_new_n113_));
  NA2        g0091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g0093(.A(new_new_n115_), .B(i_0_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  OAI210     g0095(.A0(new_new_n116_), .A1(new_new_n114_), .B0(new_new_n117_), .Y(new_new_n118_));
  INV        g0096(.A(new_new_n118_), .Y(new_new_n119_));
  NAi31      g0097(.An(new_new_n110_), .B(new_new_n119_), .C(new_new_n103_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n46_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NO2        g0107(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n86_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n47_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n109_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n98_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g0127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g0128(.A(new_new_n150_), .B(new_new_n25_), .Y(new_new_n151_));
  AN2        g0129(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g0131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n155_));
  NA2        g0133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g0135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g0138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g0139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n39_), .Y(new_new_n163_));
  NO2        g0141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g0142(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g0144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  AOI210     g0146(.A0(new_new_n168_), .A1(new_new_n151_), .B0(new_new_n143_), .Y(new_new_n169_));
  NA3        g0147(.A(new_new_n73_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n48_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  OR2        g0152(.A(new_new_n174_), .B(new_new_n171_), .Y(new_new_n175_));
  NO2        g0153(.A(i_4_), .B(i_5_), .Y(new_new_n176_));
  NAi21      g0154(.An(i_12_), .B(i_11_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n177_), .B(i_13_), .Y(new_new_n178_));
  NA3        g0156(.A(new_new_n178_), .B(new_new_n176_), .C(new_new_n83_), .Y(new_new_n179_));
  AOI210     g0157(.A0(new_new_n179_), .A1(new_new_n175_), .B0(new_new_n170_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n181_), .B(new_new_n46_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NAi31      g0161(.An(new_new_n183_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n184_));
  NA2        g0162(.A(i_3_), .B(i_5_), .Y(new_new_n185_));
  OR2        g0163(.A(new_new_n185_), .B(new_new_n174_), .Y(new_new_n186_));
  AOI210     g0164(.A0(new_new_n186_), .A1(new_new_n184_), .B0(new_new_n182_), .Y(new_new_n187_));
  NO2        g0165(.A(new_new_n73_), .B(i_5_), .Y(new_new_n188_));
  NO2        g0166(.A(i_13_), .B(i_10_), .Y(new_new_n189_));
  NA3        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n44_), .Y(new_new_n190_));
  NO2        g0168(.A(i_2_), .B(i_1_), .Y(new_new_n191_));
  NAi21      g0169(.An(i_4_), .B(i_12_), .Y(new_new_n192_));
  NO4        g0170(.A(new_new_n192_), .B(i_1_), .C(new_new_n190_), .D(new_new_n25_), .Y(new_new_n193_));
  NO3        g0171(.A(new_new_n193_), .B(new_new_n187_), .C(new_new_n180_), .Y(new_new_n194_));
  INV        g0172(.A(i_8_), .Y(new_new_n195_));
  NO2        g0173(.A(new_new_n195_), .B(i_7_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(i_6_), .Y(new_new_n197_));
  NO3        g0175(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(new_new_n113_), .Y(new_new_n199_));
  NO3        g0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n200_));
  NA3        g0178(.A(new_new_n200_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n202_));
  OAI210     g0180(.A0(new_new_n99_), .A1(i_12_), .B0(new_new_n202_), .Y(new_new_n203_));
  AOI210     g0181(.A0(new_new_n203_), .A1(new_new_n201_), .B0(new_new_n199_), .Y(new_new_n204_));
  NO2        g0182(.A(i_3_), .B(i_8_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n206_));
  NA3        g0184(.A(new_new_n206_), .B(new_new_n205_), .C(new_new_n39_), .Y(new_new_n207_));
  NO2        g0185(.A(new_new_n106_), .B(new_new_n58_), .Y(new_new_n208_));
  INV        g0186(.A(new_new_n208_), .Y(new_new_n209_));
  NO2        g0187(.A(i_13_), .B(i_9_), .Y(new_new_n210_));
  NA3        g0188(.A(new_new_n210_), .B(i_6_), .C(new_new_n195_), .Y(new_new_n211_));
  NAi21      g0189(.An(i_12_), .B(i_3_), .Y(new_new_n212_));
  NO2        g0190(.A(new_new_n44_), .B(i_5_), .Y(new_new_n213_));
  NO3        g0191(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n214_));
  NA3        g0192(.A(new_new_n214_), .B(new_new_n213_), .C(i_10_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(new_new_n211_), .B0(new_new_n209_), .B1(new_new_n207_), .Y(new_new_n216_));
  AOI210     g0194(.A0(new_new_n216_), .A1(i_7_), .B0(new_new_n204_), .Y(new_new_n217_));
  OAI220     g0195(.A0(new_new_n217_), .A1(i_4_), .B0(new_new_n197_), .B1(new_new_n194_), .Y(new_new_n218_));
  NAi21      g0196(.An(i_12_), .B(i_7_), .Y(new_new_n219_));
  NA3        g0197(.A(i_13_), .B(new_new_n195_), .C(i_10_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  NA2        g0199(.A(i_0_), .B(i_5_), .Y(new_new_n222_));
  NA2        g0200(.A(new_new_n222_), .B(new_new_n107_), .Y(new_new_n223_));
  OAI220     g0201(.A0(new_new_n223_), .A1(i_1_), .B0(new_new_n182_), .B1(new_new_n133_), .Y(new_new_n224_));
  NAi31      g0202(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n36_), .B(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n228_));
  NA3        g0206(.A(new_new_n228_), .B(new_new_n227_), .C(new_new_n226_), .Y(new_new_n229_));
  INV        g0207(.A(i_13_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n230_), .Y(new_new_n231_));
  NA3        g0209(.A(new_new_n231_), .B(new_new_n200_), .C(new_new_n198_), .Y(new_new_n232_));
  OAI210     g0210(.A0(new_new_n229_), .A1(new_new_n225_), .B0(new_new_n232_), .Y(new_new_n233_));
  AOI220     g0211(.A0(new_new_n233_), .A1(new_new_n142_), .B0(new_new_n224_), .B1(new_new_n221_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n185_), .B(i_4_), .Y(new_new_n235_));
  INV        g0213(.A(new_new_n235_), .Y(new_new_n236_));
  OR2        g0214(.A(i_8_), .B(i_7_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n237_), .B(new_new_n86_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n53_), .B(i_1_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  INV        g0218(.A(i_12_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n44_), .B(new_new_n241_), .Y(new_new_n242_));
  NO3        g0220(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(i_2_), .B(i_1_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n240_), .B(new_new_n236_), .Y(new_new_n245_));
  NO3        g0223(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_4_), .B(i_3_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n247_), .B(new_new_n75_), .Y(new_new_n248_));
  NO2        g0226(.A(i_0_), .B(i_6_), .Y(new_new_n249_));
  NOi41      g0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n250_));
  NA2        g0228(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n244_), .B(new_new_n185_), .Y(new_new_n252_));
  NAi21      g0230(.An(new_new_n251_), .B(new_new_n252_), .Y(new_new_n253_));
  INV        g0231(.A(new_new_n253_), .Y(new_new_n254_));
  AOI220     g0232(.A0(new_new_n254_), .A1(new_new_n39_), .B0(new_new_n245_), .B1(new_new_n210_), .Y(new_new_n255_));
  NO2        g0233(.A(i_11_), .B(new_new_n230_), .Y(new_new_n256_));
  NOi21      g0234(.An(i_1_), .B(i_6_), .Y(new_new_n257_));
  NAi21      g0235(.An(i_3_), .B(i_7_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n241_), .B(i_9_), .Y(new_new_n259_));
  OR4        g0237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n257_), .D(new_new_n188_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n73_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NA3        g0244(.A(new_new_n266_), .B(new_new_n263_), .C(new_new_n64_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n267_), .B(new_new_n260_), .Y(new_new_n268_));
  NA3        g0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n269_));
  INV        g0247(.A(new_new_n143_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n241_), .B(i_13_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n75_), .Y(new_new_n272_));
  AOI220     g0250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n268_), .B1(new_new_n256_), .Y(new_new_n273_));
  NO2        g0251(.A(new_new_n237_), .B(new_new_n37_), .Y(new_new_n274_));
  NA2        g0252(.A(i_12_), .B(i_6_), .Y(new_new_n275_));
  OR2        g0253(.A(i_13_), .B(i_9_), .Y(new_new_n276_));
  NO3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n48_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n247_), .B(i_2_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n277_), .C(new_new_n44_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n256_), .B(i_9_), .Y(new_new_n280_));
  NA2        g0258(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n281_));
  OAI210     g0259(.A0(new_new_n281_), .A1(new_new_n280_), .B0(new_new_n279_), .Y(new_new_n282_));
  NO3        g0260(.A(i_11_), .B(new_new_n230_), .C(new_new_n25_), .Y(new_new_n283_));
  NO2        g0261(.A(new_new_n258_), .B(i_8_), .Y(new_new_n284_));
  NO2        g0262(.A(i_6_), .B(new_new_n48_), .Y(new_new_n285_));
  NA3        g0263(.A(new_new_n285_), .B(new_new_n284_), .C(new_new_n283_), .Y(new_new_n286_));
  NO3        g0264(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n287_));
  NA3        g0265(.A(new_new_n287_), .B(new_new_n274_), .C(new_new_n231_), .Y(new_new_n288_));
  AOI210     g0266(.A0(new_new_n288_), .A1(new_new_n286_), .B0(i_1_), .Y(new_new_n289_));
  AOI210     g0267(.A0(new_new_n282_), .A1(new_new_n274_), .B0(new_new_n289_), .Y(new_new_n290_));
  NA4        g0268(.A(new_new_n290_), .B(new_new_n273_), .C(new_new_n255_), .D(new_new_n234_), .Y(new_new_n291_));
  NO3        g0269(.A(i_12_), .B(new_new_n230_), .C(new_new_n37_), .Y(new_new_n292_));
  INV        g0270(.A(new_new_n292_), .Y(new_new_n293_));
  NOi21      g0271(.An(new_new_n164_), .B(new_new_n86_), .Y(new_new_n294_));
  NO3        g0272(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n295_));
  AOI220     g0273(.A0(new_new_n295_), .A1(new_new_n198_), .B0(new_new_n294_), .B1(new_new_n239_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n296_), .B(i_7_), .Y(new_new_n297_));
  NO3        g0275(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n244_), .B(i_0_), .Y(new_new_n299_));
  AOI220     g0277(.A0(new_new_n299_), .A1(new_new_n196_), .B0(new_new_n298_), .B1(new_new_n142_), .Y(new_new_n300_));
  NA2        g0278(.A(new_new_n285_), .B(new_new_n26_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n301_), .B(new_new_n300_), .Y(new_new_n302_));
  NA2        g0280(.A(i_0_), .B(i_1_), .Y(new_new_n303_));
  NO2        g0281(.A(new_new_n303_), .B(i_2_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n59_), .B(i_6_), .Y(new_new_n305_));
  NA3        g0283(.A(new_new_n305_), .B(new_new_n304_), .C(new_new_n164_), .Y(new_new_n306_));
  OAI210     g0284(.A0(new_new_n166_), .A1(new_new_n143_), .B0(new_new_n306_), .Y(new_new_n307_));
  NO3        g0285(.A(new_new_n307_), .B(new_new_n302_), .C(new_new_n297_), .Y(new_new_n308_));
  NO2        g0286(.A(i_3_), .B(i_10_), .Y(new_new_n309_));
  NA3        g0287(.A(new_new_n309_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n310_));
  NO2        g0288(.A(i_2_), .B(new_new_n104_), .Y(new_new_n311_));
  NA2        g0289(.A(i_1_), .B(new_new_n36_), .Y(new_new_n312_));
  NOi21      g0290(.An(new_new_n222_), .B(new_new_n106_), .Y(new_new_n313_));
  NA3        g0291(.A(new_new_n313_), .B(i_1_), .C(new_new_n311_), .Y(new_new_n314_));
  AN2        g0292(.A(i_3_), .B(i_10_), .Y(new_new_n315_));
  NA4        g0293(.A(new_new_n315_), .B(new_new_n200_), .C(new_new_n178_), .D(new_new_n176_), .Y(new_new_n316_));
  NO2        g0294(.A(i_5_), .B(new_new_n37_), .Y(new_new_n317_));
  NO2        g0295(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n318_));
  OR2        g0296(.A(new_new_n314_), .B(new_new_n310_), .Y(new_new_n319_));
  OAI220     g0297(.A0(new_new_n319_), .A1(i_6_), .B0(new_new_n308_), .B1(new_new_n293_), .Y(new_new_n320_));
  NO4        g0298(.A(new_new_n320_), .B(new_new_n291_), .C(new_new_n218_), .D(new_new_n169_), .Y(new_new_n321_));
  NO3        g0299(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n322_));
  NO2        g0300(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n323_));
  NA2        g0301(.A(new_new_n299_), .B(new_new_n323_), .Y(new_new_n324_));
  NO3        g0302(.A(i_6_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n325_));
  NA2        g0303(.A(new_new_n325_), .B(new_new_n200_), .Y(new_new_n326_));
  AOI210     g0304(.A0(new_new_n326_), .A1(new_new_n324_), .B0(new_new_n171_), .Y(new_new_n327_));
  NO2        g0305(.A(i_2_), .B(i_3_), .Y(new_new_n328_));
  OR2        g0306(.A(i_0_), .B(i_5_), .Y(new_new_n329_));
  NA2        g0307(.A(new_new_n222_), .B(new_new_n329_), .Y(new_new_n330_));
  NA4        g0308(.A(new_new_n330_), .B(new_new_n238_), .C(new_new_n328_), .D(i_1_), .Y(new_new_n331_));
  NA3        g0309(.A(new_new_n299_), .B(new_new_n294_), .C(new_new_n113_), .Y(new_new_n332_));
  NAi21      g0310(.An(i_8_), .B(i_7_), .Y(new_new_n333_));
  NO2        g0311(.A(new_new_n333_), .B(i_6_), .Y(new_new_n334_));
  NO2        g0312(.A(new_new_n158_), .B(new_new_n46_), .Y(new_new_n335_));
  NA3        g0313(.A(new_new_n335_), .B(new_new_n334_), .C(new_new_n164_), .Y(new_new_n336_));
  NA3        g0314(.A(new_new_n336_), .B(new_new_n332_), .C(new_new_n331_), .Y(new_new_n337_));
  OAI210     g0315(.A0(new_new_n337_), .A1(new_new_n327_), .B0(i_4_), .Y(new_new_n338_));
  NO2        g0316(.A(i_12_), .B(i_10_), .Y(new_new_n339_));
  NOi21      g0317(.An(i_5_), .B(i_0_), .Y(new_new_n340_));
  AOI210     g0318(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n104_), .Y(new_new_n341_));
  NO4        g0319(.A(new_new_n341_), .B(new_new_n312_), .C(new_new_n340_), .D(new_new_n128_), .Y(new_new_n342_));
  NA4        g0320(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n343_));
  NA2        g0321(.A(new_new_n342_), .B(new_new_n339_), .Y(new_new_n344_));
  NO2        g0322(.A(i_6_), .B(i_8_), .Y(new_new_n345_));
  NOi21      g0323(.An(i_0_), .B(i_2_), .Y(new_new_n346_));
  AN2        g0324(.A(new_new_n346_), .B(new_new_n345_), .Y(new_new_n347_));
  NO2        g0325(.A(i_1_), .B(i_7_), .Y(new_new_n348_));
  AO220      g0326(.A0(new_new_n348_), .A1(new_new_n347_), .B0(new_new_n334_), .B1(new_new_n239_), .Y(new_new_n349_));
  NA3        g0327(.A(new_new_n349_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n350_), .B(new_new_n344_), .C(new_new_n338_), .Y(new_new_n351_));
  NO3        g0329(.A(new_new_n237_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n352_));
  NO3        g0330(.A(new_new_n333_), .B(i_2_), .C(i_1_), .Y(new_new_n353_));
  OAI210     g0331(.A0(new_new_n353_), .A1(new_new_n352_), .B0(i_6_), .Y(new_new_n354_));
  NA3        g0332(.A(new_new_n257_), .B(new_new_n311_), .C(new_new_n195_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n355_), .A1(new_new_n354_), .B0(new_new_n330_), .Y(new_new_n356_));
  NOi21      g0334(.An(new_new_n154_), .B(new_new_n107_), .Y(new_new_n357_));
  NO2        g0335(.A(new_new_n357_), .B(new_new_n124_), .Y(new_new_n358_));
  OAI210     g0336(.A0(new_new_n358_), .A1(new_new_n356_), .B0(i_3_), .Y(new_new_n359_));
  INV        g0337(.A(new_new_n84_), .Y(new_new_n360_));
  NO2        g0338(.A(new_new_n303_), .B(new_new_n81_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n132_), .Y(new_new_n362_));
  NO2        g0340(.A(new_new_n95_), .B(new_new_n195_), .Y(new_new_n363_));
  NA3        g0341(.A(new_new_n313_), .B(new_new_n363_), .C(new_new_n63_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n364_), .A1(new_new_n362_), .B0(new_new_n360_), .Y(new_new_n365_));
  NO2        g0343(.A(new_new_n195_), .B(i_9_), .Y(new_new_n366_));
  NA2        g0344(.A(new_new_n366_), .B(new_new_n208_), .Y(new_new_n367_));
  NO2        g0345(.A(new_new_n367_), .B(new_new_n46_), .Y(new_new_n368_));
  NO3        g0346(.A(new_new_n368_), .B(new_new_n365_), .C(new_new_n302_), .Y(new_new_n369_));
  AOI210     g0347(.A0(new_new_n369_), .A1(new_new_n359_), .B0(new_new_n163_), .Y(new_new_n370_));
  AOI210     g0348(.A0(new_new_n351_), .A1(new_new_n322_), .B0(new_new_n370_), .Y(new_new_n371_));
  NOi32      g0349(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n372_));
  INV        g0350(.A(new_new_n372_), .Y(new_new_n373_));
  NAi21      g0351(.An(i_0_), .B(i_6_), .Y(new_new_n374_));
  NAi21      g0352(.An(i_1_), .B(i_5_), .Y(new_new_n375_));
  NA2        g0353(.A(new_new_n375_), .B(new_new_n374_), .Y(new_new_n376_));
  NA2        g0354(.A(new_new_n376_), .B(new_new_n25_), .Y(new_new_n377_));
  OAI210     g0355(.A0(new_new_n377_), .A1(new_new_n160_), .B0(new_new_n251_), .Y(new_new_n378_));
  NAi41      g0356(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n379_));
  OAI220     g0357(.A0(new_new_n379_), .A1(new_new_n375_), .B0(new_new_n225_), .B1(new_new_n160_), .Y(new_new_n380_));
  AOI210     g0358(.A0(new_new_n379_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n381_));
  NOi32      g0359(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n382_));
  NAi21      g0360(.An(i_6_), .B(i_1_), .Y(new_new_n383_));
  NA3        g0361(.A(new_new_n383_), .B(new_new_n382_), .C(new_new_n46_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n384_), .B(i_0_), .Y(new_new_n385_));
  OR3        g0363(.A(new_new_n385_), .B(new_new_n381_), .C(new_new_n380_), .Y(new_new_n386_));
  NO2        g0364(.A(i_1_), .B(new_new_n104_), .Y(new_new_n387_));
  NAi21      g0365(.An(i_3_), .B(i_4_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n388_), .B(i_9_), .Y(new_new_n389_));
  AN2        g0367(.A(i_6_), .B(i_7_), .Y(new_new_n390_));
  OAI210     g0368(.A0(new_new_n390_), .A1(new_new_n387_), .B0(new_new_n389_), .Y(new_new_n391_));
  NA2        g0369(.A(i_2_), .B(i_7_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n388_), .B(i_10_), .Y(new_new_n393_));
  NA3        g0371(.A(new_new_n393_), .B(new_new_n392_), .C(new_new_n249_), .Y(new_new_n394_));
  AOI210     g0372(.A0(new_new_n394_), .A1(new_new_n391_), .B0(new_new_n188_), .Y(new_new_n395_));
  AOI210     g0373(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n396_));
  OAI210     g0374(.A0(new_new_n396_), .A1(new_new_n191_), .B0(new_new_n393_), .Y(new_new_n397_));
  AOI220     g0375(.A0(new_new_n393_), .A1(new_new_n348_), .B0(new_new_n243_), .B1(new_new_n191_), .Y(new_new_n398_));
  AOI210     g0376(.A0(new_new_n398_), .A1(new_new_n397_), .B0(i_5_), .Y(new_new_n399_));
  NO4        g0377(.A(new_new_n399_), .B(new_new_n395_), .C(new_new_n386_), .D(new_new_n378_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n400_), .B(new_new_n373_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n402_));
  AN2        g0380(.A(i_12_), .B(i_5_), .Y(new_new_n403_));
  NO2        g0381(.A(i_4_), .B(new_new_n26_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n404_), .B(new_new_n403_), .Y(new_new_n405_));
  NO2        g0383(.A(i_11_), .B(i_6_), .Y(new_new_n406_));
  NA3        g0384(.A(new_new_n406_), .B(new_new_n335_), .C(new_new_n230_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n405_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n247_), .B(i_5_), .Y(new_new_n409_));
  NO2        g0387(.A(i_5_), .B(i_10_), .Y(new_new_n410_));
  AOI220     g0388(.A0(new_new_n410_), .A1(new_new_n278_), .B0(new_new_n409_), .B1(new_new_n200_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n144_), .B(new_new_n45_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n412_), .B(new_new_n411_), .Y(new_new_n413_));
  OAI210     g0391(.A0(new_new_n413_), .A1(new_new_n408_), .B0(new_new_n402_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n150_), .B(new_new_n86_), .Y(new_new_n416_));
  OAI210     g0394(.A0(new_new_n416_), .A1(new_new_n408_), .B0(new_new_n415_), .Y(new_new_n417_));
  NO3        g0395(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n418_));
  NO2        g0396(.A(i_3_), .B(new_new_n104_), .Y(new_new_n419_));
  NA2        g0397(.A(new_new_n309_), .B(new_new_n75_), .Y(new_new_n420_));
  NO2        g0398(.A(i_11_), .B(i_12_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n421_), .B(new_new_n36_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n420_), .B(new_new_n422_), .Y(new_new_n423_));
  NA2        g0401(.A(new_new_n410_), .B(new_new_n241_), .Y(new_new_n424_));
  NA3        g0402(.A(new_new_n113_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(new_new_n225_), .Y(new_new_n426_));
  NAi21      g0404(.An(i_13_), .B(i_0_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(new_new_n244_), .Y(new_new_n428_));
  OAI210     g0406(.A0(new_new_n426_), .A1(new_new_n423_), .B0(new_new_n428_), .Y(new_new_n429_));
  NA3        g0407(.A(new_new_n429_), .B(new_new_n417_), .C(new_new_n414_), .Y(new_new_n430_));
  NA2        g0408(.A(new_new_n44_), .B(new_new_n230_), .Y(new_new_n431_));
  NO3        g0409(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n432_));
  NO2        g0410(.A(i_0_), .B(i_11_), .Y(new_new_n433_));
  AN2        g0411(.A(i_1_), .B(i_6_), .Y(new_new_n434_));
  NOi21      g0412(.An(i_2_), .B(i_12_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n435_), .B(new_new_n434_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(new_new_n1109_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n1113_), .B(i_4_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n437_), .B(new_new_n438_), .Y(new_new_n439_));
  NAi21      g0417(.An(i_9_), .B(i_4_), .Y(new_new_n440_));
  OR2        g0418(.A(i_13_), .B(i_10_), .Y(new_new_n441_));
  NO3        g0419(.A(new_new_n441_), .B(new_new_n117_), .C(new_new_n440_), .Y(new_new_n442_));
  NO2        g0420(.A(new_new_n174_), .B(new_new_n123_), .Y(new_new_n443_));
  OR2        g0421(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n292_), .B(new_new_n445_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n285_), .B(new_new_n214_), .Y(new_new_n447_));
  OAI220     g0425(.A0(new_new_n447_), .A1(new_new_n444_), .B0(new_new_n446_), .B1(new_new_n357_), .Y(new_new_n448_));
  INV        g0426(.A(new_new_n448_), .Y(new_new_n449_));
  AOI210     g0427(.A0(new_new_n449_), .A1(new_new_n439_), .B0(new_new_n26_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n332_), .B(new_new_n331_), .Y(new_new_n451_));
  AOI220     g0429(.A0(new_new_n305_), .A1(new_new_n295_), .B0(new_new_n299_), .B1(new_new_n323_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n452_), .B(new_new_n171_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n185_), .B(new_new_n86_), .Y(new_new_n454_));
  AOI220     g0432(.A0(new_new_n454_), .A1(new_new_n304_), .B0(new_new_n287_), .B1(new_new_n214_), .Y(new_new_n455_));
  NO2        g0433(.A(new_new_n455_), .B(i_7_), .Y(new_new_n456_));
  NO3        g0434(.A(new_new_n456_), .B(new_new_n453_), .C(new_new_n451_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n198_), .B(new_new_n99_), .Y(new_new_n458_));
  NA3        g0436(.A(new_new_n335_), .B(new_new_n164_), .C(new_new_n86_), .Y(new_new_n459_));
  AOI210     g0437(.A0(new_new_n459_), .A1(new_new_n458_), .B0(new_new_n333_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n195_), .B(i_10_), .Y(new_new_n461_));
  NA3        g0439(.A(new_new_n263_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n462_));
  NA2        g0440(.A(new_new_n305_), .B(new_new_n239_), .Y(new_new_n463_));
  OAI220     g0441(.A0(new_new_n463_), .A1(new_new_n185_), .B0(new_new_n462_), .B1(new_new_n461_), .Y(new_new_n464_));
  NO2        g0442(.A(i_3_), .B(new_new_n48_), .Y(new_new_n465_));
  NA3        g0443(.A(new_new_n348_), .B(new_new_n347_), .C(new_new_n465_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n325_), .B(new_new_n330_), .Y(new_new_n467_));
  OAI210     g0445(.A0(new_new_n467_), .A1(i_1_), .B0(new_new_n466_), .Y(new_new_n468_));
  NO3        g0446(.A(new_new_n468_), .B(new_new_n464_), .C(new_new_n460_), .Y(new_new_n469_));
  AOI210     g0447(.A0(new_new_n469_), .A1(new_new_n457_), .B0(new_new_n280_), .Y(new_new_n470_));
  NO4        g0448(.A(new_new_n470_), .B(new_new_n450_), .C(new_new_n430_), .D(new_new_n401_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n63_), .B(i_4_), .Y(new_new_n472_));
  NO2        g0450(.A(new_new_n73_), .B(i_13_), .Y(new_new_n473_));
  NO2        g0451(.A(i_10_), .B(i_9_), .Y(new_new_n474_));
  NAi21      g0452(.An(i_12_), .B(i_8_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n475_), .B(i_3_), .Y(new_new_n476_));
  NO2        g0454(.A(new_new_n46_), .B(i_4_), .Y(new_new_n477_));
  NA2        g0455(.A(new_new_n477_), .B(new_new_n107_), .Y(new_new_n478_));
  NO2        g0456(.A(new_new_n478_), .B(new_new_n207_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n318_), .B(i_0_), .Y(new_new_n480_));
  NO3        g0458(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n481_));
  NA2        g0459(.A(new_new_n275_), .B(new_new_n100_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n482_), .B(new_new_n481_), .Y(new_new_n483_));
  NA2        g0461(.A(i_8_), .B(i_9_), .Y(new_new_n484_));
  AOI210     g0462(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n485_));
  OR2        g0463(.A(new_new_n485_), .B(new_new_n484_), .Y(new_new_n486_));
  NA2        g0464(.A(new_new_n292_), .B(new_new_n208_), .Y(new_new_n487_));
  OAI220     g0465(.A0(new_new_n487_), .A1(new_new_n486_), .B0(new_new_n483_), .B1(new_new_n480_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n256_), .B(new_new_n317_), .Y(new_new_n489_));
  NO3        g0467(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n490_));
  INV        g0468(.A(new_new_n490_), .Y(new_new_n491_));
  NA3        g0469(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n492_));
  NA4        g0470(.A(new_new_n145_), .B(new_new_n115_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n493_));
  OAI220     g0471(.A0(new_new_n493_), .A1(new_new_n492_), .B0(new_new_n491_), .B1(new_new_n489_), .Y(new_new_n494_));
  NO3        g0472(.A(new_new_n494_), .B(new_new_n488_), .C(new_new_n479_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n304_), .B(new_new_n109_), .Y(new_new_n496_));
  OR2        g0474(.A(new_new_n496_), .B(new_new_n211_), .Y(new_new_n497_));
  OR2        g0475(.A(new_new_n367_), .B(new_new_n104_), .Y(new_new_n498_));
  OA220      g0476(.A0(new_new_n498_), .A1(new_new_n163_), .B0(new_new_n497_), .B1(new_new_n236_), .Y(new_new_n499_));
  NA2        g0477(.A(new_new_n99_), .B(i_13_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n454_), .B(new_new_n402_), .Y(new_new_n501_));
  NO2        g0479(.A(i_2_), .B(i_13_), .Y(new_new_n502_));
  NO2        g0480(.A(new_new_n501_), .B(new_new_n500_), .Y(new_new_n503_));
  NO3        g0481(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n504_));
  NO2        g0482(.A(i_6_), .B(i_7_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n505_), .B(new_new_n504_), .Y(new_new_n506_));
  NO2        g0484(.A(i_11_), .B(i_1_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n73_), .B(i_3_), .Y(new_new_n508_));
  OR2        g0486(.A(i_11_), .B(i_8_), .Y(new_new_n509_));
  NOi21      g0487(.An(i_2_), .B(i_7_), .Y(new_new_n510_));
  NAi31      g0488(.An(new_new_n509_), .B(new_new_n510_), .C(new_new_n508_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n441_), .B(i_6_), .Y(new_new_n512_));
  NA3        g0490(.A(new_new_n512_), .B(new_new_n472_), .C(new_new_n75_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n513_), .B(new_new_n511_), .Y(new_new_n514_));
  NO2        g0492(.A(i_3_), .B(new_new_n195_), .Y(new_new_n515_));
  NO2        g0493(.A(i_6_), .B(i_10_), .Y(new_new_n516_));
  NA3        g0494(.A(new_new_n516_), .B(new_new_n322_), .C(new_new_n515_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n517_), .B(new_new_n156_), .Y(new_new_n518_));
  NA3        g0496(.A(new_new_n250_), .B(new_new_n173_), .C(new_new_n132_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n520_));
  NO2        g0498(.A(new_new_n158_), .B(i_3_), .Y(new_new_n521_));
  NAi31      g0499(.An(new_new_n520_), .B(new_new_n521_), .C(new_new_n231_), .Y(new_new_n522_));
  NA3        g0500(.A(new_new_n415_), .B(new_new_n181_), .C(new_new_n149_), .Y(new_new_n523_));
  NA3        g0501(.A(new_new_n523_), .B(new_new_n522_), .C(new_new_n519_), .Y(new_new_n524_));
  NO4        g0502(.A(new_new_n524_), .B(new_new_n518_), .C(new_new_n514_), .D(new_new_n503_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n481_), .B(new_new_n403_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n490_), .B(new_new_n410_), .Y(new_new_n527_));
  NO2        g0505(.A(new_new_n527_), .B(new_new_n229_), .Y(new_new_n528_));
  NAi21      g0506(.An(new_new_n220_), .B(new_new_n421_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n26_), .B(i_5_), .Y(new_new_n530_));
  NO2        g0508(.A(i_0_), .B(new_new_n86_), .Y(new_new_n531_));
  NA3        g0509(.A(new_new_n531_), .B(new_new_n530_), .C(new_new_n142_), .Y(new_new_n532_));
  OR3        g0510(.A(new_new_n312_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n533_));
  NO2        g0511(.A(new_new_n533_), .B(new_new_n532_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n27_), .B(i_10_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n322_), .B(new_new_n243_), .Y(new_new_n536_));
  OAI220     g0514(.A0(new_new_n536_), .A1(new_new_n462_), .B0(new_new_n535_), .B1(new_new_n500_), .Y(new_new_n537_));
  NA4        g0515(.A(new_new_n315_), .B(new_new_n228_), .C(new_new_n73_), .D(new_new_n241_), .Y(new_new_n538_));
  NO2        g0516(.A(new_new_n538_), .B(new_new_n506_), .Y(new_new_n539_));
  NO4        g0517(.A(new_new_n539_), .B(new_new_n537_), .C(new_new_n534_), .D(new_new_n528_), .Y(new_new_n540_));
  NA4        g0518(.A(new_new_n540_), .B(new_new_n525_), .C(new_new_n499_), .D(new_new_n495_), .Y(new_new_n541_));
  NA3        g0519(.A(new_new_n315_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n542_));
  OAI210     g0520(.A0(new_new_n310_), .A1(new_new_n183_), .B0(new_new_n542_), .Y(new_new_n543_));
  AN2        g0521(.A(new_new_n295_), .B(new_new_n238_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n544_), .B(new_new_n543_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n122_), .B(new_new_n112_), .Y(new_new_n546_));
  AN2        g0524(.A(new_new_n546_), .B(new_new_n481_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n322_), .B(new_new_n165_), .Y(new_new_n548_));
  OAI210     g0526(.A0(new_new_n548_), .A1(new_new_n236_), .B0(new_new_n316_), .Y(new_new_n549_));
  AOI220     g0527(.A0(new_new_n549_), .A1(new_new_n334_), .B0(new_new_n547_), .B1(new_new_n318_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n403_), .B(new_new_n230_), .Y(new_new_n551_));
  NA2        g0529(.A(new_new_n372_), .B(new_new_n73_), .Y(new_new_n552_));
  NA2        g0530(.A(new_new_n390_), .B(new_new_n382_), .Y(new_new_n553_));
  AO210      g0531(.A0(new_new_n552_), .A1(new_new_n551_), .B0(new_new_n553_), .Y(new_new_n554_));
  NO2        g0532(.A(new_new_n36_), .B(i_8_), .Y(new_new_n555_));
  NAi41      g0533(.An(new_new_n552_), .B(new_new_n516_), .C(new_new_n555_), .D(new_new_n46_), .Y(new_new_n556_));
  INV        g0534(.A(new_new_n442_), .Y(new_new_n557_));
  NA3        g0535(.A(new_new_n557_), .B(new_new_n556_), .C(new_new_n554_), .Y(new_new_n558_));
  INV        g0536(.A(new_new_n558_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n560_));
  OAI210     g0538(.A0(i_8_), .A1(new_new_n560_), .B0(new_new_n134_), .Y(new_new_n561_));
  AOI210     g0539(.A0(new_new_n196_), .A1(i_9_), .B0(new_new_n274_), .Y(new_new_n562_));
  NO2        g0540(.A(new_new_n562_), .B(new_new_n201_), .Y(new_new_n563_));
  OR2        g0541(.A(new_new_n185_), .B(i_4_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n564_), .B(new_new_n86_), .Y(new_new_n565_));
  AOI220     g0543(.A0(new_new_n565_), .A1(new_new_n563_), .B0(new_new_n561_), .B1(new_new_n443_), .Y(new_new_n566_));
  NA4        g0544(.A(new_new_n566_), .B(new_new_n559_), .C(new_new_n550_), .D(new_new_n545_), .Y(new_new_n567_));
  NA2        g0545(.A(new_new_n409_), .B(new_new_n304_), .Y(new_new_n568_));
  NA2        g0546(.A(new_new_n170_), .B(new_new_n568_), .Y(new_new_n569_));
  NO2        g0547(.A(i_12_), .B(new_new_n195_), .Y(new_new_n570_));
  NA2        g0548(.A(new_new_n570_), .B(new_new_n230_), .Y(new_new_n571_));
  NA3        g0549(.A(new_new_n516_), .B(new_new_n176_), .C(new_new_n27_), .Y(new_new_n572_));
  NO3        g0550(.A(new_new_n572_), .B(new_new_n571_), .C(new_new_n496_), .Y(new_new_n573_));
  NOi31      g0551(.An(new_new_n325_), .B(new_new_n441_), .C(new_new_n38_), .Y(new_new_n574_));
  OAI210     g0552(.A0(new_new_n574_), .A1(new_new_n573_), .B0(new_new_n569_), .Y(new_new_n575_));
  NO2        g0553(.A(i_8_), .B(i_7_), .Y(new_new_n576_));
  OAI210     g0554(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n577_));
  NA2        g0555(.A(new_new_n577_), .B(new_new_n228_), .Y(new_new_n578_));
  AOI220     g0556(.A0(new_new_n335_), .A1(new_new_n39_), .B0(new_new_n239_), .B1(new_new_n210_), .Y(new_new_n579_));
  OAI220     g0557(.A0(new_new_n579_), .A1(new_new_n564_), .B0(new_new_n578_), .B1(new_new_n247_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n44_), .B(i_10_), .Y(new_new_n581_));
  NO2        g0559(.A(new_new_n581_), .B(i_6_), .Y(new_new_n582_));
  NA3        g0560(.A(new_new_n582_), .B(new_new_n580_), .C(new_new_n576_), .Y(new_new_n583_));
  AOI220     g0561(.A0(new_new_n454_), .A1(new_new_n335_), .B0(new_new_n252_), .B1(new_new_n249_), .Y(new_new_n584_));
  OAI220     g0562(.A0(new_new_n584_), .A1(new_new_n271_), .B0(new_new_n500_), .B1(new_new_n133_), .Y(new_new_n585_));
  NA2        g0563(.A(new_new_n585_), .B(new_new_n274_), .Y(new_new_n586_));
  NOi31      g0564(.An(new_new_n299_), .B(new_new_n310_), .C(new_new_n183_), .Y(new_new_n587_));
  NA3        g0565(.A(new_new_n315_), .B(new_new_n176_), .C(new_new_n99_), .Y(new_new_n588_));
  NO2        g0566(.A(new_new_n226_), .B(new_new_n44_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n158_), .B(i_5_), .Y(new_new_n590_));
  NA3        g0568(.A(new_new_n590_), .B(new_new_n431_), .C(new_new_n328_), .Y(new_new_n591_));
  OAI210     g0569(.A0(new_new_n591_), .A1(new_new_n589_), .B0(new_new_n588_), .Y(new_new_n592_));
  OAI210     g0570(.A0(new_new_n592_), .A1(new_new_n587_), .B0(new_new_n490_), .Y(new_new_n593_));
  NA4        g0571(.A(new_new_n593_), .B(new_new_n586_), .C(new_new_n583_), .D(new_new_n575_), .Y(new_new_n594_));
  NA3        g0572(.A(new_new_n222_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n595_));
  NA2        g0573(.A(new_new_n292_), .B(new_new_n84_), .Y(new_new_n596_));
  AOI210     g0574(.A0(new_new_n595_), .A1(new_new_n362_), .B0(new_new_n596_), .Y(new_new_n597_));
  NA2        g0575(.A(new_new_n305_), .B(new_new_n295_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n598_), .B(new_new_n175_), .Y(new_new_n599_));
  NA2        g0577(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n600_));
  NA2        g0578(.A(new_new_n474_), .B(new_new_n226_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n600_), .B(new_new_n601_), .Y(new_new_n602_));
  NA2        g0580(.A(i_0_), .B(new_new_n48_), .Y(new_new_n603_));
  NA3        g0581(.A(new_new_n570_), .B(new_new_n283_), .C(new_new_n603_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n1110_), .B(new_new_n604_), .Y(new_new_n605_));
  NO4        g0583(.A(new_new_n605_), .B(new_new_n602_), .C(new_new_n599_), .D(new_new_n597_), .Y(new_new_n606_));
  NO4        g0584(.A(new_new_n257_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n607_));
  NO3        g0585(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n608_));
  NO2        g0586(.A(new_new_n237_), .B(new_new_n36_), .Y(new_new_n609_));
  AN2        g0587(.A(new_new_n609_), .B(new_new_n608_), .Y(new_new_n610_));
  OA210      g0588(.A0(new_new_n610_), .A1(new_new_n607_), .B0(new_new_n372_), .Y(new_new_n611_));
  NO2        g0589(.A(new_new_n441_), .B(i_1_), .Y(new_new_n612_));
  NOi31      g0590(.An(new_new_n612_), .B(new_new_n482_), .C(new_new_n73_), .Y(new_new_n613_));
  AN4        g0591(.A(new_new_n613_), .B(new_new_n438_), .C(new_new_n530_), .D(i_2_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n452_), .B(new_new_n179_), .Y(new_new_n615_));
  NO3        g0593(.A(new_new_n615_), .B(new_new_n614_), .C(new_new_n611_), .Y(new_new_n616_));
  NOi21      g0594(.An(i_10_), .B(i_6_), .Y(new_new_n617_));
  NO2        g0595(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n618_));
  AOI220     g0596(.A0(new_new_n292_), .A1(new_new_n618_), .B0(new_new_n283_), .B1(new_new_n617_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n619_), .B(new_new_n480_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n325_), .B(new_new_n165_), .Y(new_new_n622_));
  AOI220     g0600(.A0(new_new_n622_), .A1(new_new_n463_), .B0(new_new_n186_), .B1(new_new_n184_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n200_), .B(new_new_n37_), .Y(new_new_n624_));
  NOi31      g0602(.An(new_new_n146_), .B(new_new_n624_), .C(new_new_n343_), .Y(new_new_n625_));
  NO3        g0603(.A(new_new_n625_), .B(new_new_n623_), .C(new_new_n620_), .Y(new_new_n626_));
  NO2        g0604(.A(new_new_n552_), .B(new_new_n398_), .Y(new_new_n627_));
  INV        g0605(.A(new_new_n328_), .Y(new_new_n628_));
  NO2        g0606(.A(i_12_), .B(new_new_n86_), .Y(new_new_n629_));
  NA3        g0607(.A(new_new_n629_), .B(new_new_n283_), .C(new_new_n603_), .Y(new_new_n630_));
  NA3        g0608(.A(new_new_n406_), .B(new_new_n292_), .C(new_new_n222_), .Y(new_new_n631_));
  AOI210     g0609(.A0(new_new_n631_), .A1(new_new_n630_), .B0(new_new_n628_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n176_), .B(i_0_), .Y(new_new_n633_));
  NO3        g0611(.A(new_new_n633_), .B(new_new_n354_), .C(new_new_n310_), .Y(new_new_n634_));
  OR2        g0612(.A(i_2_), .B(i_5_), .Y(new_new_n635_));
  OR2        g0613(.A(new_new_n635_), .B(new_new_n434_), .Y(new_new_n636_));
  AOI210     g0614(.A0(new_new_n392_), .A1(new_new_n249_), .B0(new_new_n200_), .Y(new_new_n637_));
  AOI210     g0615(.A0(new_new_n637_), .A1(new_new_n636_), .B0(new_new_n529_), .Y(new_new_n638_));
  NO4        g0616(.A(new_new_n638_), .B(new_new_n634_), .C(new_new_n632_), .D(new_new_n627_), .Y(new_new_n639_));
  NA4        g0617(.A(new_new_n639_), .B(new_new_n626_), .C(new_new_n616_), .D(new_new_n606_), .Y(new_new_n640_));
  NO4        g0618(.A(new_new_n640_), .B(new_new_n594_), .C(new_new_n567_), .D(new_new_n541_), .Y(new_new_n641_));
  NA4        g0619(.A(new_new_n641_), .B(new_new_n471_), .C(new_new_n371_), .D(new_new_n321_), .Y(men7));
  NO2        g0620(.A(new_new_n109_), .B(new_new_n92_), .Y(new_new_n643_));
  NA2        g0621(.A(new_new_n404_), .B(new_new_n643_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n516_), .B(new_new_n84_), .Y(new_new_n645_));
  OAI210     g0623(.A0(new_new_n1111_), .A1(new_new_n645_), .B0(new_new_n644_), .Y(new_new_n646_));
  NA3        g0624(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n241_), .B(i_4_), .Y(new_new_n648_));
  NA2        g0626(.A(new_new_n648_), .B(i_8_), .Y(new_new_n649_));
  AOI210     g0627(.A0(new_new_n649_), .A1(new_new_n108_), .B0(new_new_n647_), .Y(new_new_n650_));
  NA2        g0628(.A(i_2_), .B(new_new_n86_), .Y(new_new_n651_));
  OAI210     g0629(.A0(new_new_n89_), .A1(new_new_n205_), .B0(new_new_n206_), .Y(new_new_n652_));
  NO2        g0630(.A(i_7_), .B(new_new_n37_), .Y(new_new_n653_));
  NA2        g0631(.A(i_4_), .B(i_8_), .Y(new_new_n654_));
  AOI210     g0632(.A0(new_new_n654_), .A1(new_new_n315_), .B0(new_new_n653_), .Y(new_new_n655_));
  OAI220     g0633(.A0(new_new_n655_), .A1(new_new_n651_), .B0(new_new_n652_), .B1(i_13_), .Y(new_new_n656_));
  NO3        g0634(.A(new_new_n656_), .B(new_new_n650_), .C(new_new_n646_), .Y(new_new_n657_));
  AOI210     g0635(.A0(new_new_n128_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n658_));
  AOI210     g0636(.A0(new_new_n658_), .A1(new_new_n241_), .B0(new_new_n162_), .Y(new_new_n659_));
  OR2        g0637(.A(i_6_), .B(i_10_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n660_), .B(new_new_n23_), .Y(new_new_n661_));
  OR3        g0639(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n662_));
  NO3        g0640(.A(new_new_n662_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n663_));
  INV        g0641(.A(new_new_n202_), .Y(new_new_n664_));
  OR2        g0642(.A(new_new_n659_), .B(new_new_n276_), .Y(new_new_n665_));
  AOI210     g0643(.A0(new_new_n665_), .A1(new_new_n657_), .B0(new_new_n63_), .Y(new_new_n666_));
  NOi21      g0644(.An(i_11_), .B(i_7_), .Y(new_new_n667_));
  AO210      g0645(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n667_), .Y(new_new_n669_));
  NA2        g0647(.A(new_new_n669_), .B(new_new_n210_), .Y(new_new_n670_));
  NA3        g0648(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n671_));
  NAi31      g0649(.An(new_new_n671_), .B(new_new_n219_), .C(i_11_), .Y(new_new_n672_));
  AOI210     g0650(.A0(new_new_n672_), .A1(new_new_n670_), .B0(new_new_n63_), .Y(new_new_n673_));
  NO3        g0651(.A(new_new_n265_), .B(new_new_n212_), .C(i_8_), .Y(new_new_n674_));
  OAI210     g0652(.A0(new_new_n674_), .A1(new_new_n231_), .B0(new_new_n63_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n435_), .B(new_new_n31_), .Y(new_new_n676_));
  OR2        g0654(.A(new_new_n212_), .B(new_new_n109_), .Y(new_new_n677_));
  INV        g0655(.A(new_new_n676_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n63_), .B(i_9_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n679_), .B(i_4_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n680_), .B(new_new_n678_), .Y(new_new_n681_));
  NO2        g0659(.A(i_1_), .B(i_12_), .Y(new_new_n682_));
  NA3        g0660(.A(new_new_n682_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n683_));
  NA4        g0661(.A(new_new_n683_), .B(new_new_n681_), .C(new_new_n675_), .D(new_new_n398_), .Y(new_new_n684_));
  OAI210     g0662(.A0(new_new_n684_), .A1(new_new_n673_), .B0(i_6_), .Y(new_new_n685_));
  OAI210     g0663(.A0(new_new_n671_), .A1(new_new_n109_), .B0(new_new_n492_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n686_), .B(new_new_n629_), .Y(new_new_n687_));
  NO2        g0665(.A(new_new_n241_), .B(new_new_n86_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(i_11_), .Y(new_new_n689_));
  INV        g0667(.A(new_new_n687_), .Y(new_new_n690_));
  NO4        g0668(.A(new_new_n219_), .B(new_new_n128_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n691_));
  NA2        g0669(.A(new_new_n691_), .B(new_new_n679_), .Y(new_new_n692_));
  NA2        g0670(.A(new_new_n241_), .B(i_6_), .Y(new_new_n693_));
  NO3        g0671(.A(new_new_n660_), .B(new_new_n237_), .C(new_new_n23_), .Y(new_new_n694_));
  AOI210     g0672(.A0(i_1_), .A1(new_new_n266_), .B0(new_new_n694_), .Y(new_new_n695_));
  OAI210     g0673(.A0(new_new_n695_), .A1(new_new_n44_), .B0(new_new_n692_), .Y(new_new_n696_));
  NA3        g0674(.A(new_new_n576_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n697_));
  NA3        g0675(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n46_), .B(i_1_), .Y(new_new_n699_));
  NA3        g0677(.A(new_new_n699_), .B(new_new_n275_), .C(new_new_n44_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n700_), .B(new_new_n698_), .Y(new_new_n701_));
  NA3        g0679(.A(new_new_n679_), .B(new_new_n328_), .C(i_6_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n702_), .B(new_new_n23_), .Y(new_new_n703_));
  AOI210     g0681(.A0(new_new_n507_), .A1(new_new_n445_), .B0(new_new_n246_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n704_), .B(new_new_n651_), .Y(new_new_n705_));
  NAi21      g0683(.An(new_new_n697_), .B(new_new_n94_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n699_), .B(new_new_n275_), .Y(new_new_n707_));
  NO2        g0685(.A(i_11_), .B(new_new_n37_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n708_), .B(new_new_n24_), .Y(new_new_n709_));
  OAI210     g0687(.A0(new_new_n709_), .A1(new_new_n707_), .B0(new_new_n706_), .Y(new_new_n710_));
  OR4        g0688(.A(new_new_n710_), .B(new_new_n705_), .C(new_new_n703_), .D(new_new_n701_), .Y(new_new_n711_));
  NO3        g0689(.A(new_new_n711_), .B(new_new_n696_), .C(new_new_n690_), .Y(new_new_n712_));
  INV        g0690(.A(i_1_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n713_), .B(new_new_n662_), .Y(new_new_n714_));
  NO2        g0692(.A(new_new_n440_), .B(new_new_n86_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n714_), .B(new_new_n46_), .Y(new_new_n716_));
  NA2        g0694(.A(i_3_), .B(new_new_n195_), .Y(new_new_n717_));
  NO2        g0695(.A(new_new_n717_), .B(new_new_n114_), .Y(new_new_n718_));
  AN2        g0696(.A(new_new_n718_), .B(new_new_n582_), .Y(new_new_n719_));
  NO2        g0697(.A(new_new_n237_), .B(new_new_n44_), .Y(new_new_n720_));
  NO3        g0698(.A(new_new_n720_), .B(new_new_n318_), .C(new_new_n242_), .Y(new_new_n721_));
  NO2        g0699(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n722_));
  NO2        g0700(.A(new_new_n722_), .B(i_6_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n86_), .B(i_9_), .Y(new_new_n724_));
  NO2        g0702(.A(new_new_n724_), .B(new_new_n63_), .Y(new_new_n725_));
  NO2        g0703(.A(new_new_n725_), .B(new_new_n682_), .Y(new_new_n726_));
  NO4        g0704(.A(new_new_n726_), .B(new_new_n723_), .C(new_new_n721_), .D(i_4_), .Y(new_new_n727_));
  NA2        g0705(.A(i_1_), .B(i_3_), .Y(new_new_n728_));
  NO2        g0706(.A(new_new_n484_), .B(new_new_n95_), .Y(new_new_n729_));
  INV        g0707(.A(new_new_n729_), .Y(new_new_n730_));
  NO2        g0708(.A(new_new_n730_), .B(new_new_n728_), .Y(new_new_n731_));
  NO3        g0709(.A(new_new_n731_), .B(new_new_n727_), .C(new_new_n719_), .Y(new_new_n732_));
  NA4        g0710(.A(new_new_n732_), .B(new_new_n716_), .C(new_new_n712_), .D(new_new_n685_), .Y(new_new_n733_));
  NO3        g0711(.A(new_new_n509_), .B(i_3_), .C(i_7_), .Y(new_new_n734_));
  NOi21      g0712(.An(new_new_n734_), .B(i_10_), .Y(new_new_n735_));
  OA210      g0713(.A0(new_new_n735_), .A1(new_new_n250_), .B0(new_new_n86_), .Y(new_new_n736_));
  NA2        g0714(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n737_));
  NO3        g0715(.A(new_new_n510_), .B(new_new_n654_), .C(new_new_n86_), .Y(new_new_n738_));
  NA2        g0716(.A(new_new_n738_), .B(new_new_n25_), .Y(new_new_n739_));
  NA2        g0717(.A(new_new_n162_), .B(new_new_n86_), .Y(new_new_n740_));
  NA3        g0718(.A(new_new_n740_), .B(new_new_n739_), .C(new_new_n737_), .Y(new_new_n741_));
  OAI210     g0719(.A0(new_new_n741_), .A1(new_new_n736_), .B0(i_1_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n702_), .B(new_new_n475_), .Y(new_new_n743_));
  INV        g0721(.A(new_new_n743_), .Y(new_new_n744_));
  AOI210     g0722(.A0(new_new_n744_), .A1(new_new_n742_), .B0(i_13_), .Y(new_new_n745_));
  OR2        g0723(.A(i_11_), .B(i_7_), .Y(new_new_n746_));
  NA3        g0724(.A(new_new_n746_), .B(i_3_), .C(new_new_n138_), .Y(new_new_n747_));
  AOI220     g0725(.A0(new_new_n502_), .A1(new_new_n162_), .B0(new_new_n477_), .B1(new_new_n138_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n748_), .B(new_new_n747_), .Y(new_new_n749_));
  NO2        g0727(.A(new_new_n510_), .B(new_new_n24_), .Y(new_new_n750_));
  AOI210     g0728(.A0(new_new_n750_), .A1(new_new_n715_), .B0(new_new_n250_), .Y(new_new_n751_));
  OAI220     g0729(.A0(new_new_n751_), .A1(new_new_n40_), .B0(new_new_n54_), .B1(new_new_n95_), .Y(new_new_n752_));
  AOI210     g0730(.A0(new_new_n749_), .A1(new_new_n345_), .B0(new_new_n752_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n114_), .B(new_new_n109_), .Y(new_new_n754_));
  AOI220     g0732(.A0(new_new_n754_), .A1(new_new_n72_), .B0(new_new_n406_), .B1(new_new_n699_), .Y(new_new_n755_));
  NO2        g0733(.A(new_new_n755_), .B(new_new_n247_), .Y(new_new_n756_));
  AOI210     g0734(.A0(new_new_n475_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n757_));
  NOi21      g0735(.An(new_new_n757_), .B(new_new_n645_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n127_), .B(i_13_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n698_), .B(new_new_n114_), .Y(new_new_n760_));
  INV        g0738(.A(new_new_n760_), .Y(new_new_n761_));
  OAI220     g0739(.A0(new_new_n761_), .A1(new_new_n71_), .B0(new_new_n759_), .B1(new_new_n1112_), .Y(new_new_n762_));
  NO3        g0740(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n26_), .B(new_new_n195_), .Y(new_new_n764_));
  INV        g0742(.A(new_new_n763_), .Y(new_new_n765_));
  AOI220     g0743(.A0(new_new_n406_), .A1(new_new_n699_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n766_));
  OAI220     g0744(.A0(new_new_n766_), .A1(new_new_n649_), .B0(new_new_n765_), .B1(new_new_n664_), .Y(new_new_n767_));
  NO4        g0745(.A(new_new_n767_), .B(new_new_n762_), .C(new_new_n758_), .D(new_new_n756_), .Y(new_new_n768_));
  OR2        g0746(.A(i_11_), .B(i_6_), .Y(new_new_n769_));
  NA3        g0747(.A(new_new_n648_), .B(new_new_n764_), .C(i_7_), .Y(new_new_n770_));
  AOI210     g0748(.A0(new_new_n770_), .A1(new_new_n761_), .B0(new_new_n769_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n689_), .B(i_13_), .Y(new_new_n772_));
  NA2        g0750(.A(new_new_n105_), .B(new_new_n764_), .Y(new_new_n773_));
  NAi21      g0751(.An(i_11_), .B(i_12_), .Y(new_new_n774_));
  NO3        g0752(.A(new_new_n774_), .B(i_13_), .C(new_new_n86_), .Y(new_new_n775_));
  NO3        g0753(.A(new_new_n510_), .B(new_new_n629_), .C(new_new_n654_), .Y(new_new_n776_));
  AOI220     g0754(.A0(new_new_n776_), .A1(new_new_n322_), .B0(new_new_n775_), .B1(new_new_n773_), .Y(new_new_n777_));
  NA2        g0755(.A(new_new_n777_), .B(new_new_n772_), .Y(new_new_n778_));
  OAI210     g0756(.A0(new_new_n778_), .A1(new_new_n771_), .B0(new_new_n63_), .Y(new_new_n779_));
  NO2        g0757(.A(i_2_), .B(i_12_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n387_), .B(new_new_n780_), .Y(new_new_n781_));
  OAI210     g0759(.A0(i_8_), .A1(new_new_n389_), .B0(new_new_n387_), .Y(new_new_n782_));
  NO2        g0760(.A(new_new_n128_), .B(i_2_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(new_new_n682_), .Y(new_new_n784_));
  NA3        g0762(.A(new_new_n784_), .B(new_new_n782_), .C(new_new_n781_), .Y(new_new_n785_));
  NA3        g0763(.A(new_new_n785_), .B(new_new_n45_), .C(new_new_n230_), .Y(new_new_n786_));
  NA4        g0764(.A(new_new_n786_), .B(new_new_n779_), .C(new_new_n768_), .D(new_new_n753_), .Y(new_new_n787_));
  OR4        g0765(.A(new_new_n787_), .B(new_new_n745_), .C(new_new_n733_), .D(new_new_n666_), .Y(men5));
  NA3        g0766(.A(new_new_n24_), .B(new_new_n780_), .C(new_new_n109_), .Y(new_new_n789_));
  NO2        g0767(.A(new_new_n649_), .B(i_11_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n89_), .B(new_new_n790_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n791_), .B(new_new_n789_), .Y(new_new_n792_));
  NO3        g0770(.A(i_11_), .B(new_new_n241_), .C(i_13_), .Y(new_new_n793_));
  NO2        g0771(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n794_));
  NA2        g0772(.A(i_12_), .B(i_8_), .Y(new_new_n795_));
  INV        g0773(.A(new_new_n474_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n1116_), .B(new_new_n794_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n797_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n798_), .B(new_new_n792_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n173_), .Y(new_new_n800_));
  INV        g0778(.A(new_new_n250_), .Y(new_new_n801_));
  INV        g0779(.A(new_new_n476_), .Y(new_new_n802_));
  AOI210     g0780(.A0(new_new_n802_), .A1(new_new_n801_), .B0(new_new_n800_), .Y(new_new_n803_));
  NO2        g0781(.A(new_new_n484_), .B(new_new_n26_), .Y(new_new_n804_));
  NO2        g0782(.A(new_new_n804_), .B(new_new_n445_), .Y(new_new_n805_));
  INV        g0783(.A(new_new_n803_), .Y(new_new_n806_));
  INV        g0784(.A(new_new_n794_), .Y(new_new_n807_));
  INV        g0785(.A(new_new_n174_), .Y(new_new_n808_));
  NO3        g0786(.A(new_new_n668_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n809_));
  AOI210     g0787(.A0(new_new_n808_), .A1(new_new_n89_), .B0(new_new_n809_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n810_), .A1(new_new_n807_), .B0(new_new_n195_), .Y(new_new_n811_));
  OA210      g0789(.A0(new_new_n669_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n812_));
  NA2        g0790(.A(new_new_n202_), .B(new_new_n205_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n152_), .B(i_8_), .Y(new_new_n814_));
  AOI210     g0792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n392_), .Y(new_new_n815_));
  NA2        g0793(.A(new_new_n212_), .B(new_new_n148_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n816_), .B(new_new_n445_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n105_), .B(new_new_n44_), .Y(new_new_n818_));
  NA3        g0796(.A(new_new_n104_), .B(new_new_n315_), .C(new_new_n42_), .Y(new_new_n819_));
  OAI210     g0797(.A0(new_new_n819_), .A1(new_new_n818_), .B0(new_new_n817_), .Y(new_new_n820_));
  NO4        g0798(.A(new_new_n820_), .B(new_new_n815_), .C(new_new_n812_), .D(new_new_n811_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n621_), .B(new_new_n28_), .Y(new_new_n822_));
  NA2        g0800(.A(new_new_n793_), .B(new_new_n284_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n823_), .B(new_new_n822_), .Y(new_new_n824_));
  NO2        g0802(.A(new_new_n62_), .B(i_12_), .Y(new_new_n825_));
  INV        g0803(.A(new_new_n824_), .Y(new_new_n826_));
  NA4        g0804(.A(new_new_n826_), .B(new_new_n821_), .C(new_new_n806_), .D(new_new_n799_), .Y(men6));
  NO2        g0805(.A(new_new_n317_), .B(i_1_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n188_), .B(new_new_n139_), .Y(new_new_n829_));
  OAI210     g0807(.A0(new_new_n829_), .A1(new_new_n828_), .B0(new_new_n783_), .Y(new_new_n830_));
  NA4        g0808(.A(new_new_n410_), .B(new_new_n515_), .C(new_new_n71_), .D(new_new_n104_), .Y(new_new_n831_));
  INV        g0809(.A(new_new_n831_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n225_), .B(new_new_n520_), .Y(new_new_n833_));
  NO2        g0811(.A(new_new_n832_), .B(new_new_n340_), .Y(new_new_n834_));
  AO210      g0812(.A0(new_new_n834_), .A1(new_new_n830_), .B0(i_12_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n393_), .B(new_new_n348_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n735_), .B(new_new_n71_), .Y(new_new_n837_));
  NA2        g0815(.A(new_new_n837_), .B(new_new_n836_), .Y(new_new_n838_));
  INV        g0816(.A(new_new_n199_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n838_), .B(new_new_n839_), .Y(new_new_n840_));
  INV        g0818(.A(new_new_n339_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n75_), .B(new_new_n131_), .Y(new_new_n842_));
  NO2        g0820(.A(new_new_n842_), .B(new_new_n841_), .Y(new_new_n843_));
  NO3        g0821(.A(new_new_n257_), .B(new_new_n132_), .C(i_9_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n844_), .B(new_new_n825_), .Y(new_new_n845_));
  AOI210     g0823(.A0(new_new_n845_), .A1(new_new_n553_), .B0(new_new_n188_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n32_), .B(i_11_), .Y(new_new_n847_));
  NAi32      g0825(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n848_));
  AOI210     g0826(.A0(new_new_n769_), .A1(new_new_n87_), .B0(new_new_n848_), .Y(new_new_n849_));
  OAI210     g0827(.A0(new_new_n734_), .A1(new_new_n609_), .B0(new_new_n608_), .Y(new_new_n850_));
  NAi21      g0828(.An(new_new_n849_), .B(new_new_n850_), .Y(new_new_n851_));
  OR3        g0829(.A(new_new_n851_), .B(new_new_n846_), .C(new_new_n843_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n746_), .B(i_2_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n854_));
  OAI210     g0832(.A0(new_new_n854_), .A1(new_new_n434_), .B0(new_new_n377_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n855_), .B(new_new_n853_), .Y(new_new_n856_));
  AO220      g0834(.A0(new_new_n376_), .A1(new_new_n366_), .B0(new_new_n418_), .B1(i_8_), .Y(new_new_n857_));
  NA3        g0835(.A(new_new_n857_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n858_));
  OR2        g0836(.A(new_new_n669_), .B(new_new_n476_), .Y(new_new_n859_));
  NA3        g0837(.A(new_new_n859_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n860_));
  OR2        g0838(.A(new_new_n796_), .B(new_new_n36_), .Y(new_new_n861_));
  NA4        g0839(.A(new_new_n861_), .B(new_new_n860_), .C(new_new_n858_), .D(new_new_n856_), .Y(new_new_n862_));
  INV        g0840(.A(new_new_n87_), .Y(new_new_n863_));
  AOI220     g0841(.A0(new_new_n863_), .A1(new_new_n608_), .B0(new_new_n833_), .B1(new_new_n1115_), .Y(new_new_n864_));
  NA3        g0842(.A(new_new_n392_), .B(new_new_n243_), .C(new_new_n147_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n418_), .B(new_new_n70_), .Y(new_new_n866_));
  NA4        g0844(.A(new_new_n866_), .B(new_new_n865_), .C(new_new_n864_), .D(new_new_n652_), .Y(new_new_n867_));
  AO210      g0845(.A0(new_new_n555_), .A1(new_new_n46_), .B0(new_new_n88_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n868_), .B(new_new_n516_), .Y(new_new_n869_));
  AOI210     g0847(.A0(new_new_n476_), .A1(new_new_n474_), .B0(new_new_n607_), .Y(new_new_n870_));
  NO2        g0848(.A(new_new_n660_), .B(new_new_n105_), .Y(new_new_n871_));
  OAI210     g0849(.A0(new_new_n871_), .A1(new_new_n112_), .B0(new_new_n433_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n249_), .B(new_new_n46_), .Y(new_new_n873_));
  INV        g0851(.A(new_new_n636_), .Y(new_new_n874_));
  NA3        g0852(.A(new_new_n874_), .B(new_new_n339_), .C(i_7_), .Y(new_new_n875_));
  NA4        g0853(.A(new_new_n875_), .B(new_new_n872_), .C(new_new_n870_), .D(new_new_n869_), .Y(new_new_n876_));
  NO4        g0854(.A(new_new_n876_), .B(new_new_n867_), .C(new_new_n862_), .D(new_new_n852_), .Y(new_new_n877_));
  NA4        g0855(.A(new_new_n877_), .B(new_new_n840_), .C(new_new_n835_), .D(new_new_n400_), .Y(men3));
  NA2        g0856(.A(i_12_), .B(i_10_), .Y(new_new_n879_));
  NA2        g0857(.A(i_6_), .B(i_7_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n880_), .B(i_0_), .Y(new_new_n881_));
  NO2        g0859(.A(i_11_), .B(new_new_n241_), .Y(new_new_n882_));
  OAI210     g0860(.A0(new_new_n881_), .A1(new_new_n299_), .B0(new_new_n882_), .Y(new_new_n883_));
  NO2        g0861(.A(new_new_n883_), .B(new_new_n195_), .Y(new_new_n884_));
  NO3        g0862(.A(new_new_n480_), .B(new_new_n92_), .C(new_new_n44_), .Y(new_new_n885_));
  OA210      g0863(.A0(new_new_n885_), .A1(new_new_n884_), .B0(new_new_n176_), .Y(new_new_n886_));
  NA3        g0864(.A(new_new_n865_), .B(new_new_n652_), .C(new_new_n391_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n887_), .B(new_new_n39_), .Y(new_new_n888_));
  NOi21      g0866(.An(new_new_n99_), .B(new_new_n805_), .Y(new_new_n889_));
  NO3        g0867(.A(new_new_n677_), .B(new_new_n484_), .C(new_new_n131_), .Y(new_new_n890_));
  NA2        g0868(.A(new_new_n435_), .B(new_new_n45_), .Y(new_new_n891_));
  AN2        g0869(.A(new_new_n482_), .B(new_new_n55_), .Y(new_new_n892_));
  NO3        g0870(.A(new_new_n892_), .B(new_new_n890_), .C(new_new_n889_), .Y(new_new_n893_));
  AOI210     g0871(.A0(new_new_n893_), .A1(new_new_n888_), .B0(new_new_n48_), .Y(new_new_n894_));
  NO4        g0872(.A(new_new_n396_), .B(new_new_n403_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n188_), .B(new_new_n617_), .Y(new_new_n896_));
  NOi21      g0874(.An(new_new_n896_), .B(new_new_n895_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n757_), .B(new_new_n724_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n346_), .B(new_new_n465_), .Y(new_new_n899_));
  OAI220     g0877(.A0(new_new_n899_), .A1(new_new_n898_), .B0(new_new_n897_), .B1(new_new_n63_), .Y(new_new_n900_));
  NOi21      g0878(.An(i_5_), .B(i_9_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n901_), .B(new_new_n473_), .Y(new_new_n902_));
  INV        g0880(.A(new_new_n738_), .Y(new_new_n903_));
  NO3        g0881(.A(new_new_n1113_), .B(new_new_n275_), .C(new_new_n73_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n177_), .B(new_new_n148_), .Y(new_new_n905_));
  AOI210     g0883(.A0(new_new_n905_), .A1(new_new_n249_), .B0(new_new_n904_), .Y(new_new_n906_));
  OAI220     g0884(.A0(new_new_n906_), .A1(new_new_n183_), .B0(new_new_n903_), .B1(new_new_n902_), .Y(new_new_n907_));
  NO4        g0885(.A(new_new_n907_), .B(new_new_n900_), .C(new_new_n894_), .D(new_new_n886_), .Y(new_new_n908_));
  NA2        g0886(.A(new_new_n188_), .B(new_new_n24_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n722_), .B(new_new_n643_), .Y(new_new_n910_));
  NO2        g0888(.A(new_new_n910_), .B(new_new_n909_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n322_), .B(new_new_n129_), .Y(new_new_n912_));
  NAi21      g0890(.An(new_new_n163_), .B(new_new_n465_), .Y(new_new_n913_));
  OAI220     g0891(.A0(new_new_n913_), .A1(new_new_n873_), .B0(new_new_n912_), .B1(new_new_n424_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n914_), .B(new_new_n911_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n410_), .B(new_new_n303_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n916_), .B(new_new_n760_), .Y(new_new_n917_));
  NO4        g0895(.A(new_new_n635_), .B(new_new_n219_), .C(new_new_n441_), .D(new_new_n434_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n918_), .B(i_11_), .Y(new_new_n919_));
  AN2        g0897(.A(new_new_n99_), .B(new_new_n248_), .Y(new_new_n920_));
  NA2        g0898(.A(new_new_n793_), .B(new_new_n340_), .Y(new_new_n921_));
  AOI210     g0899(.A0(new_new_n516_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n922_));
  OAI220     g0900(.A0(new_new_n922_), .A1(new_new_n921_), .B0(new_new_n709_), .B1(new_new_n578_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n259_), .B(new_new_n154_), .Y(new_new_n924_));
  NA2        g0902(.A(i_0_), .B(i_10_), .Y(new_new_n925_));
  OAI210     g0903(.A0(new_new_n925_), .A1(new_new_n86_), .B0(new_new_n581_), .Y(new_new_n926_));
  NO4        g0904(.A(new_new_n114_), .B(new_new_n58_), .C(new_new_n717_), .D(i_5_), .Y(new_new_n927_));
  AO220      g0905(.A0(new_new_n927_), .A1(new_new_n926_), .B0(new_new_n924_), .B1(i_6_), .Y(new_new_n928_));
  AOI220     g0906(.A0(new_new_n346_), .A1(new_new_n101_), .B0(new_new_n188_), .B1(new_new_n84_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n612_), .B(i_4_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n191_), .B(new_new_n205_), .Y(new_new_n931_));
  OAI220     g0909(.A0(new_new_n931_), .A1(new_new_n921_), .B0(new_new_n930_), .B1(new_new_n929_), .Y(new_new_n932_));
  NO4        g0910(.A(new_new_n932_), .B(new_new_n928_), .C(new_new_n923_), .D(new_new_n920_), .Y(new_new_n933_));
  NA4        g0911(.A(new_new_n933_), .B(new_new_n919_), .C(new_new_n917_), .D(new_new_n915_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n935_));
  NA2        g0913(.A(i_11_), .B(i_9_), .Y(new_new_n936_));
  NO3        g0914(.A(i_12_), .B(new_new_n936_), .C(new_new_n651_), .Y(new_new_n937_));
  AO220      g0915(.A0(new_new_n937_), .A1(new_new_n935_), .B0(new_new_n277_), .B1(new_new_n88_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n48_), .B(i_7_), .Y(new_new_n939_));
  NAi31      g0917(.An(new_new_n272_), .B(new_new_n489_), .C(new_new_n161_), .Y(new_new_n940_));
  NO2        g0918(.A(new_new_n936_), .B(new_new_n73_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n177_), .B(i_0_), .Y(new_new_n942_));
  INV        g0920(.A(new_new_n942_), .Y(new_new_n943_));
  NA2        g0921(.A(new_new_n505_), .B(new_new_n235_), .Y(new_new_n944_));
  AOI210     g0922(.A0(new_new_n390_), .A1(new_new_n41_), .B0(new_new_n432_), .Y(new_new_n945_));
  OAI220     g0923(.A0(new_new_n945_), .A1(new_new_n902_), .B0(new_new_n944_), .B1(new_new_n943_), .Y(new_new_n946_));
  NO3        g0924(.A(new_new_n946_), .B(new_new_n940_), .C(new_new_n938_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n475_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n173_), .B(new_new_n106_), .Y(new_new_n949_));
  NOi32      g0927(.An(new_new_n948_), .Bn(new_new_n191_), .C(new_new_n949_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n653_), .A1(new_new_n340_), .B0(new_new_n248_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n951_), .B(new_new_n891_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n952_), .B(new_new_n950_), .Y(new_new_n953_));
  NOi21      g0931(.An(i_7_), .B(i_5_), .Y(new_new_n954_));
  NOi31      g0932(.An(new_new_n954_), .B(i_0_), .C(new_new_n774_), .Y(new_new_n955_));
  NA3        g0933(.A(new_new_n955_), .B(new_new_n404_), .C(i_6_), .Y(new_new_n956_));
  OA210      g0934(.A0(new_new_n949_), .A1(new_new_n553_), .B0(new_new_n956_), .Y(new_new_n957_));
  NO3        g0935(.A(new_new_n427_), .B(new_new_n379_), .C(new_new_n375_), .Y(new_new_n958_));
  NO2        g0936(.A(new_new_n269_), .B(new_new_n329_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n774_), .B(new_new_n264_), .Y(new_new_n960_));
  AOI210     g0938(.A0(new_new_n960_), .A1(new_new_n959_), .B0(new_new_n958_), .Y(new_new_n961_));
  NA4        g0939(.A(new_new_n961_), .B(new_new_n957_), .C(new_new_n953_), .D(new_new_n947_), .Y(new_new_n962_));
  NO2        g0940(.A(new_new_n909_), .B(new_new_n244_), .Y(new_new_n963_));
  AN2        g0941(.A(new_new_n345_), .B(new_new_n340_), .Y(new_new_n964_));
  AO220      g0942(.A0(new_new_n964_), .A1(new_new_n905_), .B0(new_new_n361_), .B1(new_new_n27_), .Y(new_new_n965_));
  OAI210     g0943(.A0(new_new_n965_), .A1(new_new_n963_), .B0(i_10_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n879_), .B(new_new_n328_), .Y(new_new_n967_));
  OA210      g0945(.A0(new_new_n505_), .A1(new_new_n228_), .B0(new_new_n504_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n967_), .B(new_new_n941_), .Y(new_new_n969_));
  NA3        g0947(.A(new_new_n504_), .B(new_new_n435_), .C(new_new_n45_), .Y(new_new_n970_));
  OAI210     g0948(.A0(new_new_n913_), .A1(i_7_), .B0(new_new_n970_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n262_), .B(new_new_n46_), .Y(new_new_n972_));
  NA2        g0950(.A(new_new_n941_), .B(new_new_n315_), .Y(new_new_n973_));
  OAI210     g0951(.A0(new_new_n972_), .A1(new_new_n190_), .B0(new_new_n973_), .Y(new_new_n974_));
  AOI220     g0952(.A0(new_new_n974_), .A1(new_new_n505_), .B0(new_new_n971_), .B1(new_new_n73_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n854_), .B(new_new_n402_), .C(new_new_n688_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n95_), .B(new_new_n44_), .Y(new_new_n977_));
  NO2        g0955(.A(new_new_n75_), .B(new_new_n795_), .Y(new_new_n978_));
  AOI220     g0956(.A0(new_new_n978_), .A1(new_new_n977_), .B0(new_new_n176_), .B1(new_new_n643_), .Y(new_new_n979_));
  AOI210     g0957(.A0(new_new_n979_), .A1(new_new_n976_), .B0(new_new_n47_), .Y(new_new_n980_));
  NO3        g0958(.A(new_new_n635_), .B(new_new_n374_), .C(new_new_n24_), .Y(new_new_n981_));
  AOI210     g0959(.A0(new_new_n750_), .A1(new_new_n590_), .B0(new_new_n981_), .Y(new_new_n982_));
  NAi21      g0960(.An(i_9_), .B(i_5_), .Y(new_new_n983_));
  NO2        g0961(.A(new_new_n983_), .B(new_new_n427_), .Y(new_new_n984_));
  NO2        g0962(.A(new_new_n647_), .B(new_new_n108_), .Y(new_new_n985_));
  AOI220     g0963(.A0(new_new_n985_), .A1(i_0_), .B0(new_new_n984_), .B1(new_new_n669_), .Y(new_new_n986_));
  OAI220     g0964(.A0(new_new_n986_), .A1(new_new_n86_), .B0(new_new_n982_), .B1(new_new_n174_), .Y(new_new_n987_));
  NO3        g0965(.A(new_new_n987_), .B(new_new_n980_), .C(new_new_n558_), .Y(new_new_n988_));
  NA4        g0966(.A(new_new_n988_), .B(new_new_n975_), .C(new_new_n969_), .D(new_new_n966_), .Y(new_new_n989_));
  NO3        g0967(.A(new_new_n989_), .B(new_new_n962_), .C(new_new_n934_), .Y(new_new_n990_));
  NO2        g0968(.A(i_0_), .B(new_new_n774_), .Y(new_new_n991_));
  NA2        g0969(.A(new_new_n73_), .B(new_new_n44_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n108_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n993_));
  AO220      g0971(.A0(new_new_n993_), .A1(new_new_n73_), .B0(new_new_n991_), .B1(new_new_n176_), .Y(new_new_n994_));
  NO2        g0972(.A(new_new_n737_), .B(new_new_n949_), .Y(new_new_n995_));
  AOI210     g0973(.A0(new_new_n994_), .A1(new_new_n363_), .B0(new_new_n995_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n783_), .B(new_new_n146_), .Y(new_new_n997_));
  INV        g0975(.A(new_new_n997_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n998_), .B(new_new_n724_), .C(new_new_n73_), .Y(new_new_n999_));
  NO2        g0977(.A(new_new_n850_), .B(new_new_n427_), .Y(new_new_n1000_));
  NA3        g0978(.A(new_new_n881_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n882_), .B(i_9_), .Y(new_new_n1002_));
  AOI210     g0980(.A0(new_new_n1001_), .A1(new_new_n532_), .B0(new_new_n1002_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n1003_), .B(new_new_n1000_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n1004_), .B(new_new_n999_), .C(new_new_n996_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n964_), .B(new_new_n392_), .Y(new_new_n1006_));
  AOI210     g0984(.A0(new_new_n310_), .A1(new_new_n163_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  NA2        g0985(.A(new_new_n939_), .B(new_new_n521_), .Y(new_new_n1008_));
  AOI210     g0986(.A0(i_11_), .A1(new_new_n163_), .B0(new_new_n1008_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n1009_), .B(new_new_n1007_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n925_), .B(new_new_n901_), .C(new_new_n192_), .Y(new_new_n1011_));
  AOI220     g0989(.A0(new_new_n1011_), .A1(i_11_), .B0(new_new_n613_), .B1(new_new_n75_), .Y(new_new_n1012_));
  NO3        g0990(.A(new_new_n213_), .B(new_new_n403_), .C(i_0_), .Y(new_new_n1013_));
  OAI210     g0991(.A0(new_new_n1013_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n222_), .Y(new_new_n1015_));
  OAI220     g0993(.A0(new_new_n571_), .A1(new_new_n139_), .B0(new_new_n693_), .B1(new_new_n664_), .Y(new_new_n1016_));
  NA3        g0994(.A(new_new_n1016_), .B(new_new_n419_), .C(new_new_n1015_), .Y(new_new_n1017_));
  NA4        g0995(.A(new_new_n1017_), .B(new_new_n1014_), .C(new_new_n1012_), .D(new_new_n1010_), .Y(new_new_n1018_));
  NO2        g0996(.A(new_new_n247_), .B(new_new_n95_), .Y(new_new_n1019_));
  AOI210     g0997(.A0(new_new_n1019_), .A1(new_new_n991_), .B0(new_new_n110_), .Y(new_new_n1020_));
  AOI220     g0998(.A0(new_new_n954_), .A1(new_new_n521_), .B0(new_new_n881_), .B1(new_new_n164_), .Y(new_new_n1021_));
  NA2        g0999(.A(new_new_n366_), .B(new_new_n178_), .Y(new_new_n1022_));
  OA220      g1000(.A0(new_new_n1022_), .A1(new_new_n1021_), .B0(new_new_n1020_), .B1(i_5_), .Y(new_new_n1023_));
  AOI210     g1001(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n177_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n1024_), .B(new_new_n968_), .Y(new_new_n1025_));
  NA3        g1003(.A(new_new_n661_), .B(new_new_n188_), .C(new_new_n84_), .Y(new_new_n1026_));
  NA2        g1004(.A(new_new_n1026_), .B(new_new_n588_), .Y(new_new_n1027_));
  NO3        g1005(.A(new_new_n891_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n526_), .B(new_new_n519_), .Y(new_new_n1029_));
  NO3        g1007(.A(new_new_n1029_), .B(new_new_n1028_), .C(new_new_n1027_), .Y(new_new_n1030_));
  NA3        g1008(.A(new_new_n410_), .B(new_new_n173_), .C(new_new_n172_), .Y(new_new_n1031_));
  NA3        g1009(.A(new_new_n939_), .B(new_new_n299_), .C(i_10_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n1032_), .B(new_new_n1031_), .Y(new_new_n1033_));
  NA3        g1011(.A(new_new_n410_), .B(new_new_n347_), .C(new_new_n226_), .Y(new_new_n1034_));
  INV        g1012(.A(new_new_n1034_), .Y(new_new_n1035_));
  NOi31      g1013(.An(new_new_n409_), .B(new_new_n992_), .C(new_new_n244_), .Y(new_new_n1036_));
  NO3        g1014(.A(new_new_n936_), .B(new_new_n222_), .C(new_new_n192_), .Y(new_new_n1037_));
  NO4        g1015(.A(new_new_n1037_), .B(new_new_n1036_), .C(new_new_n1035_), .D(new_new_n1033_), .Y(new_new_n1038_));
  NA4        g1016(.A(new_new_n1038_), .B(new_new_n1030_), .C(new_new_n1025_), .D(new_new_n1023_), .Y(new_new_n1039_));
  AOI210     g1017(.A0(new_new_n612_), .A1(new_new_n570_), .B0(new_new_n663_), .Y(new_new_n1040_));
  NO3        g1018(.A(new_new_n1040_), .B(new_new_n603_), .C(new_new_n360_), .Y(new_new_n1041_));
  NA3        g1019(.A(new_new_n882_), .B(new_new_n111_), .C(new_new_n124_), .Y(new_new_n1042_));
  INV        g1020(.A(new_new_n1042_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n1043_), .A1(new_new_n1114_), .B0(new_new_n1041_), .Y(new_new_n1044_));
  NA3        g1022(.A(new_new_n315_), .B(i_5_), .C(new_new_n195_), .Y(new_new_n1045_));
  NAi31      g1023(.An(new_new_n246_), .B(new_new_n1045_), .C(new_new_n247_), .Y(new_new_n1046_));
  NO4        g1024(.A(new_new_n244_), .B(new_new_n213_), .C(i_0_), .D(i_12_), .Y(new_new_n1047_));
  AOI220     g1025(.A0(new_new_n1047_), .A1(new_new_n1046_), .B0(new_new_n832_), .B1(new_new_n178_), .Y(new_new_n1048_));
  AN2        g1026(.A(new_new_n925_), .B(new_new_n154_), .Y(new_new_n1049_));
  NO4        g1027(.A(new_new_n1049_), .B(i_12_), .C(new_new_n697_), .D(new_new_n131_), .Y(new_new_n1050_));
  NA2        g1028(.A(new_new_n1050_), .B(new_new_n222_), .Y(new_new_n1051_));
  NA3        g1029(.A(new_new_n101_), .B(new_new_n617_), .C(i_11_), .Y(new_new_n1052_));
  NO2        g1030(.A(new_new_n1052_), .B(new_new_n156_), .Y(new_new_n1053_));
  NA2        g1031(.A(new_new_n954_), .B(new_new_n502_), .Y(new_new_n1054_));
  OAI220     g1032(.A0(i_7_), .A1(new_new_n1045_), .B0(new_new_n1054_), .B1(new_new_n725_), .Y(new_new_n1055_));
  AOI210     g1033(.A0(new_new_n1055_), .A1(new_new_n942_), .B0(new_new_n1053_), .Y(new_new_n1056_));
  NA4        g1034(.A(new_new_n1056_), .B(new_new_n1051_), .C(new_new_n1048_), .D(new_new_n1044_), .Y(new_new_n1057_));
  NO4        g1035(.A(new_new_n1057_), .B(new_new_n1039_), .C(new_new_n1018_), .D(new_new_n1005_), .Y(new_new_n1058_));
  OAI210     g1036(.A0(new_new_n853_), .A1(new_new_n847_), .B0(new_new_n37_), .Y(new_new_n1059_));
  NA3        g1037(.A(new_new_n948_), .B(new_new_n387_), .C(i_5_), .Y(new_new_n1060_));
  NA3        g1038(.A(new_new_n1060_), .B(new_new_n1059_), .C(new_new_n659_), .Y(new_new_n1061_));
  NA2        g1039(.A(new_new_n1061_), .B(new_new_n210_), .Y(new_new_n1062_));
  AN2        g1040(.A(new_new_n746_), .B(new_new_n388_), .Y(new_new_n1063_));
  NA2        g1041(.A(new_new_n189_), .B(new_new_n191_), .Y(new_new_n1064_));
  AO210      g1042(.A0(new_new_n1063_), .A1(new_new_n33_), .B0(new_new_n1064_), .Y(new_new_n1065_));
  OAI210     g1043(.A0(new_new_n663_), .A1(new_new_n661_), .B0(new_new_n328_), .Y(new_new_n1066_));
  NAi31      g1044(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1067_));
  NO2        g1045(.A(new_new_n70_), .B(new_new_n1067_), .Y(new_new_n1068_));
  NO2        g1046(.A(new_new_n1068_), .B(new_new_n694_), .Y(new_new_n1069_));
  NA3        g1047(.A(new_new_n1069_), .B(new_new_n1066_), .C(new_new_n1065_), .Y(new_new_n1070_));
  NO2        g1048(.A(new_new_n492_), .B(new_new_n275_), .Y(new_new_n1071_));
  NO4        g1049(.A(new_new_n237_), .B(new_new_n145_), .C(new_new_n728_), .D(new_new_n37_), .Y(new_new_n1072_));
  NO3        g1050(.A(new_new_n1072_), .B(new_new_n1071_), .C(new_new_n918_), .Y(new_new_n1073_));
  OAI210     g1051(.A0(new_new_n1052_), .A1(new_new_n148_), .B0(new_new_n1073_), .Y(new_new_n1074_));
  AOI210     g1052(.A0(new_new_n1070_), .A1(new_new_n48_), .B0(new_new_n1074_), .Y(new_new_n1075_));
  AOI210     g1053(.A0(new_new_n1075_), .A1(new_new_n1062_), .B0(new_new_n73_), .Y(new_new_n1076_));
  NO2        g1054(.A(new_new_n610_), .B(new_new_n399_), .Y(new_new_n1077_));
  NO2        g1055(.A(new_new_n1077_), .B(new_new_n800_), .Y(new_new_n1078_));
  OAI210     g1056(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n109_), .Y(new_new_n1079_));
  NA2        g1057(.A(new_new_n1079_), .B(new_new_n76_), .Y(new_new_n1080_));
  AOI210     g1058(.A0(new_new_n1024_), .A1(new_new_n939_), .B0(new_new_n955_), .Y(new_new_n1081_));
  AOI210     g1059(.A0(new_new_n1081_), .A1(new_new_n1080_), .B0(new_new_n728_), .Y(new_new_n1082_));
  NA2        g1060(.A(new_new_n269_), .B(new_new_n57_), .Y(new_new_n1083_));
  AOI220     g1061(.A0(new_new_n1083_), .A1(new_new_n76_), .B0(new_new_n361_), .B1(new_new_n261_), .Y(new_new_n1084_));
  NO2        g1062(.A(new_new_n1084_), .B(new_new_n241_), .Y(new_new_n1085_));
  NA3        g1063(.A(new_new_n99_), .B(new_new_n317_), .C(new_new_n31_), .Y(new_new_n1086_));
  INV        g1064(.A(new_new_n1086_), .Y(new_new_n1087_));
  NO3        g1065(.A(new_new_n1087_), .B(new_new_n1085_), .C(new_new_n1082_), .Y(new_new_n1088_));
  OAI210     g1066(.A0(new_new_n277_), .A1(new_new_n159_), .B0(new_new_n89_), .Y(new_new_n1089_));
  NA3        g1067(.A(new_new_n804_), .B(new_new_n299_), .C(new_new_n80_), .Y(new_new_n1090_));
  AOI210     g1068(.A0(new_new_n1090_), .A1(new_new_n1089_), .B0(i_11_), .Y(new_new_n1091_));
  NA2        g1069(.A(new_new_n654_), .B(new_new_n219_), .Y(new_new_n1092_));
  OAI210     g1070(.A0(new_new_n1092_), .A1(new_new_n948_), .B0(new_new_n210_), .Y(new_new_n1093_));
  NA2        g1071(.A(new_new_n165_), .B(i_5_), .Y(new_new_n1094_));
  AOI210     g1072(.A0(new_new_n1093_), .A1(new_new_n813_), .B0(new_new_n1094_), .Y(new_new_n1095_));
  NO3        g1073(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1096_));
  OAI210     g1074(.A0(new_new_n959_), .A1(new_new_n317_), .B0(new_new_n1096_), .Y(new_new_n1097_));
  NO2        g1075(.A(new_new_n1097_), .B(new_new_n774_), .Y(new_new_n1098_));
  NO4        g1076(.A(new_new_n983_), .B(new_new_n509_), .C(new_new_n258_), .D(new_new_n257_), .Y(new_new_n1099_));
  NO2        g1077(.A(new_new_n1099_), .B(new_new_n607_), .Y(new_new_n1100_));
  NO2        g1078(.A(new_new_n849_), .B(new_new_n380_), .Y(new_new_n1101_));
  AOI210     g1079(.A0(new_new_n1101_), .A1(new_new_n1100_), .B0(new_new_n40_), .Y(new_new_n1102_));
  NO4        g1080(.A(new_new_n1102_), .B(new_new_n1098_), .C(new_new_n1095_), .D(new_new_n1091_), .Y(new_new_n1103_));
  OAI210     g1081(.A0(new_new_n1088_), .A1(i_4_), .B0(new_new_n1103_), .Y(new_new_n1104_));
  NO3        g1082(.A(new_new_n1104_), .B(new_new_n1078_), .C(new_new_n1076_), .Y(new_new_n1105_));
  NA4        g1083(.A(new_new_n1105_), .B(new_new_n1058_), .C(new_new_n990_), .D(new_new_n908_), .Y(men4));
  INV        g1084(.A(i_5_), .Y(new_new_n1109_));
  INV        g1085(.A(new_new_n383_), .Y(new_new_n1110_));
  INV        g1086(.A(new_new_n144_), .Y(new_new_n1111_));
  INV        g1087(.A(i_1_), .Y(new_new_n1112_));
  INV        g1088(.A(i_9_), .Y(new_new_n1113_));
  INV        g1089(.A(i_5_), .Y(new_new_n1114_));
  INV        g1090(.A(i_7_), .Y(new_new_n1115_));
  INV        g1091(.A(i_3_), .Y(new_new_n1116_));
endmodule


