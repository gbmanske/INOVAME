// Benchmark "top" written by ABC on Thu Jun 20 14:00:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n135_,
    new_new_n136_, new_new_n137_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1012_, new_new_n1013_, new_new_n1014_, new_new_n1015_,
    new_new_n1016_, new_new_n1017_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(men1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA3        g031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  OAI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi31      g042(.An(new_new_n64_), .B(new_new_n62_), .C(new_new_n58_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_9_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_7_), .Y(new_new_n80_));
  NO2        g058(.A(new_new_n79_), .B(new_new_n60_), .Y(new_new_n81_));
  INV        g059(.A(i_6_), .Y(new_new_n82_));
  OR4        g060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n83_));
  INV        g061(.A(new_new_n83_), .Y(new_new_n84_));
  NO2        g062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  NO2        g063(.A(new_new_n84_), .B(new_new_n85_), .Y(new_new_n86_));
  NA2        g064(.A(new_new_n81_), .B(new_new_n86_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_10_), .Y(new_new_n88_));
  NA2        g066(.A(i_6_), .B(i_9_), .Y(new_new_n89_));
  AOI210     g067(.A0(new_new_n89_), .A1(new_new_n88_), .B0(new_new_n60_), .Y(new_new_n90_));
  NA2        g068(.A(i_2_), .B(i_6_), .Y(new_new_n91_));
  INV        g069(.A(new_new_n90_), .Y(new_new_n92_));
  AOI210     g070(.A0(new_new_n92_), .A1(new_new_n87_), .B0(new_new_n77_), .Y(new_new_n93_));
  AN3        g071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NO2        g073(.A(i_5_), .B(i_8_), .Y(new_new_n96_));
  NOi21      g074(.An(new_new_n96_), .B(new_new_n95_), .Y(new_new_n97_));
  AOI220     g075(.A0(new_new_n97_), .A1(new_new_n59_), .B0(new_new_n94_), .B1(new_new_n32_), .Y(new_new_n98_));
  INV        g076(.A(i_7_), .Y(new_new_n99_));
  NA2        g077(.A(new_new_n46_), .B(new_new_n99_), .Y(new_new_n100_));
  NO2        g078(.A(i_0_), .B(i_5_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(new_new_n82_), .Y(new_new_n102_));
  NA2        g080(.A(i_12_), .B(i_3_), .Y(new_new_n103_));
  INV        g081(.A(new_new_n103_), .Y(new_new_n104_));
  NA3        g082(.A(new_new_n104_), .B(new_new_n102_), .C(new_new_n100_), .Y(new_new_n105_));
  NAi21      g083(.An(i_7_), .B(i_11_), .Y(new_new_n106_));
  AN2        g084(.A(i_2_), .B(i_10_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n107_), .B(i_7_), .Y(new_new_n108_));
  OR2        g086(.A(new_new_n77_), .B(new_new_n55_), .Y(new_new_n109_));
  NO2        g087(.A(i_8_), .B(new_new_n99_), .Y(new_new_n110_));
  NO3        g088(.A(new_new_n110_), .B(new_new_n109_), .C(new_new_n108_), .Y(new_new_n111_));
  NA2        g089(.A(i_12_), .B(i_7_), .Y(new_new_n112_));
  NO2        g090(.A(new_new_n60_), .B(new_new_n26_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n113_), .B(i_0_), .Y(new_new_n114_));
  NA2        g092(.A(i_11_), .B(i_12_), .Y(new_new_n115_));
  OAI210     g093(.A0(new_new_n114_), .A1(new_new_n112_), .B0(new_new_n115_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n116_), .B(new_new_n111_), .Y(new_new_n117_));
  NA3        g095(.A(new_new_n117_), .B(new_new_n105_), .C(new_new_n98_), .Y(new_new_n118_));
  NOi21      g096(.An(i_1_), .B(i_5_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_11_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n121_));
  NA2        g099(.A(i_7_), .B(new_new_n25_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n122_), .B(new_new_n121_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n123_), .B(new_new_n46_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n89_), .B(new_new_n88_), .Y(new_new_n125_));
  NAi21      g103(.An(i_3_), .B(i_8_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n59_), .Y(new_new_n127_));
  NOi31      g105(.An(new_new_n127_), .B(new_new_n125_), .C(new_new_n124_), .Y(new_new_n128_));
  NO2        g106(.A(i_1_), .B(new_new_n82_), .Y(new_new_n129_));
  NO2        g107(.A(i_6_), .B(i_5_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(i_3_), .Y(new_new_n131_));
  OAI220     g109(.A0(new_new_n131_), .A1(new_new_n106_), .B0(new_new_n128_), .B1(new_new_n120_), .Y(new_new_n132_));
  NO3        g110(.A(new_new_n132_), .B(new_new_n118_), .C(new_new_n93_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n76_), .Y(men2));
  NO2        g112(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n135_));
  NA2        g113(.A(i_6_), .B(new_new_n25_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(new_new_n135_), .Y(new_new_n137_));
  NA4        g115(.A(new_new_n137_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(men0));
  AN2        g116(.A(i_8_), .B(i_7_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(i_6_), .Y(new_new_n140_));
  NO2        g118(.A(i_12_), .B(i_13_), .Y(new_new_n141_));
  NAi21      g119(.An(i_5_), .B(i_11_), .Y(new_new_n142_));
  NOi21      g120(.An(new_new_n141_), .B(new_new_n142_), .Y(new_new_n143_));
  NO2        g121(.A(i_0_), .B(i_1_), .Y(new_new_n144_));
  NA2        g122(.A(i_2_), .B(i_3_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(i_4_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(new_new_n143_), .Y(new_new_n147_));
  AN2        g125(.A(new_new_n141_), .B(new_new_n79_), .Y(new_new_n148_));
  NO2        g126(.A(new_new_n148_), .B(new_new_n27_), .Y(new_new_n149_));
  NA2        g127(.A(i_1_), .B(i_5_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n70_), .B(new_new_n46_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n36_), .Y(new_new_n152_));
  NO3        g130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  OR2        g131(.A(i_0_), .B(i_1_), .Y(new_new_n154_));
  NO3        g132(.A(new_new_n154_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n155_));
  NAi32      g133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n156_));
  NAi21      g134(.An(new_new_n156_), .B(new_new_n155_), .Y(new_new_n157_));
  NOi21      g135(.An(i_4_), .B(i_10_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n40_), .Y(new_new_n159_));
  NO2        g137(.A(i_3_), .B(i_5_), .Y(new_new_n160_));
  NO3        g138(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n161_));
  NA2        g139(.A(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  OAI210     g140(.A0(new_new_n162_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n163_), .B(new_new_n153_), .Y(new_new_n164_));
  AOI210     g142(.A0(new_new_n164_), .A1(new_new_n147_), .B0(new_new_n140_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n70_), .B(i_1_), .Y(new_new_n166_));
  NA2        g144(.A(i_3_), .B(new_new_n48_), .Y(new_new_n167_));
  NOi21      g145(.An(i_4_), .B(i_9_), .Y(new_new_n168_));
  NOi21      g146(.An(i_11_), .B(i_13_), .Y(new_new_n169_));
  NA2        g147(.A(new_new_n169_), .B(new_new_n168_), .Y(new_new_n170_));
  OR2        g148(.A(new_new_n170_), .B(new_new_n167_), .Y(new_new_n171_));
  NO2        g149(.A(i_4_), .B(i_5_), .Y(new_new_n172_));
  NAi21      g150(.An(i_12_), .B(i_11_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n173_), .B(i_13_), .Y(new_new_n174_));
  NA3        g152(.A(new_new_n174_), .B(new_new_n172_), .C(new_new_n79_), .Y(new_new_n175_));
  AOI210     g153(.A0(new_new_n175_), .A1(new_new_n171_), .B0(new_new_n166_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n70_), .B(new_new_n60_), .Y(new_new_n177_));
  INV        g155(.A(new_new_n177_), .Y(new_new_n178_));
  NA2        g156(.A(new_new_n36_), .B(i_5_), .Y(new_new_n179_));
  NAi31      g157(.An(new_new_n179_), .B(new_new_n148_), .C(i_11_), .Y(new_new_n180_));
  NA2        g158(.A(i_3_), .B(i_5_), .Y(new_new_n181_));
  OR2        g159(.A(new_new_n181_), .B(new_new_n170_), .Y(new_new_n182_));
  AOI210     g160(.A0(new_new_n182_), .A1(new_new_n180_), .B0(new_new_n178_), .Y(new_new_n183_));
  NO2        g161(.A(new_new_n70_), .B(i_5_), .Y(new_new_n184_));
  NO2        g162(.A(i_13_), .B(i_10_), .Y(new_new_n185_));
  NA3        g163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n44_), .Y(new_new_n186_));
  NO2        g164(.A(i_2_), .B(i_1_), .Y(new_new_n187_));
  NA2        g165(.A(new_new_n187_), .B(i_3_), .Y(new_new_n188_));
  NAi21      g166(.An(i_4_), .B(i_12_), .Y(new_new_n189_));
  NO4        g167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n186_), .D(new_new_n25_), .Y(new_new_n190_));
  NO3        g168(.A(new_new_n190_), .B(new_new_n183_), .C(new_new_n176_), .Y(new_new_n191_));
  INV        g169(.A(i_8_), .Y(new_new_n192_));
  NA2        g170(.A(i_8_), .B(i_6_), .Y(new_new_n193_));
  NO3        g171(.A(i_3_), .B(new_new_n82_), .C(new_new_n48_), .Y(new_new_n194_));
  NA2        g172(.A(new_new_n194_), .B(new_new_n110_), .Y(new_new_n195_));
  NO3        g173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n197_));
  NO3        g175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n198_));
  OAI210     g176(.A0(new_new_n94_), .A1(i_12_), .B0(new_new_n198_), .Y(new_new_n199_));
  AOI210     g177(.A0(new_new_n199_), .A1(new_new_n197_), .B0(new_new_n195_), .Y(new_new_n200_));
  NO2        g178(.A(i_3_), .B(i_8_), .Y(new_new_n201_));
  NO3        g179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n202_));
  NA3        g180(.A(new_new_n202_), .B(new_new_n201_), .C(new_new_n40_), .Y(new_new_n203_));
  INV        g181(.A(i_1_), .Y(new_new_n204_));
  NO2        g182(.A(i_13_), .B(i_9_), .Y(new_new_n205_));
  NA3        g183(.A(new_new_n205_), .B(i_6_), .C(new_new_n192_), .Y(new_new_n206_));
  NAi21      g184(.An(i_12_), .B(i_3_), .Y(new_new_n207_));
  OR2        g185(.A(new_new_n207_), .B(new_new_n206_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n44_), .B(i_5_), .Y(new_new_n209_));
  NO3        g187(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n210_));
  INV        g188(.A(new_new_n210_), .Y(new_new_n211_));
  OAI220     g189(.A0(new_new_n211_), .A1(new_new_n208_), .B0(new_new_n204_), .B1(new_new_n203_), .Y(new_new_n212_));
  AOI210     g190(.A0(new_new_n212_), .A1(i_7_), .B0(new_new_n200_), .Y(new_new_n213_));
  OAI220     g191(.A0(new_new_n213_), .A1(i_4_), .B0(new_new_n193_), .B1(new_new_n191_), .Y(new_new_n214_));
  NA3        g192(.A(i_13_), .B(new_new_n192_), .C(i_10_), .Y(new_new_n215_));
  NA2        g193(.A(i_0_), .B(i_5_), .Y(new_new_n216_));
  NAi31      g194(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n36_), .B(i_13_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n46_), .B(new_new_n60_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n219_), .C(new_new_n218_), .Y(new_new_n221_));
  INV        g199(.A(i_13_), .Y(new_new_n222_));
  NO2        g200(.A(i_12_), .B(new_new_n222_), .Y(new_new_n223_));
  NA3        g201(.A(new_new_n223_), .B(new_new_n196_), .C(new_new_n194_), .Y(new_new_n224_));
  OAI210     g202(.A0(new_new_n221_), .A1(new_new_n217_), .B0(new_new_n224_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n225_), .B(new_new_n139_), .Y(new_new_n226_));
  NO2        g204(.A(i_12_), .B(new_new_n37_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n181_), .B(i_4_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  OR2        g207(.A(i_8_), .B(i_7_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n230_), .B(new_new_n82_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n51_), .B(i_1_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  INV        g211(.A(i_12_), .Y(new_new_n234_));
  NO3        g212(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n235_));
  NA2        g213(.A(i_2_), .B(i_1_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n233_), .B(new_new_n229_), .Y(new_new_n237_));
  NO3        g215(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n238_));
  NAi21      g216(.An(i_4_), .B(i_3_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n72_), .Y(new_new_n240_));
  NO2        g218(.A(i_0_), .B(i_6_), .Y(new_new_n241_));
  NOi41      g219(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n242_));
  NA2        g220(.A(new_new_n242_), .B(new_new_n241_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n236_), .B(new_new_n181_), .Y(new_new_n244_));
  NAi21      g222(.An(new_new_n243_), .B(new_new_n244_), .Y(new_new_n245_));
  INV        g223(.A(new_new_n245_), .Y(new_new_n246_));
  AOI210     g224(.A0(new_new_n246_), .A1(new_new_n40_), .B0(new_new_n237_), .Y(new_new_n247_));
  NO2        g225(.A(i_11_), .B(new_new_n222_), .Y(new_new_n248_));
  NOi21      g226(.An(i_1_), .B(i_6_), .Y(new_new_n249_));
  NAi21      g227(.An(i_3_), .B(i_7_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n234_), .B(i_9_), .Y(new_new_n251_));
  OR4        g229(.A(new_new_n251_), .B(new_new_n250_), .C(new_new_n249_), .D(new_new_n184_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n70_), .B(i_5_), .Y(new_new_n254_));
  NA2        g232(.A(i_3_), .B(i_9_), .Y(new_new_n255_));
  NAi21      g233(.An(i_7_), .B(i_10_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n256_), .B(new_new_n255_), .Y(new_new_n257_));
  NA3        g235(.A(new_new_n257_), .B(new_new_n254_), .C(new_new_n61_), .Y(new_new_n258_));
  NA2        g236(.A(new_new_n258_), .B(new_new_n252_), .Y(new_new_n259_));
  NA3        g237(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n260_));
  INV        g238(.A(new_new_n140_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n234_), .B(i_13_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n262_), .B(new_new_n72_), .Y(new_new_n263_));
  AOI220     g241(.A0(new_new_n263_), .A1(new_new_n261_), .B0(new_new_n259_), .B1(new_new_n248_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n230_), .B(new_new_n37_), .Y(new_new_n265_));
  NA2        g243(.A(i_12_), .B(i_6_), .Y(new_new_n266_));
  OR2        g244(.A(i_13_), .B(i_9_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n239_), .B(i_2_), .Y(new_new_n268_));
  NA2        g246(.A(new_new_n248_), .B(i_9_), .Y(new_new_n269_));
  NA2        g247(.A(new_new_n151_), .B(new_new_n60_), .Y(new_new_n270_));
  NO3        g248(.A(i_11_), .B(new_new_n222_), .C(new_new_n25_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n250_), .B(i_8_), .Y(new_new_n272_));
  NO2        g250(.A(i_6_), .B(new_new_n48_), .Y(new_new_n273_));
  NA3        g251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n271_), .Y(new_new_n274_));
  NA3        g252(.A(i_6_), .B(new_new_n265_), .C(new_new_n223_), .Y(new_new_n275_));
  AOI210     g253(.A0(new_new_n275_), .A1(new_new_n274_), .B0(new_new_n270_), .Y(new_new_n276_));
  INV        g254(.A(new_new_n276_), .Y(new_new_n277_));
  NA4        g255(.A(new_new_n277_), .B(new_new_n264_), .C(new_new_n247_), .D(new_new_n226_), .Y(new_new_n278_));
  NO3        g256(.A(i_12_), .B(new_new_n222_), .C(new_new_n37_), .Y(new_new_n279_));
  INV        g257(.A(new_new_n279_), .Y(new_new_n280_));
  NA2        g258(.A(i_8_), .B(new_new_n99_), .Y(new_new_n281_));
  NOi21      g259(.An(new_new_n160_), .B(new_new_n82_), .Y(new_new_n282_));
  NO3        g260(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n283_));
  AOI220     g261(.A0(new_new_n283_), .A1(new_new_n194_), .B0(new_new_n282_), .B1(new_new_n232_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(new_new_n281_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n236_), .B(i_0_), .Y(new_new_n286_));
  AOI220     g264(.A0(new_new_n286_), .A1(i_8_), .B0(i_1_), .B1(new_new_n139_), .Y(new_new_n287_));
  NA2        g265(.A(new_new_n273_), .B(new_new_n26_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n288_), .B(new_new_n287_), .Y(new_new_n289_));
  NA2        g267(.A(i_0_), .B(i_1_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(i_2_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n56_), .B(i_6_), .Y(new_new_n292_));
  NA3        g270(.A(new_new_n292_), .B(new_new_n291_), .C(new_new_n160_), .Y(new_new_n293_));
  OAI210     g271(.A0(new_new_n162_), .A1(new_new_n140_), .B0(new_new_n293_), .Y(new_new_n294_));
  NO3        g272(.A(new_new_n294_), .B(new_new_n289_), .C(new_new_n285_), .Y(new_new_n295_));
  NO2        g273(.A(i_3_), .B(i_10_), .Y(new_new_n296_));
  NA3        g274(.A(new_new_n296_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n297_));
  NO2        g275(.A(i_2_), .B(new_new_n99_), .Y(new_new_n298_));
  NA2        g276(.A(i_1_), .B(new_new_n36_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n299_), .B(i_8_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n300_), .B(new_new_n298_), .Y(new_new_n301_));
  AN2        g279(.A(i_3_), .B(i_10_), .Y(new_new_n302_));
  NA4        g280(.A(new_new_n302_), .B(new_new_n196_), .C(new_new_n174_), .D(new_new_n172_), .Y(new_new_n303_));
  NO2        g281(.A(i_5_), .B(new_new_n37_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n305_));
  OR2        g283(.A(new_new_n301_), .B(new_new_n297_), .Y(new_new_n306_));
  OAI220     g284(.A0(new_new_n306_), .A1(i_6_), .B0(new_new_n295_), .B1(new_new_n280_), .Y(new_new_n307_));
  NO4        g285(.A(new_new_n307_), .B(new_new_n278_), .C(new_new_n214_), .D(new_new_n165_), .Y(new_new_n308_));
  NO3        g286(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n56_), .B(new_new_n82_), .Y(new_new_n310_));
  NO3        g288(.A(i_6_), .B(new_new_n192_), .C(i_7_), .Y(new_new_n311_));
  INV        g289(.A(new_new_n311_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n312_), .B(new_new_n167_), .Y(new_new_n313_));
  NO2        g291(.A(i_2_), .B(i_3_), .Y(new_new_n314_));
  OR2        g292(.A(i_0_), .B(i_5_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n216_), .B(new_new_n315_), .Y(new_new_n316_));
  NA4        g294(.A(new_new_n316_), .B(new_new_n231_), .C(new_new_n314_), .D(i_1_), .Y(new_new_n317_));
  NA3        g295(.A(new_new_n286_), .B(new_new_n282_), .C(new_new_n110_), .Y(new_new_n318_));
  NAi21      g296(.An(i_8_), .B(i_7_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n319_), .B(i_6_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n154_), .B(new_new_n46_), .Y(new_new_n321_));
  NA3        g299(.A(new_new_n321_), .B(new_new_n320_), .C(new_new_n160_), .Y(new_new_n322_));
  NA3        g300(.A(new_new_n322_), .B(new_new_n318_), .C(new_new_n317_), .Y(new_new_n323_));
  OAI210     g301(.A0(new_new_n323_), .A1(new_new_n313_), .B0(i_4_), .Y(new_new_n324_));
  NO2        g302(.A(i_12_), .B(i_10_), .Y(new_new_n325_));
  NOi21      g303(.An(i_5_), .B(i_0_), .Y(new_new_n326_));
  NO3        g304(.A(new_new_n299_), .B(new_new_n326_), .C(new_new_n126_), .Y(new_new_n327_));
  NA4        g305(.A(new_new_n80_), .B(new_new_n36_), .C(new_new_n82_), .D(i_8_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n327_), .B(new_new_n325_), .Y(new_new_n329_));
  NO2        g307(.A(i_6_), .B(i_8_), .Y(new_new_n330_));
  NOi21      g308(.An(i_0_), .B(i_2_), .Y(new_new_n331_));
  AN2        g309(.A(new_new_n331_), .B(new_new_n330_), .Y(new_new_n332_));
  NO2        g310(.A(i_1_), .B(i_7_), .Y(new_new_n333_));
  AO220      g311(.A0(new_new_n333_), .A1(new_new_n332_), .B0(new_new_n320_), .B1(new_new_n232_), .Y(new_new_n334_));
  NA3        g312(.A(new_new_n334_), .B(i_4_), .C(i_5_), .Y(new_new_n335_));
  NA3        g313(.A(new_new_n335_), .B(new_new_n329_), .C(new_new_n324_), .Y(new_new_n336_));
  NO3        g314(.A(new_new_n230_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n337_));
  NO3        g315(.A(new_new_n319_), .B(i_2_), .C(i_1_), .Y(new_new_n338_));
  OAI210     g316(.A0(new_new_n338_), .A1(new_new_n337_), .B0(i_6_), .Y(new_new_n339_));
  NA3        g317(.A(new_new_n249_), .B(new_new_n298_), .C(new_new_n192_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n340_), .A1(new_new_n339_), .B0(new_new_n316_), .Y(new_new_n341_));
  NOi21      g319(.An(new_new_n150_), .B(new_new_n102_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n342_), .B(new_new_n122_), .Y(new_new_n343_));
  OAI210     g321(.A0(new_new_n343_), .A1(new_new_n341_), .B0(i_3_), .Y(new_new_n344_));
  INV        g322(.A(new_new_n80_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n290_), .B(new_new_n78_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n346_), .B(new_new_n130_), .Y(new_new_n347_));
  NO2        g325(.A(new_new_n91_), .B(new_new_n192_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n348_), .B(new_new_n60_), .Y(new_new_n349_));
  AOI210     g327(.A0(new_new_n349_), .A1(new_new_n347_), .B0(new_new_n345_), .Y(new_new_n350_));
  INV        g328(.A(i_9_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n350_), .B(new_new_n289_), .Y(new_new_n352_));
  AOI210     g330(.A0(new_new_n352_), .A1(new_new_n344_), .B0(new_new_n159_), .Y(new_new_n353_));
  AOI210     g331(.A0(new_new_n336_), .A1(new_new_n309_), .B0(new_new_n353_), .Y(new_new_n354_));
  NOi32      g332(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n355_));
  INV        g333(.A(new_new_n355_), .Y(new_new_n356_));
  NAi21      g334(.An(i_1_), .B(i_5_), .Y(new_new_n357_));
  INV        g335(.A(new_new_n243_), .Y(new_new_n358_));
  NAi41      g336(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n359_));
  OAI220     g337(.A0(new_new_n359_), .A1(new_new_n357_), .B0(new_new_n217_), .B1(new_new_n156_), .Y(new_new_n360_));
  AOI210     g338(.A0(new_new_n359_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n361_));
  NOi32      g339(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n362_));
  OR2        g340(.A(new_new_n361_), .B(new_new_n360_), .Y(new_new_n363_));
  NO2        g341(.A(i_1_), .B(new_new_n99_), .Y(new_new_n364_));
  NAi21      g342(.An(i_3_), .B(i_4_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n365_), .B(i_9_), .Y(new_new_n366_));
  AN2        g344(.A(i_6_), .B(i_7_), .Y(new_new_n367_));
  OAI210     g345(.A0(new_new_n367_), .A1(new_new_n364_), .B0(new_new_n366_), .Y(new_new_n368_));
  NA2        g346(.A(i_2_), .B(i_7_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n365_), .B(i_10_), .Y(new_new_n370_));
  NA3        g348(.A(new_new_n370_), .B(new_new_n369_), .C(new_new_n241_), .Y(new_new_n371_));
  AOI210     g349(.A0(new_new_n371_), .A1(new_new_n368_), .B0(new_new_n184_), .Y(new_new_n372_));
  AOI210     g350(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n373_));
  OAI210     g351(.A0(new_new_n373_), .A1(new_new_n187_), .B0(new_new_n370_), .Y(new_new_n374_));
  AOI220     g352(.A0(new_new_n370_), .A1(new_new_n333_), .B0(new_new_n235_), .B1(new_new_n187_), .Y(new_new_n375_));
  AOI210     g353(.A0(new_new_n375_), .A1(new_new_n374_), .B0(i_5_), .Y(new_new_n376_));
  NO4        g354(.A(new_new_n376_), .B(new_new_n372_), .C(new_new_n363_), .D(new_new_n358_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n377_), .B(new_new_n356_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n379_));
  AN2        g357(.A(i_12_), .B(i_5_), .Y(new_new_n380_));
  NO2        g358(.A(i_4_), .B(new_new_n26_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n381_), .B(new_new_n380_), .Y(new_new_n382_));
  NO2        g360(.A(i_11_), .B(i_6_), .Y(new_new_n383_));
  NA3        g361(.A(new_new_n383_), .B(new_new_n321_), .C(new_new_n222_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n384_), .B(new_new_n382_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n239_), .B(i_5_), .Y(new_new_n386_));
  NO2        g364(.A(i_5_), .B(i_10_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n141_), .B(new_new_n45_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n388_), .B(new_new_n239_), .Y(new_new_n389_));
  OAI210     g367(.A0(new_new_n389_), .A1(new_new_n385_), .B0(new_new_n379_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n385_), .B(new_new_n391_), .Y(new_new_n392_));
  NO3        g370(.A(new_new_n82_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n393_));
  NA3        g371(.A(new_new_n296_), .B(new_new_n89_), .C(new_new_n52_), .Y(new_new_n394_));
  NO2        g372(.A(i_11_), .B(i_12_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n395_), .B(new_new_n36_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n394_), .B(new_new_n396_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n387_), .B(new_new_n234_), .Y(new_new_n398_));
  NA3        g376(.A(new_new_n110_), .B(i_4_), .C(i_11_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n217_), .Y(new_new_n400_));
  NAi21      g378(.An(i_13_), .B(i_0_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n401_), .B(new_new_n236_), .Y(new_new_n402_));
  OAI210     g380(.A0(new_new_n400_), .A1(new_new_n397_), .B0(new_new_n402_), .Y(new_new_n403_));
  NA3        g381(.A(new_new_n403_), .B(new_new_n392_), .C(new_new_n390_), .Y(new_new_n404_));
  NO3        g382(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n405_));
  NO2        g383(.A(i_0_), .B(i_11_), .Y(new_new_n406_));
  AN2        g384(.A(i_1_), .B(i_6_), .Y(new_new_n407_));
  NOi21      g385(.An(i_2_), .B(i_12_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n408_), .B(new_new_n407_), .Y(new_new_n409_));
  INV        g387(.A(new_new_n409_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n139_), .B(i_9_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(i_4_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n410_), .B(new_new_n412_), .Y(new_new_n413_));
  NAi21      g391(.An(i_9_), .B(i_4_), .Y(new_new_n414_));
  OR2        g392(.A(i_13_), .B(i_10_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n115_), .C(new_new_n414_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n99_), .B(new_new_n25_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n279_), .B(new_new_n417_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n273_), .B(new_new_n210_), .Y(new_new_n419_));
  OAI220     g397(.A0(new_new_n419_), .A1(new_new_n215_), .B0(new_new_n418_), .B1(new_new_n342_), .Y(new_new_n420_));
  INV        g398(.A(new_new_n420_), .Y(new_new_n421_));
  AOI210     g399(.A0(new_new_n421_), .A1(new_new_n413_), .B0(new_new_n26_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n318_), .B(new_new_n317_), .Y(new_new_n423_));
  AOI220     g401(.A0(new_new_n292_), .A1(new_new_n283_), .B0(new_new_n286_), .B1(new_new_n310_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n424_), .B(new_new_n167_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n181_), .B(new_new_n82_), .Y(new_new_n426_));
  AOI220     g404(.A0(new_new_n426_), .A1(new_new_n291_), .B0(i_6_), .B1(new_new_n210_), .Y(new_new_n427_));
  NO2        g405(.A(new_new_n427_), .B(new_new_n281_), .Y(new_new_n428_));
  NO3        g406(.A(new_new_n428_), .B(new_new_n425_), .C(new_new_n423_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n194_), .B(new_new_n94_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n321_), .B(new_new_n160_), .C(new_new_n82_), .Y(new_new_n431_));
  AOI210     g409(.A0(new_new_n431_), .A1(new_new_n430_), .B0(new_new_n319_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n192_), .B(i_10_), .Y(new_new_n433_));
  NA3        g411(.A(new_new_n254_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n292_), .B(new_new_n232_), .Y(new_new_n435_));
  OAI220     g413(.A0(new_new_n435_), .A1(new_new_n181_), .B0(new_new_n434_), .B1(new_new_n433_), .Y(new_new_n436_));
  NO2        g414(.A(i_3_), .B(new_new_n48_), .Y(new_new_n437_));
  NA3        g415(.A(new_new_n333_), .B(new_new_n332_), .C(new_new_n437_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n311_), .B(new_new_n316_), .Y(new_new_n439_));
  OAI210     g417(.A0(new_new_n439_), .A1(new_new_n188_), .B0(new_new_n438_), .Y(new_new_n440_));
  NO3        g418(.A(new_new_n440_), .B(new_new_n436_), .C(new_new_n432_), .Y(new_new_n441_));
  AOI210     g419(.A0(new_new_n441_), .A1(new_new_n429_), .B0(new_new_n269_), .Y(new_new_n442_));
  NO4        g420(.A(new_new_n442_), .B(new_new_n422_), .C(new_new_n404_), .D(new_new_n378_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n60_), .B(i_4_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n70_), .B(i_13_), .Y(new_new_n445_));
  NO2        g423(.A(i_10_), .B(i_9_), .Y(new_new_n446_));
  NAi21      g424(.An(i_12_), .B(i_8_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n447_), .B(i_3_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n46_), .B(i_4_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n449_), .B(new_new_n102_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n450_), .B(new_new_n203_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n305_), .B(i_0_), .Y(new_new_n452_));
  NO3        g430(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n266_), .B(new_new_n95_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NA2        g433(.A(i_8_), .B(i_9_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n248_), .B(new_new_n304_), .Y(new_new_n457_));
  NO3        g435(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n458_));
  INV        g436(.A(new_new_n458_), .Y(new_new_n459_));
  NA3        g437(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n460_));
  NA4        g438(.A(new_new_n142_), .B(new_new_n113_), .C(new_new_n77_), .D(new_new_n23_), .Y(new_new_n461_));
  OAI220     g439(.A0(new_new_n461_), .A1(new_new_n460_), .B0(new_new_n459_), .B1(new_new_n457_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n451_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n291_), .B(new_new_n106_), .Y(new_new_n464_));
  OR2        g442(.A(new_new_n464_), .B(new_new_n206_), .Y(new_new_n465_));
  BUFFER     g443(.A(new_new_n293_), .Y(new_new_n466_));
  OA220      g444(.A0(new_new_n466_), .A1(new_new_n159_), .B0(new_new_n465_), .B1(new_new_n229_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n94_), .B(i_13_), .Y(new_new_n468_));
  NA2        g446(.A(new_new_n426_), .B(new_new_n379_), .Y(new_new_n469_));
  NO2        g447(.A(i_2_), .B(i_13_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n471_));
  NO3        g449(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n472_));
  NO2        g450(.A(i_6_), .B(i_7_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NO2        g452(.A(i_11_), .B(i_1_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n70_), .B(i_3_), .Y(new_new_n476_));
  NOi21      g454(.An(i_2_), .B(i_7_), .Y(new_new_n477_));
  NAi31      g455(.An(i_11_), .B(new_new_n477_), .C(new_new_n476_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n415_), .B(i_6_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(new_new_n444_), .Y(new_new_n480_));
  NO2        g458(.A(new_new_n480_), .B(new_new_n478_), .Y(new_new_n481_));
  NO2        g459(.A(i_3_), .B(new_new_n192_), .Y(new_new_n482_));
  NO2        g460(.A(i_6_), .B(i_10_), .Y(new_new_n483_));
  NA4        g461(.A(new_new_n483_), .B(new_new_n309_), .C(new_new_n482_), .D(new_new_n234_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(new_new_n152_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n154_), .B(i_3_), .Y(new_new_n487_));
  NAi31      g465(.An(new_new_n486_), .B(new_new_n487_), .C(new_new_n223_), .Y(new_new_n488_));
  NA3        g466(.A(new_new_n391_), .B(new_new_n177_), .C(new_new_n146_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NO4        g468(.A(new_new_n490_), .B(new_new_n485_), .C(new_new_n481_), .D(new_new_n471_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n458_), .B(new_new_n387_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n492_), .B(new_new_n221_), .Y(new_new_n493_));
  NAi21      g471(.An(new_new_n215_), .B(new_new_n395_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n26_), .B(i_5_), .Y(new_new_n495_));
  NO2        g473(.A(i_0_), .B(new_new_n82_), .Y(new_new_n496_));
  NA3        g474(.A(new_new_n496_), .B(new_new_n495_), .C(new_new_n139_), .Y(new_new_n497_));
  OR3        g475(.A(new_new_n299_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(new_new_n497_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n27_), .B(i_10_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n309_), .B(new_new_n235_), .Y(new_new_n501_));
  OAI220     g479(.A0(new_new_n501_), .A1(new_new_n434_), .B0(new_new_n500_), .B1(new_new_n468_), .Y(new_new_n502_));
  NA4        g480(.A(new_new_n302_), .B(new_new_n220_), .C(new_new_n70_), .D(new_new_n234_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(new_new_n474_), .Y(new_new_n504_));
  NO4        g482(.A(new_new_n504_), .B(new_new_n502_), .C(new_new_n499_), .D(new_new_n493_), .Y(new_new_n505_));
  NA4        g483(.A(new_new_n505_), .B(new_new_n491_), .C(new_new_n467_), .D(new_new_n463_), .Y(new_new_n506_));
  NA3        g484(.A(new_new_n302_), .B(new_new_n174_), .C(new_new_n172_), .Y(new_new_n507_));
  OAI210     g485(.A0(new_new_n297_), .A1(new_new_n179_), .B0(new_new_n507_), .Y(new_new_n508_));
  BUFFER     g486(.A(new_new_n283_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n509_), .B(new_new_n508_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n120_), .B(new_new_n109_), .Y(new_new_n511_));
  AN2        g489(.A(new_new_n511_), .B(new_new_n453_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n309_), .B(new_new_n161_), .Y(new_new_n513_));
  OAI210     g491(.A0(new_new_n513_), .A1(new_new_n229_), .B0(new_new_n303_), .Y(new_new_n514_));
  AOI220     g492(.A0(new_new_n514_), .A1(new_new_n320_), .B0(new_new_n512_), .B1(new_new_n305_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n380_), .B(new_new_n222_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n355_), .B(new_new_n70_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n367_), .B(new_new_n362_), .Y(new_new_n518_));
  AO210      g496(.A0(new_new_n517_), .A1(new_new_n516_), .B0(new_new_n518_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n36_), .B(i_8_), .Y(new_new_n520_));
  NAi41      g498(.An(new_new_n517_), .B(new_new_n483_), .C(new_new_n520_), .D(new_new_n46_), .Y(new_new_n521_));
  AOI210     g499(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n416_), .Y(new_new_n522_));
  NA3        g500(.A(new_new_n522_), .B(new_new_n521_), .C(new_new_n519_), .Y(new_new_n523_));
  INV        g501(.A(new_new_n523_), .Y(new_new_n524_));
  NO2        g502(.A(i_7_), .B(new_new_n197_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n181_), .B(new_new_n82_), .Y(new_new_n526_));
  NA2        g504(.A(new_new_n526_), .B(new_new_n525_), .Y(new_new_n527_));
  NA4        g505(.A(new_new_n527_), .B(new_new_n524_), .C(new_new_n515_), .D(new_new_n510_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n386_), .B(new_new_n291_), .Y(new_new_n529_));
  OAI210     g507(.A0(new_new_n382_), .A1(new_new_n166_), .B0(new_new_n529_), .Y(new_new_n530_));
  NA2        g508(.A(new_new_n1016_), .B(new_new_n222_), .Y(new_new_n531_));
  NO3        g509(.A(new_new_n1014_), .B(new_new_n531_), .C(new_new_n464_), .Y(new_new_n532_));
  NOi31      g510(.An(new_new_n311_), .B(new_new_n415_), .C(new_new_n38_), .Y(new_new_n533_));
  OAI210     g511(.A0(new_new_n533_), .A1(new_new_n532_), .B0(new_new_n530_), .Y(new_new_n534_));
  NO2        g512(.A(i_8_), .B(i_7_), .Y(new_new_n535_));
  INV        g513(.A(i_5_), .Y(new_new_n536_));
  NA2        g514(.A(new_new_n536_), .B(new_new_n220_), .Y(new_new_n537_));
  AOI220     g515(.A0(new_new_n321_), .A1(new_new_n40_), .B0(new_new_n232_), .B1(new_new_n205_), .Y(new_new_n538_));
  OAI220     g516(.A0(new_new_n538_), .A1(new_new_n181_), .B0(new_new_n537_), .B1(new_new_n239_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n44_), .B(i_10_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n540_), .B(i_6_), .Y(new_new_n541_));
  NA3        g519(.A(new_new_n541_), .B(new_new_n539_), .C(new_new_n535_), .Y(new_new_n542_));
  AOI220     g520(.A0(new_new_n426_), .A1(new_new_n321_), .B0(new_new_n244_), .B1(new_new_n241_), .Y(new_new_n543_));
  OAI220     g521(.A0(new_new_n543_), .A1(new_new_n262_), .B0(new_new_n468_), .B1(new_new_n131_), .Y(new_new_n544_));
  NA2        g522(.A(new_new_n544_), .B(new_new_n265_), .Y(new_new_n545_));
  NOi21      g523(.An(new_new_n286_), .B(new_new_n297_), .Y(new_new_n546_));
  NA2        g524(.A(new_new_n546_), .B(new_new_n458_), .Y(new_new_n547_));
  NA4        g525(.A(new_new_n547_), .B(new_new_n545_), .C(new_new_n542_), .D(new_new_n534_), .Y(new_new_n548_));
  NA3        g526(.A(new_new_n216_), .B(new_new_n68_), .C(new_new_n44_), .Y(new_new_n549_));
  NA2        g527(.A(new_new_n279_), .B(new_new_n80_), .Y(new_new_n550_));
  AOI210     g528(.A0(new_new_n549_), .A1(new_new_n347_), .B0(new_new_n550_), .Y(new_new_n551_));
  NA2        g529(.A(new_new_n292_), .B(new_new_n283_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n552_), .B(new_new_n171_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n554_));
  NA2        g532(.A(new_new_n446_), .B(new_new_n218_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n554_), .B(new_new_n555_), .Y(new_new_n556_));
  NO3        g534(.A(new_new_n556_), .B(new_new_n553_), .C(new_new_n551_), .Y(new_new_n557_));
  NO4        g535(.A(new_new_n249_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n558_));
  NO3        g536(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n230_), .B(new_new_n36_), .Y(new_new_n560_));
  AN2        g538(.A(new_new_n560_), .B(new_new_n559_), .Y(new_new_n561_));
  OA210      g539(.A0(new_new_n561_), .A1(new_new_n558_), .B0(new_new_n355_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n415_), .B(i_1_), .Y(new_new_n563_));
  NOi31      g541(.An(new_new_n563_), .B(new_new_n454_), .C(new_new_n70_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n424_), .B(new_new_n175_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n565_), .B(new_new_n562_), .Y(new_new_n566_));
  NOi21      g544(.An(i_10_), .B(i_6_), .Y(new_new_n567_));
  NO2        g545(.A(new_new_n82_), .B(new_new_n25_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n569_));
  NA2        g547(.A(new_new_n311_), .B(new_new_n161_), .Y(new_new_n570_));
  AOI220     g548(.A0(new_new_n570_), .A1(new_new_n435_), .B0(new_new_n182_), .B1(new_new_n180_), .Y(new_new_n571_));
  NOi21      g549(.An(new_new_n143_), .B(new_new_n328_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n572_), .B(new_new_n571_), .Y(new_new_n573_));
  NO2        g551(.A(i_12_), .B(new_new_n82_), .Y(new_new_n574_));
  NA2        g552(.A(new_new_n172_), .B(i_0_), .Y(new_new_n575_));
  NO3        g553(.A(new_new_n575_), .B(new_new_n339_), .C(new_new_n297_), .Y(new_new_n576_));
  INV        g554(.A(new_new_n196_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n577_), .B(new_new_n494_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n578_), .B(new_new_n576_), .Y(new_new_n579_));
  NA4        g557(.A(new_new_n579_), .B(new_new_n573_), .C(new_new_n566_), .D(new_new_n557_), .Y(new_new_n580_));
  NO4        g558(.A(new_new_n580_), .B(new_new_n548_), .C(new_new_n528_), .D(new_new_n506_), .Y(new_new_n581_));
  NA4        g559(.A(new_new_n581_), .B(new_new_n443_), .C(new_new_n354_), .D(new_new_n308_), .Y(men7));
  NO2        g560(.A(new_new_n91_), .B(new_new_n52_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n106_), .B(new_new_n88_), .Y(new_new_n584_));
  NA2        g562(.A(new_new_n381_), .B(new_new_n584_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n483_), .B(new_new_n80_), .Y(new_new_n586_));
  NA2        g564(.A(i_11_), .B(new_new_n192_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n141_), .B(new_new_n587_), .Y(new_new_n588_));
  OAI210     g566(.A0(new_new_n588_), .A1(new_new_n586_), .B0(new_new_n585_), .Y(new_new_n589_));
  NA3        g567(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n234_), .B(i_4_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(i_8_), .Y(new_new_n592_));
  NO2        g570(.A(new_new_n103_), .B(new_new_n590_), .Y(new_new_n593_));
  NA2        g571(.A(i_2_), .B(new_new_n82_), .Y(new_new_n594_));
  OAI210     g572(.A0(new_new_n85_), .A1(new_new_n201_), .B0(new_new_n202_), .Y(new_new_n595_));
  NO2        g573(.A(i_7_), .B(new_new_n37_), .Y(new_new_n596_));
  NA2        g574(.A(i_4_), .B(i_8_), .Y(new_new_n597_));
  AOI210     g575(.A0(new_new_n597_), .A1(new_new_n302_), .B0(new_new_n596_), .Y(new_new_n598_));
  OAI220     g576(.A0(new_new_n598_), .A1(new_new_n594_), .B0(new_new_n595_), .B1(i_13_), .Y(new_new_n599_));
  NO4        g577(.A(new_new_n599_), .B(new_new_n593_), .C(new_new_n589_), .D(new_new_n583_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n126_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n601_));
  AOI210     g579(.A0(new_new_n601_), .A1(new_new_n234_), .B0(new_new_n158_), .Y(new_new_n602_));
  OR2        g580(.A(i_6_), .B(i_10_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n603_), .B(new_new_n23_), .Y(new_new_n604_));
  OR3        g582(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n605_));
  NO3        g583(.A(new_new_n605_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n606_));
  INV        g584(.A(new_new_n198_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n606_), .B(new_new_n604_), .Y(new_new_n608_));
  OA220      g586(.A0(new_new_n608_), .A1(i_2_), .B0(new_new_n602_), .B1(new_new_n267_), .Y(new_new_n609_));
  AOI210     g587(.A0(new_new_n609_), .A1(new_new_n600_), .B0(new_new_n60_), .Y(new_new_n610_));
  NOi21      g588(.An(i_11_), .B(i_7_), .Y(new_new_n611_));
  AO210      g589(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n611_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n205_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n614_), .B(new_new_n60_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n84_), .B(new_new_n60_), .Y(new_new_n616_));
  AO210      g594(.A0(new_new_n616_), .A1(new_new_n375_), .B0(new_new_n41_), .Y(new_new_n617_));
  NA2        g595(.A(new_new_n223_), .B(new_new_n60_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n408_), .B(new_new_n31_), .Y(new_new_n619_));
  OR2        g597(.A(new_new_n207_), .B(new_new_n106_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n619_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n60_), .B(i_9_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n622_), .B(i_4_), .Y(new_new_n623_));
  NA2        g601(.A(new_new_n623_), .B(new_new_n621_), .Y(new_new_n624_));
  NO2        g602(.A(i_1_), .B(i_12_), .Y(new_new_n625_));
  NA3        g603(.A(new_new_n625_), .B(new_new_n107_), .C(new_new_n24_), .Y(new_new_n626_));
  NA4        g604(.A(new_new_n626_), .B(new_new_n624_), .C(new_new_n618_), .D(new_new_n617_), .Y(new_new_n627_));
  OAI210     g605(.A0(new_new_n627_), .A1(new_new_n615_), .B0(i_6_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n234_), .B(new_new_n82_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(i_11_), .Y(new_new_n630_));
  INV        g608(.A(new_new_n455_), .Y(new_new_n631_));
  NO4        g609(.A(i_12_), .B(new_new_n126_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n632_), .B(new_new_n622_), .Y(new_new_n633_));
  NO3        g611(.A(new_new_n603_), .B(new_new_n230_), .C(new_new_n23_), .Y(new_new_n634_));
  AOI210     g612(.A0(i_1_), .A1(new_new_n257_), .B0(new_new_n634_), .Y(new_new_n635_));
  OAI210     g613(.A0(new_new_n635_), .A1(new_new_n44_), .B0(new_new_n633_), .Y(new_new_n636_));
  NA3        g614(.A(new_new_n535_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n135_), .B(i_9_), .Y(new_new_n638_));
  NA3        g616(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n46_), .B(i_1_), .Y(new_new_n640_));
  NA3        g618(.A(new_new_n640_), .B(new_new_n266_), .C(new_new_n44_), .Y(new_new_n641_));
  OAI220     g619(.A0(new_new_n641_), .A1(new_new_n639_), .B0(new_new_n638_), .B1(new_new_n1013_), .Y(new_new_n642_));
  NA3        g620(.A(new_new_n622_), .B(new_new_n314_), .C(i_6_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(new_new_n23_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n475_), .A1(new_new_n417_), .B0(new_new_n238_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n594_), .Y(new_new_n646_));
  NAi21      g624(.An(new_new_n637_), .B(new_new_n90_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n640_), .B(new_new_n266_), .Y(new_new_n648_));
  NO2        g626(.A(i_11_), .B(new_new_n37_), .Y(new_new_n649_));
  NA2        g627(.A(new_new_n649_), .B(new_new_n24_), .Y(new_new_n650_));
  OAI210     g628(.A0(new_new_n650_), .A1(new_new_n648_), .B0(new_new_n647_), .Y(new_new_n651_));
  OR4        g629(.A(new_new_n651_), .B(new_new_n646_), .C(new_new_n644_), .D(new_new_n642_), .Y(new_new_n652_));
  NO3        g630(.A(new_new_n652_), .B(new_new_n636_), .C(new_new_n631_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n234_), .B(new_new_n99_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n654_), .B(new_new_n611_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n414_), .B(new_new_n82_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n115_), .B(new_new_n37_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n82_), .B(i_9_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n658_), .B(new_new_n60_), .Y(new_new_n659_));
  NA2        g637(.A(i_1_), .B(i_3_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n653_), .B(new_new_n628_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n367_), .B(new_new_n366_), .Y(new_new_n662_));
  NO3        g640(.A(new_new_n477_), .B(new_new_n597_), .C(new_new_n82_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n663_), .B(new_new_n25_), .Y(new_new_n664_));
  NA3        g642(.A(new_new_n158_), .B(new_new_n80_), .C(new_new_n82_), .Y(new_new_n665_));
  NA3        g643(.A(new_new_n665_), .B(new_new_n664_), .C(new_new_n662_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n666_), .B(i_1_), .Y(new_new_n667_));
  AOI210     g645(.A0(new_new_n266_), .A1(new_new_n95_), .B0(i_1_), .Y(new_new_n668_));
  NO2        g646(.A(new_new_n365_), .B(i_2_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n669_), .B(new_new_n668_), .Y(new_new_n670_));
  AOI210     g648(.A0(new_new_n670_), .A1(new_new_n667_), .B0(i_13_), .Y(new_new_n671_));
  OR2        g649(.A(i_11_), .B(i_7_), .Y(new_new_n672_));
  NA3        g650(.A(new_new_n672_), .B(new_new_n104_), .C(new_new_n135_), .Y(new_new_n673_));
  AOI220     g651(.A0(new_new_n470_), .A1(new_new_n158_), .B0(new_new_n449_), .B1(new_new_n135_), .Y(new_new_n674_));
  OAI210     g652(.A0(new_new_n674_), .A1(new_new_n44_), .B0(new_new_n673_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n52_), .B(i_12_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n477_), .B(new_new_n24_), .Y(new_new_n677_));
  AOI220     g655(.A0(new_new_n677_), .A1(new_new_n656_), .B0(new_new_n242_), .B1(new_new_n129_), .Y(new_new_n678_));
  OAI220     g656(.A0(new_new_n678_), .A1(new_new_n41_), .B0(new_new_n1012_), .B1(new_new_n91_), .Y(new_new_n679_));
  AOI210     g657(.A0(new_new_n675_), .A1(new_new_n330_), .B0(new_new_n679_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n383_), .B(new_new_n640_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n681_), .B(new_new_n239_), .Y(new_new_n682_));
  AOI210     g660(.A0(new_new_n447_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n683_));
  NOi31      g661(.An(new_new_n683_), .B(new_new_n586_), .C(new_new_n44_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n125_), .B(i_13_), .Y(new_new_n685_));
  NO2        g663(.A(new_new_n639_), .B(new_new_n112_), .Y(new_new_n686_));
  INV        g664(.A(new_new_n686_), .Y(new_new_n687_));
  OAI220     g665(.A0(new_new_n687_), .A1(new_new_n68_), .B0(new_new_n685_), .B1(new_new_n668_), .Y(new_new_n688_));
  NO3        g666(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n99_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n26_), .B(new_new_n192_), .Y(new_new_n690_));
  INV        g668(.A(i_7_), .Y(new_new_n691_));
  INV        g669(.A(new_new_n689_), .Y(new_new_n692_));
  AOI220     g670(.A0(new_new_n383_), .A1(new_new_n640_), .B0(new_new_n90_), .B1(new_new_n100_), .Y(new_new_n693_));
  OAI220     g671(.A0(new_new_n693_), .A1(new_new_n592_), .B0(new_new_n692_), .B1(new_new_n607_), .Y(new_new_n694_));
  NO4        g672(.A(new_new_n694_), .B(new_new_n688_), .C(new_new_n684_), .D(new_new_n682_), .Y(new_new_n695_));
  OR2        g673(.A(i_11_), .B(i_6_), .Y(new_new_n696_));
  NA3        g674(.A(new_new_n591_), .B(new_new_n690_), .C(i_7_), .Y(new_new_n697_));
  AOI210     g675(.A0(new_new_n697_), .A1(new_new_n687_), .B0(new_new_n696_), .Y(new_new_n698_));
  NA3        g676(.A(new_new_n408_), .B(new_new_n596_), .C(new_new_n95_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n630_), .B(i_13_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n100_), .B(new_new_n690_), .Y(new_new_n701_));
  NAi21      g679(.An(i_11_), .B(i_12_), .Y(new_new_n702_));
  NOi41      g680(.An(new_new_n108_), .B(new_new_n702_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n703_));
  NA2        g681(.A(new_new_n703_), .B(new_new_n701_), .Y(new_new_n704_));
  NA3        g682(.A(new_new_n704_), .B(new_new_n700_), .C(new_new_n699_), .Y(new_new_n705_));
  OAI210     g683(.A0(new_new_n705_), .A1(new_new_n698_), .B0(new_new_n60_), .Y(new_new_n706_));
  NO2        g684(.A(i_2_), .B(i_12_), .Y(new_new_n707_));
  NA2        g685(.A(new_new_n364_), .B(new_new_n707_), .Y(new_new_n708_));
  NA2        g686(.A(i_8_), .B(new_new_n25_), .Y(new_new_n709_));
  NO3        g687(.A(new_new_n709_), .B(new_new_n381_), .C(new_new_n591_), .Y(new_new_n710_));
  OAI210     g688(.A0(new_new_n710_), .A1(new_new_n366_), .B0(new_new_n364_), .Y(new_new_n711_));
  NO2        g689(.A(new_new_n126_), .B(i_2_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n712_), .B(new_new_n625_), .Y(new_new_n713_));
  NA3        g691(.A(new_new_n713_), .B(new_new_n711_), .C(new_new_n708_), .Y(new_new_n714_));
  NA3        g692(.A(new_new_n714_), .B(new_new_n45_), .C(new_new_n222_), .Y(new_new_n715_));
  NA4        g693(.A(new_new_n715_), .B(new_new_n706_), .C(new_new_n695_), .D(new_new_n680_), .Y(new_new_n716_));
  OR4        g694(.A(new_new_n716_), .B(new_new_n671_), .C(new_new_n661_), .D(new_new_n610_), .Y(men5));
  NA2        g695(.A(new_new_n655_), .B(new_new_n268_), .Y(new_new_n718_));
  AN2        g696(.A(new_new_n24_), .B(i_10_), .Y(new_new_n719_));
  NA3        g697(.A(new_new_n719_), .B(new_new_n707_), .C(new_new_n106_), .Y(new_new_n720_));
  NO2        g698(.A(new_new_n592_), .B(i_11_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n85_), .B(new_new_n721_), .Y(new_new_n722_));
  NA3        g700(.A(new_new_n722_), .B(new_new_n720_), .C(new_new_n718_), .Y(new_new_n723_));
  NO3        g701(.A(i_11_), .B(new_new_n234_), .C(i_13_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n122_), .B(new_new_n23_), .Y(new_new_n725_));
  NA2        g703(.A(i_12_), .B(i_8_), .Y(new_new_n726_));
  OAI210     g704(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n726_), .Y(new_new_n727_));
  INV        g705(.A(new_new_n446_), .Y(new_new_n728_));
  AOI220     g706(.A0(new_new_n314_), .A1(new_new_n569_), .B0(new_new_n727_), .B1(new_new_n725_), .Y(new_new_n729_));
  INV        g707(.A(new_new_n729_), .Y(new_new_n730_));
  NO2        g708(.A(new_new_n730_), .B(new_new_n723_), .Y(new_new_n731_));
  INV        g709(.A(new_new_n169_), .Y(new_new_n732_));
  INV        g710(.A(new_new_n242_), .Y(new_new_n733_));
  OAI210     g711(.A0(new_new_n669_), .A1(new_new_n448_), .B0(new_new_n108_), .Y(new_new_n734_));
  AOI210     g712(.A0(new_new_n734_), .A1(new_new_n733_), .B0(new_new_n732_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n456_), .B(new_new_n26_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n736_), .B(new_new_n417_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n737_), .B(i_2_), .Y(new_new_n738_));
  INV        g716(.A(new_new_n738_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n415_), .Y(new_new_n740_));
  AOI210     g718(.A0(new_new_n740_), .A1(new_new_n739_), .B0(new_new_n735_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n189_), .B(new_new_n123_), .Y(new_new_n742_));
  OAI210     g720(.A0(new_new_n742_), .A1(new_new_n725_), .B0(i_2_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n170_), .Y(new_new_n744_));
  NO3        g722(.A(new_new_n612_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n744_), .A1(new_new_n85_), .B0(new_new_n745_), .Y(new_new_n746_));
  AOI210     g724(.A0(new_new_n746_), .A1(new_new_n743_), .B0(new_new_n192_), .Y(new_new_n747_));
  OA210      g725(.A0(new_new_n613_), .A1(new_new_n124_), .B0(i_13_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n148_), .B(new_new_n587_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n749_), .B(new_new_n369_), .Y(new_new_n750_));
  AOI210     g728(.A0(new_new_n207_), .A1(new_new_n145_), .B0(new_new_n520_), .Y(new_new_n751_));
  NA2        g729(.A(new_new_n751_), .B(new_new_n417_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n100_), .B(new_new_n44_), .Y(new_new_n753_));
  INV        g731(.A(new_new_n298_), .Y(new_new_n754_));
  NA4        g732(.A(new_new_n754_), .B(new_new_n302_), .C(new_new_n122_), .D(new_new_n42_), .Y(new_new_n755_));
  OAI210     g733(.A0(new_new_n755_), .A1(new_new_n753_), .B0(new_new_n752_), .Y(new_new_n756_));
  NO4        g734(.A(new_new_n756_), .B(new_new_n750_), .C(new_new_n748_), .D(new_new_n747_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n569_), .B(new_new_n28_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n724_), .B(new_new_n272_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n759_), .B(new_new_n758_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n59_), .B(i_12_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n761_), .B(new_new_n124_), .Y(new_new_n762_));
  NO2        g740(.A(new_new_n762_), .B(new_new_n587_), .Y(new_new_n763_));
  AOI220     g741(.A0(new_new_n763_), .A1(new_new_n36_), .B0(new_new_n760_), .B1(new_new_n46_), .Y(new_new_n764_));
  NA4        g742(.A(new_new_n764_), .B(new_new_n757_), .C(new_new_n741_), .D(new_new_n731_), .Y(men6));
  NO3        g743(.A(new_new_n253_), .B(new_new_n304_), .C(i_1_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n184_), .B(new_new_n136_), .Y(new_new_n767_));
  OAI210     g745(.A0(new_new_n767_), .A1(new_new_n766_), .B0(new_new_n712_), .Y(new_new_n768_));
  NA4        g746(.A(new_new_n387_), .B(new_new_n482_), .C(new_new_n68_), .D(new_new_n99_), .Y(new_new_n769_));
  INV        g747(.A(new_new_n769_), .Y(new_new_n770_));
  NO2        g748(.A(new_new_n217_), .B(new_new_n486_), .Y(new_new_n771_));
  NO2        g749(.A(i_11_), .B(i_9_), .Y(new_new_n772_));
  NO2        g750(.A(new_new_n770_), .B(new_new_n326_), .Y(new_new_n773_));
  AO210      g751(.A0(new_new_n773_), .A1(new_new_n768_), .B0(i_12_), .Y(new_new_n774_));
  NA2        g752(.A(new_new_n370_), .B(new_new_n333_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n574_), .B(new_new_n60_), .Y(new_new_n776_));
  BUFFER     g754(.A(new_new_n616_), .Y(new_new_n777_));
  NA3        g755(.A(new_new_n777_), .B(new_new_n776_), .C(new_new_n775_), .Y(new_new_n778_));
  INV        g756(.A(new_new_n195_), .Y(new_new_n779_));
  AOI220     g757(.A0(new_new_n779_), .A1(new_new_n772_), .B0(new_new_n778_), .B1(new_new_n70_), .Y(new_new_n780_));
  INV        g758(.A(new_new_n325_), .Y(new_new_n781_));
  NA2        g759(.A(new_new_n72_), .B(new_new_n129_), .Y(new_new_n782_));
  INV        g760(.A(new_new_n122_), .Y(new_new_n783_));
  NA2        g761(.A(new_new_n783_), .B(new_new_n46_), .Y(new_new_n784_));
  AOI210     g762(.A0(new_new_n784_), .A1(new_new_n782_), .B0(new_new_n781_), .Y(new_new_n785_));
  NO2        g763(.A(new_new_n249_), .B(i_9_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n786_), .B(new_new_n761_), .Y(new_new_n787_));
  AOI210     g765(.A0(new_new_n787_), .A1(new_new_n518_), .B0(new_new_n184_), .Y(new_new_n788_));
  NAi32      g766(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n789_));
  NO2        g767(.A(new_new_n696_), .B(new_new_n789_), .Y(new_new_n790_));
  OR3        g768(.A(new_new_n790_), .B(new_new_n788_), .C(new_new_n785_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n672_), .B(i_2_), .Y(new_new_n792_));
  NA2        g770(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n793_), .B(new_new_n407_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n794_), .B(new_new_n792_), .Y(new_new_n795_));
  OR2        g773(.A(new_new_n613_), .B(new_new_n448_), .Y(new_new_n796_));
  NA3        g774(.A(new_new_n796_), .B(new_new_n144_), .C(new_new_n66_), .Y(new_new_n797_));
  AO210      g775(.A0(new_new_n492_), .A1(new_new_n728_), .B0(new_new_n36_), .Y(new_new_n798_));
  NA3        g776(.A(new_new_n798_), .B(new_new_n797_), .C(new_new_n795_), .Y(new_new_n799_));
  OAI210     g777(.A0(new_new_n629_), .A1(i_11_), .B0(new_new_n83_), .Y(new_new_n800_));
  AOI220     g778(.A0(new_new_n800_), .A1(new_new_n559_), .B0(new_new_n771_), .B1(new_new_n691_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n393_), .B(new_new_n67_), .Y(new_new_n802_));
  NA3        g780(.A(new_new_n802_), .B(new_new_n801_), .C(new_new_n595_), .Y(new_new_n803_));
  AO210      g781(.A0(new_new_n520_), .A1(new_new_n46_), .B0(new_new_n84_), .Y(new_new_n804_));
  NA3        g782(.A(new_new_n804_), .B(new_new_n483_), .C(new_new_n216_), .Y(new_new_n805_));
  AOI210     g783(.A0(new_new_n448_), .A1(new_new_n446_), .B0(new_new_n558_), .Y(new_new_n806_));
  NA2        g784(.A(new_new_n109_), .B(new_new_n406_), .Y(new_new_n807_));
  INV        g785(.A(new_new_n241_), .Y(new_new_n808_));
  NA3        g786(.A(new_new_n807_), .B(new_new_n806_), .C(new_new_n805_), .Y(new_new_n809_));
  NO4        g787(.A(new_new_n809_), .B(new_new_n803_), .C(new_new_n799_), .D(new_new_n791_), .Y(new_new_n810_));
  NA4        g788(.A(new_new_n810_), .B(new_new_n780_), .C(new_new_n774_), .D(new_new_n377_), .Y(men3));
  NA2        g789(.A(i_6_), .B(i_7_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n812_), .B(i_0_), .Y(new_new_n813_));
  NO2        g791(.A(i_11_), .B(new_new_n234_), .Y(new_new_n814_));
  OAI210     g792(.A0(new_new_n813_), .A1(new_new_n286_), .B0(new_new_n814_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n815_), .B(new_new_n192_), .Y(new_new_n816_));
  NO3        g794(.A(new_new_n452_), .B(new_new_n88_), .C(new_new_n44_), .Y(new_new_n817_));
  OA210      g795(.A0(new_new_n817_), .A1(new_new_n816_), .B0(new_new_n172_), .Y(new_new_n818_));
  NA2        g796(.A(new_new_n595_), .B(new_new_n368_), .Y(new_new_n819_));
  NA2        g797(.A(new_new_n819_), .B(new_new_n40_), .Y(new_new_n820_));
  NO3        g798(.A(new_new_n620_), .B(new_new_n456_), .C(new_new_n129_), .Y(new_new_n821_));
  AN2        g799(.A(new_new_n454_), .B(new_new_n53_), .Y(new_new_n822_));
  NO2        g800(.A(new_new_n822_), .B(new_new_n821_), .Y(new_new_n823_));
  AOI210     g801(.A0(new_new_n823_), .A1(new_new_n820_), .B0(new_new_n48_), .Y(new_new_n824_));
  NO4        g802(.A(new_new_n373_), .B(new_new_n380_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n184_), .B(new_new_n567_), .Y(new_new_n826_));
  NOi21      g804(.An(new_new_n826_), .B(new_new_n825_), .Y(new_new_n827_));
  NO2        g805(.A(new_new_n827_), .B(new_new_n60_), .Y(new_new_n828_));
  NOi21      g806(.An(i_5_), .B(i_9_), .Y(new_new_n829_));
  NA2        g807(.A(new_new_n829_), .B(new_new_n445_), .Y(new_new_n830_));
  BUFFER     g808(.A(new_new_n266_), .Y(new_new_n831_));
  AOI210     g809(.A0(new_new_n831_), .A1(new_new_n475_), .B0(new_new_n663_), .Y(new_new_n832_));
  NO2        g810(.A(new_new_n173_), .B(new_new_n145_), .Y(new_new_n833_));
  NO2        g811(.A(new_new_n832_), .B(new_new_n830_), .Y(new_new_n834_));
  NO4        g812(.A(new_new_n834_), .B(new_new_n828_), .C(new_new_n824_), .D(new_new_n818_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n184_), .B(new_new_n24_), .Y(new_new_n836_));
  NO2        g814(.A(new_new_n657_), .B(new_new_n584_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n836_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n309_), .B(new_new_n127_), .Y(new_new_n839_));
  NAi21      g817(.An(new_new_n159_), .B(new_new_n437_), .Y(new_new_n840_));
  OAI220     g818(.A0(new_new_n840_), .A1(new_new_n808_), .B0(new_new_n839_), .B1(new_new_n398_), .Y(new_new_n841_));
  NO2        g819(.A(new_new_n841_), .B(new_new_n838_), .Y(new_new_n842_));
  NO2        g820(.A(new_new_n387_), .B(new_new_n290_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n843_), .B(new_new_n686_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n568_), .B(i_0_), .Y(new_new_n845_));
  NO3        g823(.A(new_new_n845_), .B(new_new_n382_), .C(new_new_n85_), .Y(new_new_n846_));
  INV        g824(.A(new_new_n846_), .Y(new_new_n847_));
  AN2        g825(.A(new_new_n94_), .B(new_new_n240_), .Y(new_new_n848_));
  NA2        g826(.A(new_new_n724_), .B(new_new_n326_), .Y(new_new_n849_));
  INV        g827(.A(new_new_n55_), .Y(new_new_n850_));
  OAI220     g828(.A0(new_new_n850_), .A1(new_new_n849_), .B0(new_new_n650_), .B1(new_new_n537_), .Y(new_new_n851_));
  NO2        g829(.A(new_new_n251_), .B(new_new_n150_), .Y(new_new_n852_));
  NA2        g830(.A(i_0_), .B(i_10_), .Y(new_new_n853_));
  AN2        g831(.A(new_new_n852_), .B(i_6_), .Y(new_new_n854_));
  AOI220     g832(.A0(new_new_n331_), .A1(new_new_n96_), .B0(new_new_n184_), .B1(new_new_n80_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n563_), .B(i_4_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n187_), .B(new_new_n201_), .Y(new_new_n857_));
  OAI220     g835(.A0(new_new_n857_), .A1(new_new_n849_), .B0(new_new_n856_), .B1(new_new_n855_), .Y(new_new_n858_));
  NO4        g836(.A(new_new_n858_), .B(new_new_n854_), .C(new_new_n851_), .D(new_new_n848_), .Y(new_new_n859_));
  NA4        g837(.A(new_new_n859_), .B(new_new_n847_), .C(new_new_n844_), .D(new_new_n842_), .Y(new_new_n860_));
  NO2        g838(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n861_));
  NA2        g839(.A(i_11_), .B(i_9_), .Y(new_new_n862_));
  NO3        g840(.A(i_12_), .B(new_new_n862_), .C(new_new_n594_), .Y(new_new_n863_));
  AN2        g841(.A(new_new_n863_), .B(new_new_n861_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n48_), .B(i_7_), .Y(new_new_n865_));
  NA2        g843(.A(new_new_n391_), .B(new_new_n177_), .Y(new_new_n866_));
  NA2        g844(.A(new_new_n866_), .B(new_new_n157_), .Y(new_new_n867_));
  NO2        g845(.A(new_new_n173_), .B(i_0_), .Y(new_new_n868_));
  INV        g846(.A(new_new_n868_), .Y(new_new_n869_));
  NA2        g847(.A(new_new_n473_), .B(new_new_n228_), .Y(new_new_n870_));
  INV        g848(.A(new_new_n405_), .Y(new_new_n871_));
  OAI220     g849(.A0(new_new_n871_), .A1(new_new_n830_), .B0(new_new_n870_), .B1(new_new_n869_), .Y(new_new_n872_));
  NO3        g850(.A(new_new_n872_), .B(new_new_n867_), .C(new_new_n864_), .Y(new_new_n873_));
  NA2        g851(.A(new_new_n649_), .B(new_new_n119_), .Y(new_new_n874_));
  NO2        g852(.A(i_6_), .B(new_new_n874_), .Y(new_new_n875_));
  AOI210     g853(.A0(new_new_n447_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n876_));
  NA2        g854(.A(new_new_n169_), .B(new_new_n101_), .Y(new_new_n877_));
  NOi32      g855(.An(new_new_n876_), .Bn(new_new_n187_), .C(new_new_n877_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n878_), .B(new_new_n875_), .Y(new_new_n879_));
  NOi21      g857(.An(i_7_), .B(i_5_), .Y(new_new_n880_));
  NOi31      g858(.An(new_new_n880_), .B(i_0_), .C(new_new_n702_), .Y(new_new_n881_));
  NA3        g859(.A(new_new_n881_), .B(new_new_n381_), .C(i_6_), .Y(new_new_n882_));
  OA210      g860(.A0(new_new_n877_), .A1(new_new_n518_), .B0(new_new_n882_), .Y(new_new_n883_));
  NO3        g861(.A(new_new_n401_), .B(new_new_n359_), .C(new_new_n357_), .Y(new_new_n884_));
  NO2        g862(.A(new_new_n260_), .B(new_new_n315_), .Y(new_new_n885_));
  NO2        g863(.A(new_new_n702_), .B(new_new_n255_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n886_), .A1(new_new_n885_), .B0(new_new_n884_), .Y(new_new_n887_));
  NA4        g865(.A(new_new_n887_), .B(new_new_n883_), .C(new_new_n879_), .D(new_new_n873_), .Y(new_new_n888_));
  NO2        g866(.A(new_new_n836_), .B(new_new_n236_), .Y(new_new_n889_));
  AN2        g867(.A(new_new_n330_), .B(new_new_n326_), .Y(new_new_n890_));
  AN2        g868(.A(new_new_n890_), .B(new_new_n833_), .Y(new_new_n891_));
  OAI210     g869(.A0(new_new_n891_), .A1(new_new_n889_), .B0(i_10_), .Y(new_new_n892_));
  OA210      g870(.A0(new_new_n473_), .A1(new_new_n220_), .B0(new_new_n472_), .Y(new_new_n893_));
  NA3        g871(.A(new_new_n472_), .B(new_new_n408_), .C(new_new_n45_), .Y(new_new_n894_));
  INV        g872(.A(new_new_n894_), .Y(new_new_n895_));
  NO2        g873(.A(i_3_), .B(new_new_n186_), .Y(new_new_n896_));
  AOI220     g874(.A0(new_new_n896_), .A1(new_new_n473_), .B0(new_new_n895_), .B1(new_new_n70_), .Y(new_new_n897_));
  NA3        g875(.A(new_new_n793_), .B(new_new_n379_), .C(new_new_n629_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n91_), .B(new_new_n44_), .Y(new_new_n899_));
  NO2        g877(.A(new_new_n72_), .B(new_new_n726_), .Y(new_new_n900_));
  AOI220     g878(.A0(new_new_n900_), .A1(new_new_n899_), .B0(new_new_n172_), .B1(new_new_n584_), .Y(new_new_n901_));
  AOI210     g879(.A0(new_new_n901_), .A1(new_new_n898_), .B0(new_new_n47_), .Y(new_new_n902_));
  NAi21      g880(.An(i_9_), .B(i_5_), .Y(new_new_n903_));
  NO2        g881(.A(new_new_n903_), .B(new_new_n401_), .Y(new_new_n904_));
  NO2        g882(.A(new_new_n590_), .B(new_new_n103_), .Y(new_new_n905_));
  AOI220     g883(.A0(new_new_n905_), .A1(i_0_), .B0(new_new_n904_), .B1(new_new_n613_), .Y(new_new_n906_));
  NO2        g884(.A(new_new_n906_), .B(new_new_n82_), .Y(new_new_n907_));
  NO3        g885(.A(new_new_n907_), .B(new_new_n902_), .C(new_new_n523_), .Y(new_new_n908_));
  NA3        g886(.A(new_new_n908_), .B(new_new_n897_), .C(new_new_n892_), .Y(new_new_n909_));
  NO3        g887(.A(new_new_n909_), .B(new_new_n888_), .C(new_new_n860_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n70_), .B(new_new_n44_), .Y(new_new_n911_));
  NA2        g889(.A(new_new_n853_), .B(new_new_n911_), .Y(new_new_n912_));
  NO3        g890(.A(new_new_n103_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n913_));
  AN2        g891(.A(new_new_n913_), .B(new_new_n912_), .Y(new_new_n914_));
  AOI210     g892(.A0(new_new_n776_), .A1(new_new_n662_), .B0(new_new_n877_), .Y(new_new_n915_));
  AOI210     g893(.A0(new_new_n914_), .A1(new_new_n348_), .B0(new_new_n915_), .Y(new_new_n916_));
  NA2        g894(.A(new_new_n712_), .B(new_new_n143_), .Y(new_new_n917_));
  INV        g895(.A(new_new_n917_), .Y(new_new_n918_));
  NA3        g896(.A(new_new_n918_), .B(new_new_n658_), .C(new_new_n70_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n813_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n814_), .B(i_9_), .Y(new_new_n921_));
  AOI210     g899(.A0(new_new_n920_), .A1(new_new_n497_), .B0(new_new_n921_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n241_), .B(new_new_n227_), .Y(new_new_n923_));
  AOI210     g901(.A0(new_new_n923_), .A1(new_new_n845_), .B0(new_new_n150_), .Y(new_new_n924_));
  NO2        g902(.A(new_new_n924_), .B(new_new_n922_), .Y(new_new_n925_));
  NA3        g903(.A(new_new_n925_), .B(new_new_n919_), .C(new_new_n916_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n890_), .B(new_new_n369_), .Y(new_new_n927_));
  AOI210     g905(.A0(new_new_n297_), .A1(new_new_n159_), .B0(new_new_n927_), .Y(new_new_n928_));
  NA2        g906(.A(new_new_n40_), .B(new_new_n44_), .Y(new_new_n929_));
  NA2        g907(.A(new_new_n865_), .B(new_new_n487_), .Y(new_new_n930_));
  AOI210     g908(.A0(new_new_n929_), .A1(new_new_n159_), .B0(new_new_n930_), .Y(new_new_n931_));
  NO2        g909(.A(new_new_n931_), .B(new_new_n928_), .Y(new_new_n932_));
  NO3        g910(.A(new_new_n853_), .B(new_new_n829_), .C(new_new_n189_), .Y(new_new_n933_));
  AOI220     g911(.A0(new_new_n933_), .A1(i_11_), .B0(new_new_n564_), .B1(new_new_n72_), .Y(new_new_n934_));
  NO3        g912(.A(new_new_n209_), .B(new_new_n380_), .C(i_0_), .Y(new_new_n935_));
  OAI210     g913(.A0(new_new_n935_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n936_));
  INV        g914(.A(new_new_n216_), .Y(new_new_n937_));
  NO2        g915(.A(new_new_n531_), .B(new_new_n136_), .Y(new_new_n938_));
  NA3        g916(.A(new_new_n938_), .B(new_new_n1017_), .C(new_new_n937_), .Y(new_new_n939_));
  NA4        g917(.A(new_new_n939_), .B(new_new_n936_), .C(new_new_n934_), .D(new_new_n932_), .Y(new_new_n940_));
  AOI220     g918(.A0(new_new_n880_), .A1(new_new_n487_), .B0(new_new_n813_), .B1(new_new_n160_), .Y(new_new_n941_));
  NA2        g919(.A(new_new_n351_), .B(new_new_n174_), .Y(new_new_n942_));
  OR2        g920(.A(new_new_n942_), .B(new_new_n941_), .Y(new_new_n943_));
  AOI210     g921(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n173_), .Y(new_new_n944_));
  NA2        g922(.A(new_new_n944_), .B(new_new_n893_), .Y(new_new_n945_));
  NA3        g923(.A(new_new_n387_), .B(new_new_n169_), .C(new_new_n168_), .Y(new_new_n946_));
  NA3        g924(.A(new_new_n865_), .B(new_new_n286_), .C(new_new_n227_), .Y(new_new_n947_));
  NA2        g925(.A(new_new_n947_), .B(new_new_n946_), .Y(new_new_n948_));
  NA3        g926(.A(new_new_n387_), .B(new_new_n332_), .C(new_new_n218_), .Y(new_new_n949_));
  INV        g927(.A(new_new_n949_), .Y(new_new_n950_));
  NOi31      g928(.An(new_new_n386_), .B(new_new_n911_), .C(new_new_n236_), .Y(new_new_n951_));
  NO3        g929(.A(new_new_n951_), .B(new_new_n950_), .C(new_new_n948_), .Y(new_new_n952_));
  NA3        g930(.A(new_new_n952_), .B(new_new_n945_), .C(new_new_n943_), .Y(new_new_n953_));
  NO2        g931(.A(new_new_n82_), .B(i_5_), .Y(new_new_n954_));
  NA3        g932(.A(new_new_n814_), .B(new_new_n107_), .C(new_new_n122_), .Y(new_new_n955_));
  INV        g933(.A(new_new_n955_), .Y(new_new_n956_));
  NA2        g934(.A(new_new_n956_), .B(new_new_n954_), .Y(new_new_n957_));
  NA2        g935(.A(new_new_n770_), .B(new_new_n174_), .Y(new_new_n958_));
  AN2        g936(.A(new_new_n853_), .B(new_new_n150_), .Y(new_new_n959_));
  NO4        g937(.A(new_new_n959_), .B(i_12_), .C(new_new_n637_), .D(new_new_n129_), .Y(new_new_n960_));
  NA2        g938(.A(new_new_n960_), .B(new_new_n216_), .Y(new_new_n961_));
  NA3        g939(.A(new_new_n96_), .B(new_new_n567_), .C(i_11_), .Y(new_new_n962_));
  NO2        g940(.A(new_new_n962_), .B(new_new_n152_), .Y(new_new_n963_));
  NA2        g941(.A(new_new_n880_), .B(new_new_n470_), .Y(new_new_n964_));
  NO2        g942(.A(new_new_n964_), .B(new_new_n659_), .Y(new_new_n965_));
  AOI210     g943(.A0(new_new_n965_), .A1(new_new_n868_), .B0(new_new_n963_), .Y(new_new_n966_));
  NA4        g944(.A(new_new_n966_), .B(new_new_n961_), .C(new_new_n958_), .D(new_new_n957_), .Y(new_new_n967_));
  NO4        g945(.A(new_new_n967_), .B(new_new_n953_), .C(new_new_n940_), .D(new_new_n926_), .Y(new_new_n968_));
  NA2        g946(.A(new_new_n792_), .B(new_new_n37_), .Y(new_new_n969_));
  NA3        g947(.A(new_new_n876_), .B(new_new_n364_), .C(i_5_), .Y(new_new_n970_));
  NA3        g948(.A(new_new_n970_), .B(new_new_n969_), .C(new_new_n602_), .Y(new_new_n971_));
  NA2        g949(.A(new_new_n971_), .B(new_new_n205_), .Y(new_new_n972_));
  NA2        g950(.A(new_new_n185_), .B(new_new_n187_), .Y(new_new_n973_));
  AO210      g951(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n973_), .Y(new_new_n974_));
  OAI210     g952(.A0(new_new_n606_), .A1(new_new_n604_), .B0(new_new_n314_), .Y(new_new_n975_));
  NAi31      g953(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n976_));
  AOI210     g954(.A0(new_new_n115_), .A1(new_new_n67_), .B0(new_new_n976_), .Y(new_new_n977_));
  NO2        g955(.A(new_new_n977_), .B(new_new_n634_), .Y(new_new_n978_));
  NA3        g956(.A(new_new_n978_), .B(new_new_n975_), .C(new_new_n974_), .Y(new_new_n979_));
  NO2        g957(.A(new_new_n460_), .B(new_new_n266_), .Y(new_new_n980_));
  NO4        g958(.A(new_new_n230_), .B(new_new_n142_), .C(new_new_n660_), .D(new_new_n37_), .Y(new_new_n981_));
  NO2        g959(.A(new_new_n981_), .B(new_new_n980_), .Y(new_new_n982_));
  OAI210     g960(.A0(new_new_n962_), .A1(new_new_n145_), .B0(new_new_n982_), .Y(new_new_n983_));
  AOI210     g961(.A0(new_new_n979_), .A1(new_new_n48_), .B0(new_new_n983_), .Y(new_new_n984_));
  AOI210     g962(.A0(new_new_n984_), .A1(new_new_n972_), .B0(new_new_n70_), .Y(new_new_n985_));
  NO2        g963(.A(new_new_n561_), .B(new_new_n376_), .Y(new_new_n986_));
  NO2        g964(.A(new_new_n986_), .B(new_new_n732_), .Y(new_new_n987_));
  OAI210     g965(.A0(new_new_n77_), .A1(new_new_n52_), .B0(new_new_n106_), .Y(new_new_n988_));
  NA2        g966(.A(new_new_n988_), .B(new_new_n73_), .Y(new_new_n989_));
  AOI210     g967(.A0(new_new_n944_), .A1(new_new_n865_), .B0(new_new_n881_), .Y(new_new_n990_));
  AOI210     g968(.A0(new_new_n990_), .A1(new_new_n989_), .B0(new_new_n660_), .Y(new_new_n991_));
  NA2        g969(.A(new_new_n260_), .B(new_new_n54_), .Y(new_new_n992_));
  AOI220     g970(.A0(new_new_n992_), .A1(new_new_n73_), .B0(new_new_n346_), .B1(new_new_n253_), .Y(new_new_n993_));
  NO2        g971(.A(new_new_n993_), .B(new_new_n234_), .Y(new_new_n994_));
  NA3        g972(.A(new_new_n94_), .B(new_new_n304_), .C(new_new_n31_), .Y(new_new_n995_));
  INV        g973(.A(new_new_n995_), .Y(new_new_n996_));
  NO3        g974(.A(new_new_n996_), .B(new_new_n994_), .C(new_new_n991_), .Y(new_new_n997_));
  OAI210     g975(.A0(new_new_n1015_), .A1(new_new_n876_), .B0(new_new_n205_), .Y(new_new_n998_));
  NA2        g976(.A(new_new_n161_), .B(i_5_), .Y(new_new_n999_));
  NO2        g977(.A(new_new_n998_), .B(new_new_n999_), .Y(new_new_n1000_));
  NO3        g978(.A(new_new_n56_), .B(new_new_n55_), .C(i_4_), .Y(new_new_n1001_));
  OAI210     g979(.A0(new_new_n885_), .A1(new_new_n304_), .B0(new_new_n1001_), .Y(new_new_n1002_));
  NO2        g980(.A(new_new_n1002_), .B(new_new_n702_), .Y(new_new_n1003_));
  INV        g981(.A(new_new_n360_), .Y(new_new_n1004_));
  NO2        g982(.A(new_new_n1004_), .B(new_new_n41_), .Y(new_new_n1005_));
  NO3        g983(.A(new_new_n1005_), .B(new_new_n1003_), .C(new_new_n1000_), .Y(new_new_n1006_));
  OAI210     g984(.A0(new_new_n997_), .A1(i_4_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  NO3        g985(.A(new_new_n1007_), .B(new_new_n987_), .C(new_new_n985_), .Y(new_new_n1008_));
  NA4        g986(.A(new_new_n1008_), .B(new_new_n968_), .C(new_new_n910_), .D(new_new_n835_), .Y(men4));
  INV        g987(.A(new_new_n676_), .Y(new_new_n1012_));
  INV        g988(.A(i_2_), .Y(new_new_n1013_));
  INV        g989(.A(new_new_n483_), .Y(new_new_n1014_));
  INV        g990(.A(i_12_), .Y(new_new_n1015_));
  INV        g991(.A(i_12_), .Y(new_new_n1016_));
  INV        g992(.A(i_3_), .Y(new_new_n1017_));
endmodule


