// Benchmark "top" written by ABC on Fri Jun 21 17:49:20 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n133_, new_new_n134_, new_new_n135_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1093_, new_new_n1094_, new_new_n1095_,
    new_new_n1096_, new_new_n1097_, new_new_n1098_, new_new_n1099_,
    new_new_n1100_, new_new_n1101_, new_new_n1102_, new_new_n1103_,
    new_new_n1104_, new_new_n1105_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_5_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n51_));
  NA2        g0029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g0030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NO2        g0031(.A(new_new_n53_), .B(new_new_n52_), .Y(new_new_n54_));
  OAI210     g0032(.A0(new_new_n54_), .A1(new_new_n51_), .B0(new_new_n45_), .Y(new_new_n55_));
  NA3        g0033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g0034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g0035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  OAI210     g0036(.A0(new_new_n58_), .A1(new_new_n57_), .B0(new_new_n56_), .Y(new_new_n59_));
  NA2        g0037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g0038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g0039(.A(i_1_), .Y(new_new_n62_));
  NA2        g0040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA2        g0041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi21      g0043(.An(new_new_n65_), .B(new_new_n60_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n50_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g0053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n62_), .Y(new_new_n83_));
  INV        g0061(.A(i_6_), .Y(new_new_n84_));
  OR4        g0062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n85_));
  INV        g0063(.A(new_new_n85_), .Y(new_new_n86_));
  NO2        g0064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  OAI210     g0065(.A0(new_new_n83_), .A1(new_new_n80_), .B0(new_new_n85_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n62_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n90_), .A1(new_new_n88_), .B0(new_new_n78_), .Y(new_new_n93_));
  AN3        g0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g0072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NO2        g0073(.A(i_5_), .B(i_8_), .Y(new_new_n96_));
  NA2        g0074(.A(new_new_n94_), .B(new_new_n32_), .Y(new_new_n97_));
  INV        g0075(.A(i_7_), .Y(new_new_n98_));
  NO2        g0076(.A(i_0_), .B(i_5_), .Y(new_new_n99_));
  NO2        g0077(.A(new_new_n99_), .B(new_new_n84_), .Y(new_new_n100_));
  NA2        g0078(.A(i_12_), .B(i_3_), .Y(new_new_n101_));
  INV        g0079(.A(new_new_n101_), .Y(new_new_n102_));
  NAi21      g0080(.An(i_7_), .B(i_11_), .Y(new_new_n103_));
  NO3        g0081(.A(new_new_n103_), .B(new_new_n89_), .C(new_new_n52_), .Y(new_new_n104_));
  AN2        g0082(.A(i_2_), .B(i_10_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(i_7_), .Y(new_new_n106_));
  OR2        g0084(.A(new_new_n78_), .B(new_new_n57_), .Y(new_new_n107_));
  NO2        g0085(.A(i_8_), .B(new_new_n98_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NO2        g0087(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n110_));
  NA2        g0088(.A(new_new_n110_), .B(i_0_), .Y(new_new_n111_));
  NA2        g0089(.A(i_11_), .B(i_12_), .Y(new_new_n112_));
  OAI210     g0090(.A0(new_new_n111_), .A1(new_new_n109_), .B0(new_new_n112_), .Y(new_new_n113_));
  INV        g0091(.A(new_new_n113_), .Y(new_new_n114_));
  NAi31      g0092(.An(new_new_n104_), .B(new_new_n114_), .C(new_new_n97_), .Y(new_new_n115_));
  NOi21      g0093(.An(i_1_), .B(i_5_), .Y(new_new_n116_));
  NA2        g0094(.A(new_new_n116_), .B(i_11_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n98_), .B(new_new_n37_), .Y(new_new_n118_));
  NA2        g0096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g0097(.A(new_new_n119_), .B(new_new_n118_), .Y(new_new_n120_));
  NO2        g0098(.A(new_new_n120_), .B(new_new_n46_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n122_));
  NAi21      g0100(.An(i_3_), .B(i_8_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(new_new_n61_), .Y(new_new_n124_));
  NOi31      g0102(.An(new_new_n124_), .B(new_new_n122_), .C(new_new_n121_), .Y(new_new_n125_));
  NO2        g0103(.A(i_1_), .B(new_new_n84_), .Y(new_new_n126_));
  NO2        g0104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  AO210      g0106(.A0(new_new_n128_), .A1(new_new_n47_), .B0(new_new_n126_), .Y(new_new_n129_));
  OAI220     g0107(.A0(new_new_n129_), .A1(new_new_n103_), .B0(new_new_n125_), .B1(new_new_n117_), .Y(new_new_n130_));
  NO3        g0108(.A(new_new_n130_), .B(new_new_n115_), .C(new_new_n93_), .Y(new_new_n131_));
  NA3        g0109(.A(new_new_n131_), .B(new_new_n77_), .C(new_new_n55_), .Y(men2));
  NO2        g0110(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n133_));
  NA2        g0111(.A(i_6_), .B(new_new_n25_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(new_new_n133_), .Y(new_new_n135_));
  NA4        g0113(.A(new_new_n135_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(men0));
  AN2        g0114(.A(i_8_), .B(i_7_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(i_6_), .Y(new_new_n138_));
  NO2        g0116(.A(i_12_), .B(i_13_), .Y(new_new_n139_));
  NAi21      g0117(.An(i_5_), .B(i_11_), .Y(new_new_n140_));
  NOi21      g0118(.An(new_new_n139_), .B(new_new_n140_), .Y(new_new_n141_));
  NO2        g0119(.A(i_0_), .B(i_1_), .Y(new_new_n142_));
  NA2        g0120(.A(i_2_), .B(i_3_), .Y(new_new_n143_));
  NO2        g0121(.A(new_new_n143_), .B(i_4_), .Y(new_new_n144_));
  NA3        g0122(.A(new_new_n144_), .B(new_new_n142_), .C(new_new_n141_), .Y(new_new_n145_));
  OR2        g0123(.A(new_new_n145_), .B(new_new_n25_), .Y(new_new_n146_));
  AN2        g0124(.A(new_new_n139_), .B(new_new_n81_), .Y(new_new_n147_));
  NO2        g0125(.A(new_new_n147_), .B(new_new_n27_), .Y(new_new_n148_));
  NA2        g0126(.A(i_1_), .B(i_5_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n71_), .B(new_new_n46_), .Y(new_new_n150_));
  NA2        g0128(.A(new_new_n150_), .B(new_new_n36_), .Y(new_new_n151_));
  NO3        g0129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  OR2        g0130(.A(i_0_), .B(i_1_), .Y(new_new_n153_));
  NO3        g0131(.A(new_new_n153_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n154_));
  NAi32      g0132(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n155_));
  NAi21      g0133(.An(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  NOi21      g0134(.An(i_4_), .B(i_10_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n39_), .Y(new_new_n158_));
  NO2        g0136(.A(i_3_), .B(i_5_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n160_));
  NA2        g0138(.A(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  OAI210     g0139(.A0(new_new_n161_), .A1(new_new_n158_), .B0(new_new_n156_), .Y(new_new_n162_));
  NO2        g0140(.A(new_new_n162_), .B(new_new_n152_), .Y(new_new_n163_));
  AOI210     g0141(.A0(new_new_n163_), .A1(new_new_n146_), .B0(new_new_n138_), .Y(new_new_n164_));
  NA3        g0142(.A(new_new_n71_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(i_3_), .B(new_new_n48_), .Y(new_new_n166_));
  NOi21      g0144(.An(i_4_), .B(i_9_), .Y(new_new_n167_));
  NOi21      g0145(.An(i_11_), .B(i_13_), .Y(new_new_n168_));
  NA2        g0146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  OR2        g0147(.A(new_new_n169_), .B(new_new_n166_), .Y(new_new_n170_));
  NO2        g0148(.A(i_4_), .B(i_5_), .Y(new_new_n171_));
  NAi21      g0149(.An(i_12_), .B(i_11_), .Y(new_new_n172_));
  NO2        g0150(.A(new_new_n172_), .B(i_13_), .Y(new_new_n173_));
  NA3        g0151(.A(new_new_n173_), .B(new_new_n171_), .C(new_new_n81_), .Y(new_new_n174_));
  AOI210     g0152(.A0(new_new_n174_), .A1(new_new_n170_), .B0(new_new_n165_), .Y(new_new_n175_));
  NO2        g0153(.A(new_new_n71_), .B(new_new_n62_), .Y(new_new_n176_));
  NA2        g0154(.A(new_new_n176_), .B(new_new_n46_), .Y(new_new_n177_));
  NA2        g0155(.A(new_new_n36_), .B(i_5_), .Y(new_new_n178_));
  NAi31      g0156(.An(new_new_n178_), .B(new_new_n147_), .C(i_11_), .Y(new_new_n179_));
  NA2        g0157(.A(i_3_), .B(i_5_), .Y(new_new_n180_));
  OR2        g0158(.A(new_new_n180_), .B(new_new_n169_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n179_), .B0(new_new_n177_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n71_), .B(i_5_), .Y(new_new_n183_));
  NO2        g0161(.A(i_13_), .B(i_10_), .Y(new_new_n184_));
  NA3        g0162(.A(new_new_n184_), .B(new_new_n183_), .C(new_new_n44_), .Y(new_new_n185_));
  NO2        g0163(.A(i_2_), .B(i_1_), .Y(new_new_n186_));
  NA2        g0164(.A(new_new_n186_), .B(i_3_), .Y(new_new_n187_));
  NAi21      g0165(.An(i_4_), .B(i_12_), .Y(new_new_n188_));
  NO4        g0166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n185_), .D(new_new_n25_), .Y(new_new_n189_));
  NO3        g0167(.A(new_new_n189_), .B(new_new_n182_), .C(new_new_n175_), .Y(new_new_n190_));
  INV        g0168(.A(i_8_), .Y(new_new_n191_));
  NO2        g0169(.A(new_new_n191_), .B(i_7_), .Y(new_new_n192_));
  NA2        g0170(.A(new_new_n192_), .B(i_6_), .Y(new_new_n193_));
  NO3        g0171(.A(i_3_), .B(new_new_n84_), .C(new_new_n48_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(new_new_n108_), .Y(new_new_n195_));
  NO3        g0173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n196_));
  NA3        g0174(.A(new_new_n196_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n197_));
  NO3        g0175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n198_));
  OAI210     g0176(.A0(new_new_n94_), .A1(i_12_), .B0(new_new_n198_), .Y(new_new_n199_));
  AOI210     g0177(.A0(new_new_n199_), .A1(new_new_n197_), .B0(new_new_n195_), .Y(new_new_n200_));
  NO2        g0178(.A(i_3_), .B(i_8_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n202_));
  NA3        g0180(.A(new_new_n202_), .B(new_new_n201_), .C(new_new_n39_), .Y(new_new_n203_));
  NO2        g0181(.A(new_new_n99_), .B(new_new_n57_), .Y(new_new_n204_));
  NO2        g0182(.A(i_13_), .B(i_9_), .Y(new_new_n205_));
  NA3        g0183(.A(new_new_n205_), .B(i_6_), .C(new_new_n191_), .Y(new_new_n206_));
  NAi21      g0184(.An(i_12_), .B(i_3_), .Y(new_new_n207_));
  OR2        g0185(.A(new_new_n207_), .B(new_new_n206_), .Y(new_new_n208_));
  NO2        g0186(.A(new_new_n44_), .B(i_5_), .Y(new_new_n209_));
  NA2        g0187(.A(new_new_n209_), .B(i_10_), .Y(new_new_n210_));
  OAI220     g0188(.A0(new_new_n210_), .A1(new_new_n208_), .B0(new_new_n99_), .B1(new_new_n203_), .Y(new_new_n211_));
  AOI210     g0189(.A0(new_new_n211_), .A1(i_7_), .B0(new_new_n200_), .Y(new_new_n212_));
  OAI220     g0190(.A0(new_new_n212_), .A1(i_4_), .B0(new_new_n193_), .B1(new_new_n190_), .Y(new_new_n213_));
  NAi21      g0191(.An(i_12_), .B(i_7_), .Y(new_new_n214_));
  NA3        g0192(.A(i_13_), .B(new_new_n191_), .C(i_10_), .Y(new_new_n215_));
  NO2        g0193(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n216_));
  NA2        g0194(.A(i_0_), .B(i_5_), .Y(new_new_n217_));
  NA2        g0195(.A(new_new_n217_), .B(new_new_n100_), .Y(new_new_n218_));
  OAI220     g0196(.A0(new_new_n218_), .A1(new_new_n187_), .B0(new_new_n177_), .B1(new_new_n128_), .Y(new_new_n219_));
  NAi31      g0197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n36_), .B(i_13_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n223_));
  NA3        g0201(.A(new_new_n223_), .B(new_new_n222_), .C(new_new_n221_), .Y(new_new_n224_));
  INV        g0202(.A(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(i_12_), .B(new_new_n225_), .Y(new_new_n226_));
  NA3        g0204(.A(new_new_n226_), .B(new_new_n196_), .C(new_new_n194_), .Y(new_new_n227_));
  OAI210     g0205(.A0(new_new_n224_), .A1(new_new_n220_), .B0(new_new_n227_), .Y(new_new_n228_));
  AOI220     g0206(.A0(new_new_n228_), .A1(new_new_n137_), .B0(new_new_n219_), .B1(new_new_n216_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n37_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n180_), .B(i_4_), .Y(new_new_n231_));
  OR2        g0209(.A(i_8_), .B(i_7_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n232_), .B(new_new_n84_), .Y(new_new_n233_));
  NO2        g0211(.A(new_new_n52_), .B(i_1_), .Y(new_new_n234_));
  NA2        g0212(.A(new_new_n234_), .B(new_new_n233_), .Y(new_new_n235_));
  INV        g0213(.A(i_12_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n44_), .B(new_new_n236_), .Y(new_new_n237_));
  NO3        g0215(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n238_));
  NA2        g0216(.A(i_2_), .B(i_1_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n235_), .B(new_new_n180_), .Y(new_new_n240_));
  NO3        g0218(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n241_));
  NAi21      g0219(.An(i_4_), .B(i_3_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n242_), .B(new_new_n73_), .Y(new_new_n243_));
  NO2        g0221(.A(i_0_), .B(i_6_), .Y(new_new_n244_));
  NOi41      g0222(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n245_));
  NA2        g0223(.A(new_new_n245_), .B(new_new_n244_), .Y(new_new_n246_));
  NO2        g0224(.A(new_new_n239_), .B(new_new_n180_), .Y(new_new_n247_));
  NAi21      g0225(.An(new_new_n246_), .B(new_new_n247_), .Y(new_new_n248_));
  INV        g0226(.A(new_new_n248_), .Y(new_new_n249_));
  AOI220     g0227(.A0(new_new_n249_), .A1(new_new_n39_), .B0(new_new_n240_), .B1(new_new_n205_), .Y(new_new_n250_));
  NO2        g0228(.A(i_11_), .B(new_new_n225_), .Y(new_new_n251_));
  NOi21      g0229(.An(i_1_), .B(i_6_), .Y(new_new_n252_));
  NAi21      g0230(.An(i_3_), .B(i_7_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n236_), .B(i_9_), .Y(new_new_n254_));
  OR4        g0232(.A(new_new_n254_), .B(new_new_n253_), .C(new_new_n252_), .D(new_new_n183_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n256_));
  NO2        g0234(.A(i_12_), .B(i_3_), .Y(new_new_n257_));
  NA2        g0235(.A(new_new_n71_), .B(i_5_), .Y(new_new_n258_));
  NA2        g0236(.A(i_3_), .B(i_9_), .Y(new_new_n259_));
  NAi21      g0237(.An(i_7_), .B(i_10_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  NA3        g0239(.A(new_new_n261_), .B(new_new_n258_), .C(new_new_n63_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n262_), .B(new_new_n255_), .Y(new_new_n263_));
  NA3        g0241(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n264_));
  INV        g0242(.A(new_new_n138_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n236_), .B(i_13_), .Y(new_new_n266_));
  NO2        g0244(.A(new_new_n266_), .B(new_new_n73_), .Y(new_new_n267_));
  AOI220     g0245(.A0(new_new_n267_), .A1(new_new_n265_), .B0(new_new_n263_), .B1(new_new_n251_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n232_), .B(new_new_n37_), .Y(new_new_n269_));
  NA2        g0247(.A(i_12_), .B(i_6_), .Y(new_new_n270_));
  OR2        g0248(.A(i_13_), .B(i_9_), .Y(new_new_n271_));
  NO3        g0249(.A(new_new_n271_), .B(new_new_n270_), .C(new_new_n48_), .Y(new_new_n272_));
  NO2        g0250(.A(new_new_n242_), .B(i_2_), .Y(new_new_n273_));
  NA3        g0251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n44_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n251_), .B(i_9_), .Y(new_new_n275_));
  OAI210     g0253(.A0(new_new_n71_), .A1(new_new_n275_), .B0(new_new_n274_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n150_), .B(new_new_n62_), .Y(new_new_n277_));
  NO3        g0255(.A(i_11_), .B(new_new_n225_), .C(new_new_n25_), .Y(new_new_n278_));
  NO2        g0256(.A(i_6_), .B(new_new_n48_), .Y(new_new_n279_));
  NA3        g0257(.A(new_new_n279_), .B(i_7_), .C(new_new_n278_), .Y(new_new_n280_));
  NO3        g0258(.A(new_new_n26_), .B(new_new_n84_), .C(i_5_), .Y(new_new_n281_));
  NA3        g0259(.A(new_new_n281_), .B(new_new_n269_), .C(new_new_n226_), .Y(new_new_n282_));
  AOI210     g0260(.A0(new_new_n282_), .A1(new_new_n280_), .B0(new_new_n277_), .Y(new_new_n283_));
  AOI210     g0261(.A0(new_new_n276_), .A1(new_new_n269_), .B0(new_new_n283_), .Y(new_new_n284_));
  NA4        g0262(.A(new_new_n284_), .B(new_new_n268_), .C(new_new_n250_), .D(new_new_n229_), .Y(new_new_n285_));
  NO3        g0263(.A(i_12_), .B(new_new_n225_), .C(new_new_n37_), .Y(new_new_n286_));
  INV        g0264(.A(new_new_n286_), .Y(new_new_n287_));
  NOi21      g0265(.An(new_new_n159_), .B(new_new_n84_), .Y(new_new_n288_));
  NO3        g0266(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n289_));
  AOI220     g0267(.A0(new_new_n289_), .A1(new_new_n194_), .B0(new_new_n288_), .B1(new_new_n234_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n290_), .B(i_7_), .Y(new_new_n291_));
  NO3        g0269(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n239_), .B(i_0_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n192_), .B0(new_new_n292_), .B1(new_new_n137_), .Y(new_new_n294_));
  NA2        g0272(.A(new_new_n279_), .B(new_new_n26_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(new_new_n294_), .Y(new_new_n296_));
  NA2        g0274(.A(i_0_), .B(i_1_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(i_2_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n58_), .B(i_6_), .Y(new_new_n299_));
  NA3        g0277(.A(new_new_n299_), .B(new_new_n298_), .C(new_new_n159_), .Y(new_new_n300_));
  OAI210     g0278(.A0(new_new_n161_), .A1(new_new_n138_), .B0(new_new_n300_), .Y(new_new_n301_));
  NO3        g0279(.A(new_new_n301_), .B(new_new_n296_), .C(new_new_n291_), .Y(new_new_n302_));
  NO2        g0280(.A(i_3_), .B(i_10_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n304_));
  NO2        g0282(.A(i_4_), .B(i_8_), .Y(new_new_n305_));
  NOi21      g0283(.An(new_new_n217_), .B(new_new_n99_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(new_new_n305_), .C(i_7_), .Y(new_new_n307_));
  AN2        g0285(.A(i_3_), .B(i_10_), .Y(new_new_n308_));
  NA4        g0286(.A(new_new_n308_), .B(new_new_n196_), .C(new_new_n173_), .D(new_new_n171_), .Y(new_new_n309_));
  NO2        g0287(.A(i_5_), .B(new_new_n37_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n311_));
  OR2        g0289(.A(new_new_n307_), .B(new_new_n304_), .Y(new_new_n312_));
  OAI220     g0290(.A0(new_new_n312_), .A1(i_6_), .B0(new_new_n302_), .B1(new_new_n287_), .Y(new_new_n313_));
  NO4        g0291(.A(new_new_n313_), .B(new_new_n285_), .C(new_new_n213_), .D(new_new_n164_), .Y(new_new_n314_));
  NO3        g0292(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n315_));
  NO3        g0293(.A(i_6_), .B(new_new_n191_), .C(i_7_), .Y(new_new_n316_));
  AOI210     g0294(.A0(new_new_n1104_), .A1(new_new_n239_), .B0(new_new_n166_), .Y(new_new_n317_));
  NO2        g0295(.A(i_2_), .B(i_3_), .Y(new_new_n318_));
  OR2        g0296(.A(i_0_), .B(i_5_), .Y(new_new_n319_));
  NA2        g0297(.A(new_new_n217_), .B(new_new_n319_), .Y(new_new_n320_));
  NA4        g0298(.A(new_new_n320_), .B(new_new_n233_), .C(new_new_n318_), .D(i_1_), .Y(new_new_n321_));
  NA3        g0299(.A(new_new_n293_), .B(new_new_n288_), .C(new_new_n108_), .Y(new_new_n322_));
  NAi21      g0300(.An(i_8_), .B(i_7_), .Y(new_new_n323_));
  NO2        g0301(.A(new_new_n323_), .B(i_6_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n153_), .B(new_new_n46_), .Y(new_new_n325_));
  NA3        g0303(.A(new_new_n325_), .B(new_new_n324_), .C(new_new_n159_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n322_), .C(new_new_n321_), .Y(new_new_n327_));
  OAI210     g0305(.A0(new_new_n327_), .A1(new_new_n317_), .B0(i_4_), .Y(new_new_n328_));
  NO2        g0306(.A(i_12_), .B(i_10_), .Y(new_new_n329_));
  NOi21      g0307(.An(i_5_), .B(i_0_), .Y(new_new_n330_));
  AOI210     g0308(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n98_), .Y(new_new_n331_));
  NO4        g0309(.A(new_new_n331_), .B(i_4_), .C(new_new_n330_), .D(new_new_n123_), .Y(new_new_n332_));
  NA4        g0310(.A(new_new_n82_), .B(new_new_n36_), .C(new_new_n84_), .D(i_8_), .Y(new_new_n333_));
  NA2        g0311(.A(new_new_n332_), .B(new_new_n329_), .Y(new_new_n334_));
  NO2        g0312(.A(i_6_), .B(i_8_), .Y(new_new_n335_));
  NOi21      g0313(.An(i_0_), .B(i_2_), .Y(new_new_n336_));
  AN2        g0314(.A(new_new_n336_), .B(new_new_n335_), .Y(new_new_n337_));
  NO2        g0315(.A(i_1_), .B(i_7_), .Y(new_new_n338_));
  AO220      g0316(.A0(new_new_n338_), .A1(new_new_n337_), .B0(new_new_n324_), .B1(new_new_n234_), .Y(new_new_n339_));
  NA3        g0317(.A(new_new_n339_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n340_), .B(new_new_n334_), .C(new_new_n328_), .Y(new_new_n341_));
  AOI210     g0319(.A0(i_8_), .A1(i_8_), .B0(new_new_n320_), .Y(new_new_n342_));
  NOi21      g0320(.An(new_new_n149_), .B(new_new_n100_), .Y(new_new_n343_));
  NO2        g0321(.A(new_new_n343_), .B(new_new_n119_), .Y(new_new_n344_));
  OAI210     g0322(.A0(new_new_n344_), .A1(new_new_n342_), .B0(i_3_), .Y(new_new_n345_));
  INV        g0323(.A(new_new_n82_), .Y(new_new_n346_));
  NO2        g0324(.A(new_new_n297_), .B(new_new_n79_), .Y(new_new_n347_));
  NA2        g0325(.A(new_new_n347_), .B(new_new_n127_), .Y(new_new_n348_));
  NO2        g0326(.A(new_new_n92_), .B(new_new_n191_), .Y(new_new_n349_));
  NA3        g0327(.A(new_new_n306_), .B(new_new_n349_), .C(new_new_n62_), .Y(new_new_n350_));
  AOI210     g0328(.A0(new_new_n350_), .A1(new_new_n348_), .B0(new_new_n346_), .Y(new_new_n351_));
  NO2        g0329(.A(new_new_n191_), .B(i_9_), .Y(new_new_n352_));
  NA3        g0330(.A(new_new_n352_), .B(new_new_n204_), .C(new_new_n153_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n353_), .B(new_new_n46_), .Y(new_new_n354_));
  NO3        g0332(.A(new_new_n354_), .B(new_new_n351_), .C(new_new_n296_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n355_), .A1(new_new_n345_), .B0(new_new_n158_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n341_), .A1(new_new_n315_), .B0(new_new_n356_), .Y(new_new_n357_));
  NOi32      g0335(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n358_));
  INV        g0336(.A(new_new_n358_), .Y(new_new_n359_));
  NAi21      g0337(.An(i_0_), .B(i_6_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_1_), .B(i_5_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n360_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n25_), .Y(new_new_n363_));
  OAI210     g0341(.A0(new_new_n363_), .A1(new_new_n155_), .B0(new_new_n246_), .Y(new_new_n364_));
  NAi41      g0342(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n365_));
  OAI220     g0343(.A0(new_new_n365_), .A1(new_new_n361_), .B0(new_new_n220_), .B1(new_new_n155_), .Y(new_new_n366_));
  AOI210     g0344(.A0(new_new_n365_), .A1(new_new_n155_), .B0(new_new_n153_), .Y(new_new_n367_));
  NOi32      g0345(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n368_));
  NAi21      g0346(.An(i_6_), .B(i_1_), .Y(new_new_n369_));
  NA3        g0347(.A(new_new_n369_), .B(new_new_n368_), .C(new_new_n46_), .Y(new_new_n370_));
  NO2        g0348(.A(new_new_n370_), .B(i_0_), .Y(new_new_n371_));
  OR3        g0349(.A(new_new_n371_), .B(new_new_n367_), .C(new_new_n366_), .Y(new_new_n372_));
  NO2        g0350(.A(i_1_), .B(new_new_n98_), .Y(new_new_n373_));
  NAi21      g0351(.An(i_3_), .B(i_4_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n374_), .B(i_9_), .Y(new_new_n375_));
  AN2        g0353(.A(i_6_), .B(i_7_), .Y(new_new_n376_));
  OAI210     g0354(.A0(new_new_n376_), .A1(new_new_n373_), .B0(new_new_n375_), .Y(new_new_n377_));
  NA2        g0355(.A(i_2_), .B(i_7_), .Y(new_new_n378_));
  NO2        g0356(.A(new_new_n374_), .B(i_10_), .Y(new_new_n379_));
  NA3        g0357(.A(new_new_n379_), .B(new_new_n378_), .C(new_new_n244_), .Y(new_new_n380_));
  AOI210     g0358(.A0(new_new_n380_), .A1(new_new_n377_), .B0(new_new_n183_), .Y(new_new_n381_));
  AOI210     g0359(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n382_));
  OAI210     g0360(.A0(new_new_n382_), .A1(new_new_n186_), .B0(new_new_n379_), .Y(new_new_n383_));
  AOI220     g0361(.A0(new_new_n379_), .A1(new_new_n338_), .B0(new_new_n238_), .B1(new_new_n186_), .Y(new_new_n384_));
  AOI210     g0362(.A0(new_new_n384_), .A1(new_new_n383_), .B0(i_5_), .Y(new_new_n385_));
  NO4        g0363(.A(new_new_n385_), .B(new_new_n381_), .C(new_new_n372_), .D(new_new_n364_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n386_), .B(new_new_n359_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n388_));
  AN2        g0366(.A(i_12_), .B(i_5_), .Y(new_new_n389_));
  NO2        g0367(.A(i_4_), .B(new_new_n26_), .Y(new_new_n390_));
  NA2        g0368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  NO2        g0369(.A(i_11_), .B(i_6_), .Y(new_new_n392_));
  NA3        g0370(.A(new_new_n392_), .B(new_new_n325_), .C(new_new_n225_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n393_), .B(new_new_n391_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n242_), .B(i_5_), .Y(new_new_n395_));
  NO2        g0373(.A(i_5_), .B(i_10_), .Y(new_new_n396_));
  AOI220     g0374(.A0(new_new_n396_), .A1(new_new_n273_), .B0(new_new_n395_), .B1(new_new_n196_), .Y(new_new_n397_));
  NO2        g0375(.A(i_6_), .B(new_new_n397_), .Y(new_new_n398_));
  OAI210     g0376(.A0(new_new_n398_), .A1(new_new_n394_), .B0(new_new_n388_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n145_), .B(new_new_n84_), .Y(new_new_n401_));
  OAI210     g0379(.A0(new_new_n401_), .A1(new_new_n394_), .B0(new_new_n400_), .Y(new_new_n402_));
  NO3        g0380(.A(new_new_n84_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n403_));
  NO2        g0381(.A(i_3_), .B(new_new_n98_), .Y(new_new_n404_));
  NA4        g0382(.A(new_new_n303_), .B(new_new_n90_), .C(new_new_n73_), .D(new_new_n53_), .Y(new_new_n405_));
  NO2        g0383(.A(i_11_), .B(i_12_), .Y(new_new_n406_));
  NA2        g0384(.A(new_new_n406_), .B(new_new_n36_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n405_), .B(new_new_n407_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n396_), .B(new_new_n236_), .Y(new_new_n409_));
  NA3        g0387(.A(new_new_n108_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n410_));
  OAI220     g0388(.A0(new_new_n410_), .A1(new_new_n220_), .B0(new_new_n409_), .B1(new_new_n333_), .Y(new_new_n411_));
  NAi21      g0389(.An(i_13_), .B(i_0_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n412_), .B(new_new_n239_), .Y(new_new_n413_));
  OAI210     g0391(.A0(new_new_n411_), .A1(new_new_n408_), .B0(new_new_n413_), .Y(new_new_n414_));
  NA3        g0392(.A(new_new_n414_), .B(new_new_n402_), .C(new_new_n399_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n44_), .B(new_new_n225_), .Y(new_new_n416_));
  NO3        g0394(.A(i_1_), .B(i_12_), .C(new_new_n84_), .Y(new_new_n417_));
  NO2        g0395(.A(i_0_), .B(i_11_), .Y(new_new_n418_));
  AN2        g0396(.A(i_1_), .B(i_6_), .Y(new_new_n419_));
  NOi21      g0397(.An(i_2_), .B(i_12_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n420_), .B(new_new_n419_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n421_), .B(new_new_n1095_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n137_), .B(i_9_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n423_), .B(i_4_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n422_), .B(new_new_n424_), .Y(new_new_n425_));
  NAi21      g0403(.An(i_9_), .B(i_4_), .Y(new_new_n426_));
  OR2        g0404(.A(i_13_), .B(i_10_), .Y(new_new_n427_));
  NO3        g0405(.A(new_new_n427_), .B(new_new_n112_), .C(new_new_n426_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n169_), .B(new_new_n118_), .Y(new_new_n429_));
  OR2        g0407(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n98_), .B(new_new_n25_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n286_), .B(new_new_n431_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n279_), .B(i_1_), .Y(new_new_n433_));
  OAI220     g0411(.A0(new_new_n433_), .A1(new_new_n430_), .B0(new_new_n432_), .B1(new_new_n343_), .Y(new_new_n434_));
  INV        g0412(.A(new_new_n434_), .Y(new_new_n435_));
  AOI210     g0413(.A0(new_new_n435_), .A1(new_new_n425_), .B0(new_new_n26_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n322_), .B(new_new_n321_), .Y(new_new_n437_));
  AOI220     g0415(.A0(new_new_n299_), .A1(new_new_n289_), .B0(new_new_n293_), .B1(i_6_), .Y(new_new_n438_));
  NO2        g0416(.A(new_new_n438_), .B(new_new_n166_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n180_), .B(new_new_n84_), .Y(new_new_n440_));
  AOI220     g0418(.A0(new_new_n440_), .A1(new_new_n298_), .B0(new_new_n281_), .B1(i_1_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n441_), .B(i_7_), .Y(new_new_n442_));
  NO3        g0420(.A(new_new_n442_), .B(new_new_n439_), .C(new_new_n437_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n194_), .B(new_new_n94_), .Y(new_new_n444_));
  NA3        g0422(.A(new_new_n325_), .B(new_new_n159_), .C(new_new_n84_), .Y(new_new_n445_));
  AOI210     g0423(.A0(new_new_n445_), .A1(new_new_n444_), .B0(new_new_n323_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n191_), .B(i_10_), .Y(new_new_n447_));
  NA3        g0425(.A(new_new_n258_), .B(new_new_n63_), .C(i_2_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n299_), .B(new_new_n234_), .Y(new_new_n449_));
  OAI220     g0427(.A0(new_new_n449_), .A1(new_new_n180_), .B0(new_new_n448_), .B1(new_new_n447_), .Y(new_new_n450_));
  NO2        g0428(.A(i_3_), .B(new_new_n48_), .Y(new_new_n451_));
  NA3        g0429(.A(new_new_n338_), .B(new_new_n337_), .C(new_new_n451_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n316_), .B(new_new_n320_), .Y(new_new_n453_));
  OAI210     g0431(.A0(new_new_n453_), .A1(new_new_n187_), .B0(new_new_n452_), .Y(new_new_n454_));
  NO3        g0432(.A(new_new_n454_), .B(new_new_n450_), .C(new_new_n446_), .Y(new_new_n455_));
  AOI210     g0433(.A0(new_new_n455_), .A1(new_new_n443_), .B0(new_new_n275_), .Y(new_new_n456_));
  NO4        g0434(.A(new_new_n456_), .B(new_new_n436_), .C(new_new_n415_), .D(new_new_n387_), .Y(new_new_n457_));
  NO2        g0435(.A(new_new_n71_), .B(i_13_), .Y(new_new_n458_));
  NO2        g0436(.A(i_10_), .B(i_9_), .Y(new_new_n459_));
  NAi21      g0437(.An(i_12_), .B(i_8_), .Y(new_new_n460_));
  NO2        g0438(.A(new_new_n460_), .B(i_3_), .Y(new_new_n461_));
  NO2        g0439(.A(new_new_n46_), .B(i_4_), .Y(new_new_n462_));
  NA2        g0440(.A(new_new_n462_), .B(new_new_n100_), .Y(new_new_n463_));
  NO2        g0441(.A(new_new_n463_), .B(new_new_n203_), .Y(new_new_n464_));
  NA2        g0442(.A(new_new_n311_), .B(i_0_), .Y(new_new_n465_));
  NO3        g0443(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n270_), .B(new_new_n95_), .Y(new_new_n467_));
  NA2        g0445(.A(new_new_n467_), .B(new_new_n466_), .Y(new_new_n468_));
  NA2        g0446(.A(i_8_), .B(i_9_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n286_), .B(new_new_n204_), .Y(new_new_n470_));
  OAI220     g0448(.A0(new_new_n470_), .A1(new_new_n469_), .B0(new_new_n468_), .B1(new_new_n465_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n251_), .B(new_new_n310_), .Y(new_new_n472_));
  NO3        g0450(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n473_));
  AOI210     g0451(.A0(new_new_n257_), .A1(new_new_n186_), .B0(new_new_n473_), .Y(new_new_n474_));
  NA3        g0452(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n475_));
  NA4        g0453(.A(new_new_n140_), .B(new_new_n110_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n476_));
  OAI220     g0454(.A0(new_new_n476_), .A1(new_new_n475_), .B0(new_new_n474_), .B1(new_new_n472_), .Y(new_new_n477_));
  NO3        g0455(.A(new_new_n477_), .B(new_new_n471_), .C(new_new_n464_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n298_), .B(new_new_n103_), .Y(new_new_n479_));
  OR2        g0457(.A(new_new_n479_), .B(new_new_n206_), .Y(new_new_n480_));
  OA210      g0458(.A0(new_new_n353_), .A1(new_new_n98_), .B0(new_new_n300_), .Y(new_new_n481_));
  OA220      g0459(.A0(new_new_n481_), .A1(new_new_n158_), .B0(new_new_n480_), .B1(new_new_n180_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n94_), .B(i_13_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n440_), .B(new_new_n388_), .Y(new_new_n484_));
  NO2        g0462(.A(i_2_), .B(i_13_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n484_), .B(new_new_n483_), .Y(new_new_n486_));
  NO3        g0464(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n487_));
  NO2        g0465(.A(i_6_), .B(i_7_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n488_), .B(new_new_n487_), .Y(new_new_n489_));
  OR2        g0467(.A(i_11_), .B(i_8_), .Y(new_new_n490_));
  NOi21      g0468(.An(i_2_), .B(i_7_), .Y(new_new_n491_));
  NAi31      g0469(.An(new_new_n490_), .B(new_new_n491_), .C(new_new_n1097_), .Y(new_new_n492_));
  NO2        g0470(.A(new_new_n427_), .B(i_6_), .Y(new_new_n493_));
  NA3        g0471(.A(new_new_n493_), .B(new_new_n1100_), .C(new_new_n73_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n494_), .B(new_new_n492_), .Y(new_new_n495_));
  NO2        g0473(.A(i_3_), .B(new_new_n191_), .Y(new_new_n496_));
  NO2        g0474(.A(i_6_), .B(i_10_), .Y(new_new_n497_));
  NA4        g0475(.A(new_new_n497_), .B(new_new_n315_), .C(new_new_n496_), .D(new_new_n236_), .Y(new_new_n498_));
  NO2        g0476(.A(new_new_n498_), .B(new_new_n151_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n245_), .B(new_new_n168_), .C(new_new_n127_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n501_));
  NO2        g0479(.A(new_new_n153_), .B(i_3_), .Y(new_new_n502_));
  NAi31      g0480(.An(new_new_n501_), .B(new_new_n502_), .C(new_new_n226_), .Y(new_new_n503_));
  NA3        g0481(.A(new_new_n400_), .B(new_new_n176_), .C(new_new_n144_), .Y(new_new_n504_));
  NA3        g0482(.A(new_new_n504_), .B(new_new_n503_), .C(new_new_n500_), .Y(new_new_n505_));
  NO4        g0483(.A(new_new_n505_), .B(new_new_n499_), .C(new_new_n495_), .D(new_new_n486_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n473_), .B(new_new_n396_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n507_), .B(new_new_n224_), .Y(new_new_n508_));
  NAi21      g0486(.An(new_new_n215_), .B(new_new_n406_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n26_), .B(i_5_), .Y(new_new_n510_));
  NO2        g0488(.A(i_0_), .B(new_new_n84_), .Y(new_new_n511_));
  NA3        g0489(.A(new_new_n511_), .B(new_new_n510_), .C(new_new_n137_), .Y(new_new_n512_));
  OAI220     g0490(.A0(new_new_n38_), .A1(new_new_n512_), .B0(i_0_), .B1(new_new_n509_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n27_), .B(i_10_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n315_), .B(new_new_n238_), .Y(new_new_n515_));
  OAI220     g0493(.A0(new_new_n515_), .A1(new_new_n448_), .B0(new_new_n514_), .B1(new_new_n483_), .Y(new_new_n516_));
  NA4        g0494(.A(new_new_n308_), .B(new_new_n223_), .C(new_new_n71_), .D(new_new_n236_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n517_), .B(new_new_n489_), .Y(new_new_n518_));
  NO4        g0496(.A(new_new_n518_), .B(new_new_n516_), .C(new_new_n513_), .D(new_new_n508_), .Y(new_new_n519_));
  NA4        g0497(.A(new_new_n519_), .B(new_new_n506_), .C(new_new_n482_), .D(new_new_n478_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n308_), .B(new_new_n173_), .C(new_new_n171_), .Y(new_new_n521_));
  OAI210     g0499(.A0(new_new_n304_), .A1(new_new_n178_), .B0(new_new_n521_), .Y(new_new_n522_));
  AN2        g0500(.A(new_new_n289_), .B(new_new_n233_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n523_), .B(new_new_n522_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n117_), .B(new_new_n107_), .Y(new_new_n525_));
  AO220      g0503(.A0(new_new_n525_), .A1(new_new_n466_), .B0(new_new_n428_), .B1(i_6_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n315_), .B(new_new_n160_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n527_), .A1(new_new_n180_), .B0(new_new_n309_), .Y(new_new_n528_));
  AOI220     g0506(.A0(new_new_n528_), .A1(new_new_n324_), .B0(new_new_n526_), .B1(new_new_n311_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n389_), .B(new_new_n225_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n358_), .B(new_new_n71_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n376_), .B(new_new_n368_), .Y(new_new_n532_));
  AO210      g0510(.A0(new_new_n531_), .A1(new_new_n530_), .B0(new_new_n532_), .Y(new_new_n533_));
  NO2        g0511(.A(new_new_n36_), .B(i_8_), .Y(new_new_n534_));
  NAi41      g0512(.An(new_new_n531_), .B(new_new_n497_), .C(new_new_n534_), .D(new_new_n46_), .Y(new_new_n535_));
  INV        g0513(.A(new_new_n428_), .Y(new_new_n536_));
  NA3        g0514(.A(new_new_n536_), .B(new_new_n535_), .C(new_new_n533_), .Y(new_new_n537_));
  INV        g0515(.A(new_new_n537_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n258_), .B(new_new_n63_), .Y(new_new_n539_));
  OAI210     g0517(.A0(i_8_), .A1(new_new_n539_), .B0(new_new_n129_), .Y(new_new_n540_));
  AOI210     g0518(.A0(new_new_n192_), .A1(i_9_), .B0(new_new_n269_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n541_), .B(new_new_n197_), .Y(new_new_n542_));
  AOI220     g0520(.A0(i_6_), .A1(new_new_n542_), .B0(new_new_n540_), .B1(new_new_n429_), .Y(new_new_n543_));
  NA4        g0521(.A(new_new_n543_), .B(new_new_n538_), .C(new_new_n529_), .D(new_new_n524_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n395_), .B(new_new_n298_), .Y(new_new_n545_));
  OAI210     g0523(.A0(new_new_n391_), .A1(new_new_n165_), .B0(new_new_n545_), .Y(new_new_n546_));
  NO2        g0524(.A(i_12_), .B(new_new_n191_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n547_), .B(new_new_n225_), .Y(new_new_n548_));
  NA3        g0526(.A(new_new_n497_), .B(new_new_n171_), .C(new_new_n27_), .Y(new_new_n549_));
  NO3        g0527(.A(new_new_n549_), .B(new_new_n548_), .C(new_new_n479_), .Y(new_new_n550_));
  NOi31      g0528(.An(new_new_n316_), .B(new_new_n427_), .C(new_new_n38_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n551_), .A1(new_new_n550_), .B0(new_new_n546_), .Y(new_new_n552_));
  NO2        g0530(.A(i_8_), .B(i_7_), .Y(new_new_n553_));
  OAI210     g0531(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n223_), .Y(new_new_n555_));
  AOI220     g0533(.A0(new_new_n325_), .A1(new_new_n39_), .B0(new_new_n234_), .B1(new_new_n205_), .Y(new_new_n556_));
  OAI220     g0534(.A0(new_new_n556_), .A1(new_new_n180_), .B0(new_new_n555_), .B1(new_new_n242_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n44_), .B(i_10_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n558_), .B(i_6_), .Y(new_new_n559_));
  NA3        g0537(.A(new_new_n559_), .B(new_new_n557_), .C(new_new_n553_), .Y(new_new_n560_));
  AOI220     g0538(.A0(new_new_n440_), .A1(new_new_n325_), .B0(new_new_n247_), .B1(new_new_n244_), .Y(new_new_n561_));
  OAI220     g0539(.A0(new_new_n561_), .A1(new_new_n266_), .B0(new_new_n483_), .B1(new_new_n128_), .Y(new_new_n562_));
  NA2        g0540(.A(new_new_n562_), .B(new_new_n269_), .Y(new_new_n563_));
  NOi31      g0541(.An(new_new_n293_), .B(new_new_n304_), .C(new_new_n178_), .Y(new_new_n564_));
  NA3        g0542(.A(new_new_n308_), .B(new_new_n171_), .C(new_new_n94_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n221_), .B(new_new_n44_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n153_), .B(i_5_), .Y(new_new_n567_));
  NA3        g0545(.A(new_new_n567_), .B(new_new_n416_), .C(new_new_n318_), .Y(new_new_n568_));
  OAI210     g0546(.A0(new_new_n568_), .A1(new_new_n566_), .B0(new_new_n565_), .Y(new_new_n569_));
  OAI210     g0547(.A0(new_new_n569_), .A1(new_new_n564_), .B0(new_new_n473_), .Y(new_new_n570_));
  NA4        g0548(.A(new_new_n570_), .B(new_new_n563_), .C(new_new_n560_), .D(new_new_n552_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n286_), .B(new_new_n82_), .Y(new_new_n572_));
  AOI210     g0550(.A0(i_11_), .A1(new_new_n348_), .B0(new_new_n572_), .Y(new_new_n573_));
  NA2        g0551(.A(new_new_n299_), .B(new_new_n289_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n574_), .B(new_new_n170_), .Y(new_new_n575_));
  NA2        g0553(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n459_), .B(new_new_n221_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n576_), .B(new_new_n577_), .Y(new_new_n578_));
  NA2        g0556(.A(i_0_), .B(new_new_n48_), .Y(new_new_n579_));
  NA3        g0557(.A(new_new_n547_), .B(new_new_n278_), .C(new_new_n579_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n1101_), .B(new_new_n580_), .Y(new_new_n581_));
  NO4        g0559(.A(new_new_n581_), .B(new_new_n578_), .C(new_new_n575_), .D(new_new_n573_), .Y(new_new_n582_));
  NO4        g0560(.A(new_new_n252_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n583_));
  NO3        g0561(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n232_), .B(new_new_n36_), .Y(new_new_n585_));
  AN2        g0563(.A(new_new_n585_), .B(new_new_n584_), .Y(new_new_n586_));
  OA210      g0564(.A0(new_new_n586_), .A1(new_new_n583_), .B0(new_new_n358_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n427_), .B(i_1_), .Y(new_new_n588_));
  NOi31      g0566(.An(new_new_n588_), .B(new_new_n467_), .C(new_new_n71_), .Y(new_new_n589_));
  AN4        g0567(.A(new_new_n589_), .B(new_new_n424_), .C(new_new_n510_), .D(i_2_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n438_), .B(new_new_n174_), .Y(new_new_n591_));
  NO3        g0569(.A(new_new_n591_), .B(new_new_n590_), .C(new_new_n587_), .Y(new_new_n592_));
  NOi21      g0570(.An(i_10_), .B(i_6_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n84_), .B(new_new_n25_), .Y(new_new_n594_));
  AOI220     g0572(.A0(new_new_n286_), .A1(new_new_n594_), .B0(new_new_n278_), .B1(new_new_n593_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n595_), .B(new_new_n465_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n597_));
  NA2        g0575(.A(new_new_n316_), .B(new_new_n160_), .Y(new_new_n598_));
  AOI220     g0576(.A0(new_new_n598_), .A1(new_new_n449_), .B0(new_new_n181_), .B1(new_new_n179_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n196_), .B(new_new_n37_), .Y(new_new_n600_));
  NOi31      g0578(.An(new_new_n141_), .B(new_new_n600_), .C(new_new_n333_), .Y(new_new_n601_));
  NO3        g0579(.A(new_new_n601_), .B(new_new_n599_), .C(new_new_n596_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n531_), .B(new_new_n384_), .Y(new_new_n603_));
  INV        g0581(.A(new_new_n318_), .Y(new_new_n604_));
  NO2        g0582(.A(i_12_), .B(new_new_n84_), .Y(new_new_n605_));
  NA3        g0583(.A(new_new_n605_), .B(new_new_n278_), .C(new_new_n579_), .Y(new_new_n606_));
  NA3        g0584(.A(new_new_n392_), .B(new_new_n286_), .C(new_new_n217_), .Y(new_new_n607_));
  AOI210     g0585(.A0(new_new_n607_), .A1(new_new_n606_), .B0(new_new_n604_), .Y(new_new_n608_));
  NA2        g0586(.A(new_new_n171_), .B(i_0_), .Y(new_new_n609_));
  NO3        g0587(.A(new_new_n609_), .B(i_8_), .C(new_new_n304_), .Y(new_new_n610_));
  OR2        g0588(.A(i_2_), .B(i_5_), .Y(new_new_n611_));
  OR2        g0589(.A(new_new_n611_), .B(new_new_n419_), .Y(new_new_n612_));
  AOI210     g0590(.A0(i_0_), .A1(new_new_n612_), .B0(new_new_n509_), .Y(new_new_n613_));
  NO4        g0591(.A(new_new_n613_), .B(new_new_n610_), .C(new_new_n608_), .D(new_new_n603_), .Y(new_new_n614_));
  NA4        g0592(.A(new_new_n614_), .B(new_new_n602_), .C(new_new_n592_), .D(new_new_n582_), .Y(new_new_n615_));
  NO4        g0593(.A(new_new_n615_), .B(new_new_n571_), .C(new_new_n544_), .D(new_new_n520_), .Y(new_new_n616_));
  NA4        g0594(.A(new_new_n616_), .B(new_new_n457_), .C(new_new_n357_), .D(new_new_n314_), .Y(men7));
  NO2        g0595(.A(new_new_n103_), .B(new_new_n89_), .Y(new_new_n618_));
  NA2        g0596(.A(new_new_n390_), .B(new_new_n618_), .Y(new_new_n619_));
  NA2        g0597(.A(new_new_n497_), .B(new_new_n82_), .Y(new_new_n620_));
  NA2        g0598(.A(i_11_), .B(new_new_n191_), .Y(new_new_n621_));
  OAI210     g0599(.A0(new_new_n1102_), .A1(new_new_n620_), .B0(new_new_n619_), .Y(new_new_n622_));
  NA3        g0600(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n236_), .B(i_4_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n624_), .B(i_8_), .Y(new_new_n625_));
  AOI210     g0603(.A0(new_new_n625_), .A1(new_new_n101_), .B0(new_new_n623_), .Y(new_new_n626_));
  NA2        g0604(.A(i_2_), .B(new_new_n84_), .Y(new_new_n627_));
  OAI210     g0605(.A0(new_new_n87_), .A1(new_new_n201_), .B0(new_new_n202_), .Y(new_new_n628_));
  NO2        g0606(.A(i_7_), .B(new_new_n37_), .Y(new_new_n629_));
  NA2        g0607(.A(i_4_), .B(i_8_), .Y(new_new_n630_));
  AOI210     g0608(.A0(new_new_n630_), .A1(new_new_n308_), .B0(new_new_n629_), .Y(new_new_n631_));
  OAI220     g0609(.A0(new_new_n631_), .A1(new_new_n627_), .B0(new_new_n628_), .B1(i_13_), .Y(new_new_n632_));
  NO3        g0610(.A(new_new_n632_), .B(new_new_n626_), .C(new_new_n622_), .Y(new_new_n633_));
  AOI210     g0611(.A0(new_new_n123_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n634_));
  AOI210     g0612(.A0(new_new_n634_), .A1(new_new_n236_), .B0(new_new_n157_), .Y(new_new_n635_));
  OR2        g0613(.A(i_6_), .B(i_10_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n636_), .B(new_new_n23_), .Y(new_new_n637_));
  OR3        g0615(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n638_));
  NO3        g0616(.A(new_new_n638_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n639_));
  INV        g0617(.A(new_new_n198_), .Y(new_new_n640_));
  NO2        g0618(.A(new_new_n639_), .B(new_new_n637_), .Y(new_new_n641_));
  OA220      g0619(.A0(new_new_n641_), .A1(new_new_n604_), .B0(new_new_n635_), .B1(new_new_n271_), .Y(new_new_n642_));
  AOI210     g0620(.A0(new_new_n642_), .A1(new_new_n633_), .B0(new_new_n62_), .Y(new_new_n643_));
  NOi21      g0621(.An(i_11_), .B(i_7_), .Y(new_new_n644_));
  AO210      g0622(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n645_), .B(new_new_n644_), .Y(new_new_n646_));
  NA3        g0624(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n647_));
  NAi31      g0625(.An(new_new_n647_), .B(new_new_n214_), .C(i_11_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n648_), .B(new_new_n62_), .Y(new_new_n649_));
  AO210      g0627(.A0(new_new_n85_), .A1(new_new_n384_), .B0(new_new_n40_), .Y(new_new_n650_));
  NO3        g0628(.A(new_new_n260_), .B(new_new_n207_), .C(new_new_n621_), .Y(new_new_n651_));
  OAI210     g0629(.A0(new_new_n651_), .A1(new_new_n226_), .B0(new_new_n62_), .Y(new_new_n652_));
  NA2        g0630(.A(new_new_n420_), .B(new_new_n31_), .Y(new_new_n653_));
  OR2        g0631(.A(new_new_n207_), .B(new_new_n103_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n654_), .B(new_new_n653_), .Y(new_new_n655_));
  NO2        g0633(.A(new_new_n62_), .B(i_9_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n62_), .B(new_new_n655_), .Y(new_new_n657_));
  NO2        g0635(.A(i_1_), .B(i_12_), .Y(new_new_n658_));
  NA3        g0636(.A(new_new_n658_), .B(new_new_n105_), .C(new_new_n24_), .Y(new_new_n659_));
  NA4        g0637(.A(new_new_n659_), .B(new_new_n657_), .C(new_new_n652_), .D(new_new_n650_), .Y(new_new_n660_));
  OAI210     g0638(.A0(new_new_n660_), .A1(new_new_n649_), .B0(i_6_), .Y(new_new_n661_));
  OAI210     g0639(.A0(new_new_n647_), .A1(new_new_n103_), .B0(new_new_n475_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(new_new_n605_), .Y(new_new_n663_));
  NO2        g0641(.A(i_6_), .B(i_11_), .Y(new_new_n664_));
  NA3        g0642(.A(new_new_n663_), .B(new_new_n536_), .C(new_new_n468_), .Y(new_new_n665_));
  NO4        g0643(.A(new_new_n214_), .B(new_new_n123_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n666_));
  NA2        g0644(.A(new_new_n666_), .B(new_new_n656_), .Y(new_new_n667_));
  NO3        g0645(.A(new_new_n636_), .B(new_new_n232_), .C(new_new_n23_), .Y(new_new_n668_));
  AOI210     g0646(.A0(i_1_), .A1(new_new_n261_), .B0(new_new_n668_), .Y(new_new_n669_));
  OAI210     g0647(.A0(new_new_n669_), .A1(new_new_n44_), .B0(new_new_n667_), .Y(new_new_n670_));
  NA3        g0648(.A(new_new_n553_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n671_));
  NA2        g0649(.A(new_new_n133_), .B(i_9_), .Y(new_new_n672_));
  NA3        g0650(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n46_), .B(i_1_), .Y(new_new_n674_));
  NA3        g0652(.A(new_new_n674_), .B(new_new_n270_), .C(new_new_n44_), .Y(new_new_n675_));
  OAI220     g0653(.A0(new_new_n675_), .A1(new_new_n673_), .B0(new_new_n672_), .B1(new_new_n1094_), .Y(new_new_n676_));
  NA3        g0654(.A(new_new_n656_), .B(new_new_n318_), .C(i_6_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n677_), .B(new_new_n23_), .Y(new_new_n678_));
  NAi21      g0656(.An(new_new_n671_), .B(new_new_n91_), .Y(new_new_n679_));
  NA2        g0657(.A(new_new_n674_), .B(new_new_n270_), .Y(new_new_n680_));
  NO2        g0658(.A(i_11_), .B(new_new_n37_), .Y(new_new_n681_));
  NA2        g0659(.A(new_new_n681_), .B(new_new_n24_), .Y(new_new_n682_));
  OAI210     g0660(.A0(new_new_n682_), .A1(new_new_n680_), .B0(new_new_n679_), .Y(new_new_n683_));
  OR3        g0661(.A(new_new_n683_), .B(new_new_n678_), .C(new_new_n676_), .Y(new_new_n684_));
  NO3        g0662(.A(new_new_n684_), .B(new_new_n670_), .C(new_new_n665_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n236_), .B(new_new_n98_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n686_), .B(new_new_n644_), .Y(new_new_n687_));
  NO2        g0665(.A(new_new_n426_), .B(new_new_n84_), .Y(new_new_n688_));
  NA2        g0666(.A(i_3_), .B(new_new_n191_), .Y(new_new_n689_));
  AN2        g0667(.A(new_new_n1105_), .B(new_new_n559_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n232_), .B(new_new_n44_), .Y(new_new_n691_));
  NO3        g0669(.A(new_new_n691_), .B(new_new_n311_), .C(new_new_n237_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n112_), .B(new_new_n37_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n693_), .B(i_6_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n84_), .B(i_9_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n62_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n658_), .Y(new_new_n697_));
  NO4        g0675(.A(new_new_n697_), .B(new_new_n694_), .C(new_new_n692_), .D(i_4_), .Y(new_new_n698_));
  NA2        g0676(.A(i_1_), .B(i_3_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n469_), .B(new_new_n92_), .Y(new_new_n700_));
  AOI210     g0678(.A0(new_new_n691_), .A1(new_new_n593_), .B0(new_new_n700_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n701_), .B(new_new_n699_), .Y(new_new_n702_));
  NO3        g0680(.A(new_new_n702_), .B(new_new_n698_), .C(new_new_n690_), .Y(new_new_n703_));
  NA3        g0681(.A(new_new_n703_), .B(new_new_n685_), .C(new_new_n661_), .Y(new_new_n704_));
  NO3        g0682(.A(new_new_n490_), .B(i_3_), .C(i_7_), .Y(new_new_n705_));
  OA210      g0683(.A0(new_new_n705_), .A1(new_new_n245_), .B0(new_new_n84_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n707_));
  NA3        g0685(.A(new_new_n497_), .B(new_new_n534_), .C(new_new_n46_), .Y(new_new_n708_));
  NO3        g0686(.A(new_new_n491_), .B(new_new_n630_), .C(new_new_n84_), .Y(new_new_n709_));
  NA2        g0687(.A(new_new_n709_), .B(new_new_n25_), .Y(new_new_n710_));
  NA3        g0688(.A(new_new_n157_), .B(new_new_n82_), .C(new_new_n84_), .Y(new_new_n711_));
  NA4        g0689(.A(new_new_n711_), .B(new_new_n710_), .C(new_new_n708_), .D(new_new_n707_), .Y(new_new_n712_));
  OAI210     g0690(.A0(new_new_n712_), .A1(new_new_n706_), .B0(i_1_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n374_), .B(i_2_), .Y(new_new_n714_));
  AOI210     g0692(.A0(new_new_n677_), .A1(new_new_n713_), .B0(i_13_), .Y(new_new_n715_));
  OR2        g0693(.A(i_11_), .B(i_7_), .Y(new_new_n716_));
  NA3        g0694(.A(new_new_n716_), .B(new_new_n102_), .C(new_new_n133_), .Y(new_new_n717_));
  AOI220     g0695(.A0(new_new_n485_), .A1(new_new_n157_), .B0(new_new_n462_), .B1(new_new_n133_), .Y(new_new_n718_));
  OAI210     g0696(.A0(new_new_n718_), .A1(new_new_n44_), .B0(new_new_n717_), .Y(new_new_n719_));
  AOI210     g0697(.A0(new_new_n673_), .A1(new_new_n53_), .B0(i_12_), .Y(new_new_n720_));
  NO2        g0698(.A(new_new_n491_), .B(new_new_n24_), .Y(new_new_n721_));
  AOI220     g0699(.A0(new_new_n721_), .A1(new_new_n688_), .B0(new_new_n245_), .B1(new_new_n126_), .Y(new_new_n722_));
  OAI220     g0700(.A0(new_new_n722_), .A1(new_new_n40_), .B0(new_new_n1093_), .B1(new_new_n92_), .Y(new_new_n723_));
  AOI210     g0701(.A0(new_new_n719_), .A1(new_new_n335_), .B0(new_new_n723_), .Y(new_new_n724_));
  NA2        g0702(.A(new_new_n109_), .B(new_new_n103_), .Y(new_new_n725_));
  AOI220     g0703(.A0(new_new_n725_), .A1(new_new_n70_), .B0(new_new_n392_), .B1(new_new_n674_), .Y(new_new_n726_));
  NO2        g0704(.A(new_new_n726_), .B(new_new_n242_), .Y(new_new_n727_));
  AOI210     g0705(.A0(new_new_n460_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n728_));
  NOi31      g0706(.An(new_new_n728_), .B(new_new_n620_), .C(new_new_n44_), .Y(new_new_n729_));
  NA2        g0707(.A(new_new_n122_), .B(i_13_), .Y(new_new_n730_));
  NO2        g0708(.A(new_new_n673_), .B(new_new_n109_), .Y(new_new_n731_));
  INV        g0709(.A(new_new_n731_), .Y(new_new_n732_));
  OAI220     g0710(.A0(new_new_n732_), .A1(new_new_n69_), .B0(new_new_n730_), .B1(new_new_n1099_), .Y(new_new_n733_));
  NO3        g0711(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n98_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n26_), .B(new_new_n191_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(i_7_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n491_), .B(new_new_n236_), .C(new_new_n84_), .Y(new_new_n737_));
  AOI210     g0715(.A0(new_new_n737_), .A1(new_new_n736_), .B0(new_new_n734_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n392_), .A1(new_new_n674_), .B0(new_new_n91_), .B1(i_2_), .Y(new_new_n739_));
  OAI220     g0717(.A0(new_new_n739_), .A1(new_new_n625_), .B0(new_new_n738_), .B1(new_new_n640_), .Y(new_new_n740_));
  NO4        g0718(.A(new_new_n740_), .B(new_new_n733_), .C(new_new_n729_), .D(new_new_n727_), .Y(new_new_n741_));
  OR2        g0719(.A(i_11_), .B(i_6_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n624_), .B(new_new_n735_), .C(i_7_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n743_), .A1(new_new_n732_), .B0(new_new_n742_), .Y(new_new_n744_));
  NA2        g0722(.A(new_new_n664_), .B(i_13_), .Y(new_new_n745_));
  NA2        g0723(.A(i_2_), .B(new_new_n735_), .Y(new_new_n746_));
  NAi21      g0724(.An(i_11_), .B(i_12_), .Y(new_new_n747_));
  NOi41      g0725(.An(new_new_n106_), .B(new_new_n747_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n748_));
  NO3        g0726(.A(new_new_n491_), .B(new_new_n605_), .C(new_new_n630_), .Y(new_new_n749_));
  AOI220     g0727(.A0(new_new_n749_), .A1(new_new_n315_), .B0(new_new_n748_), .B1(new_new_n746_), .Y(new_new_n750_));
  NA2        g0728(.A(new_new_n750_), .B(new_new_n745_), .Y(new_new_n751_));
  OAI210     g0729(.A0(new_new_n751_), .A1(new_new_n744_), .B0(new_new_n62_), .Y(new_new_n752_));
  NO2        g0730(.A(i_2_), .B(i_12_), .Y(new_new_n753_));
  OAI210     g0731(.A0(new_new_n634_), .A1(new_new_n373_), .B0(new_new_n753_), .Y(new_new_n754_));
  NA2        g0732(.A(i_8_), .B(new_new_n25_), .Y(new_new_n755_));
  NO3        g0733(.A(new_new_n755_), .B(new_new_n390_), .C(new_new_n624_), .Y(new_new_n756_));
  OAI210     g0734(.A0(new_new_n756_), .A1(new_new_n375_), .B0(new_new_n373_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n123_), .B(i_2_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n758_), .B(new_new_n658_), .Y(new_new_n759_));
  NA3        g0737(.A(new_new_n759_), .B(new_new_n757_), .C(new_new_n754_), .Y(new_new_n760_));
  NA3        g0738(.A(new_new_n760_), .B(new_new_n45_), .C(new_new_n225_), .Y(new_new_n761_));
  NA4        g0739(.A(new_new_n761_), .B(new_new_n752_), .C(new_new_n741_), .D(new_new_n724_), .Y(new_new_n762_));
  OR4        g0740(.A(new_new_n762_), .B(new_new_n715_), .C(new_new_n704_), .D(new_new_n643_), .Y(men5));
  AOI210     g0741(.A0(new_new_n687_), .A1(new_new_n273_), .B0(new_new_n429_), .Y(new_new_n764_));
  AO210      g0742(.A0(new_new_n24_), .A1(i_10_), .B0(new_new_n251_), .Y(new_new_n765_));
  NA3        g0743(.A(new_new_n765_), .B(new_new_n753_), .C(new_new_n103_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n764_), .C(new_new_n536_), .Y(new_new_n767_));
  NO3        g0745(.A(i_11_), .B(new_new_n236_), .C(i_13_), .Y(new_new_n768_));
  NO2        g0746(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n769_));
  NA2        g0747(.A(i_12_), .B(i_8_), .Y(new_new_n770_));
  INV        g0748(.A(new_new_n459_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n318_), .B(new_new_n597_), .Y(new_new_n772_));
  INV        g0750(.A(new_new_n772_), .Y(new_new_n773_));
  NO2        g0751(.A(new_new_n773_), .B(new_new_n767_), .Y(new_new_n774_));
  INV        g0752(.A(new_new_n168_), .Y(new_new_n775_));
  OAI210     g0753(.A0(new_new_n714_), .A1(new_new_n461_), .B0(new_new_n106_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n776_), .B(new_new_n775_), .Y(new_new_n777_));
  NO2        g0755(.A(new_new_n469_), .B(new_new_n26_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n778_), .B(new_new_n431_), .Y(new_new_n779_));
  NA2        g0757(.A(new_new_n779_), .B(i_2_), .Y(new_new_n780_));
  INV        g0758(.A(new_new_n780_), .Y(new_new_n781_));
  AOI210     g0759(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n427_), .Y(new_new_n782_));
  AOI210     g0760(.A0(new_new_n782_), .A1(new_new_n781_), .B0(new_new_n777_), .Y(new_new_n783_));
  NO2        g0761(.A(new_new_n188_), .B(new_new_n120_), .Y(new_new_n784_));
  OAI210     g0762(.A0(new_new_n784_), .A1(new_new_n769_), .B0(i_2_), .Y(new_new_n785_));
  INV        g0763(.A(new_new_n169_), .Y(new_new_n786_));
  NO3        g0764(.A(new_new_n645_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n787_));
  AOI210     g0765(.A0(new_new_n786_), .A1(new_new_n87_), .B0(new_new_n787_), .Y(new_new_n788_));
  AOI210     g0766(.A0(new_new_n788_), .A1(new_new_n785_), .B0(new_new_n191_), .Y(new_new_n789_));
  OA210      g0767(.A0(new_new_n646_), .A1(new_new_n121_), .B0(i_13_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n198_), .B(new_new_n201_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n147_), .B(new_new_n621_), .Y(new_new_n792_));
  AOI210     g0770(.A0(new_new_n792_), .A1(new_new_n791_), .B0(new_new_n378_), .Y(new_new_n793_));
  AOI210     g0771(.A0(new_new_n207_), .A1(new_new_n143_), .B0(new_new_n534_), .Y(new_new_n794_));
  OAI210     g0772(.A0(new_new_n794_), .A1(new_new_n226_), .B0(new_new_n431_), .Y(new_new_n795_));
  NA3        g0773(.A(new_new_n308_), .B(new_new_n119_), .C(new_new_n42_), .Y(new_new_n796_));
  OAI210     g0774(.A0(new_new_n796_), .A1(new_new_n46_), .B0(new_new_n795_), .Y(new_new_n797_));
  NO4        g0775(.A(new_new_n797_), .B(new_new_n793_), .C(new_new_n790_), .D(new_new_n789_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n61_), .B(i_12_), .Y(new_new_n799_));
  NO2        g0777(.A(new_new_n799_), .B(new_new_n121_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n800_), .B(new_new_n621_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n801_), .B(new_new_n36_), .Y(new_new_n802_));
  NA4        g0780(.A(new_new_n802_), .B(new_new_n798_), .C(new_new_n783_), .D(new_new_n774_), .Y(men6));
  NO3        g0781(.A(new_new_n256_), .B(new_new_n310_), .C(i_1_), .Y(new_new_n804_));
  NO2        g0782(.A(new_new_n183_), .B(new_new_n134_), .Y(new_new_n805_));
  OAI210     g0783(.A0(new_new_n805_), .A1(new_new_n804_), .B0(new_new_n758_), .Y(new_new_n806_));
  NA4        g0784(.A(new_new_n396_), .B(new_new_n496_), .C(new_new_n69_), .D(new_new_n98_), .Y(new_new_n807_));
  INV        g0785(.A(new_new_n807_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n220_), .B(new_new_n501_), .Y(new_new_n809_));
  NO2        g0787(.A(i_11_), .B(i_9_), .Y(new_new_n810_));
  NO3        g0788(.A(new_new_n809_), .B(new_new_n808_), .C(new_new_n330_), .Y(new_new_n811_));
  AO210      g0789(.A0(new_new_n811_), .A1(new_new_n806_), .B0(i_12_), .Y(new_new_n812_));
  NA2        g0790(.A(new_new_n379_), .B(new_new_n338_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n605_), .B(new_new_n62_), .Y(new_new_n814_));
  NA2        g0792(.A(new_new_n705_), .B(new_new_n69_), .Y(new_new_n815_));
  NA4        g0793(.A(new_new_n85_), .B(new_new_n815_), .C(new_new_n814_), .D(new_new_n813_), .Y(new_new_n816_));
  INV        g0794(.A(new_new_n195_), .Y(new_new_n817_));
  AOI220     g0795(.A0(new_new_n817_), .A1(new_new_n810_), .B0(new_new_n816_), .B1(new_new_n71_), .Y(new_new_n818_));
  INV        g0796(.A(new_new_n329_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n73_), .B(new_new_n126_), .Y(new_new_n820_));
  INV        g0798(.A(new_new_n119_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n821_), .B(new_new_n46_), .Y(new_new_n822_));
  AOI210     g0800(.A0(new_new_n822_), .A1(new_new_n820_), .B0(new_new_n819_), .Y(new_new_n823_));
  NO3        g0801(.A(new_new_n252_), .B(new_new_n127_), .C(i_9_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n824_), .B(new_new_n799_), .Y(new_new_n825_));
  AOI210     g0803(.A0(new_new_n825_), .A1(new_new_n532_), .B0(new_new_n183_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n32_), .B(i_11_), .Y(new_new_n827_));
  NA3        g0805(.A(new_new_n827_), .B(new_new_n488_), .C(new_new_n396_), .Y(new_new_n828_));
  OAI210     g0806(.A0(new_new_n705_), .A1(new_new_n585_), .B0(new_new_n584_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n829_), .B(new_new_n828_), .Y(new_new_n830_));
  OR3        g0808(.A(new_new_n830_), .B(new_new_n826_), .C(new_new_n823_), .Y(new_new_n831_));
  NO2        g0809(.A(new_new_n716_), .B(i_2_), .Y(new_new_n832_));
  NA2        g0810(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n833_));
  NA2        g0811(.A(new_new_n1103_), .B(new_new_n832_), .Y(new_new_n834_));
  AO220      g0812(.A0(new_new_n362_), .A1(new_new_n352_), .B0(new_new_n403_), .B1(new_new_n621_), .Y(new_new_n835_));
  NA3        g0813(.A(new_new_n835_), .B(new_new_n257_), .C(i_7_), .Y(new_new_n836_));
  OR2        g0814(.A(new_new_n646_), .B(new_new_n461_), .Y(new_new_n837_));
  NA3        g0815(.A(new_new_n837_), .B(new_new_n142_), .C(new_new_n67_), .Y(new_new_n838_));
  AO210      g0816(.A0(new_new_n507_), .A1(new_new_n771_), .B0(new_new_n36_), .Y(new_new_n839_));
  NA4        g0817(.A(new_new_n839_), .B(new_new_n838_), .C(new_new_n836_), .D(new_new_n834_), .Y(new_new_n840_));
  OAI210     g0818(.A0(i_6_), .A1(i_11_), .B0(new_new_n85_), .Y(new_new_n841_));
  AOI220     g0819(.A0(new_new_n841_), .A1(new_new_n584_), .B0(new_new_n809_), .B1(new_new_n736_), .Y(new_new_n842_));
  NA3        g0820(.A(new_new_n378_), .B(new_new_n238_), .C(new_new_n142_), .Y(new_new_n843_));
  OAI210     g0821(.A0(new_new_n403_), .A1(new_new_n202_), .B0(new_new_n68_), .Y(new_new_n844_));
  NA4        g0822(.A(new_new_n844_), .B(new_new_n843_), .C(new_new_n842_), .D(new_new_n628_), .Y(new_new_n845_));
  AO210      g0823(.A0(new_new_n534_), .A1(new_new_n46_), .B0(new_new_n86_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n846_), .B(new_new_n497_), .C(new_new_n217_), .Y(new_new_n847_));
  AOI210     g0825(.A0(new_new_n461_), .A1(new_new_n459_), .B0(new_new_n583_), .Y(new_new_n848_));
  NO2        g0826(.A(new_new_n636_), .B(i_2_), .Y(new_new_n849_));
  OAI210     g0827(.A0(new_new_n849_), .A1(new_new_n107_), .B0(new_new_n418_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n244_), .B(new_new_n46_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n851_), .B(new_new_n612_), .Y(new_new_n852_));
  NA3        g0830(.A(new_new_n852_), .B(new_new_n329_), .C(i_7_), .Y(new_new_n853_));
  NA4        g0831(.A(new_new_n853_), .B(new_new_n850_), .C(new_new_n848_), .D(new_new_n847_), .Y(new_new_n854_));
  NO4        g0832(.A(new_new_n854_), .B(new_new_n845_), .C(new_new_n840_), .D(new_new_n831_), .Y(new_new_n855_));
  NA4        g0833(.A(new_new_n855_), .B(new_new_n818_), .C(new_new_n812_), .D(new_new_n386_), .Y(men3));
  NA2        g0834(.A(i_12_), .B(i_10_), .Y(new_new_n857_));
  NA2        g0835(.A(i_6_), .B(i_7_), .Y(new_new_n858_));
  NO2        g0836(.A(new_new_n858_), .B(i_0_), .Y(new_new_n859_));
  NO2        g0837(.A(i_11_), .B(new_new_n236_), .Y(new_new_n860_));
  OAI210     g0838(.A0(new_new_n859_), .A1(new_new_n293_), .B0(new_new_n860_), .Y(new_new_n861_));
  NO2        g0839(.A(new_new_n861_), .B(new_new_n191_), .Y(new_new_n862_));
  NO3        g0840(.A(new_new_n465_), .B(new_new_n89_), .C(new_new_n44_), .Y(new_new_n863_));
  OA210      g0841(.A0(new_new_n863_), .A1(new_new_n862_), .B0(new_new_n171_), .Y(new_new_n864_));
  NA3        g0842(.A(new_new_n843_), .B(new_new_n628_), .C(new_new_n377_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n865_), .B(new_new_n39_), .Y(new_new_n866_));
  NOi21      g0844(.An(new_new_n94_), .B(new_new_n779_), .Y(new_new_n867_));
  NO3        g0845(.A(new_new_n654_), .B(new_new_n469_), .C(new_new_n126_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n420_), .B(new_new_n45_), .Y(new_new_n869_));
  AN2        g0847(.A(new_new_n467_), .B(new_new_n54_), .Y(new_new_n870_));
  NO3        g0848(.A(new_new_n870_), .B(new_new_n868_), .C(new_new_n867_), .Y(new_new_n871_));
  AOI210     g0849(.A0(new_new_n871_), .A1(new_new_n866_), .B0(new_new_n48_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n183_), .B(new_new_n593_), .Y(new_new_n873_));
  NA2        g0851(.A(new_new_n728_), .B(new_new_n695_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n336_), .B(new_new_n451_), .Y(new_new_n875_));
  OAI220     g0853(.A0(new_new_n875_), .A1(new_new_n874_), .B0(new_new_n873_), .B1(new_new_n62_), .Y(new_new_n876_));
  NOi21      g0854(.An(i_5_), .B(i_9_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n877_), .B(new_new_n458_), .Y(new_new_n878_));
  INV        g0856(.A(new_new_n709_), .Y(new_new_n879_));
  NO3        g0857(.A(new_new_n423_), .B(new_new_n270_), .C(new_new_n71_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n172_), .B(new_new_n143_), .Y(new_new_n881_));
  AOI210     g0859(.A0(new_new_n881_), .A1(new_new_n244_), .B0(new_new_n880_), .Y(new_new_n882_));
  OAI220     g0860(.A0(new_new_n882_), .A1(new_new_n178_), .B0(new_new_n879_), .B1(new_new_n878_), .Y(new_new_n883_));
  NO4        g0861(.A(new_new_n883_), .B(new_new_n876_), .C(new_new_n872_), .D(new_new_n864_), .Y(new_new_n884_));
  NOi21      g0862(.An(i_0_), .B(i_10_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n183_), .B(new_new_n24_), .Y(new_new_n886_));
  NO2        g0864(.A(new_new_n693_), .B(new_new_n618_), .Y(new_new_n887_));
  NO2        g0865(.A(new_new_n887_), .B(new_new_n886_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n315_), .B(new_new_n124_), .Y(new_new_n889_));
  NAi21      g0867(.An(new_new_n158_), .B(new_new_n451_), .Y(new_new_n890_));
  OAI220     g0868(.A0(new_new_n890_), .A1(new_new_n851_), .B0(new_new_n889_), .B1(new_new_n409_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n891_), .B(new_new_n888_), .Y(new_new_n892_));
  NO2        g0870(.A(new_new_n396_), .B(new_new_n297_), .Y(new_new_n893_));
  NA2        g0871(.A(new_new_n893_), .B(new_new_n731_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n594_), .B(i_0_), .Y(new_new_n895_));
  NO3        g0873(.A(new_new_n895_), .B(new_new_n391_), .C(new_new_n87_), .Y(new_new_n896_));
  NO4        g0874(.A(new_new_n611_), .B(new_new_n214_), .C(new_new_n427_), .D(new_new_n419_), .Y(new_new_n897_));
  AOI210     g0875(.A0(new_new_n897_), .A1(i_11_), .B0(new_new_n896_), .Y(new_new_n898_));
  INV        g0876(.A(new_new_n488_), .Y(new_new_n899_));
  AN2        g0877(.A(new_new_n94_), .B(new_new_n243_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n768_), .B(new_new_n330_), .Y(new_new_n901_));
  AOI210     g0879(.A0(new_new_n497_), .A1(new_new_n87_), .B0(new_new_n57_), .Y(new_new_n902_));
  OAI220     g0880(.A0(new_new_n902_), .A1(new_new_n901_), .B0(new_new_n682_), .B1(new_new_n555_), .Y(new_new_n903_));
  NO2        g0881(.A(new_new_n254_), .B(new_new_n149_), .Y(new_new_n904_));
  NA2        g0882(.A(i_0_), .B(i_10_), .Y(new_new_n905_));
  OAI210     g0883(.A0(new_new_n905_), .A1(new_new_n84_), .B0(new_new_n558_), .Y(new_new_n906_));
  NO4        g0884(.A(new_new_n109_), .B(new_new_n57_), .C(new_new_n689_), .D(i_5_), .Y(new_new_n907_));
  AO220      g0885(.A0(new_new_n907_), .A1(new_new_n906_), .B0(new_new_n904_), .B1(i_6_), .Y(new_new_n908_));
  AOI220     g0886(.A0(new_new_n336_), .A1(new_new_n96_), .B0(new_new_n183_), .B1(new_new_n82_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n588_), .B(i_4_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n186_), .B(new_new_n201_), .Y(new_new_n911_));
  OAI220     g0889(.A0(new_new_n911_), .A1(new_new_n901_), .B0(new_new_n910_), .B1(new_new_n909_), .Y(new_new_n912_));
  NO4        g0890(.A(new_new_n912_), .B(new_new_n908_), .C(new_new_n903_), .D(new_new_n900_), .Y(new_new_n913_));
  NA4        g0891(.A(new_new_n913_), .B(new_new_n898_), .C(new_new_n894_), .D(new_new_n892_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n915_));
  NA2        g0893(.A(i_11_), .B(i_9_), .Y(new_new_n916_));
  NO3        g0894(.A(i_12_), .B(new_new_n916_), .C(new_new_n627_), .Y(new_new_n917_));
  AO220      g0895(.A0(new_new_n917_), .A1(new_new_n915_), .B0(new_new_n272_), .B1(new_new_n86_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n48_), .B(i_7_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n916_), .B(new_new_n71_), .Y(new_new_n920_));
  NO2        g0898(.A(new_new_n172_), .B(i_0_), .Y(new_new_n921_));
  INV        g0899(.A(new_new_n921_), .Y(new_new_n922_));
  NA2        g0900(.A(new_new_n488_), .B(new_new_n231_), .Y(new_new_n923_));
  AOI210     g0901(.A0(new_new_n376_), .A1(new_new_n41_), .B0(new_new_n417_), .Y(new_new_n924_));
  OAI220     g0902(.A0(new_new_n924_), .A1(new_new_n878_), .B0(new_new_n923_), .B1(new_new_n922_), .Y(new_new_n925_));
  NO2        g0903(.A(new_new_n925_), .B(new_new_n918_), .Y(new_new_n926_));
  AOI210     g0904(.A0(new_new_n460_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n927_));
  NA2        g0905(.A(new_new_n168_), .B(new_new_n99_), .Y(new_new_n928_));
  NOi32      g0906(.An(new_new_n927_), .Bn(new_new_n186_), .C(new_new_n928_), .Y(new_new_n929_));
  AOI210     g0907(.A0(new_new_n629_), .A1(new_new_n330_), .B0(new_new_n243_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n930_), .B(new_new_n869_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n931_), .B(new_new_n929_), .Y(new_new_n932_));
  NOi21      g0910(.An(i_7_), .B(i_5_), .Y(new_new_n933_));
  NOi31      g0911(.An(new_new_n933_), .B(new_new_n885_), .C(new_new_n747_), .Y(new_new_n934_));
  NA3        g0912(.A(new_new_n934_), .B(new_new_n390_), .C(i_6_), .Y(new_new_n935_));
  OA210      g0913(.A0(new_new_n928_), .A1(new_new_n532_), .B0(new_new_n935_), .Y(new_new_n936_));
  NO3        g0914(.A(new_new_n412_), .B(new_new_n365_), .C(new_new_n361_), .Y(new_new_n937_));
  INV        g0915(.A(new_new_n319_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n747_), .B(new_new_n259_), .Y(new_new_n939_));
  AOI210     g0917(.A0(new_new_n939_), .A1(new_new_n938_), .B0(new_new_n937_), .Y(new_new_n940_));
  NA4        g0918(.A(new_new_n940_), .B(new_new_n936_), .C(new_new_n932_), .D(new_new_n926_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n886_), .B(new_new_n239_), .Y(new_new_n942_));
  AN2        g0920(.A(new_new_n335_), .B(new_new_n330_), .Y(new_new_n943_));
  AO220      g0921(.A0(new_new_n943_), .A1(new_new_n881_), .B0(new_new_n347_), .B1(new_new_n27_), .Y(new_new_n944_));
  OAI210     g0922(.A0(new_new_n944_), .A1(new_new_n942_), .B0(i_10_), .Y(new_new_n945_));
  INV        g0923(.A(new_new_n857_), .Y(new_new_n946_));
  OA210      g0924(.A0(new_new_n488_), .A1(new_new_n223_), .B0(new_new_n487_), .Y(new_new_n947_));
  OAI210     g0925(.A0(new_new_n947_), .A1(new_new_n946_), .B0(new_new_n920_), .Y(new_new_n948_));
  NA3        g0926(.A(new_new_n487_), .B(new_new_n420_), .C(new_new_n45_), .Y(new_new_n949_));
  OAI210     g0927(.A0(new_new_n890_), .A1(new_new_n899_), .B0(new_new_n949_), .Y(new_new_n950_));
  NO2        g0928(.A(new_new_n257_), .B(new_new_n46_), .Y(new_new_n951_));
  NA2        g0929(.A(new_new_n920_), .B(new_new_n308_), .Y(new_new_n952_));
  OAI210     g0930(.A0(new_new_n951_), .A1(new_new_n185_), .B0(new_new_n952_), .Y(new_new_n953_));
  AOI220     g0931(.A0(new_new_n953_), .A1(new_new_n488_), .B0(new_new_n950_), .B1(new_new_n71_), .Y(new_new_n954_));
  NA3        g0932(.A(new_new_n833_), .B(new_new_n388_), .C(i_6_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n92_), .B(new_new_n44_), .Y(new_new_n956_));
  NO2        g0934(.A(new_new_n73_), .B(new_new_n770_), .Y(new_new_n957_));
  AOI220     g0935(.A0(new_new_n957_), .A1(new_new_n956_), .B0(new_new_n171_), .B1(new_new_n618_), .Y(new_new_n958_));
  AOI210     g0936(.A0(new_new_n958_), .A1(new_new_n955_), .B0(new_new_n47_), .Y(new_new_n959_));
  NO3        g0937(.A(new_new_n611_), .B(new_new_n360_), .C(new_new_n24_), .Y(new_new_n960_));
  AOI210     g0938(.A0(new_new_n721_), .A1(new_new_n567_), .B0(new_new_n960_), .Y(new_new_n961_));
  NAi21      g0939(.An(i_9_), .B(i_5_), .Y(new_new_n962_));
  NO2        g0940(.A(new_new_n962_), .B(new_new_n412_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n623_), .B(new_new_n101_), .Y(new_new_n964_));
  AOI220     g0942(.A0(new_new_n964_), .A1(i_0_), .B0(new_new_n963_), .B1(new_new_n646_), .Y(new_new_n965_));
  OAI220     g0943(.A0(new_new_n965_), .A1(new_new_n84_), .B0(new_new_n961_), .B1(new_new_n169_), .Y(new_new_n966_));
  NO3        g0944(.A(new_new_n966_), .B(new_new_n959_), .C(new_new_n537_), .Y(new_new_n967_));
  NA4        g0945(.A(new_new_n967_), .B(new_new_n954_), .C(new_new_n948_), .D(new_new_n945_), .Y(new_new_n968_));
  NO3        g0946(.A(new_new_n968_), .B(new_new_n941_), .C(new_new_n914_), .Y(new_new_n969_));
  NO2        g0947(.A(new_new_n885_), .B(new_new_n747_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n71_), .B(new_new_n44_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n905_), .B(new_new_n971_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n101_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n973_));
  AO220      g0951(.A0(new_new_n973_), .A1(new_new_n972_), .B0(new_new_n970_), .B1(new_new_n171_), .Y(new_new_n974_));
  AOI210     g0952(.A0(new_new_n814_), .A1(new_new_n707_), .B0(new_new_n928_), .Y(new_new_n975_));
  AOI210     g0953(.A0(new_new_n974_), .A1(new_new_n349_), .B0(new_new_n975_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n758_), .B(new_new_n141_), .Y(new_new_n977_));
  INV        g0955(.A(new_new_n977_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n978_), .B(new_new_n695_), .C(new_new_n71_), .Y(new_new_n979_));
  NO2        g0957(.A(new_new_n829_), .B(new_new_n412_), .Y(new_new_n980_));
  NA3        g0958(.A(new_new_n859_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n860_), .B(i_9_), .Y(new_new_n982_));
  AOI210     g0960(.A0(new_new_n981_), .A1(new_new_n512_), .B0(new_new_n982_), .Y(new_new_n983_));
  OAI210     g0961(.A0(new_new_n244_), .A1(i_9_), .B0(new_new_n230_), .Y(new_new_n984_));
  AOI210     g0962(.A0(new_new_n984_), .A1(new_new_n895_), .B0(new_new_n149_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n985_), .B(new_new_n983_), .C(new_new_n980_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n986_), .B(new_new_n979_), .C(new_new_n976_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n943_), .B(new_new_n378_), .Y(new_new_n988_));
  AOI210     g0966(.A0(new_new_n304_), .A1(new_new_n158_), .B0(new_new_n988_), .Y(new_new_n989_));
  NA2        g0967(.A(new_new_n39_), .B(new_new_n44_), .Y(new_new_n990_));
  NA2        g0968(.A(new_new_n919_), .B(new_new_n502_), .Y(new_new_n991_));
  AOI210     g0969(.A0(new_new_n990_), .A1(new_new_n158_), .B0(new_new_n991_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n992_), .B(new_new_n989_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n905_), .B(new_new_n877_), .C(new_new_n188_), .Y(new_new_n994_));
  AOI220     g0972(.A0(new_new_n994_), .A1(i_11_), .B0(new_new_n589_), .B1(new_new_n73_), .Y(new_new_n995_));
  NO3        g0973(.A(new_new_n209_), .B(new_new_n389_), .C(i_0_), .Y(new_new_n996_));
  OAI210     g0974(.A0(new_new_n996_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n997_));
  INV        g0975(.A(new_new_n217_), .Y(new_new_n998_));
  OAI220     g0976(.A0(new_new_n548_), .A1(new_new_n134_), .B0(new_new_n1098_), .B1(new_new_n640_), .Y(new_new_n999_));
  NA3        g0977(.A(new_new_n999_), .B(new_new_n404_), .C(new_new_n998_), .Y(new_new_n1000_));
  NA4        g0978(.A(new_new_n1000_), .B(new_new_n997_), .C(new_new_n995_), .D(new_new_n993_), .Y(new_new_n1001_));
  NO2        g0979(.A(new_new_n242_), .B(new_new_n92_), .Y(new_new_n1002_));
  AOI210     g0980(.A0(new_new_n1002_), .A1(new_new_n970_), .B0(new_new_n104_), .Y(new_new_n1003_));
  AOI220     g0981(.A0(new_new_n933_), .A1(new_new_n502_), .B0(new_new_n859_), .B1(new_new_n159_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n352_), .B(new_new_n173_), .Y(new_new_n1005_));
  OA220      g0983(.A0(new_new_n1005_), .A1(new_new_n1004_), .B0(new_new_n1003_), .B1(i_5_), .Y(new_new_n1006_));
  AOI210     g0984(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n172_), .Y(new_new_n1007_));
  NA2        g0985(.A(new_new_n1007_), .B(new_new_n947_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n637_), .B(new_new_n183_), .C(new_new_n82_), .Y(new_new_n1009_));
  NA2        g0987(.A(new_new_n1009_), .B(new_new_n565_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n869_), .B(new_new_n53_), .C(new_new_n48_), .Y(new_new_n1011_));
  NO3        g0989(.A(new_new_n1096_), .B(new_new_n1011_), .C(new_new_n1010_), .Y(new_new_n1012_));
  NA3        g0990(.A(new_new_n396_), .B(new_new_n168_), .C(new_new_n167_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n919_), .B(new_new_n293_), .C(new_new_n230_), .Y(new_new_n1014_));
  NA2        g0992(.A(new_new_n1014_), .B(new_new_n1013_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n396_), .B(new_new_n337_), .C(new_new_n221_), .Y(new_new_n1016_));
  OAI210     g0994(.A0(new_new_n873_), .A1(new_new_n671_), .B0(new_new_n1016_), .Y(new_new_n1017_));
  NOi31      g0995(.An(new_new_n395_), .B(new_new_n971_), .C(new_new_n239_), .Y(new_new_n1018_));
  NO3        g0996(.A(new_new_n916_), .B(new_new_n217_), .C(new_new_n188_), .Y(new_new_n1019_));
  NO4        g0997(.A(new_new_n1019_), .B(new_new_n1018_), .C(new_new_n1017_), .D(new_new_n1015_), .Y(new_new_n1020_));
  NA4        g0998(.A(new_new_n1020_), .B(new_new_n1012_), .C(new_new_n1008_), .D(new_new_n1006_), .Y(new_new_n1021_));
  AOI210     g0999(.A0(new_new_n588_), .A1(new_new_n547_), .B0(new_new_n639_), .Y(new_new_n1022_));
  NO3        g1000(.A(new_new_n1022_), .B(new_new_n579_), .C(new_new_n346_), .Y(new_new_n1023_));
  NO2        g1001(.A(new_new_n84_), .B(i_5_), .Y(new_new_n1024_));
  NA3        g1002(.A(new_new_n860_), .B(new_new_n105_), .C(new_new_n119_), .Y(new_new_n1025_));
  INV        g1003(.A(new_new_n1025_), .Y(new_new_n1026_));
  AOI210     g1004(.A0(new_new_n1026_), .A1(new_new_n1024_), .B0(new_new_n1023_), .Y(new_new_n1027_));
  NA3        g1005(.A(new_new_n308_), .B(i_5_), .C(new_new_n191_), .Y(new_new_n1028_));
  NAi31      g1006(.An(new_new_n241_), .B(new_new_n1028_), .C(new_new_n242_), .Y(new_new_n1029_));
  NO4        g1007(.A(new_new_n239_), .B(new_new_n209_), .C(i_0_), .D(i_12_), .Y(new_new_n1030_));
  AOI220     g1008(.A0(new_new_n1030_), .A1(new_new_n1029_), .B0(new_new_n808_), .B1(new_new_n173_), .Y(new_new_n1031_));
  AN2        g1009(.A(new_new_n905_), .B(new_new_n149_), .Y(new_new_n1032_));
  NO4        g1010(.A(new_new_n1032_), .B(i_12_), .C(new_new_n671_), .D(new_new_n126_), .Y(new_new_n1033_));
  NA2        g1011(.A(new_new_n1033_), .B(new_new_n217_), .Y(new_new_n1034_));
  NA3        g1012(.A(new_new_n96_), .B(new_new_n593_), .C(i_11_), .Y(new_new_n1035_));
  NO2        g1013(.A(new_new_n1035_), .B(new_new_n151_), .Y(new_new_n1036_));
  NA2        g1014(.A(new_new_n933_), .B(new_new_n485_), .Y(new_new_n1037_));
  NA2        g1015(.A(new_new_n63_), .B(new_new_n98_), .Y(new_new_n1038_));
  OAI220     g1016(.A0(new_new_n1038_), .A1(new_new_n1028_), .B0(new_new_n1037_), .B1(new_new_n696_), .Y(new_new_n1039_));
  AOI210     g1017(.A0(new_new_n1039_), .A1(new_new_n921_), .B0(new_new_n1036_), .Y(new_new_n1040_));
  NA4        g1018(.A(new_new_n1040_), .B(new_new_n1034_), .C(new_new_n1031_), .D(new_new_n1027_), .Y(new_new_n1041_));
  NO4        g1019(.A(new_new_n1041_), .B(new_new_n1021_), .C(new_new_n1001_), .D(new_new_n987_), .Y(new_new_n1042_));
  OAI210     g1020(.A0(new_new_n832_), .A1(new_new_n827_), .B0(new_new_n37_), .Y(new_new_n1043_));
  NA3        g1021(.A(new_new_n927_), .B(new_new_n373_), .C(i_5_), .Y(new_new_n1044_));
  NA3        g1022(.A(new_new_n1044_), .B(new_new_n1043_), .C(new_new_n635_), .Y(new_new_n1045_));
  NA2        g1023(.A(new_new_n1045_), .B(new_new_n205_), .Y(new_new_n1046_));
  AN2        g1024(.A(new_new_n716_), .B(new_new_n374_), .Y(new_new_n1047_));
  NA2        g1025(.A(new_new_n184_), .B(new_new_n186_), .Y(new_new_n1048_));
  AO210      g1026(.A0(new_new_n1047_), .A1(new_new_n33_), .B0(new_new_n1048_), .Y(new_new_n1049_));
  OAI210     g1027(.A0(new_new_n639_), .A1(new_new_n637_), .B0(new_new_n318_), .Y(new_new_n1050_));
  NAi31      g1028(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1051_));
  AOI210     g1029(.A0(new_new_n112_), .A1(new_new_n68_), .B0(new_new_n1051_), .Y(new_new_n1052_));
  NO2        g1030(.A(new_new_n1052_), .B(new_new_n668_), .Y(new_new_n1053_));
  NA3        g1031(.A(new_new_n1053_), .B(new_new_n1050_), .C(new_new_n1049_), .Y(new_new_n1054_));
  NO2        g1032(.A(new_new_n475_), .B(new_new_n270_), .Y(new_new_n1055_));
  NO4        g1033(.A(new_new_n232_), .B(new_new_n140_), .C(new_new_n699_), .D(new_new_n37_), .Y(new_new_n1056_));
  NO3        g1034(.A(new_new_n1056_), .B(new_new_n1055_), .C(new_new_n897_), .Y(new_new_n1057_));
  OAI210     g1035(.A0(new_new_n1035_), .A1(new_new_n143_), .B0(new_new_n1057_), .Y(new_new_n1058_));
  AOI210     g1036(.A0(new_new_n1054_), .A1(new_new_n48_), .B0(new_new_n1058_), .Y(new_new_n1059_));
  AOI210     g1037(.A0(new_new_n1059_), .A1(new_new_n1046_), .B0(new_new_n71_), .Y(new_new_n1060_));
  NO2        g1038(.A(new_new_n586_), .B(new_new_n385_), .Y(new_new_n1061_));
  NO2        g1039(.A(new_new_n1061_), .B(new_new_n775_), .Y(new_new_n1062_));
  OAI210     g1040(.A0(new_new_n78_), .A1(new_new_n53_), .B0(new_new_n103_), .Y(new_new_n1063_));
  NA2        g1041(.A(new_new_n1063_), .B(new_new_n74_), .Y(new_new_n1064_));
  AOI210     g1042(.A0(new_new_n1007_), .A1(new_new_n919_), .B0(new_new_n934_), .Y(new_new_n1065_));
  AOI210     g1043(.A0(new_new_n1065_), .A1(new_new_n1064_), .B0(new_new_n699_), .Y(new_new_n1066_));
  NA2        g1044(.A(new_new_n264_), .B(new_new_n56_), .Y(new_new_n1067_));
  AOI220     g1045(.A0(new_new_n1067_), .A1(new_new_n74_), .B0(new_new_n347_), .B1(new_new_n256_), .Y(new_new_n1068_));
  NO2        g1046(.A(new_new_n1068_), .B(new_new_n236_), .Y(new_new_n1069_));
  NA3        g1047(.A(new_new_n94_), .B(new_new_n310_), .C(new_new_n31_), .Y(new_new_n1070_));
  INV        g1048(.A(new_new_n1070_), .Y(new_new_n1071_));
  NO3        g1049(.A(new_new_n1071_), .B(new_new_n1069_), .C(new_new_n1066_), .Y(new_new_n1072_));
  OAI210     g1050(.A0(new_new_n272_), .A1(new_new_n154_), .B0(new_new_n87_), .Y(new_new_n1073_));
  NA3        g1051(.A(new_new_n778_), .B(new_new_n293_), .C(new_new_n78_), .Y(new_new_n1074_));
  AOI210     g1052(.A0(new_new_n1074_), .A1(new_new_n1073_), .B0(i_11_), .Y(new_new_n1075_));
  NA2        g1053(.A(new_new_n630_), .B(new_new_n214_), .Y(new_new_n1076_));
  OAI210     g1054(.A0(new_new_n1076_), .A1(new_new_n927_), .B0(new_new_n205_), .Y(new_new_n1077_));
  NA2        g1055(.A(new_new_n160_), .B(i_5_), .Y(new_new_n1078_));
  AOI210     g1056(.A0(new_new_n1077_), .A1(new_new_n791_), .B0(new_new_n1078_), .Y(new_new_n1079_));
  NO3        g1057(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n1080_));
  OAI210     g1058(.A0(new_new_n938_), .A1(new_new_n310_), .B0(new_new_n1080_), .Y(new_new_n1081_));
  NO2        g1059(.A(new_new_n1081_), .B(new_new_n747_), .Y(new_new_n1082_));
  NO4        g1060(.A(new_new_n962_), .B(new_new_n490_), .C(new_new_n253_), .D(new_new_n252_), .Y(new_new_n1083_));
  NO2        g1061(.A(new_new_n1083_), .B(new_new_n583_), .Y(new_new_n1084_));
  INV        g1062(.A(new_new_n366_), .Y(new_new_n1085_));
  AOI210     g1063(.A0(new_new_n1085_), .A1(new_new_n1084_), .B0(new_new_n40_), .Y(new_new_n1086_));
  NO4        g1064(.A(new_new_n1086_), .B(new_new_n1082_), .C(new_new_n1079_), .D(new_new_n1075_), .Y(new_new_n1087_));
  OAI210     g1065(.A0(new_new_n1072_), .A1(i_4_), .B0(new_new_n1087_), .Y(new_new_n1088_));
  NO3        g1066(.A(new_new_n1088_), .B(new_new_n1062_), .C(new_new_n1060_), .Y(new_new_n1089_));
  NA4        g1067(.A(new_new_n1089_), .B(new_new_n1042_), .C(new_new_n969_), .D(new_new_n884_), .Y(men4));
  INV        g1068(.A(new_new_n720_), .Y(new_new_n1093_));
  INV        g1069(.A(i_2_), .Y(new_new_n1094_));
  INV        g1070(.A(i_5_), .Y(new_new_n1095_));
  INV        g1071(.A(new_new_n500_), .Y(new_new_n1096_));
  INV        g1072(.A(i_3_), .Y(new_new_n1097_));
  INV        g1073(.A(i_6_), .Y(new_new_n1098_));
  INV        g1074(.A(i_1_), .Y(new_new_n1099_));
  INV        g1075(.A(i_4_), .Y(new_new_n1100_));
  INV        g1076(.A(new_new_n369_), .Y(new_new_n1101_));
  INV        g1077(.A(new_new_n139_), .Y(new_new_n1102_));
  INV        g1078(.A(new_new_n833_), .Y(new_new_n1103_));
  INV        g1079(.A(new_new_n196_), .Y(new_new_n1104_));
  INV        g1080(.A(new_new_n109_), .Y(new_new_n1105_));
endmodule


