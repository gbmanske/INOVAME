library verilog;
use verilog.vl_types.all;
entity tb_ex4 is
end tb_ex4;
