// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n126_, new_new_n127_,
    new_new_n128_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n640_, new_new_n641_, new_new_n642_,
    new_new_n643_, new_new_n644_, new_new_n645_, new_new_n646_,
    new_new_n647_, new_new_n648_, new_new_n649_, new_new_n650_,
    new_new_n651_, new_new_n652_, new_new_n653_, new_new_n654_,
    new_new_n655_, new_new_n656_, new_new_n657_, new_new_n658_,
    new_new_n659_, new_new_n660_, new_new_n661_, new_new_n662_,
    new_new_n663_, new_new_n664_, new_new_n665_, new_new_n666_,
    new_new_n667_, new_new_n668_, new_new_n669_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n679_,
    new_new_n680_, new_new_n681_, new_new_n682_, new_new_n683_,
    new_new_n684_, new_new_n685_, new_new_n686_, new_new_n687_,
    new_new_n688_, new_new_n689_, new_new_n690_, new_new_n691_,
    new_new_n692_, new_new_n693_, new_new_n694_, new_new_n695_,
    new_new_n696_, new_new_n697_, new_new_n698_, new_new_n699_,
    new_new_n700_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n712_, new_new_n713_, new_new_n714_, new_new_n715_,
    new_new_n716_, new_new_n717_, new_new_n718_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n901_, new_new_n902_, new_new_n903_,
    new_new_n904_, new_new_n905_, new_new_n906_, new_new_n907_,
    new_new_n908_, new_new_n909_, new_new_n910_, new_new_n911_,
    new_new_n912_, new_new_n913_, new_new_n914_, new_new_n915_,
    new_new_n916_, new_new_n917_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NO3        g015(.A(i_11_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NA2        g026(.A(i_0_), .B(i_2_), .Y(new_new_n49_));
  NA2        g027(.A(i_7_), .B(i_9_), .Y(new_new_n50_));
  NA3        g028(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n51_));
  NO2        g029(.A(i_1_), .B(i_6_), .Y(new_new_n52_));
  NA2        g030(.A(i_8_), .B(i_7_), .Y(new_new_n53_));
  OAI210     g031(.A0(new_new_n53_), .A1(new_new_n52_), .B0(new_new_n51_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n54_), .B(i_12_), .Y(new_new_n55_));
  NAi21      g033(.An(i_2_), .B(i_7_), .Y(new_new_n56_));
  INV        g034(.A(i_1_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_6_), .Y(new_new_n58_));
  NA3        g036(.A(new_new_n58_), .B(new_new_n56_), .C(new_new_n31_), .Y(new_new_n59_));
  NA2        g037(.A(i_1_), .B(i_10_), .Y(new_new_n60_));
  NO2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NAi31      g039(.An(new_new_n61_), .B(new_new_n59_), .C(new_new_n55_), .Y(new_new_n62_));
  AOI210     g040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_6_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(new_new_n25_), .Y(new_new_n65_));
  INV        g043(.A(i_0_), .Y(new_new_n66_));
  NAi21      g044(.An(i_5_), .B(i_10_), .Y(new_new_n67_));
  NA2        g045(.A(i_5_), .B(i_9_), .Y(new_new_n68_));
  AOI210     g046(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n66_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n65_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n69_), .A1(new_new_n62_), .B0(i_0_), .Y(new_new_n71_));
  NA2        g049(.A(i_12_), .B(i_5_), .Y(new_new_n72_));
  NA2        g050(.A(i_2_), .B(i_8_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n52_), .Y(new_new_n74_));
  NO2        g052(.A(i_3_), .B(i_9_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_7_), .Y(new_new_n76_));
  INV        g054(.A(i_6_), .Y(new_new_n77_));
  OR4        g055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n78_));
  INV        g056(.A(new_new_n78_), .Y(new_new_n79_));
  NO2        g057(.A(i_2_), .B(i_7_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n74_), .Y(new_new_n81_));
  NAi21      g059(.An(i_6_), .B(i_10_), .Y(new_new_n82_));
  NA2        g060(.A(i_6_), .B(i_9_), .Y(new_new_n83_));
  AOI210     g061(.A0(new_new_n83_), .A1(new_new_n82_), .B0(new_new_n57_), .Y(new_new_n84_));
  NA2        g062(.A(i_2_), .B(i_6_), .Y(new_new_n85_));
  INV        g063(.A(new_new_n84_), .Y(new_new_n86_));
  AOI210     g064(.A0(new_new_n86_), .A1(new_new_n81_), .B0(new_new_n72_), .Y(new_new_n87_));
  AN3        g065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_11_), .Y(new_new_n89_));
  NO2        g067(.A(i_5_), .B(i_8_), .Y(new_new_n90_));
  NOi21      g068(.An(new_new_n90_), .B(new_new_n89_), .Y(new_new_n91_));
  AOI220     g069(.A0(new_new_n91_), .A1(new_new_n56_), .B0(new_new_n88_), .B1(new_new_n32_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n46_), .B(new_new_n93_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NA2        g073(.A(i_12_), .B(i_3_), .Y(new_new_n96_));
  INV        g074(.A(new_new_n96_), .Y(new_new_n97_));
  NA3        g075(.A(new_new_n97_), .B(i_6_), .C(new_new_n94_), .Y(new_new_n98_));
  NAi21      g076(.An(i_7_), .B(i_11_), .Y(new_new_n99_));
  NO3        g077(.A(new_new_n99_), .B(new_new_n82_), .C(new_new_n49_), .Y(new_new_n100_));
  AN2        g078(.A(i_2_), .B(i_10_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(i_7_), .Y(new_new_n102_));
  OR2        g080(.A(new_new_n72_), .B(new_new_n52_), .Y(new_new_n103_));
  NO2        g081(.A(i_8_), .B(new_new_n93_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n103_), .C(new_new_n102_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_7_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n57_), .B(new_new_n26_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n107_), .B(i_0_), .Y(new_new_n108_));
  NA2        g086(.A(i_11_), .B(i_12_), .Y(new_new_n109_));
  OAI210     g087(.A0(new_new_n108_), .A1(new_new_n106_), .B0(new_new_n109_), .Y(new_new_n110_));
  NO2        g088(.A(new_new_n110_), .B(new_new_n105_), .Y(new_new_n111_));
  NAi41      g089(.An(new_new_n100_), .B(new_new_n111_), .C(new_new_n98_), .D(new_new_n92_), .Y(new_new_n112_));
  NOi21      g090(.An(i_1_), .B(i_5_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n113_), .B(i_11_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n115_));
  NA2        g093(.A(i_7_), .B(new_new_n25_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(new_new_n115_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n83_), .B(new_new_n82_), .Y(new_new_n118_));
  NAi21      g096(.An(i_3_), .B(i_8_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n56_), .Y(new_new_n120_));
  NOi21      g098(.An(new_new_n120_), .B(new_new_n118_), .Y(new_new_n121_));
  NO2        g099(.A(i_1_), .B(new_new_n77_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n121_), .B(new_new_n114_), .Y(new_new_n123_));
  NO3        g101(.A(new_new_n123_), .B(new_new_n112_), .C(new_new_n87_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(new_new_n71_), .Y(mai2));
  NO2        g103(.A(new_new_n57_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g104(.A(i_6_), .B(new_new_n25_), .Y(new_new_n127_));
  INV        g105(.A(new_new_n126_), .Y(new_new_n128_));
  NA3        g106(.A(new_new_n128_), .B(new_new_n70_), .C(new_new_n30_), .Y(mai0));
  AN2        g107(.A(i_8_), .B(i_7_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(i_6_), .Y(new_new_n131_));
  NO2        g109(.A(i_12_), .B(i_13_), .Y(new_new_n132_));
  NAi21      g110(.An(i_5_), .B(i_11_), .Y(new_new_n133_));
  NOi21      g111(.An(new_new_n132_), .B(new_new_n133_), .Y(new_new_n134_));
  NO2        g112(.A(i_0_), .B(i_1_), .Y(new_new_n135_));
  NA2        g113(.A(i_2_), .B(i_3_), .Y(new_new_n136_));
  NO2        g114(.A(new_new_n136_), .B(i_4_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n137_), .B(new_new_n134_), .Y(new_new_n138_));
  NA2        g116(.A(i_1_), .B(i_5_), .Y(new_new_n139_));
  NO3        g117(.A(i_4_), .B(new_new_n139_), .C(new_new_n26_), .Y(new_new_n140_));
  OR2        g118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NO3        g119(.A(new_new_n141_), .B(new_new_n72_), .C(i_13_), .Y(new_new_n142_));
  NAi32      g120(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n143_));
  NAi21      g121(.An(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NOi21      g122(.An(i_4_), .B(i_10_), .Y(new_new_n145_));
  NA2        g123(.A(new_new_n145_), .B(new_new_n39_), .Y(new_new_n146_));
  NO2        g124(.A(i_3_), .B(i_5_), .Y(new_new_n147_));
  NO3        g125(.A(new_new_n66_), .B(i_2_), .C(i_1_), .Y(new_new_n148_));
  NO2        g126(.A(new_new_n913_), .B(new_new_n140_), .Y(new_new_n149_));
  AOI210     g127(.A0(new_new_n149_), .A1(new_new_n138_), .B0(new_new_n131_), .Y(new_new_n150_));
  NA3        g128(.A(new_new_n66_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n151_));
  NOi21      g129(.An(i_4_), .B(i_9_), .Y(new_new_n152_));
  NOi21      g130(.An(i_11_), .B(i_13_), .Y(new_new_n153_));
  NA2        g131(.A(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  BUFFER     g132(.A(new_new_n154_), .Y(new_new_n155_));
  NO2        g133(.A(i_4_), .B(i_5_), .Y(new_new_n156_));
  NAi21      g134(.An(i_12_), .B(i_11_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(i_13_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n156_), .Y(new_new_n159_));
  AOI210     g137(.A0(new_new_n159_), .A1(new_new_n155_), .B0(new_new_n151_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n66_), .B(new_new_n57_), .Y(new_new_n161_));
  NA2        g139(.A(new_new_n36_), .B(i_5_), .Y(new_new_n162_));
  NAi31      g140(.An(new_new_n162_), .B(new_new_n75_), .C(i_11_), .Y(new_new_n163_));
  NA2        g141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  OR2        g142(.A(new_new_n164_), .B(new_new_n154_), .Y(new_new_n165_));
  AOI210     g143(.A0(new_new_n165_), .A1(new_new_n163_), .B0(new_new_n57_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n66_), .B(i_5_), .Y(new_new_n167_));
  NO2        g145(.A(i_13_), .B(i_10_), .Y(new_new_n168_));
  NA3        g146(.A(new_new_n168_), .B(new_new_n167_), .C(new_new_n44_), .Y(new_new_n169_));
  NO2        g147(.A(i_2_), .B(i_1_), .Y(new_new_n170_));
  NAi21      g148(.An(i_4_), .B(i_12_), .Y(new_new_n171_));
  NO3        g149(.A(new_new_n171_), .B(new_new_n909_), .C(new_new_n169_), .Y(new_new_n172_));
  NO3        g150(.A(new_new_n172_), .B(new_new_n166_), .C(new_new_n160_), .Y(new_new_n173_));
  INV        g151(.A(i_8_), .Y(new_new_n174_));
  NA2        g152(.A(i_8_), .B(i_6_), .Y(new_new_n175_));
  NO3        g153(.A(i_3_), .B(new_new_n77_), .C(new_new_n48_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n176_), .B(new_new_n104_), .Y(new_new_n177_));
  NO3        g155(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n178_));
  NA3        g156(.A(new_new_n178_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n179_));
  NO3        g157(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n180_));
  AOI210     g158(.A0(i_9_), .A1(new_new_n179_), .B0(new_new_n177_), .Y(new_new_n181_));
  NO2        g159(.A(i_3_), .B(i_8_), .Y(new_new_n182_));
  NO3        g160(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n183_));
  NA3        g161(.A(new_new_n183_), .B(new_new_n182_), .C(new_new_n39_), .Y(new_new_n184_));
  NO2        g162(.A(i_13_), .B(i_9_), .Y(new_new_n185_));
  NAi21      g163(.An(i_12_), .B(i_3_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n44_), .B(i_5_), .Y(new_new_n187_));
  NO3        g165(.A(i_0_), .B(i_2_), .C(new_new_n57_), .Y(new_new_n188_));
  NA3        g166(.A(new_new_n188_), .B(new_new_n187_), .C(i_10_), .Y(new_new_n189_));
  OAI220     g167(.A0(new_new_n189_), .A1(i_13_), .B0(new_new_n52_), .B1(new_new_n184_), .Y(new_new_n190_));
  AOI210     g168(.A0(new_new_n190_), .A1(i_7_), .B0(new_new_n181_), .Y(new_new_n191_));
  OAI220     g169(.A0(new_new_n191_), .A1(i_4_), .B0(new_new_n175_), .B1(new_new_n173_), .Y(new_new_n192_));
  NAi21      g170(.An(i_12_), .B(i_7_), .Y(new_new_n193_));
  NA3        g171(.A(i_13_), .B(new_new_n174_), .C(i_10_), .Y(new_new_n194_));
  NA2        g172(.A(i_0_), .B(i_5_), .Y(new_new_n195_));
  NAi31      g173(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n36_), .B(i_13_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n66_), .B(new_new_n26_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n46_), .B(new_new_n57_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(new_new_n198_), .C(new_new_n197_), .Y(new_new_n200_));
  INV        g178(.A(i_13_), .Y(new_new_n201_));
  NO2        g179(.A(i_12_), .B(new_new_n201_), .Y(new_new_n202_));
  NA2        g180(.A(new_new_n914_), .B(new_new_n130_), .Y(new_new_n203_));
  NO2        g181(.A(i_12_), .B(new_new_n37_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n164_), .B(i_4_), .Y(new_new_n205_));
  NA2        g183(.A(new_new_n205_), .B(new_new_n204_), .Y(new_new_n206_));
  OR2        g184(.A(i_8_), .B(i_7_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n49_), .B(i_1_), .Y(new_new_n208_));
  INV        g186(.A(i_12_), .Y(new_new_n209_));
  NO3        g187(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n210_));
  NA2        g188(.A(i_2_), .B(i_1_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n49_), .B(new_new_n206_), .Y(new_new_n212_));
  NO3        g190(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n213_));
  NAi21      g191(.An(i_4_), .B(i_3_), .Y(new_new_n214_));
  NO2        g192(.A(i_0_), .B(i_6_), .Y(new_new_n215_));
  NOi41      g193(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  AOI210     g195(.A0(new_new_n905_), .A1(new_new_n39_), .B0(new_new_n212_), .Y(new_new_n218_));
  NO2        g196(.A(i_11_), .B(new_new_n201_), .Y(new_new_n219_));
  NOi21      g197(.An(i_1_), .B(i_6_), .Y(new_new_n220_));
  NAi21      g198(.An(i_3_), .B(i_7_), .Y(new_new_n221_));
  NO2        g199(.A(i_12_), .B(i_3_), .Y(new_new_n222_));
  NA2        g200(.A(new_new_n66_), .B(i_5_), .Y(new_new_n223_));
  NA2        g201(.A(i_3_), .B(i_9_), .Y(new_new_n224_));
  NA3        g202(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n917_), .B(new_new_n68_), .Y(new_new_n226_));
  NA2        g204(.A(new_new_n226_), .B(new_new_n130_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n207_), .B(new_new_n37_), .Y(new_new_n228_));
  NA2        g206(.A(i_12_), .B(i_6_), .Y(new_new_n229_));
  OR2        g207(.A(i_13_), .B(i_9_), .Y(new_new_n230_));
  NO3        g208(.A(new_new_n230_), .B(new_new_n229_), .C(new_new_n48_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n214_), .B(i_2_), .Y(new_new_n232_));
  NA3        g210(.A(new_new_n232_), .B(new_new_n231_), .C(new_new_n44_), .Y(new_new_n233_));
  NA2        g211(.A(new_new_n219_), .B(i_9_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n223_), .B(new_new_n58_), .Y(new_new_n235_));
  OAI210     g213(.A0(new_new_n235_), .A1(new_new_n234_), .B0(new_new_n233_), .Y(new_new_n236_));
  NO2        g214(.A(i_11_), .B(new_new_n201_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n221_), .B(i_8_), .Y(new_new_n238_));
  NO2        g216(.A(i_6_), .B(new_new_n48_), .Y(new_new_n239_));
  NA3        g217(.A(i_3_), .B(new_new_n228_), .C(new_new_n202_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n240_), .B(new_new_n908_), .Y(new_new_n241_));
  AOI210     g219(.A0(new_new_n236_), .A1(new_new_n228_), .B0(new_new_n241_), .Y(new_new_n242_));
  NA4        g220(.A(new_new_n242_), .B(new_new_n227_), .C(new_new_n218_), .D(new_new_n203_), .Y(new_new_n243_));
  NO3        g221(.A(i_12_), .B(new_new_n201_), .C(new_new_n37_), .Y(new_new_n244_));
  INV        g222(.A(new_new_n244_), .Y(new_new_n245_));
  NA2        g223(.A(i_8_), .B(new_new_n93_), .Y(new_new_n246_));
  NO3        g224(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n211_), .B(i_0_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n239_), .B(new_new_n26_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n249_), .B(new_new_n906_), .Y(new_new_n250_));
  NA2        g228(.A(i_0_), .B(i_1_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n251_), .B(i_2_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n53_), .B(i_6_), .Y(new_new_n253_));
  NA3        g231(.A(new_new_n253_), .B(new_new_n252_), .C(new_new_n147_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n131_), .B(new_new_n254_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n255_), .B(new_new_n250_), .Y(new_new_n256_));
  NO2        g234(.A(i_3_), .B(i_10_), .Y(new_new_n257_));
  NA3        g235(.A(new_new_n257_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n258_));
  NO2        g236(.A(i_2_), .B(new_new_n93_), .Y(new_new_n259_));
  NA2        g237(.A(i_1_), .B(new_new_n36_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n260_), .B(i_8_), .Y(new_new_n261_));
  INV        g239(.A(new_new_n261_), .Y(new_new_n262_));
  AN2        g240(.A(i_3_), .B(i_10_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n263_), .B(new_new_n158_), .C(new_new_n156_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n265_));
  OR2        g243(.A(new_new_n262_), .B(new_new_n258_), .Y(new_new_n266_));
  OAI220     g244(.A0(new_new_n266_), .A1(i_6_), .B0(new_new_n256_), .B1(new_new_n245_), .Y(new_new_n267_));
  NO4        g245(.A(new_new_n267_), .B(new_new_n243_), .C(new_new_n192_), .D(new_new_n150_), .Y(new_new_n268_));
  NO3        g246(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n53_), .B(new_new_n77_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n248_), .B(new_new_n270_), .Y(new_new_n271_));
  NO3        g249(.A(i_6_), .B(new_new_n174_), .C(i_7_), .Y(new_new_n272_));
  NA2        g250(.A(new_new_n912_), .B(new_new_n271_), .Y(new_new_n273_));
  NO2        g251(.A(i_2_), .B(i_3_), .Y(new_new_n274_));
  OR2        g252(.A(i_0_), .B(i_5_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n195_), .B(new_new_n275_), .Y(new_new_n276_));
  NA4        g254(.A(new_new_n276_), .B(i_6_), .C(new_new_n274_), .D(i_1_), .Y(new_new_n277_));
  NA2        g255(.A(new_new_n248_), .B(new_new_n147_), .Y(new_new_n278_));
  NAi21      g256(.An(i_8_), .B(i_7_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(i_6_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n141_), .B(new_new_n46_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n281_), .B(new_new_n280_), .Y(new_new_n282_));
  NA3        g260(.A(new_new_n282_), .B(new_new_n278_), .C(new_new_n277_), .Y(new_new_n283_));
  OAI210     g261(.A0(new_new_n283_), .A1(new_new_n273_), .B0(i_4_), .Y(new_new_n284_));
  NO2        g262(.A(i_12_), .B(i_10_), .Y(new_new_n285_));
  NOi21      g263(.An(i_5_), .B(i_0_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n260_), .B(new_new_n119_), .Y(new_new_n287_));
  NA4        g265(.A(new_new_n76_), .B(new_new_n36_), .C(new_new_n77_), .D(i_8_), .Y(new_new_n288_));
  NA2        g266(.A(new_new_n287_), .B(new_new_n285_), .Y(new_new_n289_));
  NO2        g267(.A(i_6_), .B(i_8_), .Y(new_new_n290_));
  NOi21      g268(.An(i_0_), .B(i_2_), .Y(new_new_n291_));
  AN2        g269(.A(new_new_n291_), .B(new_new_n290_), .Y(new_new_n292_));
  NO2        g270(.A(i_1_), .B(i_7_), .Y(new_new_n293_));
  AO220      g271(.A0(new_new_n293_), .A1(new_new_n292_), .B0(new_new_n280_), .B1(new_new_n208_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n294_), .B(new_new_n41_), .Y(new_new_n295_));
  NA3        g273(.A(new_new_n295_), .B(new_new_n289_), .C(new_new_n284_), .Y(new_new_n296_));
  NO3        g274(.A(new_new_n207_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n297_));
  NO3        g275(.A(new_new_n279_), .B(i_2_), .C(i_1_), .Y(new_new_n298_));
  OAI210     g276(.A0(new_new_n298_), .A1(new_new_n297_), .B0(i_6_), .Y(new_new_n299_));
  NA2        g277(.A(new_new_n259_), .B(new_new_n174_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n300_), .B(new_new_n299_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n301_), .B(i_3_), .Y(new_new_n302_));
  INV        g280(.A(new_new_n76_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n85_), .B(new_new_n174_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n73_), .B(new_new_n303_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n174_), .B(i_9_), .Y(new_new_n306_));
  INV        g284(.A(new_new_n306_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n305_), .B(new_new_n250_), .Y(new_new_n308_));
  AOI210     g286(.A0(new_new_n308_), .A1(new_new_n302_), .B0(new_new_n146_), .Y(new_new_n309_));
  AOI210     g287(.A0(new_new_n296_), .A1(new_new_n269_), .B0(new_new_n309_), .Y(new_new_n310_));
  NOi32      g288(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n311_));
  INV        g289(.A(new_new_n311_), .Y(new_new_n312_));
  NAi21      g290(.An(i_0_), .B(i_6_), .Y(new_new_n313_));
  NAi21      g291(.An(i_1_), .B(i_5_), .Y(new_new_n314_));
  NA2        g292(.A(new_new_n314_), .B(new_new_n313_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n315_), .B(new_new_n25_), .Y(new_new_n316_));
  OAI210     g294(.A0(new_new_n316_), .A1(new_new_n143_), .B0(new_new_n217_), .Y(new_new_n317_));
  NAi41      g295(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n318_));
  OAI220     g296(.A0(new_new_n318_), .A1(new_new_n314_), .B0(new_new_n196_), .B1(new_new_n143_), .Y(new_new_n319_));
  AOI210     g297(.A0(new_new_n318_), .A1(new_new_n143_), .B0(new_new_n141_), .Y(new_new_n320_));
  NOi32      g298(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n321_));
  NAi21      g299(.An(i_6_), .B(i_1_), .Y(new_new_n322_));
  NA3        g300(.A(new_new_n322_), .B(new_new_n321_), .C(new_new_n46_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n323_), .B(i_0_), .Y(new_new_n324_));
  OR3        g302(.A(new_new_n324_), .B(new_new_n320_), .C(new_new_n319_), .Y(new_new_n325_));
  NO2        g303(.A(i_1_), .B(new_new_n93_), .Y(new_new_n326_));
  NAi21      g304(.An(i_3_), .B(i_4_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(i_9_), .Y(new_new_n328_));
  AN2        g306(.A(i_6_), .B(i_7_), .Y(new_new_n329_));
  NA2        g307(.A(i_2_), .B(i_7_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n327_), .B(i_10_), .Y(new_new_n331_));
  NA3        g309(.A(new_new_n331_), .B(new_new_n330_), .C(new_new_n215_), .Y(new_new_n332_));
  INV        g310(.A(new_new_n332_), .Y(new_new_n333_));
  AOI210     g311(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n334_));
  OAI210     g312(.A0(new_new_n334_), .A1(new_new_n170_), .B0(new_new_n331_), .Y(new_new_n335_));
  AOI220     g313(.A0(new_new_n331_), .A1(new_new_n293_), .B0(new_new_n210_), .B1(new_new_n170_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n336_), .A1(new_new_n335_), .B0(i_5_), .Y(new_new_n337_));
  NO4        g315(.A(new_new_n337_), .B(new_new_n333_), .C(new_new_n325_), .D(new_new_n317_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n338_), .B(new_new_n312_), .Y(new_new_n339_));
  INV        g317(.A(new_new_n53_), .Y(new_new_n340_));
  AN2        g318(.A(i_12_), .B(i_5_), .Y(new_new_n341_));
  NO2        g319(.A(i_4_), .B(new_new_n26_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NO2        g321(.A(i_11_), .B(i_6_), .Y(new_new_n344_));
  INV        g322(.A(new_new_n343_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n214_), .B(i_5_), .Y(new_new_n346_));
  NO2        g324(.A(i_5_), .B(i_10_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n132_), .B(new_new_n45_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n214_), .Y(new_new_n349_));
  OAI210     g327(.A0(new_new_n349_), .A1(new_new_n345_), .B0(new_new_n340_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n351_));
  NO3        g329(.A(new_new_n77_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n347_), .B(new_new_n209_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n41_), .B(i_11_), .Y(new_new_n354_));
  OAI220     g332(.A0(new_new_n354_), .A1(new_new_n196_), .B0(new_new_n353_), .B1(new_new_n288_), .Y(new_new_n355_));
  NAi21      g333(.An(i_13_), .B(i_0_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n355_), .B(i_0_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n357_), .B(new_new_n350_), .Y(new_new_n358_));
  NO2        g336(.A(i_0_), .B(i_11_), .Y(new_new_n359_));
  NOi21      g337(.An(i_2_), .B(i_12_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n130_), .B(i_9_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(i_4_), .Y(new_new_n362_));
  OR2        g340(.A(i_13_), .B(i_10_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n154_), .B(new_new_n115_), .Y(new_new_n364_));
  OR2        g342(.A(new_new_n194_), .B(new_new_n193_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n365_), .B(new_new_n26_), .Y(new_new_n367_));
  INV        g345(.A(new_new_n277_), .Y(new_new_n368_));
  AOI220     g346(.A0(new_new_n253_), .A1(new_new_n247_), .B0(new_new_n248_), .B1(new_new_n270_), .Y(new_new_n369_));
  INV        g347(.A(new_new_n369_), .Y(new_new_n370_));
  NO2        g348(.A(i_2_), .B(new_new_n246_), .Y(new_new_n371_));
  NO3        g349(.A(new_new_n371_), .B(new_new_n370_), .C(new_new_n368_), .Y(new_new_n372_));
  NO2        g350(.A(i_3_), .B(new_new_n279_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n253_), .B(new_new_n208_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n292_), .B(new_new_n373_), .Y(new_new_n375_));
  AOI210     g353(.A0(new_new_n375_), .A1(new_new_n372_), .B0(new_new_n234_), .Y(new_new_n376_));
  NO4        g354(.A(new_new_n376_), .B(new_new_n367_), .C(new_new_n358_), .D(new_new_n339_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n57_), .B(i_4_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n378_), .B(i_2_), .Y(new_new_n379_));
  NO2        g357(.A(i_10_), .B(i_9_), .Y(new_new_n380_));
  NAi21      g358(.An(i_12_), .B(i_8_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n381_), .B(i_3_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n382_), .B(new_new_n380_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n46_), .B(i_4_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n384_), .B(i_6_), .Y(new_new_n385_));
  OAI220     g363(.A0(new_new_n385_), .A1(new_new_n184_), .B0(new_new_n383_), .B1(new_new_n379_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n265_), .B(i_0_), .Y(new_new_n387_));
  NO3        g365(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n229_), .B(new_new_n89_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n389_), .B(new_new_n388_), .Y(new_new_n390_));
  NA2        g368(.A(i_8_), .B(i_9_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n390_), .B(new_new_n387_), .Y(new_new_n392_));
  NO3        g370(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n393_));
  NA3        g371(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n392_), .B(new_new_n386_), .Y(new_new_n395_));
  OR2        g373(.A(new_new_n251_), .B(i_13_), .Y(new_new_n396_));
  OA210      g374(.A0(new_new_n307_), .A1(new_new_n93_), .B0(new_new_n254_), .Y(new_new_n397_));
  OA220      g375(.A0(new_new_n397_), .A1(new_new_n146_), .B0(new_new_n396_), .B1(new_new_n206_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n88_), .B(i_13_), .Y(new_new_n399_));
  NO2        g377(.A(i_2_), .B(i_13_), .Y(new_new_n400_));
  NA3        g378(.A(new_new_n400_), .B(new_new_n145_), .C(new_new_n91_), .Y(new_new_n401_));
  NO3        g379(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n402_));
  NO2        g380(.A(i_6_), .B(i_7_), .Y(new_new_n403_));
  NO2        g381(.A(i_11_), .B(i_1_), .Y(new_new_n404_));
  OR2        g382(.A(i_11_), .B(i_8_), .Y(new_new_n405_));
  NOi21      g383(.An(i_2_), .B(i_7_), .Y(new_new_n406_));
  NAi21      g384(.An(new_new_n405_), .B(new_new_n406_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n363_), .B(i_6_), .Y(new_new_n408_));
  NA3        g386(.A(new_new_n408_), .B(new_new_n378_), .C(new_new_n68_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n407_), .Y(new_new_n410_));
  NO2        g388(.A(i_3_), .B(new_new_n174_), .Y(new_new_n411_));
  NO2        g389(.A(i_6_), .B(i_10_), .Y(new_new_n412_));
  NA3        g390(.A(new_new_n412_), .B(new_new_n269_), .C(new_new_n411_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n413_), .B(i_4_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n141_), .B(i_3_), .Y(new_new_n415_));
  NA3        g393(.A(new_new_n351_), .B(new_new_n161_), .C(new_new_n137_), .Y(new_new_n416_));
  INV        g394(.A(new_new_n416_), .Y(new_new_n417_));
  NO3        g395(.A(new_new_n417_), .B(new_new_n414_), .C(new_new_n410_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n393_), .B(new_new_n347_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n419_), .B(new_new_n200_), .Y(new_new_n420_));
  NO2        g398(.A(i_0_), .B(new_new_n77_), .Y(new_new_n421_));
  NA3        g399(.A(new_new_n421_), .B(new_new_n907_), .C(new_new_n130_), .Y(new_new_n422_));
  OR3        g400(.A(new_new_n260_), .B(i_11_), .C(new_new_n46_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n423_), .B(new_new_n422_), .Y(new_new_n424_));
  NA3        g402(.A(new_new_n263_), .B(new_new_n199_), .C(new_new_n66_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(i_4_), .Y(new_new_n426_));
  NO3        g404(.A(new_new_n426_), .B(new_new_n424_), .C(new_new_n420_), .Y(new_new_n427_));
  NA4        g405(.A(new_new_n427_), .B(new_new_n418_), .C(new_new_n398_), .D(new_new_n395_), .Y(new_new_n428_));
  NA3        g406(.A(new_new_n263_), .B(new_new_n158_), .C(new_new_n156_), .Y(new_new_n429_));
  INV        g407(.A(new_new_n429_), .Y(new_new_n430_));
  BUFFER     g408(.A(new_new_n247_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n431_), .B(new_new_n430_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n114_), .B(new_new_n103_), .Y(new_new_n433_));
  AN2        g411(.A(new_new_n433_), .B(new_new_n388_), .Y(new_new_n434_));
  OAI210     g412(.A0(new_new_n44_), .A1(new_new_n206_), .B0(new_new_n264_), .Y(new_new_n435_));
  AOI220     g413(.A0(new_new_n435_), .A1(new_new_n280_), .B0(new_new_n434_), .B1(new_new_n265_), .Y(new_new_n436_));
  NA3        g414(.A(new_new_n378_), .B(new_new_n182_), .C(i_2_), .Y(new_new_n437_));
  INV        g415(.A(new_new_n437_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n311_), .B(new_new_n66_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n329_), .B(new_new_n321_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n36_), .B(i_8_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n38_), .B(i_13_), .Y(new_new_n442_));
  INV        g420(.A(new_new_n442_), .Y(new_new_n443_));
  AOI210     g421(.A0(new_new_n438_), .A1(new_new_n183_), .B0(new_new_n443_), .Y(new_new_n444_));
  NO2        g422(.A(i_7_), .B(new_new_n179_), .Y(new_new_n445_));
  OR2        g423(.A(new_new_n164_), .B(i_4_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n446_), .B(new_new_n77_), .Y(new_new_n447_));
  AOI220     g425(.A0(new_new_n447_), .A1(new_new_n445_), .B0(new_new_n223_), .B1(new_new_n364_), .Y(new_new_n448_));
  NA4        g426(.A(new_new_n448_), .B(new_new_n444_), .C(new_new_n436_), .D(new_new_n432_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n346_), .B(new_new_n252_), .Y(new_new_n450_));
  OAI210     g428(.A0(new_new_n343_), .A1(new_new_n151_), .B0(new_new_n450_), .Y(new_new_n451_));
  NO2        g429(.A(i_12_), .B(new_new_n174_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n452_), .B(new_new_n201_), .Y(new_new_n453_));
  NO2        g431(.A(i_6_), .B(new_new_n453_), .Y(new_new_n454_));
  NOi21      g432(.An(new_new_n272_), .B(i_11_), .Y(new_new_n455_));
  OAI210     g433(.A0(new_new_n455_), .A1(new_new_n454_), .B0(new_new_n451_), .Y(new_new_n456_));
  NO2        g434(.A(i_8_), .B(i_7_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n46_), .B(new_new_n446_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n915_), .B(i_6_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n459_), .B(new_new_n458_), .Y(new_new_n460_));
  INV        g438(.A(new_new_n399_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n461_), .B(new_new_n228_), .Y(new_new_n462_));
  NA3        g440(.A(new_new_n263_), .B(new_new_n156_), .C(new_new_n88_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n197_), .B(new_new_n44_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n141_), .B(i_5_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n465_), .B(new_new_n274_), .Y(new_new_n466_));
  OAI210     g444(.A0(new_new_n466_), .A1(new_new_n464_), .B0(new_new_n463_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n467_), .B(new_new_n393_), .Y(new_new_n468_));
  NA4        g446(.A(new_new_n468_), .B(new_new_n462_), .C(new_new_n460_), .D(new_new_n456_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n244_), .B(new_new_n76_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n73_), .B(new_new_n470_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n253_), .B(new_new_n247_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n155_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n199_), .B(new_new_n198_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n380_), .B(new_new_n197_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n474_), .B(new_new_n475_), .Y(new_new_n476_));
  AOI210     g454(.A0(new_new_n322_), .A1(new_new_n46_), .B0(new_new_n326_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n452_), .B(new_new_n237_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n477_), .B(new_new_n478_), .Y(new_new_n479_));
  NO4        g457(.A(new_new_n479_), .B(new_new_n476_), .C(new_new_n473_), .D(new_new_n471_), .Y(new_new_n480_));
  NO4        g458(.A(new_new_n220_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n481_));
  NO3        g459(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n482_));
  NO2        g460(.A(new_new_n207_), .B(new_new_n36_), .Y(new_new_n483_));
  AN2        g461(.A(new_new_n483_), .B(new_new_n482_), .Y(new_new_n484_));
  OA210      g462(.A0(new_new_n484_), .A1(new_new_n481_), .B0(new_new_n311_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n363_), .B(i_1_), .Y(new_new_n486_));
  NOi31      g464(.An(new_new_n486_), .B(new_new_n389_), .C(new_new_n66_), .Y(new_new_n487_));
  AN2        g465(.A(new_new_n487_), .B(new_new_n362_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n369_), .B(new_new_n159_), .Y(new_new_n489_));
  NO3        g467(.A(new_new_n489_), .B(new_new_n488_), .C(new_new_n485_), .Y(new_new_n490_));
  NOi21      g468(.An(i_10_), .B(i_6_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n77_), .B(new_new_n25_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n237_), .B(new_new_n491_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n493_), .B(new_new_n387_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n106_), .B(new_new_n23_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n272_), .B(new_new_n148_), .Y(new_new_n496_));
  AOI220     g474(.A0(new_new_n496_), .A1(new_new_n374_), .B0(new_new_n165_), .B1(new_new_n163_), .Y(new_new_n497_));
  NOi21      g475(.An(new_new_n134_), .B(new_new_n288_), .Y(new_new_n498_));
  NO3        g476(.A(new_new_n498_), .B(new_new_n497_), .C(new_new_n494_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n439_), .B(new_new_n336_), .Y(new_new_n500_));
  INV        g478(.A(new_new_n274_), .Y(new_new_n501_));
  NO2        g479(.A(i_12_), .B(new_new_n77_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n502_), .B(new_new_n237_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(new_new_n501_), .Y(new_new_n504_));
  NO3        g482(.A(i_4_), .B(new_new_n299_), .C(new_new_n258_), .Y(new_new_n505_));
  NO3        g483(.A(new_new_n505_), .B(new_new_n504_), .C(new_new_n500_), .Y(new_new_n506_));
  NA4        g484(.A(new_new_n506_), .B(new_new_n499_), .C(new_new_n490_), .D(new_new_n480_), .Y(new_new_n507_));
  NO4        g485(.A(new_new_n507_), .B(new_new_n469_), .C(new_new_n449_), .D(new_new_n428_), .Y(new_new_n508_));
  NA4        g486(.A(new_new_n508_), .B(new_new_n377_), .C(new_new_n310_), .D(new_new_n268_), .Y(mai7));
  NO2        g487(.A(new_new_n85_), .B(new_new_n50_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n99_), .B(new_new_n82_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n342_), .B(new_new_n511_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n412_), .B(new_new_n76_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n132_), .B(i_8_), .Y(new_new_n514_));
  OAI210     g492(.A0(new_new_n514_), .A1(new_new_n513_), .B0(new_new_n512_), .Y(new_new_n515_));
  NA3        g493(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n209_), .B(i_4_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n517_), .B(i_8_), .Y(new_new_n518_));
  NA2        g496(.A(i_2_), .B(new_new_n77_), .Y(new_new_n519_));
  NO2        g497(.A(i_7_), .B(new_new_n37_), .Y(new_new_n520_));
  NA2        g498(.A(i_4_), .B(i_8_), .Y(new_new_n521_));
  AOI210     g499(.A0(new_new_n521_), .A1(new_new_n263_), .B0(new_new_n520_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n522_), .B(new_new_n519_), .Y(new_new_n523_));
  NO3        g501(.A(new_new_n523_), .B(new_new_n515_), .C(new_new_n510_), .Y(new_new_n524_));
  AOI210     g502(.A0(new_new_n119_), .A1(new_new_n56_), .B0(i_10_), .Y(new_new_n525_));
  AOI210     g503(.A0(new_new_n525_), .A1(new_new_n209_), .B0(new_new_n145_), .Y(new_new_n526_));
  OR2        g504(.A(i_6_), .B(i_10_), .Y(new_new_n527_));
  NO2        g505(.A(new_new_n527_), .B(new_new_n23_), .Y(new_new_n528_));
  OR3        g506(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n529_));
  NO3        g507(.A(new_new_n529_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n530_));
  INV        g508(.A(new_new_n180_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n530_), .B(new_new_n528_), .Y(new_new_n532_));
  OA220      g510(.A0(new_new_n532_), .A1(new_new_n501_), .B0(new_new_n526_), .B1(new_new_n230_), .Y(new_new_n533_));
  AOI210     g511(.A0(new_new_n533_), .A1(new_new_n524_), .B0(new_new_n57_), .Y(new_new_n534_));
  NOi21      g512(.An(i_11_), .B(i_7_), .Y(new_new_n535_));
  AO210      g513(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n536_), .B(new_new_n535_), .Y(new_new_n537_));
  NA3        g515(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n538_));
  NAi21      g516(.An(new_new_n538_), .B(i_11_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n539_), .B(new_new_n57_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n541_));
  AO210      g519(.A0(new_new_n541_), .A1(new_new_n336_), .B0(new_new_n40_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n360_), .B(new_new_n31_), .Y(new_new_n543_));
  OR2        g521(.A(new_new_n186_), .B(new_new_n99_), .Y(new_new_n544_));
  NA2        g522(.A(new_new_n544_), .B(new_new_n543_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n57_), .B(i_9_), .Y(new_new_n546_));
  NA2        g524(.A(new_new_n57_), .B(new_new_n545_), .Y(new_new_n547_));
  NO2        g525(.A(i_1_), .B(i_12_), .Y(new_new_n548_));
  NA2        g526(.A(new_new_n547_), .B(new_new_n542_), .Y(new_new_n549_));
  OAI210     g527(.A0(new_new_n549_), .A1(new_new_n540_), .B0(i_6_), .Y(new_new_n550_));
  NO2        g528(.A(i_6_), .B(i_11_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n390_), .Y(new_new_n552_));
  NO4        g530(.A(new_new_n193_), .B(new_new_n119_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n209_), .B(i_6_), .Y(new_new_n554_));
  NA3        g532(.A(new_new_n457_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n555_));
  NA2        g533(.A(new_new_n126_), .B(i_9_), .Y(new_new_n556_));
  NA3        g534(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n46_), .B(i_1_), .Y(new_new_n558_));
  NA3        g536(.A(new_new_n558_), .B(new_new_n229_), .C(new_new_n44_), .Y(new_new_n559_));
  OAI220     g537(.A0(new_new_n559_), .A1(new_new_n557_), .B0(new_new_n556_), .B1(new_new_n901_), .Y(new_new_n560_));
  NA3        g538(.A(new_new_n546_), .B(new_new_n274_), .C(i_6_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n561_), .B(new_new_n23_), .Y(new_new_n562_));
  AOI210     g540(.A0(new_new_n404_), .A1(new_new_n366_), .B0(new_new_n213_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n563_), .B(new_new_n519_), .Y(new_new_n564_));
  NAi21      g542(.An(new_new_n555_), .B(new_new_n84_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n558_), .B(new_new_n229_), .Y(new_new_n566_));
  NO2        g544(.A(i_11_), .B(new_new_n37_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n567_), .B(new_new_n24_), .Y(new_new_n568_));
  OAI210     g546(.A0(new_new_n568_), .A1(new_new_n566_), .B0(new_new_n565_), .Y(new_new_n569_));
  OR4        g547(.A(new_new_n569_), .B(new_new_n564_), .C(new_new_n562_), .D(new_new_n560_), .Y(new_new_n570_));
  NO3        g548(.A(new_new_n570_), .B(new_new_n553_), .C(new_new_n552_), .Y(new_new_n571_));
  NA2        g549(.A(i_3_), .B(new_new_n174_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n572_), .B(new_new_n106_), .Y(new_new_n573_));
  AN2        g551(.A(new_new_n573_), .B(new_new_n459_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n207_), .B(new_new_n44_), .Y(new_new_n575_));
  NO2        g553(.A(new_new_n77_), .B(i_9_), .Y(new_new_n576_));
  NA2        g554(.A(i_1_), .B(i_3_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n391_), .B(new_new_n85_), .Y(new_new_n578_));
  AOI210     g556(.A0(new_new_n575_), .A1(new_new_n491_), .B0(new_new_n578_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n579_), .B(new_new_n577_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n580_), .B(new_new_n574_), .Y(new_new_n581_));
  NA3        g559(.A(new_new_n581_), .B(new_new_n571_), .C(new_new_n550_), .Y(new_new_n582_));
  NO3        g560(.A(new_new_n405_), .B(i_3_), .C(i_7_), .Y(new_new_n583_));
  NOi21      g561(.An(new_new_n583_), .B(i_10_), .Y(new_new_n584_));
  OA210      g562(.A0(new_new_n584_), .A1(new_new_n216_), .B0(new_new_n77_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n329_), .B(new_new_n328_), .Y(new_new_n586_));
  NA3        g564(.A(new_new_n412_), .B(new_new_n441_), .C(new_new_n46_), .Y(new_new_n587_));
  NO3        g565(.A(new_new_n406_), .B(new_new_n521_), .C(new_new_n77_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(new_new_n25_), .Y(new_new_n589_));
  NA3        g567(.A(new_new_n145_), .B(new_new_n76_), .C(new_new_n77_), .Y(new_new_n590_));
  NA4        g568(.A(new_new_n590_), .B(new_new_n589_), .C(new_new_n587_), .D(new_new_n586_), .Y(new_new_n591_));
  OAI210     g569(.A0(new_new_n591_), .A1(new_new_n585_), .B0(i_1_), .Y(new_new_n592_));
  AOI210     g570(.A0(new_new_n229_), .A1(new_new_n89_), .B0(i_1_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n327_), .B(i_2_), .Y(new_new_n594_));
  NA2        g572(.A(new_new_n594_), .B(new_new_n593_), .Y(new_new_n595_));
  OAI210     g573(.A0(new_new_n561_), .A1(new_new_n381_), .B0(new_new_n595_), .Y(new_new_n596_));
  INV        g574(.A(new_new_n596_), .Y(new_new_n597_));
  AOI210     g575(.A0(new_new_n597_), .A1(new_new_n592_), .B0(i_13_), .Y(new_new_n598_));
  OR2        g576(.A(i_11_), .B(i_7_), .Y(new_new_n599_));
  AOI220     g577(.A0(new_new_n400_), .A1(new_new_n145_), .B0(new_new_n384_), .B1(new_new_n126_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n600_), .B(new_new_n44_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n216_), .B(new_new_n122_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n602_), .B(new_new_n40_), .Y(new_new_n603_));
  AOI210     g581(.A0(new_new_n601_), .A1(new_new_n290_), .B0(new_new_n603_), .Y(new_new_n604_));
  AOI220     g582(.A0(i_7_), .A1(new_new_n65_), .B0(new_new_n344_), .B1(new_new_n558_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n605_), .B(new_new_n214_), .Y(new_new_n606_));
  AOI210     g584(.A0(new_new_n381_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n607_));
  NOi31      g585(.An(new_new_n607_), .B(new_new_n513_), .C(new_new_n44_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n118_), .B(i_13_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n557_), .B(new_new_n106_), .Y(new_new_n610_));
  INV        g588(.A(new_new_n610_), .Y(new_new_n611_));
  OAI220     g589(.A0(new_new_n611_), .A1(new_new_n64_), .B0(new_new_n609_), .B1(new_new_n593_), .Y(new_new_n612_));
  NO3        g590(.A(new_new_n64_), .B(new_new_n32_), .C(new_new_n93_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n26_), .B(new_new_n174_), .Y(new_new_n614_));
  NA2        g592(.A(new_new_n614_), .B(i_7_), .Y(new_new_n615_));
  NO3        g593(.A(new_new_n406_), .B(new_new_n209_), .C(new_new_n77_), .Y(new_new_n616_));
  AOI210     g594(.A0(new_new_n616_), .A1(new_new_n615_), .B0(new_new_n613_), .Y(new_new_n617_));
  NA2        g595(.A(new_new_n84_), .B(new_new_n94_), .Y(new_new_n618_));
  OAI220     g596(.A0(new_new_n618_), .A1(new_new_n518_), .B0(new_new_n617_), .B1(new_new_n531_), .Y(new_new_n619_));
  NO4        g597(.A(new_new_n619_), .B(new_new_n612_), .C(new_new_n608_), .D(new_new_n606_), .Y(new_new_n620_));
  OR2        g598(.A(i_11_), .B(i_6_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n517_), .B(new_new_n614_), .C(i_7_), .Y(new_new_n622_));
  AOI210     g600(.A0(new_new_n622_), .A1(new_new_n611_), .B0(new_new_n621_), .Y(new_new_n623_));
  NA3        g601(.A(new_new_n360_), .B(new_new_n520_), .C(new_new_n89_), .Y(new_new_n624_));
  NA2        g602(.A(new_new_n551_), .B(i_13_), .Y(new_new_n625_));
  NA2        g603(.A(new_new_n94_), .B(new_new_n614_), .Y(new_new_n626_));
  NAi21      g604(.An(i_11_), .B(i_12_), .Y(new_new_n627_));
  NOi41      g605(.An(new_new_n102_), .B(new_new_n627_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n628_));
  AOI220     g606(.A0(new_new_n910_), .A1(new_new_n269_), .B0(new_new_n628_), .B1(new_new_n626_), .Y(new_new_n629_));
  NA3        g607(.A(new_new_n629_), .B(new_new_n625_), .C(new_new_n624_), .Y(new_new_n630_));
  OAI210     g608(.A0(new_new_n630_), .A1(new_new_n623_), .B0(new_new_n57_), .Y(new_new_n631_));
  NO2        g609(.A(i_2_), .B(i_12_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n209_), .B(new_new_n326_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n119_), .B(i_2_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n634_), .B(new_new_n548_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n635_), .B(new_new_n633_), .Y(new_new_n636_));
  NA3        g614(.A(new_new_n636_), .B(new_new_n45_), .C(new_new_n201_), .Y(new_new_n637_));
  NA4        g615(.A(new_new_n637_), .B(new_new_n631_), .C(new_new_n620_), .D(new_new_n604_), .Y(new_new_n638_));
  OR4        g616(.A(new_new_n638_), .B(new_new_n598_), .C(new_new_n582_), .D(new_new_n534_), .Y(mai5));
  AN2        g617(.A(new_new_n24_), .B(i_10_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n640_), .B(new_new_n632_), .Y(new_new_n641_));
  NO2        g619(.A(new_new_n518_), .B(i_11_), .Y(new_new_n642_));
  NA2        g620(.A(new_new_n80_), .B(new_new_n642_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n643_), .B(new_new_n641_), .Y(new_new_n644_));
  NO3        g622(.A(i_11_), .B(new_new_n209_), .C(i_13_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n646_));
  NA2        g624(.A(i_12_), .B(i_8_), .Y(new_new_n647_));
  INV        g625(.A(new_new_n380_), .Y(new_new_n648_));
  NA2        g626(.A(new_new_n274_), .B(new_new_n495_), .Y(new_new_n649_));
  INV        g627(.A(new_new_n649_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n650_), .B(new_new_n644_), .Y(new_new_n651_));
  INV        g629(.A(new_new_n153_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n594_), .B(new_new_n102_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n653_), .B(new_new_n652_), .Y(new_new_n654_));
  INV        g632(.A(new_new_n366_), .Y(new_new_n655_));
  NA2        g633(.A(new_new_n655_), .B(i_2_), .Y(new_new_n656_));
  INV        g634(.A(new_new_n656_), .Y(new_new_n657_));
  AOI210     g635(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n363_), .Y(new_new_n658_));
  AOI210     g636(.A0(new_new_n658_), .A1(new_new_n657_), .B0(new_new_n654_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n171_), .B(new_new_n117_), .Y(new_new_n660_));
  OAI210     g638(.A0(new_new_n660_), .A1(new_new_n646_), .B0(i_2_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n153_), .B(new_new_n80_), .Y(new_new_n662_));
  AOI210     g640(.A0(new_new_n662_), .A1(new_new_n661_), .B0(new_new_n174_), .Y(new_new_n663_));
  AN2        g641(.A(new_new_n537_), .B(i_13_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n180_), .B(new_new_n182_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n75_), .B(i_8_), .Y(new_new_n666_));
  AOI210     g644(.A0(new_new_n666_), .A1(new_new_n665_), .B0(new_new_n330_), .Y(new_new_n667_));
  AOI210     g645(.A0(new_new_n186_), .A1(new_new_n136_), .B0(new_new_n441_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n668_), .B(new_new_n366_), .Y(new_new_n669_));
  INV        g647(.A(new_new_n259_), .Y(new_new_n670_));
  NA4        g648(.A(new_new_n670_), .B(new_new_n263_), .C(new_new_n116_), .D(new_new_n42_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n671_), .B(new_new_n669_), .Y(new_new_n672_));
  NO4        g650(.A(new_new_n672_), .B(new_new_n667_), .C(new_new_n664_), .D(new_new_n663_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n495_), .B(new_new_n28_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n645_), .B(new_new_n238_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n675_), .B(new_new_n674_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n676_), .B(new_new_n46_), .Y(new_new_n677_));
  NA4        g655(.A(new_new_n677_), .B(new_new_n673_), .C(new_new_n659_), .D(new_new_n651_), .Y(mai6));
  NO2        g656(.A(i_9_), .B(i_1_), .Y(new_new_n679_));
  INV        g657(.A(new_new_n127_), .Y(new_new_n680_));
  OAI210     g658(.A0(new_new_n680_), .A1(new_new_n679_), .B0(new_new_n634_), .Y(new_new_n681_));
  NA4        g659(.A(new_new_n347_), .B(new_new_n411_), .C(new_new_n64_), .D(new_new_n93_), .Y(new_new_n682_));
  INV        g660(.A(new_new_n682_), .Y(new_new_n683_));
  NO2        g661(.A(i_11_), .B(i_9_), .Y(new_new_n684_));
  NO2        g662(.A(new_new_n683_), .B(new_new_n286_), .Y(new_new_n685_));
  AO210      g663(.A0(new_new_n685_), .A1(new_new_n681_), .B0(i_12_), .Y(new_new_n686_));
  NA2        g664(.A(new_new_n331_), .B(new_new_n293_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n502_), .B(new_new_n57_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n584_), .B(new_new_n64_), .Y(new_new_n689_));
  NA4        g667(.A(new_new_n541_), .B(new_new_n689_), .C(new_new_n688_), .D(new_new_n687_), .Y(new_new_n690_));
  INV        g668(.A(new_new_n177_), .Y(new_new_n691_));
  AOI220     g669(.A0(new_new_n691_), .A1(new_new_n684_), .B0(new_new_n690_), .B1(new_new_n66_), .Y(new_new_n692_));
  INV        g670(.A(new_new_n285_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n68_), .B(new_new_n122_), .Y(new_new_n694_));
  NA2        g672(.A(new_new_n25_), .B(new_new_n46_), .Y(new_new_n695_));
  AOI210     g673(.A0(new_new_n695_), .A1(new_new_n694_), .B0(new_new_n693_), .Y(new_new_n696_));
  NO2        g674(.A(new_new_n32_), .B(i_11_), .Y(new_new_n697_));
  NA3        g675(.A(new_new_n697_), .B(new_new_n403_), .C(new_new_n347_), .Y(new_new_n698_));
  NAi32      g676(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n699_));
  AOI210     g677(.A0(new_new_n621_), .A1(new_new_n78_), .B0(new_new_n699_), .Y(new_new_n700_));
  OAI210     g678(.A0(new_new_n583_), .A1(new_new_n483_), .B0(new_new_n482_), .Y(new_new_n701_));
  NAi31      g679(.An(new_new_n700_), .B(new_new_n701_), .C(new_new_n698_), .Y(new_new_n702_));
  OR2        g680(.A(new_new_n702_), .B(new_new_n696_), .Y(new_new_n703_));
  NO2        g681(.A(new_new_n599_), .B(i_2_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n916_), .B(new_new_n704_), .Y(new_new_n705_));
  AO220      g683(.A0(new_new_n315_), .A1(new_new_n306_), .B0(new_new_n352_), .B1(i_8_), .Y(new_new_n706_));
  NA3        g684(.A(new_new_n706_), .B(new_new_n222_), .C(i_7_), .Y(new_new_n707_));
  OR2        g685(.A(new_new_n537_), .B(new_new_n382_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n708_), .B(new_new_n135_), .Y(new_new_n709_));
  OR2        g687(.A(new_new_n648_), .B(new_new_n36_), .Y(new_new_n710_));
  NA4        g688(.A(new_new_n710_), .B(new_new_n709_), .C(new_new_n707_), .D(new_new_n705_), .Y(new_new_n711_));
  OAI210     g689(.A0(i_6_), .A1(i_11_), .B0(new_new_n78_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n712_), .B(new_new_n482_), .Y(new_new_n713_));
  NA3        g691(.A(new_new_n330_), .B(new_new_n210_), .C(new_new_n135_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n352_), .B(new_new_n63_), .Y(new_new_n715_));
  NA3        g693(.A(new_new_n715_), .B(new_new_n714_), .C(new_new_n713_), .Y(new_new_n716_));
  AO210      g694(.A0(new_new_n441_), .A1(new_new_n46_), .B0(new_new_n79_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n717_), .B(new_new_n412_), .Y(new_new_n718_));
  AOI210     g696(.A0(new_new_n382_), .A1(new_new_n380_), .B0(new_new_n481_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n103_), .B(new_new_n359_), .Y(new_new_n720_));
  NA3        g698(.A(new_new_n720_), .B(new_new_n719_), .C(new_new_n718_), .Y(new_new_n721_));
  NO4        g699(.A(new_new_n721_), .B(new_new_n716_), .C(new_new_n711_), .D(new_new_n703_), .Y(new_new_n722_));
  NA4        g700(.A(new_new_n722_), .B(new_new_n692_), .C(new_new_n686_), .D(new_new_n338_), .Y(mai3));
  NA2        g701(.A(i_6_), .B(i_7_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n724_), .B(i_0_), .Y(new_new_n725_));
  NO2        g703(.A(i_11_), .B(new_new_n209_), .Y(new_new_n726_));
  OAI210     g704(.A0(new_new_n725_), .A1(new_new_n248_), .B0(new_new_n726_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n727_), .B(new_new_n174_), .Y(new_new_n728_));
  NO3        g706(.A(new_new_n387_), .B(new_new_n82_), .C(new_new_n44_), .Y(new_new_n729_));
  OA210      g707(.A0(new_new_n729_), .A1(new_new_n728_), .B0(new_new_n156_), .Y(new_new_n730_));
  INV        g708(.A(new_new_n714_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n731_), .B(new_new_n39_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n544_), .B(new_new_n391_), .Y(new_new_n733_));
  AOI210     g711(.A0(new_new_n902_), .A1(new_new_n732_), .B0(new_new_n48_), .Y(new_new_n734_));
  NA2        g712(.A(new_new_n607_), .B(new_new_n576_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n291_), .B(i_5_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n736_), .B(new_new_n735_), .Y(new_new_n737_));
  NOi21      g715(.An(i_5_), .B(i_9_), .Y(new_new_n738_));
  NA2        g716(.A(new_new_n738_), .B(i_0_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n229_), .A1(new_new_n404_), .B0(new_new_n588_), .Y(new_new_n740_));
  NO2        g718(.A(new_new_n157_), .B(new_new_n136_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n741_), .B(new_new_n215_), .Y(new_new_n742_));
  OAI220     g720(.A0(new_new_n742_), .A1(new_new_n162_), .B0(new_new_n740_), .B1(new_new_n739_), .Y(new_new_n743_));
  NO4        g721(.A(new_new_n743_), .B(new_new_n737_), .C(new_new_n734_), .D(new_new_n730_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n167_), .B(new_new_n24_), .Y(new_new_n745_));
  NO2        g723(.A(new_new_n37_), .B(new_new_n745_), .Y(new_new_n746_));
  NA2        g724(.A(new_new_n269_), .B(new_new_n120_), .Y(new_new_n747_));
  NAi21      g725(.An(new_new_n146_), .B(i_5_), .Y(new_new_n748_));
  NO2        g726(.A(new_new_n747_), .B(new_new_n353_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n749_), .B(new_new_n746_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n492_), .B(i_0_), .Y(new_new_n751_));
  NO3        g729(.A(new_new_n751_), .B(new_new_n343_), .C(new_new_n80_), .Y(new_new_n752_));
  INV        g730(.A(new_new_n752_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n645_), .B(new_new_n286_), .Y(new_new_n754_));
  OAI220     g732(.A0(i_6_), .A1(new_new_n754_), .B0(new_new_n568_), .B1(new_new_n57_), .Y(new_new_n755_));
  NO4        g733(.A(new_new_n106_), .B(new_new_n52_), .C(new_new_n572_), .D(i_5_), .Y(new_new_n756_));
  AN2        g734(.A(new_new_n756_), .B(i_10_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n167_), .B(new_new_n76_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n486_), .B(i_4_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n170_), .B(new_new_n182_), .Y(new_new_n760_));
  OAI220     g738(.A0(new_new_n760_), .A1(new_new_n754_), .B0(new_new_n759_), .B1(new_new_n758_), .Y(new_new_n761_));
  NO3        g739(.A(new_new_n761_), .B(new_new_n757_), .C(new_new_n755_), .Y(new_new_n762_));
  NA3        g740(.A(new_new_n762_), .B(new_new_n753_), .C(new_new_n750_), .Y(new_new_n763_));
  NA2        g741(.A(i_11_), .B(i_9_), .Y(new_new_n764_));
  NO3        g742(.A(i_12_), .B(new_new_n764_), .C(new_new_n519_), .Y(new_new_n765_));
  AN2        g743(.A(new_new_n765_), .B(i_10_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n48_), .B(i_7_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n351_), .B(new_new_n161_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n768_), .B(new_new_n144_), .Y(new_new_n769_));
  NO2        g747(.A(new_new_n157_), .B(i_0_), .Y(new_new_n770_));
  NA2        g748(.A(new_new_n403_), .B(new_new_n205_), .Y(new_new_n771_));
  NA2        g749(.A(new_new_n329_), .B(new_new_n41_), .Y(new_new_n772_));
  OAI220     g750(.A0(new_new_n772_), .A1(new_new_n739_), .B0(new_new_n771_), .B1(new_new_n157_), .Y(new_new_n773_));
  NO3        g751(.A(new_new_n773_), .B(new_new_n769_), .C(new_new_n766_), .Y(new_new_n774_));
  NA2        g752(.A(new_new_n567_), .B(new_new_n113_), .Y(new_new_n775_));
  NO2        g753(.A(i_6_), .B(new_new_n775_), .Y(new_new_n776_));
  AOI210     g754(.A0(new_new_n381_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n153_), .B(new_new_n95_), .Y(new_new_n778_));
  NOi32      g756(.An(new_new_n777_), .Bn(new_new_n170_), .C(new_new_n778_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n520_), .B(new_new_n286_), .Y(new_new_n780_));
  NO2        g758(.A(new_new_n780_), .B(i_12_), .Y(new_new_n781_));
  NO3        g759(.A(new_new_n781_), .B(new_new_n779_), .C(new_new_n776_), .Y(new_new_n782_));
  NOi21      g760(.An(i_7_), .B(i_5_), .Y(new_new_n783_));
  NOi31      g761(.An(new_new_n783_), .B(i_0_), .C(new_new_n627_), .Y(new_new_n784_));
  NA3        g762(.A(new_new_n784_), .B(new_new_n342_), .C(i_6_), .Y(new_new_n785_));
  OA210      g763(.A0(new_new_n778_), .A1(new_new_n440_), .B0(new_new_n785_), .Y(new_new_n786_));
  NO3        g764(.A(new_new_n356_), .B(new_new_n318_), .C(new_new_n314_), .Y(new_new_n787_));
  NO2        g765(.A(new_new_n225_), .B(new_new_n275_), .Y(new_new_n788_));
  NO2        g766(.A(new_new_n627_), .B(new_new_n224_), .Y(new_new_n789_));
  AOI210     g767(.A0(new_new_n789_), .A1(new_new_n788_), .B0(new_new_n787_), .Y(new_new_n790_));
  NA4        g768(.A(new_new_n790_), .B(new_new_n786_), .C(new_new_n782_), .D(new_new_n774_), .Y(new_new_n791_));
  AN2        g769(.A(new_new_n290_), .B(new_new_n741_), .Y(new_new_n792_));
  NA2        g770(.A(new_new_n792_), .B(i_10_), .Y(new_new_n793_));
  NA3        g771(.A(new_new_n402_), .B(new_new_n360_), .C(new_new_n45_), .Y(new_new_n794_));
  OAI210     g772(.A0(new_new_n748_), .A1(i_6_), .B0(new_new_n794_), .Y(new_new_n795_));
  NA2        g773(.A(i_9_), .B(new_new_n263_), .Y(new_new_n796_));
  NA2        g774(.A(new_new_n169_), .B(new_new_n796_), .Y(new_new_n797_));
  AOI220     g775(.A0(new_new_n797_), .A1(new_new_n403_), .B0(new_new_n795_), .B1(new_new_n66_), .Y(new_new_n798_));
  NO2        g776(.A(new_new_n68_), .B(new_new_n647_), .Y(new_new_n799_));
  AOI210     g777(.A0(new_new_n156_), .A1(new_new_n511_), .B0(new_new_n799_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n47_), .Y(new_new_n801_));
  NO3        g779(.A(i_5_), .B(new_new_n313_), .C(new_new_n24_), .Y(new_new_n802_));
  NO2        g780(.A(new_new_n465_), .B(new_new_n802_), .Y(new_new_n803_));
  NAi21      g781(.An(i_9_), .B(i_5_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n804_), .B(new_new_n356_), .Y(new_new_n805_));
  NO2        g783(.A(new_new_n516_), .B(new_new_n96_), .Y(new_new_n806_));
  AOI220     g784(.A0(new_new_n806_), .A1(i_0_), .B0(new_new_n805_), .B1(new_new_n537_), .Y(new_new_n807_));
  OAI220     g785(.A0(new_new_n807_), .A1(new_new_n77_), .B0(new_new_n803_), .B1(new_new_n154_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n808_), .B(new_new_n801_), .Y(new_new_n809_));
  NA3        g787(.A(new_new_n809_), .B(new_new_n798_), .C(new_new_n793_), .Y(new_new_n810_));
  NO3        g788(.A(new_new_n810_), .B(new_new_n791_), .C(new_new_n763_), .Y(new_new_n811_));
  NO2        g789(.A(i_0_), .B(new_new_n627_), .Y(new_new_n812_));
  INV        g790(.A(i_0_), .Y(new_new_n813_));
  NO2        g791(.A(i_5_), .B(new_new_n25_), .Y(new_new_n814_));
  AO220      g792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n812_), .B1(new_new_n156_), .Y(new_new_n815_));
  AOI210     g793(.A0(new_new_n688_), .A1(new_new_n586_), .B0(new_new_n778_), .Y(new_new_n816_));
  AOI210     g794(.A0(new_new_n815_), .A1(new_new_n304_), .B0(new_new_n816_), .Y(new_new_n817_));
  NA3        g795(.A(new_new_n134_), .B(new_new_n576_), .C(new_new_n66_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n701_), .B(new_new_n356_), .Y(new_new_n819_));
  NA3        g797(.A(new_new_n725_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n726_), .B(i_9_), .Y(new_new_n821_));
  AOI210     g799(.A0(new_new_n820_), .A1(new_new_n422_), .B0(new_new_n821_), .Y(new_new_n822_));
  OAI210     g800(.A0(new_new_n215_), .A1(i_9_), .B0(new_new_n204_), .Y(new_new_n823_));
  AOI210     g801(.A0(new_new_n823_), .A1(new_new_n751_), .B0(new_new_n139_), .Y(new_new_n824_));
  NO3        g802(.A(new_new_n824_), .B(new_new_n822_), .C(new_new_n819_), .Y(new_new_n825_));
  NA3        g803(.A(new_new_n825_), .B(new_new_n818_), .C(new_new_n817_), .Y(new_new_n826_));
  NA3        g804(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n767_), .B(new_new_n415_), .Y(new_new_n828_));
  AOI210     g806(.A0(new_new_n827_), .A1(new_new_n146_), .B0(new_new_n828_), .Y(new_new_n829_));
  INV        g807(.A(new_new_n829_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n487_), .B(new_new_n68_), .Y(new_new_n831_));
  NO3        g809(.A(new_new_n187_), .B(new_new_n341_), .C(i_0_), .Y(new_new_n832_));
  OAI210     g810(.A0(new_new_n832_), .A1(new_new_n69_), .B0(i_13_), .Y(new_new_n833_));
  INV        g811(.A(new_new_n195_), .Y(new_new_n834_));
  OAI220     g812(.A0(new_new_n453_), .A1(new_new_n127_), .B0(new_new_n554_), .B1(new_new_n531_), .Y(new_new_n835_));
  NA3        g813(.A(new_new_n835_), .B(i_7_), .C(new_new_n834_), .Y(new_new_n836_));
  NA4        g814(.A(new_new_n836_), .B(new_new_n833_), .C(new_new_n831_), .D(new_new_n830_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n214_), .B(new_new_n85_), .Y(new_new_n838_));
  AOI210     g816(.A0(new_new_n838_), .A1(new_new_n812_), .B0(new_new_n100_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n783_), .B(new_new_n415_), .Y(new_new_n840_));
  NA2        g818(.A(new_new_n306_), .B(new_new_n158_), .Y(new_new_n841_));
  OA220      g819(.A0(new_new_n841_), .A1(new_new_n840_), .B0(new_new_n839_), .B1(i_5_), .Y(new_new_n842_));
  AOI210     g820(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n157_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n843_), .B(new_new_n402_), .Y(new_new_n844_));
  NA3        g822(.A(new_new_n347_), .B(new_new_n292_), .C(new_new_n197_), .Y(new_new_n845_));
  INV        g823(.A(new_new_n845_), .Y(new_new_n846_));
  NOi31      g824(.An(new_new_n346_), .B(i_0_), .C(new_new_n211_), .Y(new_new_n847_));
  NO3        g825(.A(new_new_n764_), .B(new_new_n195_), .C(new_new_n171_), .Y(new_new_n848_));
  NO3        g826(.A(new_new_n848_), .B(new_new_n847_), .C(new_new_n846_), .Y(new_new_n849_));
  NA4        g827(.A(new_new_n849_), .B(new_new_n401_), .C(new_new_n844_), .D(new_new_n842_), .Y(new_new_n850_));
  NA3        g828(.A(new_new_n263_), .B(i_5_), .C(new_new_n174_), .Y(new_new_n851_));
  NA2        g829(.A(new_new_n851_), .B(new_new_n214_), .Y(new_new_n852_));
  NO3        g830(.A(new_new_n211_), .B(i_0_), .C(i_12_), .Y(new_new_n853_));
  AOI220     g831(.A0(new_new_n853_), .A1(new_new_n852_), .B0(new_new_n683_), .B1(new_new_n158_), .Y(new_new_n854_));
  NO3        g832(.A(new_new_n911_), .B(i_12_), .C(new_new_n555_), .Y(new_new_n855_));
  INV        g833(.A(new_new_n855_), .Y(new_new_n856_));
  NA3        g834(.A(new_new_n90_), .B(new_new_n491_), .C(i_11_), .Y(new_new_n857_));
  NA2        g835(.A(new_new_n783_), .B(new_new_n400_), .Y(new_new_n858_));
  NO2        g836(.A(new_new_n858_), .B(i_1_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n859_), .B(new_new_n770_), .Y(new_new_n860_));
  NA3        g838(.A(new_new_n860_), .B(new_new_n856_), .C(new_new_n854_), .Y(new_new_n861_));
  NO4        g839(.A(new_new_n861_), .B(new_new_n850_), .C(new_new_n837_), .D(new_new_n826_), .Y(new_new_n862_));
  OAI210     g840(.A0(new_new_n704_), .A1(new_new_n697_), .B0(new_new_n37_), .Y(new_new_n863_));
  NA3        g841(.A(new_new_n777_), .B(new_new_n326_), .C(i_5_), .Y(new_new_n864_));
  NA3        g842(.A(new_new_n864_), .B(new_new_n863_), .C(new_new_n526_), .Y(new_new_n865_));
  NA2        g843(.A(new_new_n865_), .B(new_new_n185_), .Y(new_new_n866_));
  NA2        g844(.A(new_new_n168_), .B(new_new_n170_), .Y(new_new_n867_));
  OR2        g845(.A(i_11_), .B(new_new_n867_), .Y(new_new_n868_));
  OAI210     g846(.A0(new_new_n530_), .A1(new_new_n528_), .B0(new_new_n274_), .Y(new_new_n869_));
  NA2        g847(.A(new_new_n869_), .B(new_new_n868_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n394_), .B(new_new_n229_), .Y(new_new_n871_));
  INV        g849(.A(new_new_n871_), .Y(new_new_n872_));
  NA2        g850(.A(new_new_n857_), .B(new_new_n872_), .Y(new_new_n873_));
  AOI210     g851(.A0(new_new_n870_), .A1(new_new_n48_), .B0(new_new_n873_), .Y(new_new_n874_));
  AOI210     g852(.A0(new_new_n874_), .A1(new_new_n866_), .B0(new_new_n66_), .Y(new_new_n875_));
  NO2        g853(.A(new_new_n484_), .B(new_new_n337_), .Y(new_new_n876_));
  NO2        g854(.A(new_new_n876_), .B(new_new_n652_), .Y(new_new_n877_));
  INV        g855(.A(new_new_n69_), .Y(new_new_n878_));
  AOI210     g856(.A0(new_new_n843_), .A1(new_new_n767_), .B0(new_new_n784_), .Y(new_new_n879_));
  AOI210     g857(.A0(new_new_n879_), .A1(new_new_n878_), .B0(new_new_n577_), .Y(new_new_n880_));
  NA2        g858(.A(i_8_), .B(new_new_n69_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n881_), .B(new_new_n209_), .Y(new_new_n882_));
  NO2        g860(.A(new_new_n882_), .B(new_new_n880_), .Y(new_new_n883_));
  OAI210     g861(.A0(new_new_n231_), .A1(new_new_n142_), .B0(new_new_n80_), .Y(new_new_n884_));
  NO2        g862(.A(new_new_n884_), .B(i_11_), .Y(new_new_n885_));
  OAI210     g863(.A0(new_new_n903_), .A1(new_new_n777_), .B0(new_new_n185_), .Y(new_new_n886_));
  NA2        g864(.A(new_new_n148_), .B(i_5_), .Y(new_new_n887_));
  AOI210     g865(.A0(new_new_n886_), .A1(new_new_n665_), .B0(new_new_n887_), .Y(new_new_n888_));
  NA2        g866(.A(new_new_n788_), .B(new_new_n904_), .Y(new_new_n889_));
  NO2        g867(.A(new_new_n889_), .B(new_new_n627_), .Y(new_new_n890_));
  NO3        g868(.A(new_new_n804_), .B(new_new_n405_), .C(new_new_n221_), .Y(new_new_n891_));
  NO2        g869(.A(new_new_n891_), .B(new_new_n481_), .Y(new_new_n892_));
  INV        g870(.A(new_new_n319_), .Y(new_new_n893_));
  AOI210     g871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n40_), .Y(new_new_n894_));
  NO4        g872(.A(new_new_n894_), .B(new_new_n890_), .C(new_new_n888_), .D(new_new_n885_), .Y(new_new_n895_));
  OAI210     g873(.A0(new_new_n883_), .A1(i_4_), .B0(new_new_n895_), .Y(new_new_n896_));
  NO3        g874(.A(new_new_n896_), .B(new_new_n877_), .C(new_new_n875_), .Y(new_new_n897_));
  NA4        g875(.A(new_new_n897_), .B(new_new_n862_), .C(new_new_n811_), .D(new_new_n744_), .Y(mai4));
  INV        g876(.A(i_2_), .Y(new_new_n901_));
  INV        g877(.A(new_new_n733_), .Y(new_new_n902_));
  INV        g878(.A(i_12_), .Y(new_new_n903_));
  INV        g879(.A(i_4_), .Y(new_new_n904_));
  INV        g880(.A(new_new_n217_), .Y(new_new_n905_));
  INV        g881(.A(new_new_n130_), .Y(new_new_n906_));
  INV        g882(.A(i_5_), .Y(new_new_n907_));
  INV        g883(.A(i_2_), .Y(new_new_n908_));
  INV        g884(.A(i_3_), .Y(new_new_n909_));
  INV        g885(.A(new_new_n521_), .Y(new_new_n910_));
  INV        g886(.A(i_10_), .Y(new_new_n911_));
  INV        g887(.A(new_new_n178_), .Y(new_new_n912_));
  INV        g888(.A(new_new_n143_), .Y(new_new_n913_));
  INV        g889(.A(new_new_n196_), .Y(new_new_n914_));
  INV        g890(.A(i_10_), .Y(new_new_n915_));
  INV        g891(.A(i_5_), .Y(new_new_n916_));
  INV        g892(.A(i_13_), .Y(new_new_n917_));
endmodule


