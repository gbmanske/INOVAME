// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n141_, new_new_n143_,
    new_new_n144_, new_new_n145_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1058_, new_new_n1059_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g0068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g0069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g0070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g0071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g0073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g0074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g0076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g0078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g0079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g0080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g0081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g0082(.A(i_7_), .Y(new_new_n105_));
  NA2        g0083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g0084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g0085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g0087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g0088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g0089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n93_), .C(new_new_n54_), .Y(new_new_n113_));
  AN2        g0091(.A(i_2_), .B(i_10_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n114_), .B(i_7_), .Y(new_new_n115_));
  OR2        g0093(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n116_));
  NO2        g0094(.A(i_8_), .B(new_new_n105_), .Y(new_new_n117_));
  NO3        g0095(.A(new_new_n117_), .B(new_new_n116_), .C(new_new_n115_), .Y(new_new_n118_));
  NA2        g0096(.A(i_12_), .B(i_7_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n120_), .B(i_0_), .Y(new_new_n121_));
  NA2        g0099(.A(i_11_), .B(i_12_), .Y(new_new_n122_));
  OAI210     g0100(.A0(new_new_n121_), .A1(new_new_n119_), .B0(new_new_n122_), .Y(new_new_n123_));
  NO2        g0101(.A(new_new_n123_), .B(new_new_n118_), .Y(new_new_n124_));
  NAi41      g0102(.An(new_new_n113_), .B(new_new_n124_), .C(new_new_n111_), .D(new_new_n104_), .Y(new_new_n125_));
  NOi21      g0103(.An(i_1_), .B(i_5_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(i_11_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n128_));
  NA2        g0106(.A(i_7_), .B(new_new_n25_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n128_), .Y(new_new_n130_));
  NO2        g0108(.A(new_new_n130_), .B(new_new_n47_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n132_));
  NAi21      g0110(.An(i_3_), .B(i_8_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(new_new_n63_), .Y(new_new_n134_));
  NOi31      g0112(.An(new_new_n134_), .B(new_new_n132_), .C(new_new_n131_), .Y(new_new_n135_));
  NO2        g0113(.A(i_1_), .B(new_new_n87_), .Y(new_new_n136_));
  NO2        g0114(.A(i_6_), .B(i_5_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(i_3_), .Y(new_new_n138_));
  AO210      g0116(.A0(new_new_n138_), .A1(new_new_n48_), .B0(new_new_n136_), .Y(new_new_n139_));
  OAI220     g0117(.A0(new_new_n139_), .A1(new_new_n112_), .B0(new_new_n135_), .B1(new_new_n127_), .Y(new_new_n140_));
  NO3        g0118(.A(new_new_n140_), .B(new_new_n125_), .C(new_new_n99_), .Y(new_new_n141_));
  NA3        g0119(.A(new_new_n141_), .B(new_new_n80_), .C(new_new_n57_), .Y(men2));
  NO2        g0120(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n143_));
  NA2        g0121(.A(i_6_), .B(new_new_n25_), .Y(new_new_n144_));
  NA2        g0122(.A(new_new_n144_), .B(new_new_n143_), .Y(new_new_n145_));
  NA4        g0123(.A(new_new_n145_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(men0));
  AN2        g0124(.A(i_8_), .B(i_7_), .Y(new_new_n147_));
  NA2        g0125(.A(new_new_n147_), .B(i_6_), .Y(new_new_n148_));
  NO2        g0126(.A(i_12_), .B(i_13_), .Y(new_new_n149_));
  NAi21      g0127(.An(i_5_), .B(i_11_), .Y(new_new_n150_));
  NOi21      g0128(.An(new_new_n149_), .B(new_new_n150_), .Y(new_new_n151_));
  NO2        g0129(.A(i_0_), .B(i_1_), .Y(new_new_n152_));
  NA2        g0130(.A(i_2_), .B(i_3_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(i_4_), .Y(new_new_n154_));
  NA3        g0132(.A(new_new_n154_), .B(new_new_n152_), .C(new_new_n151_), .Y(new_new_n155_));
  OR2        g0133(.A(new_new_n155_), .B(new_new_n25_), .Y(new_new_n156_));
  AN2        g0134(.A(new_new_n149_), .B(new_new_n84_), .Y(new_new_n157_));
  NO2        g0135(.A(new_new_n157_), .B(new_new_n27_), .Y(new_new_n158_));
  NA2        g0136(.A(i_1_), .B(i_5_), .Y(new_new_n159_));
  NO2        g0137(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n160_));
  NA2        g0138(.A(new_new_n160_), .B(new_new_n36_), .Y(new_new_n161_));
  NO3        g0139(.A(new_new_n161_), .B(new_new_n159_), .C(new_new_n158_), .Y(new_new_n162_));
  OR2        g0140(.A(i_0_), .B(i_1_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n163_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n164_));
  NAi32      g0142(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n165_));
  NAi21      g0143(.An(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  NOi21      g0144(.An(i_4_), .B(i_10_), .Y(new_new_n167_));
  NA2        g0145(.A(new_new_n167_), .B(new_new_n40_), .Y(new_new_n168_));
  NO2        g0146(.A(i_3_), .B(i_5_), .Y(new_new_n169_));
  NO3        g0147(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n170_));
  INV        g0148(.A(new_new_n162_), .Y(new_new_n171_));
  AOI210     g0149(.A0(new_new_n171_), .A1(new_new_n156_), .B0(new_new_n148_), .Y(new_new_n172_));
  NA3        g0150(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n173_));
  NA2        g0151(.A(i_3_), .B(new_new_n49_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_4_), .B(i_9_), .Y(new_new_n175_));
  NOi21      g0153(.An(i_11_), .B(i_13_), .Y(new_new_n176_));
  NA2        g0154(.A(new_new_n176_), .B(new_new_n175_), .Y(new_new_n177_));
  NO2        g0155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g0156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n84_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n173_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n183_), .B(new_new_n47_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n36_), .B(i_5_), .Y(new_new_n185_));
  NAi31      g0163(.An(new_new_n185_), .B(new_new_n157_), .C(i_11_), .Y(new_new_n186_));
  NA2        g0164(.A(i_3_), .B(i_5_), .Y(new_new_n187_));
  OR2        g0165(.A(new_new_n187_), .B(new_new_n177_), .Y(new_new_n188_));
  AOI210     g0166(.A0(new_new_n188_), .A1(new_new_n186_), .B0(new_new_n184_), .Y(new_new_n189_));
  NO2        g0167(.A(new_new_n74_), .B(i_5_), .Y(new_new_n190_));
  NO2        g0168(.A(i_13_), .B(i_10_), .Y(new_new_n191_));
  NA3        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n45_), .Y(new_new_n192_));
  NO2        g0170(.A(i_2_), .B(i_1_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_3_), .Y(new_new_n194_));
  NAi21      g0172(.An(i_4_), .B(i_12_), .Y(new_new_n195_));
  NO4        g0173(.A(new_new_n195_), .B(new_new_n194_), .C(new_new_n192_), .D(new_new_n25_), .Y(new_new_n196_));
  NO3        g0174(.A(new_new_n196_), .B(new_new_n189_), .C(new_new_n182_), .Y(new_new_n197_));
  INV        g0175(.A(i_8_), .Y(new_new_n198_));
  NO2        g0176(.A(new_new_n198_), .B(i_7_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(i_6_), .Y(new_new_n200_));
  NO3        g0178(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n201_));
  NA2        g0179(.A(new_new_n201_), .B(new_new_n117_), .Y(new_new_n202_));
  NO3        g0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n205_));
  OAI210     g0183(.A0(new_new_n100_), .A1(i_12_), .B0(new_new_n205_), .Y(new_new_n206_));
  AOI210     g0184(.A0(new_new_n206_), .A1(new_new_n204_), .B0(new_new_n202_), .Y(new_new_n207_));
  NO2        g0185(.A(i_3_), .B(i_8_), .Y(new_new_n208_));
  NO3        g0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(new_new_n208_), .C(new_new_n40_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n211_));
  INV        g0189(.A(new_new_n211_), .Y(new_new_n212_));
  NO2        g0190(.A(i_13_), .B(i_9_), .Y(new_new_n213_));
  NA3        g0191(.A(new_new_n213_), .B(i_6_), .C(new_new_n198_), .Y(new_new_n214_));
  NAi21      g0192(.An(i_12_), .B(i_3_), .Y(new_new_n215_));
  OR2        g0193(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n45_), .B(i_5_), .Y(new_new_n217_));
  NO3        g0195(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n218_));
  NA3        g0196(.A(new_new_n218_), .B(new_new_n217_), .C(i_10_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n219_), .A1(new_new_n216_), .B0(new_new_n212_), .B1(new_new_n210_), .Y(new_new_n220_));
  AOI210     g0198(.A0(new_new_n220_), .A1(i_7_), .B0(new_new_n207_), .Y(new_new_n221_));
  OAI220     g0199(.A0(new_new_n221_), .A1(i_4_), .B0(new_new_n200_), .B1(new_new_n197_), .Y(new_new_n222_));
  NAi21      g0200(.An(i_12_), .B(i_7_), .Y(new_new_n223_));
  NA3        g0201(.A(i_13_), .B(new_new_n198_), .C(i_10_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  NA2        g0203(.A(i_0_), .B(i_5_), .Y(new_new_n226_));
  NA2        g0204(.A(new_new_n226_), .B(new_new_n108_), .Y(new_new_n227_));
  OAI220     g0205(.A0(new_new_n227_), .A1(new_new_n194_), .B0(new_new_n184_), .B1(new_new_n138_), .Y(new_new_n228_));
  NAi31      g0206(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n36_), .B(i_13_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n232_));
  NA3        g0210(.A(new_new_n232_), .B(new_new_n231_), .C(new_new_n230_), .Y(new_new_n233_));
  INV        g0211(.A(i_13_), .Y(new_new_n234_));
  NO2        g0212(.A(i_12_), .B(new_new_n234_), .Y(new_new_n235_));
  NA3        g0213(.A(new_new_n235_), .B(new_new_n203_), .C(new_new_n201_), .Y(new_new_n236_));
  OAI210     g0214(.A0(new_new_n233_), .A1(new_new_n229_), .B0(new_new_n236_), .Y(new_new_n237_));
  AOI220     g0215(.A0(new_new_n237_), .A1(new_new_n147_), .B0(new_new_n228_), .B1(new_new_n225_), .Y(new_new_n238_));
  NO2        g0216(.A(i_12_), .B(new_new_n37_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n187_), .B(i_4_), .Y(new_new_n240_));
  NA2        g0218(.A(new_new_n240_), .B(new_new_n239_), .Y(new_new_n241_));
  OR2        g0219(.A(i_8_), .B(i_7_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n242_), .B(new_new_n87_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n54_), .B(i_1_), .Y(new_new_n244_));
  INV        g0222(.A(i_12_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n45_), .B(new_new_n245_), .Y(new_new_n246_));
  NO3        g0224(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(i_2_), .B(i_1_), .Y(new_new_n248_));
  NO3        g0226(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n249_));
  NAi21      g0227(.An(i_4_), .B(i_3_), .Y(new_new_n250_));
  NO2        g0228(.A(new_new_n250_), .B(new_new_n76_), .Y(new_new_n251_));
  NO2        g0229(.A(i_0_), .B(i_6_), .Y(new_new_n252_));
  NOi41      g0230(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n253_), .B(new_new_n252_), .Y(new_new_n254_));
  NO2        g0232(.A(new_new_n248_), .B(new_new_n187_), .Y(new_new_n255_));
  NAi21      g0233(.An(new_new_n254_), .B(new_new_n255_), .Y(new_new_n256_));
  INV        g0234(.A(new_new_n256_), .Y(new_new_n257_));
  NA2        g0235(.A(new_new_n257_), .B(new_new_n40_), .Y(new_new_n258_));
  NO2        g0236(.A(i_11_), .B(new_new_n234_), .Y(new_new_n259_));
  NOi21      g0237(.An(i_1_), .B(i_6_), .Y(new_new_n260_));
  NAi21      g0238(.An(i_3_), .B(i_7_), .Y(new_new_n261_));
  NA2        g0239(.A(new_new_n245_), .B(i_9_), .Y(new_new_n262_));
  OR4        g0240(.A(new_new_n262_), .B(new_new_n261_), .C(new_new_n260_), .D(new_new_n190_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n264_));
  NO2        g0242(.A(i_12_), .B(i_3_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n74_), .B(i_5_), .Y(new_new_n266_));
  NA2        g0244(.A(i_3_), .B(i_9_), .Y(new_new_n267_));
  NAi21      g0245(.An(i_7_), .B(i_10_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n268_), .B(new_new_n267_), .Y(new_new_n269_));
  NA3        g0247(.A(new_new_n269_), .B(new_new_n266_), .C(new_new_n65_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n270_), .B(new_new_n263_), .Y(new_new_n271_));
  NA3        g0249(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n272_));
  INV        g0250(.A(new_new_n148_), .Y(new_new_n273_));
  NA2        g0251(.A(new_new_n245_), .B(i_13_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n274_), .B(new_new_n76_), .Y(new_new_n275_));
  AOI220     g0253(.A0(new_new_n275_), .A1(new_new_n273_), .B0(new_new_n271_), .B1(new_new_n259_), .Y(new_new_n276_));
  NO2        g0254(.A(new_new_n242_), .B(new_new_n37_), .Y(new_new_n277_));
  NA2        g0255(.A(i_12_), .B(i_6_), .Y(new_new_n278_));
  OR2        g0256(.A(i_13_), .B(i_9_), .Y(new_new_n279_));
  NO3        g0257(.A(new_new_n279_), .B(new_new_n278_), .C(new_new_n49_), .Y(new_new_n280_));
  NO2        g0258(.A(new_new_n250_), .B(i_2_), .Y(new_new_n281_));
  NA3        g0259(.A(new_new_n281_), .B(new_new_n280_), .C(new_new_n45_), .Y(new_new_n282_));
  NA2        g0260(.A(new_new_n259_), .B(i_9_), .Y(new_new_n283_));
  NA2        g0261(.A(new_new_n266_), .B(new_new_n65_), .Y(new_new_n284_));
  OAI210     g0262(.A0(new_new_n284_), .A1(new_new_n283_), .B0(new_new_n282_), .Y(new_new_n285_));
  NA2        g0263(.A(new_new_n160_), .B(new_new_n64_), .Y(new_new_n286_));
  NO3        g0264(.A(i_11_), .B(new_new_n234_), .C(new_new_n25_), .Y(new_new_n287_));
  NO2        g0265(.A(new_new_n261_), .B(i_8_), .Y(new_new_n288_));
  NO2        g0266(.A(i_6_), .B(new_new_n49_), .Y(new_new_n289_));
  NA3        g0267(.A(new_new_n289_), .B(new_new_n288_), .C(new_new_n287_), .Y(new_new_n290_));
  NO3        g0268(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n291_));
  NA3        g0269(.A(new_new_n291_), .B(new_new_n277_), .C(new_new_n235_), .Y(new_new_n292_));
  AOI210     g0270(.A0(new_new_n292_), .A1(new_new_n290_), .B0(new_new_n286_), .Y(new_new_n293_));
  AOI210     g0271(.A0(new_new_n285_), .A1(new_new_n277_), .B0(new_new_n293_), .Y(new_new_n294_));
  NA4        g0272(.A(new_new_n294_), .B(new_new_n276_), .C(new_new_n258_), .D(new_new_n238_), .Y(new_new_n295_));
  NO3        g0273(.A(i_12_), .B(new_new_n234_), .C(new_new_n37_), .Y(new_new_n296_));
  NO3        g0274(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n248_), .B(i_0_), .Y(new_new_n298_));
  NA2        g0276(.A(i_0_), .B(i_1_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(i_2_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n60_), .B(i_6_), .Y(new_new_n301_));
  NA3        g0279(.A(new_new_n301_), .B(new_new_n300_), .C(new_new_n169_), .Y(new_new_n302_));
  NO2        g0280(.A(i_3_), .B(i_10_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n304_));
  NO2        g0282(.A(i_2_), .B(new_new_n105_), .Y(new_new_n305_));
  NA2        g0283(.A(i_1_), .B(new_new_n36_), .Y(new_new_n306_));
  NO2        g0284(.A(new_new_n306_), .B(i_8_), .Y(new_new_n307_));
  NOi21      g0285(.An(new_new_n226_), .B(new_new_n107_), .Y(new_new_n308_));
  NA3        g0286(.A(new_new_n308_), .B(new_new_n307_), .C(new_new_n305_), .Y(new_new_n309_));
  AN2        g0287(.A(i_3_), .B(i_10_), .Y(new_new_n310_));
  NA4        g0288(.A(new_new_n310_), .B(new_new_n203_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n311_));
  NO2        g0289(.A(i_5_), .B(new_new_n37_), .Y(new_new_n312_));
  NO2        g0290(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n313_));
  OR2        g0291(.A(new_new_n309_), .B(new_new_n304_), .Y(new_new_n314_));
  NO2        g0292(.A(new_new_n314_), .B(i_6_), .Y(new_new_n315_));
  NO4        g0293(.A(new_new_n315_), .B(new_new_n295_), .C(new_new_n222_), .D(new_new_n172_), .Y(new_new_n316_));
  NO3        g0294(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n317_));
  NO2        g0295(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n318_));
  NO3        g0296(.A(i_6_), .B(new_new_n198_), .C(i_7_), .Y(new_new_n319_));
  NO2        g0297(.A(i_2_), .B(i_3_), .Y(new_new_n320_));
  OR2        g0298(.A(i_0_), .B(i_5_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n226_), .B(new_new_n321_), .Y(new_new_n322_));
  NA4        g0300(.A(new_new_n322_), .B(new_new_n243_), .C(new_new_n320_), .D(i_1_), .Y(new_new_n323_));
  NAi21      g0301(.An(i_8_), .B(i_7_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n324_), .B(i_6_), .Y(new_new_n325_));
  NO2        g0303(.A(new_new_n163_), .B(new_new_n47_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n325_), .C(new_new_n169_), .Y(new_new_n327_));
  NA2        g0305(.A(new_new_n327_), .B(new_new_n323_), .Y(new_new_n328_));
  NA2        g0306(.A(new_new_n328_), .B(i_4_), .Y(new_new_n329_));
  NO2        g0307(.A(i_12_), .B(i_10_), .Y(new_new_n330_));
  NOi21      g0308(.An(i_5_), .B(i_0_), .Y(new_new_n331_));
  NA4        g0309(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n332_));
  NO2        g0310(.A(i_6_), .B(i_8_), .Y(new_new_n333_));
  NOi21      g0311(.An(i_0_), .B(i_2_), .Y(new_new_n334_));
  AN2        g0312(.A(new_new_n334_), .B(new_new_n333_), .Y(new_new_n335_));
  NO2        g0313(.A(i_1_), .B(i_7_), .Y(new_new_n336_));
  AO220      g0314(.A0(new_new_n336_), .A1(new_new_n335_), .B0(new_new_n325_), .B1(new_new_n244_), .Y(new_new_n337_));
  NA3        g0315(.A(new_new_n337_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n338_), .B(new_new_n329_), .Y(new_new_n339_));
  NO3        g0317(.A(new_new_n242_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n340_));
  NO3        g0318(.A(new_new_n324_), .B(i_2_), .C(i_1_), .Y(new_new_n341_));
  OAI210     g0319(.A0(new_new_n341_), .A1(new_new_n340_), .B0(i_6_), .Y(new_new_n342_));
  NA3        g0320(.A(new_new_n260_), .B(new_new_n305_), .C(new_new_n198_), .Y(new_new_n343_));
  AOI210     g0321(.A0(new_new_n343_), .A1(new_new_n342_), .B0(new_new_n322_), .Y(new_new_n344_));
  INV        g0322(.A(new_new_n108_), .Y(new_new_n345_));
  NA2        g0323(.A(new_new_n344_), .B(i_3_), .Y(new_new_n346_));
  INV        g0324(.A(new_new_n85_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n299_), .B(new_new_n82_), .Y(new_new_n348_));
  NA2        g0326(.A(new_new_n348_), .B(new_new_n137_), .Y(new_new_n349_));
  NO2        g0327(.A(new_new_n96_), .B(new_new_n198_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n308_), .B(new_new_n350_), .C(new_new_n64_), .Y(new_new_n351_));
  AOI210     g0329(.A0(new_new_n351_), .A1(new_new_n349_), .B0(new_new_n347_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n198_), .B(i_9_), .Y(new_new_n353_));
  NA2        g0331(.A(new_new_n353_), .B(new_new_n211_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n354_), .B(new_new_n47_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n355_), .B(new_new_n352_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n356_), .A1(new_new_n346_), .B0(new_new_n168_), .Y(new_new_n357_));
  AOI210     g0335(.A0(new_new_n339_), .A1(new_new_n317_), .B0(new_new_n357_), .Y(new_new_n358_));
  NOi32      g0336(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n359_));
  INV        g0337(.A(new_new_n359_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_0_), .B(i_6_), .Y(new_new_n361_));
  NAi21      g0339(.An(i_1_), .B(i_5_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n361_), .Y(new_new_n363_));
  NA2        g0341(.A(new_new_n363_), .B(new_new_n25_), .Y(new_new_n364_));
  OAI210     g0342(.A0(new_new_n364_), .A1(new_new_n165_), .B0(new_new_n254_), .Y(new_new_n365_));
  NAi41      g0343(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n366_));
  AOI210     g0344(.A0(new_new_n366_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n367_));
  NOi32      g0345(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n368_));
  NAi21      g0346(.An(i_6_), .B(i_1_), .Y(new_new_n369_));
  NO2        g0347(.A(i_1_), .B(new_new_n105_), .Y(new_new_n370_));
  NAi21      g0348(.An(i_3_), .B(i_4_), .Y(new_new_n371_));
  NO2        g0349(.A(new_new_n371_), .B(i_9_), .Y(new_new_n372_));
  AN2        g0350(.A(i_6_), .B(i_7_), .Y(new_new_n373_));
  OAI210     g0351(.A0(new_new_n373_), .A1(new_new_n370_), .B0(new_new_n372_), .Y(new_new_n374_));
  NA2        g0352(.A(i_2_), .B(i_7_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n371_), .B(i_10_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n374_), .B(new_new_n190_), .Y(new_new_n377_));
  AOI210     g0355(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n378_));
  OAI210     g0356(.A0(new_new_n378_), .A1(new_new_n193_), .B0(new_new_n376_), .Y(new_new_n379_));
  AOI220     g0357(.A0(new_new_n376_), .A1(new_new_n336_), .B0(new_new_n247_), .B1(new_new_n193_), .Y(new_new_n380_));
  AOI210     g0358(.A0(new_new_n380_), .A1(new_new_n379_), .B0(i_5_), .Y(new_new_n381_));
  NO4        g0359(.A(new_new_n381_), .B(new_new_n377_), .C(new_new_n367_), .D(new_new_n365_), .Y(new_new_n382_));
  NO2        g0360(.A(new_new_n382_), .B(new_new_n360_), .Y(new_new_n383_));
  AN2        g0361(.A(i_12_), .B(i_5_), .Y(new_new_n384_));
  NA2        g0362(.A(i_3_), .B(new_new_n384_), .Y(new_new_n385_));
  NO2        g0363(.A(i_11_), .B(i_6_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n250_), .B(i_5_), .Y(new_new_n387_));
  NO2        g0365(.A(i_5_), .B(i_10_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n389_));
  NO3        g0367(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n390_));
  NO2        g0368(.A(i_3_), .B(new_new_n105_), .Y(new_new_n391_));
  NO2        g0369(.A(i_11_), .B(i_12_), .Y(new_new_n392_));
  NA2        g0370(.A(new_new_n388_), .B(new_new_n245_), .Y(new_new_n393_));
  NA3        g0371(.A(new_new_n117_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n394_));
  OAI220     g0372(.A0(new_new_n394_), .A1(new_new_n229_), .B0(new_new_n393_), .B1(new_new_n332_), .Y(new_new_n395_));
  NAi21      g0373(.An(i_13_), .B(i_0_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n396_), .B(new_new_n248_), .Y(new_new_n397_));
  NA2        g0375(.A(new_new_n395_), .B(new_new_n397_), .Y(new_new_n398_));
  INV        g0376(.A(new_new_n398_), .Y(new_new_n399_));
  NO3        g0377(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n400_));
  NO2        g0378(.A(i_0_), .B(i_11_), .Y(new_new_n401_));
  INV        g0379(.A(i_5_), .Y(new_new_n402_));
  AN2        g0380(.A(i_1_), .B(i_6_), .Y(new_new_n403_));
  NOi21      g0381(.An(i_2_), .B(i_12_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n404_), .B(new_new_n403_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n405_), .B(new_new_n402_), .Y(new_new_n406_));
  NA2        g0384(.A(new_new_n147_), .B(i_9_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(i_4_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n406_), .B(new_new_n408_), .Y(new_new_n409_));
  NAi21      g0387(.An(i_9_), .B(i_4_), .Y(new_new_n410_));
  OR2        g0388(.A(i_13_), .B(i_10_), .Y(new_new_n411_));
  NO3        g0389(.A(new_new_n411_), .B(new_new_n122_), .C(new_new_n410_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n177_), .B(new_new_n128_), .Y(new_new_n413_));
  OR2        g0391(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n296_), .B(new_new_n415_), .Y(new_new_n416_));
  NA2        g0394(.A(new_new_n289_), .B(new_new_n218_), .Y(new_new_n417_));
  OAI220     g0395(.A0(new_new_n417_), .A1(new_new_n414_), .B0(new_new_n416_), .B1(new_new_n345_), .Y(new_new_n418_));
  INV        g0396(.A(new_new_n418_), .Y(new_new_n419_));
  AOI210     g0397(.A0(new_new_n419_), .A1(new_new_n409_), .B0(new_new_n26_), .Y(new_new_n420_));
  INV        g0398(.A(new_new_n323_), .Y(new_new_n421_));
  AOI220     g0399(.A0(new_new_n301_), .A1(new_new_n297_), .B0(new_new_n298_), .B1(new_new_n318_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n422_), .B(new_new_n174_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n423_), .B(new_new_n421_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n198_), .B(i_10_), .Y(new_new_n425_));
  NA3        g0403(.A(new_new_n266_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n301_), .B(new_new_n244_), .Y(new_new_n427_));
  OAI220     g0405(.A0(new_new_n427_), .A1(new_new_n187_), .B0(new_new_n426_), .B1(new_new_n425_), .Y(new_new_n428_));
  NO2        g0406(.A(i_3_), .B(new_new_n49_), .Y(new_new_n429_));
  INV        g0407(.A(new_new_n428_), .Y(new_new_n430_));
  AOI210     g0408(.A0(new_new_n430_), .A1(new_new_n424_), .B0(new_new_n283_), .Y(new_new_n431_));
  NO4        g0409(.A(new_new_n431_), .B(new_new_n420_), .C(new_new_n399_), .D(new_new_n383_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n64_), .B(i_4_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n74_), .B(i_13_), .Y(new_new_n434_));
  NA3        g0412(.A(new_new_n434_), .B(new_new_n433_), .C(i_2_), .Y(new_new_n435_));
  NO2        g0413(.A(i_10_), .B(i_9_), .Y(new_new_n436_));
  NAi21      g0414(.An(i_12_), .B(i_8_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n437_), .B(i_3_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n438_), .B(new_new_n436_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n47_), .B(i_4_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n440_), .B(new_new_n108_), .Y(new_new_n441_));
  OAI220     g0419(.A0(new_new_n441_), .A1(new_new_n210_), .B0(new_new_n439_), .B1(new_new_n435_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n313_), .B(i_0_), .Y(new_new_n443_));
  NO3        g0421(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n278_), .B(new_new_n101_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n445_), .B(new_new_n444_), .Y(new_new_n446_));
  NA2        g0424(.A(i_8_), .B(i_9_), .Y(new_new_n447_));
  AOI210     g0425(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n448_));
  OR2        g0426(.A(new_new_n448_), .B(new_new_n447_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n296_), .B(new_new_n211_), .Y(new_new_n450_));
  OAI220     g0428(.A0(new_new_n450_), .A1(new_new_n449_), .B0(new_new_n446_), .B1(new_new_n443_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n259_), .B(new_new_n312_), .Y(new_new_n452_));
  NO3        g0430(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n453_));
  INV        g0431(.A(new_new_n453_), .Y(new_new_n454_));
  NA3        g0432(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n455_));
  NA4        g0433(.A(new_new_n150_), .B(new_new_n120_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n456_));
  OAI220     g0434(.A0(new_new_n456_), .A1(new_new_n455_), .B0(new_new_n454_), .B1(new_new_n452_), .Y(new_new_n457_));
  NO3        g0435(.A(new_new_n457_), .B(new_new_n451_), .C(new_new_n442_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n300_), .B(new_new_n112_), .Y(new_new_n459_));
  OR2        g0437(.A(new_new_n459_), .B(new_new_n214_), .Y(new_new_n460_));
  OA210      g0438(.A0(new_new_n354_), .A1(new_new_n105_), .B0(new_new_n302_), .Y(new_new_n461_));
  OA220      g0439(.A0(new_new_n461_), .A1(new_new_n168_), .B0(new_new_n460_), .B1(new_new_n241_), .Y(new_new_n462_));
  NA2        g0440(.A(new_new_n100_), .B(i_13_), .Y(new_new_n463_));
  NO2        g0441(.A(i_2_), .B(i_13_), .Y(new_new_n464_));
  NO3        g0442(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n465_));
  NO2        g0443(.A(i_6_), .B(i_7_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n466_), .B(new_new_n465_), .Y(new_new_n467_));
  NO2        g0445(.A(i_11_), .B(i_1_), .Y(new_new_n468_));
  NO2        g0446(.A(new_new_n74_), .B(i_3_), .Y(new_new_n469_));
  OR2        g0447(.A(i_11_), .B(i_8_), .Y(new_new_n470_));
  NOi21      g0448(.An(i_2_), .B(i_7_), .Y(new_new_n471_));
  NAi31      g0449(.An(new_new_n470_), .B(new_new_n471_), .C(new_new_n469_), .Y(new_new_n472_));
  NO2        g0450(.A(new_new_n411_), .B(i_6_), .Y(new_new_n473_));
  NA3        g0451(.A(new_new_n473_), .B(new_new_n433_), .C(new_new_n76_), .Y(new_new_n474_));
  NO2        g0452(.A(new_new_n474_), .B(new_new_n472_), .Y(new_new_n475_));
  NO2        g0453(.A(i_3_), .B(new_new_n198_), .Y(new_new_n476_));
  NO2        g0454(.A(i_6_), .B(i_10_), .Y(new_new_n477_));
  NA4        g0455(.A(new_new_n477_), .B(new_new_n317_), .C(new_new_n476_), .D(new_new_n245_), .Y(new_new_n478_));
  NO2        g0456(.A(new_new_n478_), .B(new_new_n161_), .Y(new_new_n479_));
  NA3        g0457(.A(new_new_n253_), .B(new_new_n176_), .C(new_new_n137_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n163_), .B(i_3_), .Y(new_new_n482_));
  NAi31      g0460(.An(new_new_n481_), .B(new_new_n482_), .C(new_new_n235_), .Y(new_new_n483_));
  NA3        g0461(.A(new_new_n389_), .B(new_new_n183_), .C(new_new_n154_), .Y(new_new_n484_));
  NA3        g0462(.A(new_new_n484_), .B(new_new_n483_), .C(new_new_n480_), .Y(new_new_n485_));
  NO3        g0463(.A(new_new_n485_), .B(new_new_n479_), .C(new_new_n475_), .Y(new_new_n486_));
  NA2        g0464(.A(new_new_n444_), .B(new_new_n384_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n453_), .B(new_new_n388_), .Y(new_new_n488_));
  NO2        g0466(.A(new_new_n488_), .B(new_new_n233_), .Y(new_new_n489_));
  NAi21      g0467(.An(new_new_n224_), .B(new_new_n392_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n26_), .B(i_5_), .Y(new_new_n491_));
  NO2        g0469(.A(i_0_), .B(new_new_n87_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n492_), .B(new_new_n491_), .C(new_new_n147_), .Y(new_new_n493_));
  OR3        g0471(.A(new_new_n306_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n27_), .B(i_10_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n317_), .B(new_new_n247_), .Y(new_new_n497_));
  OAI220     g0475(.A0(new_new_n497_), .A1(new_new_n426_), .B0(new_new_n496_), .B1(new_new_n463_), .Y(new_new_n498_));
  NA4        g0476(.A(new_new_n310_), .B(new_new_n232_), .C(new_new_n74_), .D(new_new_n245_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n499_), .B(new_new_n467_), .Y(new_new_n500_));
  NO4        g0478(.A(new_new_n500_), .B(new_new_n498_), .C(new_new_n495_), .D(new_new_n489_), .Y(new_new_n501_));
  NA4        g0479(.A(new_new_n501_), .B(new_new_n486_), .C(new_new_n462_), .D(new_new_n458_), .Y(new_new_n502_));
  NA3        g0480(.A(new_new_n310_), .B(new_new_n180_), .C(new_new_n178_), .Y(new_new_n503_));
  OAI210     g0481(.A0(new_new_n304_), .A1(new_new_n185_), .B0(new_new_n503_), .Y(new_new_n504_));
  AN2        g0482(.A(new_new_n297_), .B(new_new_n243_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n505_), .B(new_new_n504_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n127_), .B(new_new_n116_), .Y(new_new_n507_));
  AN2        g0485(.A(new_new_n507_), .B(new_new_n444_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n317_), .B(new_new_n170_), .Y(new_new_n509_));
  OAI210     g0487(.A0(new_new_n509_), .A1(new_new_n241_), .B0(new_new_n311_), .Y(new_new_n510_));
  AOI220     g0488(.A0(new_new_n510_), .A1(new_new_n325_), .B0(new_new_n508_), .B1(new_new_n313_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n384_), .B(new_new_n234_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n359_), .B(new_new_n74_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n373_), .B(new_new_n368_), .Y(new_new_n514_));
  OR2        g0492(.A(new_new_n512_), .B(new_new_n514_), .Y(new_new_n515_));
  NO2        g0493(.A(new_new_n36_), .B(i_8_), .Y(new_new_n516_));
  NAi41      g0494(.An(new_new_n513_), .B(new_new_n477_), .C(new_new_n516_), .D(new_new_n47_), .Y(new_new_n517_));
  AOI210     g0495(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n412_), .Y(new_new_n518_));
  NA3        g0496(.A(new_new_n518_), .B(new_new_n517_), .C(new_new_n515_), .Y(new_new_n519_));
  INV        g0497(.A(new_new_n519_), .Y(new_new_n520_));
  INV        g0498(.A(new_new_n139_), .Y(new_new_n521_));
  NO2        g0499(.A(i_7_), .B(new_new_n204_), .Y(new_new_n522_));
  OR2        g0500(.A(new_new_n187_), .B(i_4_), .Y(new_new_n523_));
  NO2        g0501(.A(new_new_n523_), .B(new_new_n87_), .Y(new_new_n524_));
  AOI220     g0502(.A0(new_new_n524_), .A1(new_new_n522_), .B0(new_new_n521_), .B1(new_new_n413_), .Y(new_new_n525_));
  NA4        g0503(.A(new_new_n525_), .B(new_new_n520_), .C(new_new_n511_), .D(new_new_n506_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n387_), .B(new_new_n300_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n385_), .A1(new_new_n173_), .B0(new_new_n527_), .Y(new_new_n528_));
  NO2        g0506(.A(i_12_), .B(new_new_n198_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n529_), .B(new_new_n234_), .Y(new_new_n530_));
  NO3        g0508(.A(new_new_n1059_), .B(new_new_n530_), .C(new_new_n459_), .Y(new_new_n531_));
  NOi31      g0509(.An(new_new_n319_), .B(new_new_n411_), .C(new_new_n38_), .Y(new_new_n532_));
  OAI210     g0510(.A0(new_new_n532_), .A1(new_new_n531_), .B0(new_new_n528_), .Y(new_new_n533_));
  NO2        g0511(.A(i_8_), .B(i_7_), .Y(new_new_n534_));
  OAI210     g0512(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n535_), .B(new_new_n232_), .Y(new_new_n536_));
  AOI220     g0514(.A0(new_new_n326_), .A1(new_new_n40_), .B0(new_new_n244_), .B1(new_new_n213_), .Y(new_new_n537_));
  OAI220     g0515(.A0(new_new_n537_), .A1(new_new_n523_), .B0(new_new_n536_), .B1(new_new_n250_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n45_), .B(i_10_), .Y(new_new_n539_));
  NO2        g0517(.A(new_new_n539_), .B(i_6_), .Y(new_new_n540_));
  NA3        g0518(.A(new_new_n540_), .B(new_new_n538_), .C(new_new_n534_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n463_), .B(new_new_n138_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n542_), .B(new_new_n277_), .Y(new_new_n543_));
  NOi31      g0521(.An(new_new_n298_), .B(new_new_n304_), .C(new_new_n185_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n544_), .B(new_new_n453_), .Y(new_new_n545_));
  NA4        g0523(.A(new_new_n545_), .B(new_new_n543_), .C(new_new_n541_), .D(new_new_n533_), .Y(new_new_n546_));
  NA3        g0524(.A(new_new_n226_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n296_), .B(new_new_n85_), .Y(new_new_n548_));
  AOI210     g0526(.A0(new_new_n547_), .A1(new_new_n349_), .B0(new_new_n548_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n436_), .B(new_new_n230_), .Y(new_new_n551_));
  NO2        g0529(.A(new_new_n550_), .B(new_new_n551_), .Y(new_new_n552_));
  AOI210     g0530(.A0(new_new_n369_), .A1(new_new_n47_), .B0(new_new_n370_), .Y(new_new_n553_));
  NA2        g0531(.A(i_0_), .B(new_new_n49_), .Y(new_new_n554_));
  NA3        g0532(.A(new_new_n529_), .B(new_new_n287_), .C(new_new_n554_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n553_), .B(new_new_n555_), .Y(new_new_n556_));
  NO3        g0534(.A(new_new_n556_), .B(new_new_n552_), .C(new_new_n549_), .Y(new_new_n557_));
  NO4        g0535(.A(new_new_n260_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n558_));
  NO3        g0536(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n242_), .B(new_new_n36_), .Y(new_new_n560_));
  AN2        g0538(.A(new_new_n560_), .B(new_new_n559_), .Y(new_new_n561_));
  OA210      g0539(.A0(new_new_n561_), .A1(new_new_n558_), .B0(new_new_n359_), .Y(new_new_n562_));
  NO2        g0540(.A(new_new_n411_), .B(i_1_), .Y(new_new_n563_));
  NOi31      g0541(.An(new_new_n563_), .B(new_new_n445_), .C(new_new_n74_), .Y(new_new_n564_));
  AN4        g0542(.A(new_new_n564_), .B(new_new_n408_), .C(new_new_n491_), .D(i_2_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n422_), .B(new_new_n181_), .Y(new_new_n566_));
  NO3        g0544(.A(new_new_n566_), .B(new_new_n565_), .C(new_new_n562_), .Y(new_new_n567_));
  NOi21      g0545(.An(i_10_), .B(i_6_), .Y(new_new_n568_));
  NO2        g0546(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n569_));
  AOI220     g0547(.A0(new_new_n296_), .A1(new_new_n569_), .B0(new_new_n287_), .B1(new_new_n568_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n570_), .B(new_new_n443_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n572_));
  NA2        g0550(.A(new_new_n319_), .B(new_new_n170_), .Y(new_new_n573_));
  AOI220     g0551(.A0(new_new_n573_), .A1(new_new_n427_), .B0(new_new_n188_), .B1(new_new_n186_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n203_), .B(new_new_n37_), .Y(new_new_n575_));
  NOi31      g0553(.An(new_new_n151_), .B(new_new_n575_), .C(new_new_n332_), .Y(new_new_n576_));
  NO3        g0554(.A(new_new_n576_), .B(new_new_n574_), .C(new_new_n571_), .Y(new_new_n577_));
  INV        g0555(.A(new_new_n320_), .Y(new_new_n578_));
  NO2        g0556(.A(i_12_), .B(new_new_n87_), .Y(new_new_n579_));
  NA3        g0557(.A(new_new_n579_), .B(new_new_n287_), .C(new_new_n554_), .Y(new_new_n580_));
  NA3        g0558(.A(new_new_n386_), .B(new_new_n296_), .C(new_new_n226_), .Y(new_new_n581_));
  AOI210     g0559(.A0(new_new_n581_), .A1(new_new_n580_), .B0(new_new_n578_), .Y(new_new_n582_));
  NA2        g0560(.A(new_new_n178_), .B(i_0_), .Y(new_new_n583_));
  NO3        g0561(.A(new_new_n583_), .B(new_new_n342_), .C(new_new_n304_), .Y(new_new_n584_));
  OR2        g0562(.A(i_2_), .B(i_5_), .Y(new_new_n585_));
  OR2        g0563(.A(new_new_n585_), .B(new_new_n403_), .Y(new_new_n586_));
  AOI210     g0564(.A0(new_new_n375_), .A1(new_new_n252_), .B0(new_new_n203_), .Y(new_new_n587_));
  AOI210     g0565(.A0(new_new_n587_), .A1(new_new_n586_), .B0(new_new_n490_), .Y(new_new_n588_));
  NO3        g0566(.A(new_new_n588_), .B(new_new_n584_), .C(new_new_n582_), .Y(new_new_n589_));
  NA4        g0567(.A(new_new_n589_), .B(new_new_n577_), .C(new_new_n567_), .D(new_new_n557_), .Y(new_new_n590_));
  NO4        g0568(.A(new_new_n590_), .B(new_new_n546_), .C(new_new_n526_), .D(new_new_n502_), .Y(new_new_n591_));
  NA4        g0569(.A(new_new_n591_), .B(new_new_n432_), .C(new_new_n358_), .D(new_new_n316_), .Y(men7));
  NO2        g0570(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n593_));
  NA2        g0571(.A(new_new_n477_), .B(new_new_n85_), .Y(new_new_n594_));
  NA2        g0572(.A(i_11_), .B(new_new_n198_), .Y(new_new_n595_));
  NA3        g0573(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n245_), .B(i_4_), .Y(new_new_n597_));
  NA2        g0575(.A(new_new_n597_), .B(i_8_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n109_), .B(new_new_n596_), .Y(new_new_n599_));
  NA2        g0577(.A(i_2_), .B(new_new_n87_), .Y(new_new_n600_));
  OAI210     g0578(.A0(new_new_n90_), .A1(new_new_n208_), .B0(new_new_n209_), .Y(new_new_n601_));
  NO2        g0579(.A(i_7_), .B(new_new_n37_), .Y(new_new_n602_));
  NA2        g0580(.A(i_4_), .B(i_8_), .Y(new_new_n603_));
  AOI210     g0581(.A0(new_new_n603_), .A1(new_new_n310_), .B0(new_new_n602_), .Y(new_new_n604_));
  OAI220     g0582(.A0(new_new_n604_), .A1(new_new_n600_), .B0(new_new_n601_), .B1(i_13_), .Y(new_new_n605_));
  NO3        g0583(.A(new_new_n605_), .B(new_new_n599_), .C(new_new_n593_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n133_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n607_));
  AOI210     g0585(.A0(new_new_n607_), .A1(new_new_n245_), .B0(new_new_n167_), .Y(new_new_n608_));
  OR2        g0586(.A(i_6_), .B(i_10_), .Y(new_new_n609_));
  NO2        g0587(.A(new_new_n609_), .B(new_new_n23_), .Y(new_new_n610_));
  OR3        g0588(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n611_));
  NO3        g0589(.A(new_new_n611_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n612_));
  INV        g0590(.A(new_new_n205_), .Y(new_new_n613_));
  NO2        g0591(.A(new_new_n612_), .B(new_new_n610_), .Y(new_new_n614_));
  OA220      g0592(.A0(new_new_n614_), .A1(new_new_n578_), .B0(new_new_n608_), .B1(new_new_n279_), .Y(new_new_n615_));
  AOI210     g0593(.A0(new_new_n615_), .A1(new_new_n606_), .B0(new_new_n64_), .Y(new_new_n616_));
  NOi21      g0594(.An(i_11_), .B(i_7_), .Y(new_new_n617_));
  AO210      g0595(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n618_), .B(new_new_n617_), .Y(new_new_n619_));
  NA2        g0597(.A(new_new_n619_), .B(new_new_n213_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n620_), .B(new_new_n64_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n622_));
  AO210      g0600(.A0(new_new_n622_), .A1(new_new_n380_), .B0(new_new_n41_), .Y(new_new_n623_));
  NO3        g0601(.A(new_new_n268_), .B(new_new_n215_), .C(new_new_n595_), .Y(new_new_n624_));
  OAI210     g0602(.A0(new_new_n624_), .A1(new_new_n235_), .B0(new_new_n64_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n404_), .B(new_new_n31_), .Y(new_new_n626_));
  OR2        g0604(.A(new_new_n215_), .B(new_new_n112_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n627_), .B(new_new_n626_), .Y(new_new_n628_));
  NO2        g0606(.A(new_new_n64_), .B(i_9_), .Y(new_new_n629_));
  NO2        g0607(.A(new_new_n629_), .B(i_4_), .Y(new_new_n630_));
  NA2        g0608(.A(new_new_n630_), .B(new_new_n628_), .Y(new_new_n631_));
  NO2        g0609(.A(i_1_), .B(i_12_), .Y(new_new_n632_));
  NA3        g0610(.A(new_new_n631_), .B(new_new_n625_), .C(new_new_n623_), .Y(new_new_n633_));
  OAI210     g0611(.A0(new_new_n633_), .A1(new_new_n621_), .B0(i_6_), .Y(new_new_n634_));
  NO2        g0612(.A(i_6_), .B(i_11_), .Y(new_new_n635_));
  INV        g0613(.A(new_new_n446_), .Y(new_new_n636_));
  NO4        g0614(.A(new_new_n223_), .B(new_new_n133_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n637_));
  NA2        g0615(.A(new_new_n637_), .B(new_new_n629_), .Y(new_new_n638_));
  NA2        g0616(.A(new_new_n245_), .B(i_6_), .Y(new_new_n639_));
  NO3        g0617(.A(new_new_n609_), .B(new_new_n242_), .C(new_new_n23_), .Y(new_new_n640_));
  AOI210     g0618(.A0(i_1_), .A1(new_new_n269_), .B0(new_new_n640_), .Y(new_new_n641_));
  OAI210     g0619(.A0(new_new_n641_), .A1(new_new_n45_), .B0(new_new_n638_), .Y(new_new_n642_));
  NA3        g0620(.A(new_new_n534_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n643_));
  INV        g0621(.A(i_2_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n143_), .B(i_9_), .Y(new_new_n645_));
  NA3        g0623(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n47_), .B(i_1_), .Y(new_new_n647_));
  NA3        g0625(.A(new_new_n647_), .B(new_new_n278_), .C(new_new_n45_), .Y(new_new_n648_));
  OAI220     g0626(.A0(new_new_n648_), .A1(new_new_n646_), .B0(new_new_n645_), .B1(new_new_n644_), .Y(new_new_n649_));
  NA3        g0627(.A(new_new_n629_), .B(new_new_n320_), .C(i_6_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n650_), .B(new_new_n23_), .Y(new_new_n651_));
  AOI210     g0629(.A0(new_new_n468_), .A1(new_new_n415_), .B0(new_new_n249_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n600_), .Y(new_new_n653_));
  NAi21      g0631(.An(new_new_n643_), .B(new_new_n95_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n647_), .B(new_new_n278_), .Y(new_new_n655_));
  NO2        g0633(.A(i_11_), .B(new_new_n37_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n656_), .B(new_new_n24_), .Y(new_new_n657_));
  OAI210     g0635(.A0(new_new_n657_), .A1(new_new_n655_), .B0(new_new_n654_), .Y(new_new_n658_));
  OR4        g0636(.A(new_new_n658_), .B(new_new_n653_), .C(new_new_n651_), .D(new_new_n649_), .Y(new_new_n659_));
  NO3        g0637(.A(new_new_n659_), .B(new_new_n642_), .C(new_new_n636_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n245_), .B(new_new_n105_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n617_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(i_1_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n663_), .B(new_new_n611_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n410_), .B(new_new_n87_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n664_), .B(new_new_n47_), .Y(new_new_n666_));
  NA2        g0644(.A(i_3_), .B(new_new_n198_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n667_), .B(new_new_n119_), .Y(new_new_n668_));
  AN2        g0646(.A(new_new_n668_), .B(new_new_n540_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n242_), .B(new_new_n45_), .Y(new_new_n670_));
  NO3        g0648(.A(new_new_n670_), .B(new_new_n313_), .C(new_new_n246_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n122_), .B(new_new_n37_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n672_), .B(i_6_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n87_), .B(i_9_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n64_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n675_), .B(new_new_n632_), .Y(new_new_n676_));
  NO4        g0654(.A(new_new_n676_), .B(new_new_n673_), .C(new_new_n671_), .D(i_4_), .Y(new_new_n677_));
  NA2        g0655(.A(i_1_), .B(i_3_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n447_), .B(new_new_n96_), .Y(new_new_n679_));
  AOI210     g0657(.A0(new_new_n670_), .A1(new_new_n568_), .B0(new_new_n679_), .Y(new_new_n680_));
  NO2        g0658(.A(new_new_n680_), .B(new_new_n678_), .Y(new_new_n681_));
  NO3        g0659(.A(new_new_n681_), .B(new_new_n677_), .C(new_new_n669_), .Y(new_new_n682_));
  NA4        g0660(.A(new_new_n682_), .B(new_new_n666_), .C(new_new_n660_), .D(new_new_n634_), .Y(new_new_n683_));
  NO3        g0661(.A(new_new_n470_), .B(i_3_), .C(i_7_), .Y(new_new_n684_));
  NOi21      g0662(.An(new_new_n684_), .B(i_10_), .Y(new_new_n685_));
  OA210      g0663(.A0(new_new_n685_), .A1(new_new_n253_), .B0(new_new_n87_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n373_), .B(new_new_n372_), .Y(new_new_n687_));
  NA3        g0665(.A(new_new_n477_), .B(new_new_n516_), .C(new_new_n47_), .Y(new_new_n688_));
  NA3        g0666(.A(new_new_n167_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n689_));
  NA3        g0667(.A(new_new_n689_), .B(new_new_n688_), .C(new_new_n687_), .Y(new_new_n690_));
  OAI210     g0668(.A0(new_new_n690_), .A1(new_new_n686_), .B0(i_1_), .Y(new_new_n691_));
  AOI210     g0669(.A0(new_new_n278_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n371_), .B(i_2_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n693_), .B(new_new_n692_), .Y(new_new_n694_));
  OAI210     g0672(.A0(new_new_n650_), .A1(new_new_n437_), .B0(new_new_n694_), .Y(new_new_n695_));
  INV        g0673(.A(new_new_n695_), .Y(new_new_n696_));
  AOI210     g0674(.A0(new_new_n696_), .A1(new_new_n691_), .B0(i_13_), .Y(new_new_n697_));
  OR2        g0675(.A(i_11_), .B(i_7_), .Y(new_new_n698_));
  NA3        g0676(.A(new_new_n698_), .B(new_new_n110_), .C(new_new_n143_), .Y(new_new_n699_));
  AOI220     g0677(.A0(new_new_n464_), .A1(new_new_n167_), .B0(new_new_n440_), .B1(new_new_n143_), .Y(new_new_n700_));
  OAI210     g0678(.A0(new_new_n700_), .A1(new_new_n45_), .B0(new_new_n699_), .Y(new_new_n701_));
  AOI210     g0679(.A0(new_new_n646_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n471_), .B(new_new_n24_), .Y(new_new_n703_));
  AOI220     g0681(.A0(new_new_n703_), .A1(new_new_n665_), .B0(new_new_n253_), .B1(new_new_n136_), .Y(new_new_n704_));
  OAI220     g0682(.A0(new_new_n704_), .A1(new_new_n41_), .B0(new_new_n1058_), .B1(new_new_n96_), .Y(new_new_n705_));
  AOI210     g0683(.A0(new_new_n701_), .A1(new_new_n333_), .B0(new_new_n705_), .Y(new_new_n706_));
  INV        g0684(.A(new_new_n119_), .Y(new_new_n707_));
  AOI220     g0685(.A0(new_new_n707_), .A1(new_new_n73_), .B0(new_new_n386_), .B1(new_new_n647_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n708_), .B(new_new_n250_), .Y(new_new_n709_));
  AOI210     g0687(.A0(new_new_n437_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n710_));
  NOi31      g0688(.An(new_new_n710_), .B(new_new_n594_), .C(new_new_n45_), .Y(new_new_n711_));
  NA2        g0689(.A(new_new_n132_), .B(i_13_), .Y(new_new_n712_));
  NO2        g0690(.A(new_new_n646_), .B(new_new_n119_), .Y(new_new_n713_));
  INV        g0691(.A(new_new_n713_), .Y(new_new_n714_));
  OAI220     g0692(.A0(new_new_n714_), .A1(new_new_n72_), .B0(new_new_n712_), .B1(new_new_n692_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n26_), .B(new_new_n198_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n716_), .B(i_7_), .Y(new_new_n717_));
  NO3        g0695(.A(new_new_n471_), .B(new_new_n245_), .C(new_new_n87_), .Y(new_new_n718_));
  NA2        g0696(.A(new_new_n718_), .B(new_new_n717_), .Y(new_new_n719_));
  AOI220     g0697(.A0(new_new_n386_), .A1(new_new_n647_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n720_));
  OAI220     g0698(.A0(new_new_n720_), .A1(new_new_n598_), .B0(new_new_n719_), .B1(new_new_n613_), .Y(new_new_n721_));
  NO4        g0699(.A(new_new_n721_), .B(new_new_n715_), .C(new_new_n711_), .D(new_new_n709_), .Y(new_new_n722_));
  OR2        g0700(.A(i_11_), .B(i_6_), .Y(new_new_n723_));
  NA3        g0701(.A(new_new_n597_), .B(new_new_n716_), .C(i_7_), .Y(new_new_n724_));
  AOI210     g0702(.A0(new_new_n724_), .A1(new_new_n714_), .B0(new_new_n723_), .Y(new_new_n725_));
  NA3        g0703(.A(new_new_n404_), .B(new_new_n602_), .C(new_new_n101_), .Y(new_new_n726_));
  NA2        g0704(.A(new_new_n635_), .B(i_13_), .Y(new_new_n727_));
  NA2        g0705(.A(new_new_n106_), .B(new_new_n716_), .Y(new_new_n728_));
  NAi21      g0706(.An(i_11_), .B(i_12_), .Y(new_new_n729_));
  NOi41      g0707(.An(new_new_n115_), .B(new_new_n729_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n730_));
  NO3        g0708(.A(new_new_n471_), .B(new_new_n579_), .C(new_new_n603_), .Y(new_new_n731_));
  AOI220     g0709(.A0(new_new_n731_), .A1(new_new_n317_), .B0(new_new_n730_), .B1(new_new_n728_), .Y(new_new_n732_));
  NA3        g0710(.A(new_new_n732_), .B(new_new_n727_), .C(new_new_n726_), .Y(new_new_n733_));
  OAI210     g0711(.A0(new_new_n733_), .A1(new_new_n725_), .B0(new_new_n64_), .Y(new_new_n734_));
  NO2        g0712(.A(i_2_), .B(i_12_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n370_), .B(new_new_n735_), .Y(new_new_n736_));
  NA2        g0714(.A(i_8_), .B(new_new_n25_), .Y(new_new_n737_));
  NO3        g0715(.A(new_new_n737_), .B(i_3_), .C(new_new_n597_), .Y(new_new_n738_));
  OAI210     g0716(.A0(new_new_n738_), .A1(new_new_n372_), .B0(new_new_n370_), .Y(new_new_n739_));
  NO2        g0717(.A(new_new_n133_), .B(i_2_), .Y(new_new_n740_));
  NA2        g0718(.A(new_new_n740_), .B(new_new_n632_), .Y(new_new_n741_));
  NA3        g0719(.A(new_new_n741_), .B(new_new_n739_), .C(new_new_n736_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n742_), .B(new_new_n46_), .C(new_new_n234_), .Y(new_new_n743_));
  NA4        g0721(.A(new_new_n743_), .B(new_new_n734_), .C(new_new_n722_), .D(new_new_n706_), .Y(new_new_n744_));
  OR4        g0722(.A(new_new_n744_), .B(new_new_n697_), .C(new_new_n683_), .D(new_new_n616_), .Y(men5));
  NA2        g0723(.A(new_new_n662_), .B(new_new_n281_), .Y(new_new_n746_));
  AN2        g0724(.A(new_new_n24_), .B(i_10_), .Y(new_new_n747_));
  NA3        g0725(.A(new_new_n747_), .B(new_new_n735_), .C(new_new_n112_), .Y(new_new_n748_));
  NO2        g0726(.A(new_new_n598_), .B(i_11_), .Y(new_new_n749_));
  NA2        g0727(.A(new_new_n90_), .B(new_new_n749_), .Y(new_new_n750_));
  NA3        g0728(.A(new_new_n750_), .B(new_new_n748_), .C(new_new_n746_), .Y(new_new_n751_));
  NO3        g0729(.A(i_11_), .B(new_new_n245_), .C(i_13_), .Y(new_new_n752_));
  NO2        g0730(.A(new_new_n129_), .B(new_new_n23_), .Y(new_new_n753_));
  NA2        g0731(.A(i_12_), .B(i_8_), .Y(new_new_n754_));
  OAI210     g0732(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n754_), .Y(new_new_n755_));
  INV        g0733(.A(new_new_n436_), .Y(new_new_n756_));
  AOI220     g0734(.A0(new_new_n320_), .A1(new_new_n572_), .B0(new_new_n755_), .B1(new_new_n753_), .Y(new_new_n757_));
  INV        g0735(.A(new_new_n757_), .Y(new_new_n758_));
  NO2        g0736(.A(new_new_n758_), .B(new_new_n751_), .Y(new_new_n759_));
  INV        g0737(.A(new_new_n176_), .Y(new_new_n760_));
  INV        g0738(.A(new_new_n253_), .Y(new_new_n761_));
  OAI210     g0739(.A0(new_new_n693_), .A1(new_new_n438_), .B0(new_new_n115_), .Y(new_new_n762_));
  AOI210     g0740(.A0(new_new_n762_), .A1(new_new_n761_), .B0(new_new_n760_), .Y(new_new_n763_));
  NO2        g0741(.A(new_new_n447_), .B(new_new_n26_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n764_), .B(new_new_n415_), .Y(new_new_n765_));
  NA2        g0743(.A(new_new_n765_), .B(i_2_), .Y(new_new_n766_));
  INV        g0744(.A(new_new_n766_), .Y(new_new_n767_));
  AOI210     g0745(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n411_), .Y(new_new_n768_));
  AOI210     g0746(.A0(new_new_n768_), .A1(new_new_n767_), .B0(new_new_n763_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n195_), .B(new_new_n130_), .Y(new_new_n770_));
  OAI210     g0748(.A0(new_new_n770_), .A1(new_new_n753_), .B0(i_2_), .Y(new_new_n771_));
  INV        g0749(.A(new_new_n177_), .Y(new_new_n772_));
  NO3        g0750(.A(new_new_n618_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n772_), .A1(new_new_n90_), .B0(new_new_n773_), .Y(new_new_n774_));
  AOI210     g0752(.A0(new_new_n774_), .A1(new_new_n771_), .B0(new_new_n198_), .Y(new_new_n775_));
  OA210      g0753(.A0(new_new_n619_), .A1(new_new_n131_), .B0(i_13_), .Y(new_new_n776_));
  NA2        g0754(.A(new_new_n205_), .B(new_new_n208_), .Y(new_new_n777_));
  NA2        g0755(.A(new_new_n157_), .B(new_new_n595_), .Y(new_new_n778_));
  AOI210     g0756(.A0(new_new_n778_), .A1(new_new_n777_), .B0(new_new_n375_), .Y(new_new_n779_));
  AOI210     g0757(.A0(new_new_n215_), .A1(new_new_n153_), .B0(new_new_n516_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n780_), .B(new_new_n415_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n782_));
  INV        g0760(.A(new_new_n305_), .Y(new_new_n783_));
  NA4        g0761(.A(new_new_n783_), .B(new_new_n310_), .C(new_new_n129_), .D(new_new_n43_), .Y(new_new_n784_));
  OAI210     g0762(.A0(new_new_n784_), .A1(new_new_n782_), .B0(new_new_n781_), .Y(new_new_n785_));
  NO4        g0763(.A(new_new_n785_), .B(new_new_n779_), .C(new_new_n776_), .D(new_new_n775_), .Y(new_new_n786_));
  NA2        g0764(.A(new_new_n572_), .B(new_new_n28_), .Y(new_new_n787_));
  NA2        g0765(.A(new_new_n752_), .B(new_new_n288_), .Y(new_new_n788_));
  NA2        g0766(.A(new_new_n788_), .B(new_new_n787_), .Y(new_new_n789_));
  NO2        g0767(.A(new_new_n63_), .B(i_12_), .Y(new_new_n790_));
  NO2        g0768(.A(new_new_n790_), .B(new_new_n131_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n791_), .B(new_new_n595_), .Y(new_new_n792_));
  AOI220     g0770(.A0(new_new_n792_), .A1(new_new_n36_), .B0(new_new_n789_), .B1(new_new_n47_), .Y(new_new_n793_));
  NA4        g0771(.A(new_new_n793_), .B(new_new_n786_), .C(new_new_n769_), .D(new_new_n759_), .Y(men6));
  NO3        g0772(.A(new_new_n264_), .B(new_new_n312_), .C(i_1_), .Y(new_new_n795_));
  NO2        g0773(.A(new_new_n190_), .B(new_new_n144_), .Y(new_new_n796_));
  OAI210     g0774(.A0(new_new_n796_), .A1(new_new_n795_), .B0(new_new_n740_), .Y(new_new_n797_));
  NA4        g0775(.A(new_new_n388_), .B(new_new_n476_), .C(new_new_n72_), .D(new_new_n105_), .Y(new_new_n798_));
  INV        g0776(.A(new_new_n798_), .Y(new_new_n799_));
  NO2        g0777(.A(new_new_n229_), .B(new_new_n481_), .Y(new_new_n800_));
  NO2        g0778(.A(i_11_), .B(i_9_), .Y(new_new_n801_));
  NO2        g0779(.A(new_new_n799_), .B(new_new_n331_), .Y(new_new_n802_));
  AO210      g0780(.A0(new_new_n802_), .A1(new_new_n797_), .B0(i_12_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n376_), .B(new_new_n336_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n579_), .B(new_new_n64_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n685_), .B(new_new_n72_), .Y(new_new_n806_));
  BUFFER     g0784(.A(new_new_n622_), .Y(new_new_n807_));
  NA4        g0785(.A(new_new_n807_), .B(new_new_n806_), .C(new_new_n805_), .D(new_new_n804_), .Y(new_new_n808_));
  INV        g0786(.A(new_new_n202_), .Y(new_new_n809_));
  AOI220     g0787(.A0(new_new_n809_), .A1(new_new_n801_), .B0(new_new_n808_), .B1(new_new_n74_), .Y(new_new_n810_));
  INV        g0788(.A(new_new_n330_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n76_), .B(new_new_n136_), .Y(new_new_n812_));
  INV        g0790(.A(new_new_n129_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n813_), .B(new_new_n47_), .Y(new_new_n814_));
  AOI210     g0792(.A0(new_new_n814_), .A1(new_new_n812_), .B0(new_new_n811_), .Y(new_new_n815_));
  NO3        g0793(.A(new_new_n260_), .B(new_new_n137_), .C(i_9_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n816_), .B(new_new_n790_), .Y(new_new_n817_));
  AOI210     g0795(.A0(new_new_n817_), .A1(new_new_n514_), .B0(new_new_n190_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n32_), .B(i_11_), .Y(new_new_n819_));
  NA3        g0797(.A(new_new_n819_), .B(new_new_n466_), .C(new_new_n388_), .Y(new_new_n820_));
  NAi32      g0798(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n723_), .B(new_new_n821_), .Y(new_new_n822_));
  OAI210     g0800(.A0(new_new_n684_), .A1(new_new_n560_), .B0(new_new_n559_), .Y(new_new_n823_));
  NAi31      g0801(.An(new_new_n822_), .B(new_new_n823_), .C(new_new_n820_), .Y(new_new_n824_));
  OR3        g0802(.A(new_new_n824_), .B(new_new_n818_), .C(new_new_n815_), .Y(new_new_n825_));
  NO2        g0803(.A(new_new_n698_), .B(i_2_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n827_), .B(new_new_n403_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n828_), .B(new_new_n826_), .Y(new_new_n829_));
  AO220      g0807(.A0(new_new_n363_), .A1(new_new_n353_), .B0(new_new_n390_), .B1(new_new_n595_), .Y(new_new_n830_));
  NA3        g0808(.A(new_new_n830_), .B(new_new_n265_), .C(i_7_), .Y(new_new_n831_));
  OR2        g0809(.A(new_new_n619_), .B(new_new_n438_), .Y(new_new_n832_));
  NA3        g0810(.A(new_new_n832_), .B(new_new_n152_), .C(new_new_n70_), .Y(new_new_n833_));
  AO210      g0811(.A0(new_new_n488_), .A1(new_new_n756_), .B0(new_new_n36_), .Y(new_new_n834_));
  NA4        g0812(.A(new_new_n834_), .B(new_new_n833_), .C(new_new_n831_), .D(new_new_n829_), .Y(new_new_n835_));
  NO2        g0813(.A(i_6_), .B(i_11_), .Y(new_new_n836_));
  AOI220     g0814(.A0(new_new_n836_), .A1(new_new_n559_), .B0(new_new_n800_), .B1(new_new_n717_), .Y(new_new_n837_));
  NA2        g0815(.A(new_new_n390_), .B(new_new_n71_), .Y(new_new_n838_));
  NA3        g0816(.A(new_new_n838_), .B(new_new_n837_), .C(new_new_n601_), .Y(new_new_n839_));
  AO210      g0817(.A0(new_new_n516_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n840_));
  NA3        g0818(.A(new_new_n840_), .B(new_new_n477_), .C(new_new_n226_), .Y(new_new_n841_));
  AOI210     g0819(.A0(new_new_n438_), .A1(new_new_n436_), .B0(new_new_n558_), .Y(new_new_n842_));
  NO2        g0820(.A(new_new_n609_), .B(new_new_n106_), .Y(new_new_n843_));
  OAI210     g0821(.A0(new_new_n843_), .A1(new_new_n116_), .B0(new_new_n401_), .Y(new_new_n844_));
  INV        g0822(.A(new_new_n586_), .Y(new_new_n845_));
  NA3        g0823(.A(new_new_n845_), .B(new_new_n330_), .C(i_7_), .Y(new_new_n846_));
  NA4        g0824(.A(new_new_n846_), .B(new_new_n844_), .C(new_new_n842_), .D(new_new_n841_), .Y(new_new_n847_));
  NO4        g0825(.A(new_new_n847_), .B(new_new_n839_), .C(new_new_n835_), .D(new_new_n825_), .Y(new_new_n848_));
  NA4        g0826(.A(new_new_n848_), .B(new_new_n810_), .C(new_new_n803_), .D(new_new_n382_), .Y(men3));
  NA2        g0827(.A(i_12_), .B(i_10_), .Y(new_new_n850_));
  NA2        g0828(.A(i_6_), .B(i_7_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n851_), .B(i_0_), .Y(new_new_n852_));
  NO2        g0830(.A(i_11_), .B(new_new_n245_), .Y(new_new_n853_));
  OAI210     g0831(.A0(new_new_n852_), .A1(new_new_n298_), .B0(new_new_n853_), .Y(new_new_n854_));
  NO2        g0832(.A(new_new_n854_), .B(new_new_n198_), .Y(new_new_n855_));
  NO3        g0833(.A(new_new_n443_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n856_));
  OA210      g0834(.A0(new_new_n856_), .A1(new_new_n855_), .B0(new_new_n178_), .Y(new_new_n857_));
  NA2        g0835(.A(new_new_n601_), .B(new_new_n374_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n858_), .B(new_new_n40_), .Y(new_new_n859_));
  NOi21      g0837(.An(new_new_n100_), .B(new_new_n765_), .Y(new_new_n860_));
  NO3        g0838(.A(new_new_n627_), .B(new_new_n447_), .C(new_new_n136_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n404_), .B(new_new_n46_), .Y(new_new_n862_));
  AN2        g0840(.A(new_new_n445_), .B(new_new_n56_), .Y(new_new_n863_));
  NO3        g0841(.A(new_new_n863_), .B(new_new_n861_), .C(new_new_n860_), .Y(new_new_n864_));
  AOI210     g0842(.A0(new_new_n864_), .A1(new_new_n859_), .B0(new_new_n49_), .Y(new_new_n865_));
  NO4        g0843(.A(new_new_n378_), .B(new_new_n384_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n190_), .B(new_new_n568_), .Y(new_new_n867_));
  NOi21      g0845(.An(new_new_n867_), .B(new_new_n866_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n710_), .B(new_new_n674_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n334_), .B(new_new_n429_), .Y(new_new_n870_));
  OAI220     g0848(.A0(new_new_n870_), .A1(new_new_n869_), .B0(new_new_n868_), .B1(new_new_n64_), .Y(new_new_n871_));
  NOi21      g0849(.An(i_5_), .B(i_9_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n872_), .B(new_new_n434_), .Y(new_new_n873_));
  BUFFER     g0851(.A(new_new_n278_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n874_), .B(new_new_n468_), .Y(new_new_n875_));
  NO3        g0853(.A(new_new_n407_), .B(new_new_n278_), .C(new_new_n74_), .Y(new_new_n876_));
  NO2        g0854(.A(new_new_n179_), .B(new_new_n153_), .Y(new_new_n877_));
  AOI210     g0855(.A0(new_new_n877_), .A1(new_new_n252_), .B0(new_new_n876_), .Y(new_new_n878_));
  OAI220     g0856(.A0(new_new_n878_), .A1(new_new_n185_), .B0(new_new_n875_), .B1(new_new_n873_), .Y(new_new_n879_));
  NO4        g0857(.A(new_new_n879_), .B(new_new_n871_), .C(new_new_n865_), .D(new_new_n857_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n190_), .B(new_new_n24_), .Y(new_new_n881_));
  NO2        g0859(.A(new_new_n388_), .B(new_new_n299_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n882_), .B(new_new_n713_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n569_), .B(i_0_), .Y(new_new_n884_));
  NO3        g0862(.A(new_new_n884_), .B(new_new_n385_), .C(new_new_n90_), .Y(new_new_n885_));
  NO4        g0863(.A(new_new_n585_), .B(new_new_n223_), .C(new_new_n411_), .D(new_new_n403_), .Y(new_new_n886_));
  AOI210     g0864(.A0(new_new_n886_), .A1(i_11_), .B0(new_new_n885_), .Y(new_new_n887_));
  AN2        g0865(.A(new_new_n100_), .B(new_new_n251_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n752_), .B(new_new_n331_), .Y(new_new_n889_));
  AOI210     g0867(.A0(new_new_n477_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n890_));
  OAI220     g0868(.A0(new_new_n890_), .A1(new_new_n889_), .B0(new_new_n657_), .B1(new_new_n536_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n262_), .B(new_new_n159_), .Y(new_new_n892_));
  NA2        g0870(.A(i_0_), .B(i_10_), .Y(new_new_n893_));
  INV        g0871(.A(new_new_n539_), .Y(new_new_n894_));
  NO4        g0872(.A(new_new_n119_), .B(new_new_n59_), .C(new_new_n667_), .D(i_5_), .Y(new_new_n895_));
  AO220      g0873(.A0(new_new_n895_), .A1(new_new_n894_), .B0(new_new_n892_), .B1(i_6_), .Y(new_new_n896_));
  AOI220     g0874(.A0(new_new_n334_), .A1(new_new_n102_), .B0(new_new_n190_), .B1(new_new_n85_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n563_), .B(i_4_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n193_), .B(new_new_n208_), .Y(new_new_n899_));
  OAI220     g0877(.A0(new_new_n899_), .A1(new_new_n889_), .B0(new_new_n898_), .B1(new_new_n897_), .Y(new_new_n900_));
  NO4        g0878(.A(new_new_n900_), .B(new_new_n896_), .C(new_new_n891_), .D(new_new_n888_), .Y(new_new_n901_));
  NA3        g0879(.A(new_new_n901_), .B(new_new_n887_), .C(new_new_n883_), .Y(new_new_n902_));
  NA2        g0880(.A(i_11_), .B(i_9_), .Y(new_new_n903_));
  NO2        g0881(.A(new_new_n49_), .B(i_7_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n389_), .B(new_new_n183_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n905_), .B(new_new_n166_), .Y(new_new_n906_));
  NO2        g0884(.A(new_new_n903_), .B(new_new_n74_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n179_), .B(i_0_), .Y(new_new_n908_));
  AOI210     g0886(.A0(new_new_n373_), .A1(new_new_n42_), .B0(new_new_n400_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n909_), .B(new_new_n873_), .Y(new_new_n910_));
  NO2        g0888(.A(new_new_n910_), .B(new_new_n906_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n656_), .B(new_new_n126_), .Y(new_new_n912_));
  NO2        g0890(.A(i_6_), .B(new_new_n912_), .Y(new_new_n913_));
  AOI210     g0891(.A0(new_new_n437_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n914_));
  NA2        g0892(.A(new_new_n176_), .B(new_new_n107_), .Y(new_new_n915_));
  NOi32      g0893(.An(new_new_n914_), .Bn(new_new_n193_), .C(new_new_n915_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n602_), .B(new_new_n331_), .Y(new_new_n917_));
  NO2        g0895(.A(new_new_n917_), .B(new_new_n862_), .Y(new_new_n918_));
  NO3        g0896(.A(new_new_n918_), .B(new_new_n916_), .C(new_new_n913_), .Y(new_new_n919_));
  NOi21      g0897(.An(i_7_), .B(i_5_), .Y(new_new_n920_));
  NOi31      g0898(.An(new_new_n920_), .B(i_0_), .C(new_new_n729_), .Y(new_new_n921_));
  NO3        g0899(.A(new_new_n396_), .B(new_new_n366_), .C(new_new_n362_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n272_), .B(new_new_n321_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n729_), .B(new_new_n267_), .Y(new_new_n924_));
  AOI210     g0902(.A0(new_new_n924_), .A1(new_new_n923_), .B0(new_new_n922_), .Y(new_new_n925_));
  NA3        g0903(.A(new_new_n925_), .B(new_new_n919_), .C(new_new_n911_), .Y(new_new_n926_));
  NO2        g0904(.A(new_new_n881_), .B(new_new_n248_), .Y(new_new_n927_));
  AN2        g0905(.A(new_new_n333_), .B(new_new_n331_), .Y(new_new_n928_));
  AN2        g0906(.A(new_new_n928_), .B(new_new_n877_), .Y(new_new_n929_));
  OAI210     g0907(.A0(new_new_n929_), .A1(new_new_n927_), .B0(i_10_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n850_), .B(new_new_n320_), .Y(new_new_n931_));
  OA210      g0909(.A0(new_new_n466_), .A1(new_new_n232_), .B0(new_new_n465_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n931_), .B(new_new_n907_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n265_), .B(new_new_n47_), .Y(new_new_n934_));
  NA2        g0912(.A(new_new_n907_), .B(new_new_n310_), .Y(new_new_n935_));
  OAI210     g0913(.A0(new_new_n934_), .A1(new_new_n192_), .B0(new_new_n935_), .Y(new_new_n936_));
  NA2        g0914(.A(new_new_n936_), .B(new_new_n466_), .Y(new_new_n937_));
  NO3        g0915(.A(new_new_n585_), .B(new_new_n361_), .C(new_new_n24_), .Y(new_new_n938_));
  INV        g0916(.A(new_new_n938_), .Y(new_new_n939_));
  NAi21      g0917(.An(i_9_), .B(i_5_), .Y(new_new_n940_));
  NO2        g0918(.A(new_new_n940_), .B(new_new_n396_), .Y(new_new_n941_));
  NA2        g0919(.A(new_new_n941_), .B(new_new_n619_), .Y(new_new_n942_));
  OAI220     g0920(.A0(new_new_n942_), .A1(new_new_n87_), .B0(new_new_n939_), .B1(new_new_n177_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n943_), .B(new_new_n519_), .Y(new_new_n944_));
  NA4        g0922(.A(new_new_n944_), .B(new_new_n937_), .C(new_new_n933_), .D(new_new_n930_), .Y(new_new_n945_));
  NO3        g0923(.A(new_new_n945_), .B(new_new_n926_), .C(new_new_n902_), .Y(new_new_n946_));
  NO2        g0924(.A(i_0_), .B(new_new_n729_), .Y(new_new_n947_));
  NA2        g0925(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n948_));
  INV        g0926(.A(new_new_n948_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n950_));
  AO220      g0928(.A0(new_new_n950_), .A1(new_new_n949_), .B0(new_new_n947_), .B1(new_new_n178_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n805_), .A1(new_new_n687_), .B0(new_new_n915_), .Y(new_new_n952_));
  AOI210     g0930(.A0(new_new_n951_), .A1(new_new_n350_), .B0(new_new_n952_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n740_), .B(new_new_n151_), .Y(new_new_n954_));
  INV        g0932(.A(new_new_n954_), .Y(new_new_n955_));
  NA3        g0933(.A(new_new_n955_), .B(new_new_n674_), .C(new_new_n74_), .Y(new_new_n956_));
  NO2        g0934(.A(new_new_n823_), .B(new_new_n396_), .Y(new_new_n957_));
  NA3        g0935(.A(new_new_n852_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n958_));
  NA2        g0936(.A(new_new_n853_), .B(i_9_), .Y(new_new_n959_));
  AOI210     g0937(.A0(new_new_n958_), .A1(new_new_n493_), .B0(new_new_n959_), .Y(new_new_n960_));
  OAI210     g0938(.A0(new_new_n252_), .A1(i_9_), .B0(new_new_n239_), .Y(new_new_n961_));
  AOI210     g0939(.A0(new_new_n961_), .A1(new_new_n884_), .B0(new_new_n159_), .Y(new_new_n962_));
  NO3        g0940(.A(new_new_n962_), .B(new_new_n960_), .C(new_new_n957_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n963_), .B(new_new_n956_), .C(new_new_n953_), .Y(new_new_n964_));
  NA2        g0942(.A(new_new_n928_), .B(new_new_n375_), .Y(new_new_n965_));
  AOI210     g0943(.A0(new_new_n304_), .A1(new_new_n168_), .B0(new_new_n965_), .Y(new_new_n966_));
  NA3        g0944(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n967_));
  NA2        g0945(.A(new_new_n904_), .B(new_new_n482_), .Y(new_new_n968_));
  AOI210     g0946(.A0(new_new_n967_), .A1(new_new_n168_), .B0(new_new_n968_), .Y(new_new_n969_));
  NO2        g0947(.A(new_new_n969_), .B(new_new_n966_), .Y(new_new_n970_));
  NO3        g0948(.A(new_new_n893_), .B(new_new_n872_), .C(new_new_n195_), .Y(new_new_n971_));
  AOI220     g0949(.A0(new_new_n971_), .A1(i_11_), .B0(new_new_n564_), .B1(new_new_n76_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n217_), .B(new_new_n384_), .C(i_0_), .Y(new_new_n973_));
  OAI210     g0951(.A0(new_new_n973_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n974_));
  INV        g0952(.A(new_new_n226_), .Y(new_new_n975_));
  OAI220     g0953(.A0(new_new_n530_), .A1(new_new_n144_), .B0(new_new_n639_), .B1(new_new_n613_), .Y(new_new_n976_));
  NA3        g0954(.A(new_new_n976_), .B(new_new_n391_), .C(new_new_n975_), .Y(new_new_n977_));
  NA4        g0955(.A(new_new_n977_), .B(new_new_n974_), .C(new_new_n972_), .D(new_new_n970_), .Y(new_new_n978_));
  NO2        g0956(.A(new_new_n250_), .B(new_new_n96_), .Y(new_new_n979_));
  AOI210     g0957(.A0(new_new_n979_), .A1(new_new_n947_), .B0(new_new_n113_), .Y(new_new_n980_));
  AOI220     g0958(.A0(new_new_n920_), .A1(new_new_n482_), .B0(new_new_n852_), .B1(new_new_n169_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n353_), .B(new_new_n180_), .Y(new_new_n982_));
  OA220      g0960(.A0(new_new_n982_), .A1(new_new_n981_), .B0(new_new_n980_), .B1(i_5_), .Y(new_new_n983_));
  AOI210     g0961(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n984_));
  NA2        g0962(.A(new_new_n984_), .B(new_new_n932_), .Y(new_new_n985_));
  NA3        g0963(.A(new_new_n610_), .B(new_new_n190_), .C(new_new_n85_), .Y(new_new_n986_));
  INV        g0964(.A(new_new_n986_), .Y(new_new_n987_));
  NO3        g0965(.A(new_new_n862_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n487_), .B(new_new_n480_), .Y(new_new_n989_));
  NO3        g0967(.A(new_new_n989_), .B(new_new_n988_), .C(new_new_n987_), .Y(new_new_n990_));
  NA3        g0968(.A(new_new_n388_), .B(new_new_n176_), .C(new_new_n175_), .Y(new_new_n991_));
  NA3        g0969(.A(new_new_n904_), .B(new_new_n298_), .C(new_new_n239_), .Y(new_new_n992_));
  NA2        g0970(.A(new_new_n992_), .B(new_new_n991_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n903_), .B(new_new_n226_), .C(new_new_n195_), .Y(new_new_n994_));
  NO2        g0972(.A(new_new_n994_), .B(new_new_n993_), .Y(new_new_n995_));
  NA4        g0973(.A(new_new_n995_), .B(new_new_n990_), .C(new_new_n985_), .D(new_new_n983_), .Y(new_new_n996_));
  INV        g0974(.A(new_new_n612_), .Y(new_new_n997_));
  NO3        g0975(.A(new_new_n997_), .B(new_new_n554_), .C(new_new_n347_), .Y(new_new_n998_));
  NO2        g0976(.A(new_new_n87_), .B(i_5_), .Y(new_new_n999_));
  NA3        g0977(.A(new_new_n853_), .B(new_new_n114_), .C(new_new_n129_), .Y(new_new_n1000_));
  INV        g0978(.A(new_new_n1000_), .Y(new_new_n1001_));
  AOI210     g0979(.A0(new_new_n1001_), .A1(new_new_n999_), .B0(new_new_n998_), .Y(new_new_n1002_));
  NAi21      g0980(.An(new_new_n249_), .B(new_new_n250_), .Y(new_new_n1003_));
  NO4        g0981(.A(new_new_n248_), .B(new_new_n217_), .C(i_0_), .D(i_12_), .Y(new_new_n1004_));
  AOI220     g0982(.A0(new_new_n1004_), .A1(new_new_n1003_), .B0(new_new_n799_), .B1(new_new_n180_), .Y(new_new_n1005_));
  AN2        g0983(.A(new_new_n893_), .B(new_new_n159_), .Y(new_new_n1006_));
  NO4        g0984(.A(new_new_n1006_), .B(i_12_), .C(new_new_n643_), .D(new_new_n136_), .Y(new_new_n1007_));
  NA2        g0985(.A(new_new_n1007_), .B(new_new_n226_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n102_), .B(new_new_n568_), .C(i_11_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n1009_), .B(new_new_n161_), .Y(new_new_n1010_));
  NA2        g0988(.A(new_new_n920_), .B(new_new_n464_), .Y(new_new_n1011_));
  NO2        g0989(.A(new_new_n1011_), .B(new_new_n675_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1012_), .A1(new_new_n908_), .B0(new_new_n1010_), .Y(new_new_n1013_));
  NA4        g0991(.A(new_new_n1013_), .B(new_new_n1008_), .C(new_new_n1005_), .D(new_new_n1002_), .Y(new_new_n1014_));
  NO4        g0992(.A(new_new_n1014_), .B(new_new_n996_), .C(new_new_n978_), .D(new_new_n964_), .Y(new_new_n1015_));
  OAI210     g0993(.A0(new_new_n826_), .A1(new_new_n819_), .B0(new_new_n37_), .Y(new_new_n1016_));
  NA3        g0994(.A(new_new_n914_), .B(new_new_n370_), .C(i_5_), .Y(new_new_n1017_));
  NA3        g0995(.A(new_new_n1017_), .B(new_new_n1016_), .C(new_new_n608_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n1018_), .B(new_new_n213_), .Y(new_new_n1019_));
  OAI210     g0997(.A0(new_new_n612_), .A1(new_new_n610_), .B0(new_new_n320_), .Y(new_new_n1020_));
  NAi31      g0998(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1021_));
  AOI210     g0999(.A0(new_new_n122_), .A1(new_new_n71_), .B0(new_new_n1021_), .Y(new_new_n1022_));
  NO2        g1000(.A(new_new_n1022_), .B(new_new_n640_), .Y(new_new_n1023_));
  NA2        g1001(.A(new_new_n1023_), .B(new_new_n1020_), .Y(new_new_n1024_));
  NO4        g1002(.A(new_new_n242_), .B(new_new_n150_), .C(new_new_n678_), .D(new_new_n37_), .Y(new_new_n1025_));
  NO2        g1003(.A(new_new_n1025_), .B(new_new_n886_), .Y(new_new_n1026_));
  OAI210     g1004(.A0(new_new_n1009_), .A1(new_new_n153_), .B0(new_new_n1026_), .Y(new_new_n1027_));
  AOI210     g1005(.A0(new_new_n1024_), .A1(new_new_n49_), .B0(new_new_n1027_), .Y(new_new_n1028_));
  AOI210     g1006(.A0(new_new_n1028_), .A1(new_new_n1019_), .B0(new_new_n74_), .Y(new_new_n1029_));
  NO2        g1007(.A(new_new_n561_), .B(new_new_n381_), .Y(new_new_n1030_));
  NO2        g1008(.A(new_new_n1030_), .B(new_new_n760_), .Y(new_new_n1031_));
  OAI210     g1009(.A0(new_new_n81_), .A1(new_new_n55_), .B0(new_new_n112_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n1032_), .B(new_new_n77_), .Y(new_new_n1033_));
  AOI210     g1011(.A0(new_new_n984_), .A1(new_new_n904_), .B0(new_new_n921_), .Y(new_new_n1034_));
  AOI210     g1012(.A0(new_new_n1034_), .A1(new_new_n1033_), .B0(new_new_n678_), .Y(new_new_n1035_));
  NA2        g1013(.A(new_new_n272_), .B(new_new_n58_), .Y(new_new_n1036_));
  AOI220     g1014(.A0(new_new_n1036_), .A1(new_new_n77_), .B0(new_new_n348_), .B1(new_new_n264_), .Y(new_new_n1037_));
  NO2        g1015(.A(new_new_n1037_), .B(new_new_n245_), .Y(new_new_n1038_));
  NA3        g1016(.A(new_new_n100_), .B(new_new_n312_), .C(new_new_n31_), .Y(new_new_n1039_));
  INV        g1017(.A(new_new_n1039_), .Y(new_new_n1040_));
  NO3        g1018(.A(new_new_n1040_), .B(new_new_n1038_), .C(new_new_n1035_), .Y(new_new_n1041_));
  OAI210     g1019(.A0(new_new_n280_), .A1(new_new_n164_), .B0(new_new_n90_), .Y(new_new_n1042_));
  NA3        g1020(.A(new_new_n764_), .B(new_new_n298_), .C(new_new_n81_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n1043_), .A1(new_new_n1042_), .B0(i_11_), .Y(new_new_n1044_));
  NA2        g1022(.A(new_new_n603_), .B(new_new_n223_), .Y(new_new_n1045_));
  OAI210     g1023(.A0(new_new_n1045_), .A1(new_new_n914_), .B0(new_new_n213_), .Y(new_new_n1046_));
  NA2        g1024(.A(new_new_n170_), .B(i_5_), .Y(new_new_n1047_));
  NO2        g1025(.A(new_new_n1046_), .B(new_new_n1047_), .Y(new_new_n1048_));
  NO4        g1026(.A(new_new_n940_), .B(new_new_n470_), .C(new_new_n261_), .D(new_new_n260_), .Y(new_new_n1049_));
  NO2        g1027(.A(new_new_n1049_), .B(new_new_n558_), .Y(new_new_n1050_));
  NO2        g1028(.A(new_new_n1050_), .B(new_new_n41_), .Y(new_new_n1051_));
  NO3        g1029(.A(new_new_n1051_), .B(new_new_n1048_), .C(new_new_n1044_), .Y(new_new_n1052_));
  OAI210     g1030(.A0(new_new_n1041_), .A1(i_4_), .B0(new_new_n1052_), .Y(new_new_n1053_));
  NO3        g1031(.A(new_new_n1053_), .B(new_new_n1031_), .C(new_new_n1029_), .Y(new_new_n1054_));
  NA4        g1032(.A(new_new_n1054_), .B(new_new_n1015_), .C(new_new_n946_), .D(new_new_n880_), .Y(men4));
  INV        g1033(.A(new_new_n702_), .Y(new_new_n1058_));
  INV        g1034(.A(new_new_n477_), .Y(new_new_n1059_));
endmodule


