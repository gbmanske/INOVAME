//Benchmark atmr_alu4_1266_0.125

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n129_, ori_ori_n130_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n962_, mai_mai_n963_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NOi21      o016(.An(i_12_), .B(i_13_), .Y(ori_ori_n39_));
  INV        o017(.A(ori_ori_n39_), .Y(ori_ori_n40_));
  NAi31      o018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n41_));
  INV        o019(.A(ori_ori_n35_), .Y(ori1));
  INV        o020(.A(i_11_), .Y(ori_ori_n43_));
  NO2        o021(.A(ori_ori_n43_), .B(i_6_), .Y(ori_ori_n44_));
  INV        o022(.A(i_2_), .Y(ori_ori_n45_));
  NA2        o023(.A(i_0_), .B(i_3_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_5_), .A1(ori_ori_n46_), .B0(ori_ori_n45_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_0_), .B(i_2_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NA2        o031(.A(ori_ori_n50_), .B(ori_ori_n44_), .Y(ori_ori_n54_));
  NO2        o032(.A(i_1_), .B(i_6_), .Y(ori_ori_n55_));
  NA2        o033(.A(i_8_), .B(i_7_), .Y(ori_ori_n56_));
  NAi21      o034(.An(i_2_), .B(i_7_), .Y(ori_ori_n57_));
  INV        o035(.A(i_1_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(i_6_), .Y(ori_ori_n59_));
  NA3        o037(.A(ori_ori_n59_), .B(ori_ori_n57_), .C(ori_ori_n31_), .Y(ori_ori_n60_));
  NA2        o038(.A(i_1_), .B(i_10_), .Y(ori_ori_n61_));
  NO2        o039(.A(ori_ori_n61_), .B(i_6_), .Y(ori_ori_n62_));
  NAi21      o040(.An(ori_ori_n62_), .B(ori_ori_n60_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n64_));
  AOI210     o042(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_1_), .B(i_6_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(ori_ori_n25_), .Y(ori_ori_n67_));
  INV        o045(.A(i_0_), .Y(ori_ori_n68_));
  NAi21      o046(.An(i_5_), .B(i_10_), .Y(ori_ori_n69_));
  NA2        o047(.A(i_5_), .B(i_9_), .Y(ori_ori_n70_));
  AOI210     o048(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n68_), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n71_), .B(ori_ori_n67_), .Y(ori_ori_n72_));
  INV        o050(.A(ori_ori_n72_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n73_), .A1(ori_ori_n63_), .B0(i_0_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_12_), .B(i_5_), .Y(ori_ori_n75_));
  INV        o053(.A(i_8_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n55_), .Y(ori_ori_n77_));
  INV        o055(.A(i_3_), .Y(ori_ori_n78_));
  NO2        o056(.A(i_3_), .B(i_7_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n78_), .B(ori_ori_n58_), .Y(ori_ori_n80_));
  INV        o058(.A(i_6_), .Y(ori_ori_n81_));
  OR4        o059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n82_));
  INV        o060(.A(ori_ori_n82_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_2_), .B(i_7_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n84_), .Y(ori_ori_n85_));
  OAI210     o063(.A0(ori_ori_n80_), .A1(ori_ori_n77_), .B0(ori_ori_n85_), .Y(ori_ori_n86_));
  NAi21      o064(.An(i_6_), .B(i_10_), .Y(ori_ori_n87_));
  NA2        o065(.A(i_6_), .B(i_9_), .Y(ori_ori_n88_));
  AOI210     o066(.A0(ori_ori_n88_), .A1(ori_ori_n87_), .B0(ori_ori_n58_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_2_), .B(i_6_), .Y(ori_ori_n90_));
  NO3        o068(.A(ori_ori_n90_), .B(ori_ori_n48_), .C(ori_ori_n25_), .Y(ori_ori_n91_));
  NO2        o069(.A(ori_ori_n91_), .B(ori_ori_n89_), .Y(ori_ori_n92_));
  AOI210     o070(.A0(ori_ori_n92_), .A1(ori_ori_n86_), .B0(ori_ori_n75_), .Y(ori_ori_n93_));
  AN3        o071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n94_));
  NAi21      o072(.An(i_6_), .B(i_11_), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n94_), .B(ori_ori_n32_), .Y(ori_ori_n96_));
  INV        o074(.A(i_7_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n45_), .B(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o076(.A(i_0_), .B(i_5_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n81_), .Y(ori_ori_n100_));
  NA2        o078(.A(i_12_), .B(i_3_), .Y(ori_ori_n101_));
  INV        o079(.A(ori_ori_n101_), .Y(ori_ori_n102_));
  NA3        o080(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n98_), .Y(ori_ori_n103_));
  NAi21      o081(.An(i_7_), .B(i_11_), .Y(ori_ori_n104_));
  NO3        o082(.A(ori_ori_n104_), .B(ori_ori_n87_), .C(ori_ori_n51_), .Y(ori_ori_n105_));
  AN2        o083(.A(i_2_), .B(i_10_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(i_7_), .Y(ori_ori_n107_));
  OR2        o085(.A(ori_ori_n75_), .B(ori_ori_n55_), .Y(ori_ori_n108_));
  NA2        o086(.A(i_12_), .B(i_7_), .Y(ori_ori_n109_));
  NA2        o087(.A(i_11_), .B(i_12_), .Y(ori_ori_n110_));
  NAi41      o088(.An(ori_ori_n105_), .B(ori_ori_n110_), .C(ori_ori_n103_), .D(ori_ori_n96_), .Y(ori_ori_n111_));
  NOi21      o089(.An(i_1_), .B(i_5_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(i_11_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n97_), .B(ori_ori_n37_), .Y(ori_ori_n114_));
  NA2        o092(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n115_));
  NA2        o093(.A(ori_ori_n115_), .B(ori_ori_n114_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n45_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n88_), .B(ori_ori_n87_), .Y(ori_ori_n118_));
  NAi21      o096(.An(i_3_), .B(i_8_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(ori_ori_n57_), .Y(ori_ori_n120_));
  NOi31      o098(.An(ori_ori_n120_), .B(ori_ori_n118_), .C(ori_ori_n117_), .Y(ori_ori_n121_));
  NO2        o099(.A(i_1_), .B(ori_ori_n81_), .Y(ori_ori_n122_));
  NO2        o100(.A(i_6_), .B(i_5_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(i_3_), .Y(ori_ori_n124_));
  AO210      o102(.A0(ori_ori_n124_), .A1(ori_ori_n46_), .B0(ori_ori_n122_), .Y(ori_ori_n125_));
  OAI220     o103(.A0(ori_ori_n125_), .A1(ori_ori_n104_), .B0(ori_ori_n121_), .B1(ori_ori_n113_), .Y(ori_ori_n126_));
  NO3        o104(.A(ori_ori_n126_), .B(ori_ori_n111_), .C(ori_ori_n93_), .Y(ori_ori_n127_));
  NA3        o105(.A(ori_ori_n127_), .B(ori_ori_n74_), .C(ori_ori_n54_), .Y(ori2));
  NO2        o106(.A(ori_ori_n58_), .B(ori_ori_n37_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n764_), .B(ori_ori_n129_), .Y(ori_ori_n130_));
  NA4        o108(.A(ori_ori_n130_), .B(ori_ori_n72_), .C(ori_ori_n64_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o109(.A(i_12_), .B(i_13_), .Y(ori_ori_n132_));
  NAi21      o110(.An(i_5_), .B(i_11_), .Y(ori_ori_n133_));
  NOi21      o111(.An(ori_ori_n132_), .B(ori_ori_n133_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_0_), .B(i_1_), .Y(ori_ori_n135_));
  NA2        o113(.A(i_2_), .B(i_3_), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n136_), .B(i_4_), .Y(ori_ori_n137_));
  NA3        o115(.A(ori_ori_n137_), .B(ori_ori_n135_), .C(ori_ori_n134_), .Y(ori_ori_n138_));
  NA2        o116(.A(i_1_), .B(i_5_), .Y(ori_ori_n139_));
  OR2        o117(.A(i_0_), .B(i_1_), .Y(ori_ori_n140_));
  NAi32      o118(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n141_));
  NOi21      o119(.An(i_4_), .B(i_10_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n142_), .B(ori_ori_n39_), .Y(ori_ori_n143_));
  NOi21      o121(.An(i_4_), .B(i_9_), .Y(ori_ori_n144_));
  NOi21      o122(.An(i_11_), .B(i_13_), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n145_), .B(ori_ori_n144_), .Y(ori_ori_n146_));
  NO2        o124(.A(i_4_), .B(i_5_), .Y(ori_ori_n147_));
  NAi21      o125(.An(i_12_), .B(i_11_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n148_), .B(i_13_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n68_), .B(ori_ori_n58_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n68_), .B(i_5_), .Y(ori_ori_n151_));
  NO2        o129(.A(i_13_), .B(i_10_), .Y(ori_ori_n152_));
  NA3        o130(.A(ori_ori_n152_), .B(ori_ori_n151_), .C(ori_ori_n43_), .Y(ori_ori_n153_));
  NO2        o131(.A(i_2_), .B(i_1_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n154_), .B(i_3_), .Y(ori_ori_n155_));
  NAi21      o133(.An(i_4_), .B(i_12_), .Y(ori_ori_n156_));
  INV        o134(.A(i_8_), .Y(ori_ori_n157_));
  NO3        o135(.A(i_3_), .B(ori_ori_n81_), .C(ori_ori_n47_), .Y(ori_ori_n158_));
  NA2        o136(.A(ori_ori_n158_), .B(ori_ori_n766_), .Y(ori_ori_n159_));
  NO3        o137(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n160_));
  NO3        o138(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n161_));
  NA2        o139(.A(i_12_), .B(ori_ori_n161_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n162_), .B(ori_ori_n159_), .Y(ori_ori_n163_));
  NO2        o141(.A(i_3_), .B(i_8_), .Y(ori_ori_n164_));
  NO3        o142(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n165_));
  NA3        o143(.A(ori_ori_n165_), .B(ori_ori_n164_), .C(ori_ori_n39_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n99_), .B(ori_ori_n55_), .Y(ori_ori_n167_));
  NO2        o145(.A(i_13_), .B(i_9_), .Y(ori_ori_n168_));
  NAi21      o146(.An(i_12_), .B(i_3_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n43_), .B(i_5_), .Y(ori_ori_n170_));
  INV        o148(.A(ori_ori_n163_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n171_), .B(i_4_), .Y(ori_ori_n172_));
  NAi21      o150(.An(i_12_), .B(i_7_), .Y(ori_ori_n173_));
  NA3        o151(.A(i_13_), .B(ori_ori_n157_), .C(i_10_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n174_), .B(ori_ori_n173_), .Y(ori_ori_n175_));
  NA2        o153(.A(i_0_), .B(i_5_), .Y(ori_ori_n176_));
  OAI220     o154(.A0(ori_ori_n81_), .A1(ori_ori_n155_), .B0(i_2_), .B1(ori_ori_n124_), .Y(ori_ori_n177_));
  NAi31      o155(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n45_), .B(ori_ori_n58_), .Y(ori_ori_n180_));
  NA3        o158(.A(ori_ori_n180_), .B(i_3_), .C(ori_ori_n179_), .Y(ori_ori_n181_));
  INV        o159(.A(i_13_), .Y(ori_ori_n182_));
  NO2        o160(.A(i_12_), .B(ori_ori_n182_), .Y(ori_ori_n183_));
  NA3        o161(.A(ori_ori_n183_), .B(ori_ori_n160_), .C(ori_ori_n158_), .Y(ori_ori_n184_));
  OAI210     o162(.A0(ori_ori_n181_), .A1(ori_ori_n178_), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  AOI220     o163(.A0(ori_ori_n185_), .A1(i_7_), .B0(ori_ori_n177_), .B1(ori_ori_n175_), .Y(ori_ori_n186_));
  NO2        o164(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n187_));
  OR2        o165(.A(i_8_), .B(i_7_), .Y(ori_ori_n188_));
  INV        o166(.A(i_12_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n43_), .B(ori_ori_n189_), .Y(ori_ori_n190_));
  NO3        o168(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n191_));
  NA2        o169(.A(i_2_), .B(i_1_), .Y(ori_ori_n192_));
  NO3        o170(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n193_));
  NAi21      o171(.An(i_4_), .B(i_3_), .Y(ori_ori_n194_));
  NO2        o172(.A(i_0_), .B(i_6_), .Y(ori_ori_n195_));
  NOi41      o173(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n196_));
  NO2        o174(.A(i_11_), .B(ori_ori_n182_), .Y(ori_ori_n197_));
  NOi21      o175(.An(i_1_), .B(i_6_), .Y(ori_ori_n198_));
  NAi21      o176(.An(i_3_), .B(i_7_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n189_), .B(i_9_), .Y(ori_ori_n200_));
  OR4        o178(.A(ori_ori_n200_), .B(ori_ori_n199_), .C(ori_ori_n198_), .D(ori_ori_n151_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n68_), .B(i_5_), .Y(ori_ori_n202_));
  NA2        o180(.A(i_3_), .B(i_9_), .Y(ori_ori_n203_));
  NAi21      o181(.An(i_7_), .B(i_10_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(ori_ori_n203_), .Y(ori_ori_n205_));
  NA3        o183(.A(ori_ori_n205_), .B(ori_ori_n202_), .C(ori_ori_n59_), .Y(ori_ori_n206_));
  NA2        o184(.A(ori_ori_n206_), .B(ori_ori_n201_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n189_), .B(i_13_), .Y(ori_ori_n208_));
  NA2        o186(.A(ori_ori_n207_), .B(ori_ori_n197_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n188_), .B(ori_ori_n37_), .Y(ori_ori_n210_));
  NA2        o188(.A(i_12_), .B(i_6_), .Y(ori_ori_n211_));
  OR2        o189(.A(i_13_), .B(i_9_), .Y(ori_ori_n212_));
  NO3        o190(.A(ori_ori_n212_), .B(ori_ori_n211_), .C(ori_ori_n47_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n194_), .B(i_2_), .Y(ori_ori_n214_));
  NA3        o192(.A(ori_ori_n214_), .B(ori_ori_n213_), .C(ori_ori_n43_), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n197_), .B(i_9_), .Y(ori_ori_n216_));
  NA2        o194(.A(ori_ori_n202_), .B(ori_ori_n59_), .Y(ori_ori_n217_));
  OAI210     o195(.A0(ori_ori_n217_), .A1(ori_ori_n216_), .B0(ori_ori_n215_), .Y(ori_ori_n218_));
  NO3        o196(.A(i_11_), .B(ori_ori_n182_), .C(ori_ori_n25_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n218_), .B(ori_ori_n210_), .Y(ori_ori_n220_));
  NA3        o198(.A(ori_ori_n220_), .B(ori_ori_n209_), .C(ori_ori_n186_), .Y(ori_ori_n221_));
  NO3        o199(.A(i_12_), .B(ori_ori_n182_), .C(ori_ori_n37_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n192_), .B(i_0_), .Y(ori_ori_n223_));
  NO2        o201(.A(i_3_), .B(i_10_), .Y(ori_ori_n224_));
  NO2        o202(.A(i_2_), .B(ori_ori_n97_), .Y(ori_ori_n225_));
  AN2        o203(.A(i_3_), .B(i_10_), .Y(ori_ori_n226_));
  NO2        o204(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n45_), .B(ori_ori_n26_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n221_), .B(ori_ori_n172_), .Y(ori_ori_n229_));
  NO3        o207(.A(ori_ori_n43_), .B(i_13_), .C(i_9_), .Y(ori_ori_n230_));
  NO2        o208(.A(i_2_), .B(i_3_), .Y(ori_ori_n231_));
  OR2        o209(.A(i_0_), .B(i_5_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n176_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n140_), .B(ori_ori_n45_), .Y(ori_ori_n234_));
  NO2        o212(.A(i_12_), .B(i_10_), .Y(ori_ori_n235_));
  NOi21      o213(.An(i_5_), .B(i_0_), .Y(ori_ori_n236_));
  NO2        o214(.A(i_2_), .B(ori_ori_n97_), .Y(ori_ori_n237_));
  NO4        o215(.A(ori_ori_n237_), .B(i_4_), .C(ori_ori_n236_), .D(ori_ori_n119_), .Y(ori_ori_n238_));
  NA4        o216(.A(ori_ori_n79_), .B(ori_ori_n36_), .C(ori_ori_n81_), .D(i_8_), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n238_), .B(ori_ori_n235_), .Y(ori_ori_n240_));
  NO2        o218(.A(i_6_), .B(i_8_), .Y(ori_ori_n241_));
  NO2        o219(.A(i_1_), .B(i_7_), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n240_), .Y(ori_ori_n243_));
  NA3        o221(.A(ori_ori_n198_), .B(ori_ori_n225_), .C(ori_ori_n157_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n157_), .B(i_9_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n245_), .B(ori_ori_n167_), .Y(ori_ori_n246_));
  NO2        o224(.A(ori_ori_n244_), .B(ori_ori_n143_), .Y(ori_ori_n247_));
  AOI210     o225(.A0(ori_ori_n243_), .A1(ori_ori_n230_), .B0(ori_ori_n247_), .Y(ori_ori_n248_));
  NOi32      o226(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n249_));
  INV        o227(.A(ori_ori_n249_), .Y(ori_ori_n250_));
  NAi21      o228(.An(i_1_), .B(i_5_), .Y(ori_ori_n251_));
  NAi41      o229(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n252_));
  OAI220     o230(.A0(ori_ori_n252_), .A1(ori_ori_n251_), .B0(ori_ori_n178_), .B1(ori_ori_n141_), .Y(ori_ori_n253_));
  AOI210     o231(.A0(ori_ori_n252_), .A1(ori_ori_n141_), .B0(ori_ori_n140_), .Y(ori_ori_n254_));
  NOi32      o232(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n255_));
  NAi21      o233(.An(i_6_), .B(i_1_), .Y(ori_ori_n256_));
  NA3        o234(.A(ori_ori_n256_), .B(ori_ori_n255_), .C(ori_ori_n45_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n257_), .B(i_0_), .Y(ori_ori_n258_));
  OR3        o236(.A(ori_ori_n258_), .B(ori_ori_n254_), .C(ori_ori_n253_), .Y(ori_ori_n259_));
  NO2        o237(.A(i_1_), .B(ori_ori_n97_), .Y(ori_ori_n260_));
  NAi21      o238(.An(i_3_), .B(i_4_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n261_), .B(i_9_), .Y(ori_ori_n262_));
  AN2        o240(.A(i_6_), .B(i_7_), .Y(ori_ori_n263_));
  OAI210     o241(.A0(ori_ori_n263_), .A1(ori_ori_n260_), .B0(ori_ori_n262_), .Y(ori_ori_n264_));
  NA2        o242(.A(i_2_), .B(i_7_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n261_), .B(i_10_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n264_), .B(ori_ori_n151_), .Y(ori_ori_n267_));
  AOI210     o245(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n268_));
  OAI210     o246(.A0(ori_ori_n268_), .A1(ori_ori_n154_), .B0(ori_ori_n266_), .Y(ori_ori_n269_));
  AOI220     o247(.A0(ori_ori_n266_), .A1(ori_ori_n242_), .B0(ori_ori_n191_), .B1(ori_ori_n154_), .Y(ori_ori_n270_));
  AOI210     o248(.A0(ori_ori_n270_), .A1(ori_ori_n269_), .B0(i_5_), .Y(ori_ori_n271_));
  NO3        o249(.A(ori_ori_n271_), .B(ori_ori_n267_), .C(ori_ori_n259_), .Y(ori_ori_n272_));
  NO2        o250(.A(ori_ori_n272_), .B(ori_ori_n250_), .Y(ori_ori_n273_));
  NO2        o251(.A(ori_ori_n56_), .B(ori_ori_n25_), .Y(ori_ori_n274_));
  AN2        o252(.A(i_12_), .B(i_5_), .Y(ori_ori_n275_));
  NO2        o253(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n276_), .B(ori_ori_n275_), .Y(ori_ori_n277_));
  NO2        o255(.A(i_11_), .B(i_6_), .Y(ori_ori_n278_));
  NA3        o256(.A(ori_ori_n278_), .B(ori_ori_n234_), .C(ori_ori_n182_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n279_), .B(ori_ori_n277_), .Y(ori_ori_n280_));
  NO2        o258(.A(i_5_), .B(i_10_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n281_), .B(ori_ori_n214_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n132_), .B(ori_ori_n44_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n283_), .B(ori_ori_n282_), .Y(ori_ori_n284_));
  OAI210     o262(.A0(ori_ori_n284_), .A1(ori_ori_n280_), .B0(ori_ori_n274_), .Y(ori_ori_n285_));
  NO2        o263(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n286_));
  NO2        o264(.A(ori_ori_n138_), .B(ori_ori_n81_), .Y(ori_ori_n287_));
  OAI210     o265(.A0(ori_ori_n287_), .A1(ori_ori_n280_), .B0(ori_ori_n286_), .Y(ori_ori_n288_));
  NA3        o266(.A(ori_ori_n224_), .B(ori_ori_n88_), .C(ori_ori_n70_), .Y(ori_ori_n289_));
  NO2        o267(.A(i_11_), .B(i_12_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n290_), .B(ori_ori_n36_), .Y(ori_ori_n291_));
  NO2        o269(.A(ori_ori_n289_), .B(ori_ori_n291_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n281_), .B(ori_ori_n189_), .Y(ori_ori_n293_));
  NAi21      o271(.An(i_13_), .B(i_0_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n294_), .B(ori_ori_n192_), .Y(ori_ori_n295_));
  NA2        o273(.A(ori_ori_n292_), .B(ori_ori_n295_), .Y(ori_ori_n296_));
  NA3        o274(.A(ori_ori_n296_), .B(ori_ori_n288_), .C(ori_ori_n285_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n43_), .B(ori_ori_n182_), .Y(ori_ori_n298_));
  NO2        o276(.A(i_0_), .B(i_11_), .Y(ori_ori_n299_));
  NOi21      o277(.An(i_2_), .B(i_12_), .Y(ori_ori_n300_));
  NAi21      o278(.An(i_9_), .B(i_4_), .Y(ori_ori_n301_));
  OR2        o279(.A(i_13_), .B(i_10_), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n146_), .B(ori_ori_n114_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n97_), .B(ori_ori_n25_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n157_), .B(i_10_), .Y(ori_ori_n305_));
  NA3        o283(.A(ori_ori_n202_), .B(ori_ori_n59_), .C(i_2_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n306_), .B(ori_ori_n305_), .Y(ori_ori_n307_));
  NA2        o285(.A(i_8_), .B(ori_ori_n233_), .Y(ori_ori_n308_));
  NO2        o286(.A(ori_ori_n308_), .B(ori_ori_n155_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n309_), .B(ori_ori_n307_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n310_), .B(ori_ori_n216_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n311_), .B(ori_ori_n297_), .C(ori_ori_n273_), .Y(ori_ori_n312_));
  NO2        o290(.A(i_10_), .B(i_9_), .Y(ori_ori_n313_));
  NAi21      o291(.An(i_12_), .B(i_8_), .Y(ori_ori_n314_));
  NO2        o292(.A(ori_ori_n314_), .B(i_3_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n45_), .B(i_4_), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n316_), .B(ori_ori_n100_), .Y(ori_ori_n317_));
  NO2        o295(.A(ori_ori_n317_), .B(ori_ori_n166_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n228_), .B(i_0_), .Y(ori_ori_n319_));
  NO3        o297(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n320_));
  NA2        o298(.A(ori_ori_n211_), .B(ori_ori_n95_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n321_), .B(ori_ori_n320_), .Y(ori_ori_n322_));
  NA2        o300(.A(i_8_), .B(i_9_), .Y(ori_ori_n323_));
  NO2        o301(.A(i_7_), .B(i_2_), .Y(ori_ori_n324_));
  OR2        o302(.A(ori_ori_n324_), .B(ori_ori_n323_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n222_), .B(ori_ori_n167_), .Y(ori_ori_n326_));
  OAI220     o304(.A0(ori_ori_n326_), .A1(ori_ori_n325_), .B0(ori_ori_n322_), .B1(ori_ori_n319_), .Y(ori_ori_n327_));
  NO3        o305(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n328_));
  NO2        o306(.A(ori_ori_n327_), .B(ori_ori_n318_), .Y(ori_ori_n329_));
  BUFFER     o307(.A(ori_ori_n246_), .Y(ori_ori_n330_));
  OR2        o308(.A(ori_ori_n330_), .B(ori_ori_n143_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n94_), .B(i_13_), .Y(ori_ori_n332_));
  NA2        o310(.A(i_5_), .B(ori_ori_n274_), .Y(ori_ori_n333_));
  NO2        o311(.A(i_2_), .B(i_13_), .Y(ori_ori_n334_));
  NO2        o312(.A(ori_ori_n333_), .B(ori_ori_n332_), .Y(ori_ori_n335_));
  NO3        o313(.A(i_4_), .B(ori_ori_n47_), .C(i_8_), .Y(ori_ori_n336_));
  NO2        o314(.A(i_6_), .B(i_7_), .Y(ori_ori_n337_));
  NO2        o315(.A(i_11_), .B(i_1_), .Y(ori_ori_n338_));
  NO2        o316(.A(i_3_), .B(ori_ori_n157_), .Y(ori_ori_n339_));
  NO2        o317(.A(i_6_), .B(i_10_), .Y(ori_ori_n340_));
  NA3        o318(.A(ori_ori_n196_), .B(ori_ori_n145_), .C(ori_ori_n123_), .Y(ori_ori_n341_));
  NA3        o319(.A(ori_ori_n286_), .B(ori_ori_n150_), .C(ori_ori_n137_), .Y(ori_ori_n342_));
  NA2        o320(.A(ori_ori_n342_), .B(ori_ori_n341_), .Y(ori_ori_n343_));
  NO2        o321(.A(ori_ori_n343_), .B(ori_ori_n335_), .Y(ori_ori_n344_));
  NA2        o322(.A(ori_ori_n320_), .B(ori_ori_n275_), .Y(ori_ori_n345_));
  NA2        o323(.A(ori_ori_n328_), .B(ori_ori_n281_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n346_), .B(ori_ori_n181_), .Y(ori_ori_n347_));
  NAi21      o325(.An(ori_ori_n174_), .B(ori_ori_n290_), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n242_), .B(ori_ori_n176_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n349_), .B(ori_ori_n348_), .Y(ori_ori_n350_));
  NA2        o328(.A(ori_ori_n230_), .B(ori_ori_n191_), .Y(ori_ori_n351_));
  NO2        o329(.A(ori_ori_n351_), .B(ori_ori_n306_), .Y(ori_ori_n352_));
  NO3        o330(.A(ori_ori_n352_), .B(ori_ori_n350_), .C(ori_ori_n347_), .Y(ori_ori_n353_));
  NA4        o331(.A(ori_ori_n353_), .B(ori_ori_n344_), .C(ori_ori_n331_), .D(ori_ori_n329_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n113_), .B(ori_ori_n108_), .Y(ori_ori_n355_));
  AN2        o333(.A(ori_ori_n355_), .B(ori_ori_n320_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(ori_ori_n228_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n275_), .B(ori_ori_n182_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n249_), .B(ori_ori_n68_), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n263_), .B(ori_ori_n255_), .Y(ori_ori_n360_));
  OR2        o338(.A(ori_ori_n358_), .B(ori_ori_n360_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n362_));
  INV        o340(.A(ori_ori_n361_), .Y(ori_ori_n363_));
  NA2        o341(.A(ori_ori_n202_), .B(ori_ori_n59_), .Y(ori_ori_n364_));
  OAI210     o342(.A0(i_8_), .A1(ori_ori_n364_), .B0(ori_ori_n125_), .Y(ori_ori_n365_));
  NA2        o343(.A(ori_ori_n365_), .B(ori_ori_n303_), .Y(ori_ori_n366_));
  NA3        o344(.A(ori_ori_n366_), .B(ori_ori_n361_), .C(ori_ori_n357_), .Y(ori_ori_n367_));
  NO2        o345(.A(i_12_), .B(ori_ori_n157_), .Y(ori_ori_n368_));
  NO2        o346(.A(i_8_), .B(i_7_), .Y(ori_ori_n369_));
  NA2        o347(.A(ori_ori_n43_), .B(i_10_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n370_), .B(i_6_), .Y(ori_ori_n371_));
  AOI220     o349(.A0(i_5_), .A1(ori_ori_n234_), .B0(i_2_), .B1(ori_ori_n195_), .Y(ori_ori_n372_));
  OAI220     o350(.A0(ori_ori_n372_), .A1(ori_ori_n208_), .B0(ori_ori_n332_), .B1(ori_ori_n124_), .Y(ori_ori_n373_));
  NA2        o351(.A(ori_ori_n373_), .B(ori_ori_n210_), .Y(ori_ori_n374_));
  NA3        o352(.A(ori_ori_n226_), .B(ori_ori_n147_), .C(ori_ori_n94_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n140_), .B(i_5_), .Y(ori_ori_n376_));
  NA3        o354(.A(ori_ori_n376_), .B(ori_ori_n298_), .C(ori_ori_n231_), .Y(ori_ori_n377_));
  NA2        o355(.A(ori_ori_n377_), .B(ori_ori_n375_), .Y(ori_ori_n378_));
  NA2        o356(.A(ori_ori_n378_), .B(ori_ori_n328_), .Y(ori_ori_n379_));
  NA2        o357(.A(ori_ori_n379_), .B(ori_ori_n374_), .Y(ori_ori_n380_));
  AOI210     o358(.A0(ori_ori_n256_), .A1(ori_ori_n45_), .B0(ori_ori_n260_), .Y(ori_ori_n381_));
  NA2        o359(.A(i_0_), .B(ori_ori_n47_), .Y(ori_ori_n382_));
  NA3        o360(.A(ori_ori_n368_), .B(ori_ori_n219_), .C(ori_ori_n382_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n381_), .B(ori_ori_n383_), .Y(ori_ori_n384_));
  INV        o362(.A(ori_ori_n384_), .Y(ori_ori_n385_));
  NO4        o363(.A(ori_ori_n198_), .B(ori_ori_n41_), .C(i_2_), .D(ori_ori_n47_), .Y(ori_ori_n386_));
  NO3        o364(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n387_));
  NOi21      o365(.An(i_10_), .B(i_6_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n81_), .B(ori_ori_n25_), .Y(ori_ori_n389_));
  AOI220     o367(.A0(ori_ori_n222_), .A1(ori_ori_n389_), .B0(ori_ori_n219_), .B1(ori_ori_n388_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n390_), .B(ori_ori_n319_), .Y(ori_ori_n391_));
  NO2        o369(.A(ori_ori_n109_), .B(ori_ori_n23_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n160_), .B(ori_ori_n37_), .Y(ori_ori_n393_));
  NOi31      o371(.An(ori_ori_n134_), .B(ori_ori_n393_), .C(ori_ori_n239_), .Y(ori_ori_n394_));
  NO2        o372(.A(ori_ori_n394_), .B(ori_ori_n391_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n359_), .B(ori_ori_n270_), .Y(ori_ori_n396_));
  INV        o374(.A(ori_ori_n231_), .Y(ori_ori_n397_));
  NO2        o375(.A(i_12_), .B(ori_ori_n81_), .Y(ori_ori_n398_));
  NA3        o376(.A(ori_ori_n398_), .B(ori_ori_n219_), .C(ori_ori_n382_), .Y(ori_ori_n399_));
  NA3        o377(.A(ori_ori_n278_), .B(ori_ori_n222_), .C(ori_ori_n176_), .Y(ori_ori_n400_));
  AOI210     o378(.A0(ori_ori_n400_), .A1(ori_ori_n399_), .B0(ori_ori_n397_), .Y(ori_ori_n401_));
  OR2        o379(.A(i_2_), .B(i_5_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n265_), .B(ori_ori_n195_), .Y(ori_ori_n403_));
  NO2        o381(.A(ori_ori_n403_), .B(ori_ori_n348_), .Y(ori_ori_n404_));
  NO3        o382(.A(ori_ori_n404_), .B(ori_ori_n401_), .C(ori_ori_n396_), .Y(ori_ori_n405_));
  NA3        o383(.A(ori_ori_n405_), .B(ori_ori_n395_), .C(ori_ori_n385_), .Y(ori_ori_n406_));
  NO4        o384(.A(ori_ori_n406_), .B(ori_ori_n380_), .C(ori_ori_n367_), .D(ori_ori_n354_), .Y(ori_ori_n407_));
  NA4        o385(.A(ori_ori_n407_), .B(ori_ori_n312_), .C(ori_ori_n248_), .D(ori_ori_n229_), .Y(ori7));
  NO2        o386(.A(ori_ori_n104_), .B(ori_ori_n87_), .Y(ori_ori_n409_));
  NA2        o387(.A(ori_ori_n276_), .B(ori_ori_n409_), .Y(ori_ori_n410_));
  NA2        o388(.A(ori_ori_n340_), .B(ori_ori_n79_), .Y(ori_ori_n411_));
  NA2        o389(.A(i_11_), .B(ori_ori_n157_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n132_), .B(ori_ori_n412_), .Y(ori_ori_n413_));
  OAI210     o391(.A0(ori_ori_n413_), .A1(ori_ori_n411_), .B0(ori_ori_n410_), .Y(ori_ori_n414_));
  NO2        o392(.A(ori_ori_n189_), .B(i_4_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(i_8_), .Y(ori_ori_n416_));
  NA2        o394(.A(i_2_), .B(ori_ori_n81_), .Y(ori_ori_n417_));
  OAI210     o395(.A0(ori_ori_n84_), .A1(ori_ori_n164_), .B0(ori_ori_n165_), .Y(ori_ori_n418_));
  NO2        o396(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n419_));
  NO2        o397(.A(ori_ori_n418_), .B(i_13_), .Y(ori_ori_n420_));
  NO2        o398(.A(ori_ori_n420_), .B(ori_ori_n414_), .Y(ori_ori_n421_));
  AOI210     o399(.A0(ori_ori_n119_), .A1(ori_ori_n57_), .B0(i_10_), .Y(ori_ori_n422_));
  AOI210     o400(.A0(ori_ori_n422_), .A1(ori_ori_n189_), .B0(ori_ori_n142_), .Y(ori_ori_n423_));
  OR2        o401(.A(i_6_), .B(i_10_), .Y(ori_ori_n424_));
  INV        o402(.A(ori_ori_n161_), .Y(ori_ori_n425_));
  OR2        o403(.A(ori_ori_n423_), .B(ori_ori_n212_), .Y(ori_ori_n426_));
  AOI210     o404(.A0(ori_ori_n426_), .A1(ori_ori_n421_), .B0(ori_ori_n58_), .Y(ori_ori_n427_));
  NOi21      o405(.An(i_11_), .B(i_7_), .Y(ori_ori_n428_));
  AO210      o406(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n429_));
  NO2        o407(.A(ori_ori_n429_), .B(ori_ori_n428_), .Y(ori_ori_n430_));
  NA2        o408(.A(ori_ori_n430_), .B(ori_ori_n168_), .Y(ori_ori_n431_));
  NA3        o409(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n432_));
  NAi21      o410(.An(ori_ori_n432_), .B(i_11_), .Y(ori_ori_n433_));
  AOI210     o411(.A0(ori_ori_n433_), .A1(ori_ori_n431_), .B0(ori_ori_n58_), .Y(ori_ori_n434_));
  NA2        o412(.A(ori_ori_n83_), .B(ori_ori_n58_), .Y(ori_ori_n435_));
  AO210      o413(.A0(ori_ori_n435_), .A1(ori_ori_n270_), .B0(ori_ori_n40_), .Y(ori_ori_n436_));
  NO3        o414(.A(ori_ori_n204_), .B(ori_ori_n169_), .C(ori_ori_n412_), .Y(ori_ori_n437_));
  OAI210     o415(.A0(ori_ori_n437_), .A1(ori_ori_n183_), .B0(ori_ori_n58_), .Y(ori_ori_n438_));
  NO2        o416(.A(ori_ori_n58_), .B(i_9_), .Y(ori_ori_n439_));
  NO2        o417(.A(i_1_), .B(i_12_), .Y(ori_ori_n440_));
  NA3        o418(.A(ori_ori_n440_), .B(ori_ori_n106_), .C(ori_ori_n24_), .Y(ori_ori_n441_));
  BUFFER     o419(.A(ori_ori_n441_), .Y(ori_ori_n442_));
  NA3        o420(.A(ori_ori_n442_), .B(ori_ori_n438_), .C(ori_ori_n436_), .Y(ori_ori_n443_));
  OAI210     o421(.A0(ori_ori_n443_), .A1(ori_ori_n434_), .B0(i_6_), .Y(ori_ori_n444_));
  NO2        o422(.A(ori_ori_n432_), .B(ori_ori_n104_), .Y(ori_ori_n445_));
  NA2        o423(.A(ori_ori_n445_), .B(ori_ori_n398_), .Y(ori_ori_n446_));
  NO2        o424(.A(i_6_), .B(i_11_), .Y(ori_ori_n447_));
  NA2        o425(.A(ori_ori_n446_), .B(ori_ori_n322_), .Y(ori_ori_n448_));
  NO3        o426(.A(ori_ori_n424_), .B(ori_ori_n188_), .C(ori_ori_n23_), .Y(ori_ori_n449_));
  AOI210     o427(.A0(i_1_), .A1(ori_ori_n205_), .B0(ori_ori_n449_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n450_), .B(ori_ori_n43_), .Y(ori_ori_n451_));
  NA3        o429(.A(ori_ori_n369_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n452_));
  INV        o430(.A(i_2_), .Y(ori_ori_n453_));
  NA2        o431(.A(ori_ori_n129_), .B(i_9_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n45_), .B(i_1_), .Y(ori_ori_n455_));
  NO2        o433(.A(ori_ori_n454_), .B(ori_ori_n453_), .Y(ori_ori_n456_));
  NA3        o434(.A(ori_ori_n439_), .B(ori_ori_n231_), .C(i_6_), .Y(ori_ori_n457_));
  NO2        o435(.A(ori_ori_n457_), .B(ori_ori_n23_), .Y(ori_ori_n458_));
  AOI210     o436(.A0(ori_ori_n338_), .A1(ori_ori_n304_), .B0(ori_ori_n193_), .Y(ori_ori_n459_));
  NO2        o437(.A(ori_ori_n459_), .B(ori_ori_n417_), .Y(ori_ori_n460_));
  NAi21      o438(.An(ori_ori_n452_), .B(ori_ori_n89_), .Y(ori_ori_n461_));
  NA2        o439(.A(ori_ori_n455_), .B(ori_ori_n211_), .Y(ori_ori_n462_));
  NO2        o440(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n463_), .B(ori_ori_n24_), .Y(ori_ori_n464_));
  OAI210     o442(.A0(ori_ori_n464_), .A1(ori_ori_n462_), .B0(ori_ori_n461_), .Y(ori_ori_n465_));
  OR4        o443(.A(ori_ori_n465_), .B(ori_ori_n460_), .C(ori_ori_n458_), .D(ori_ori_n456_), .Y(ori_ori_n466_));
  NO3        o444(.A(ori_ori_n466_), .B(ori_ori_n451_), .C(ori_ori_n448_), .Y(ori_ori_n467_));
  NO2        o445(.A(i_12_), .B(ori_ori_n428_), .Y(ori_ori_n468_));
  NO2        o446(.A(ori_ori_n301_), .B(ori_ori_n81_), .Y(ori_ori_n469_));
  NA2        o447(.A(i_3_), .B(ori_ori_n157_), .Y(ori_ori_n470_));
  NO2        o448(.A(ori_ori_n470_), .B(ori_ori_n109_), .Y(ori_ori_n471_));
  AN2        o449(.A(ori_ori_n471_), .B(ori_ori_n371_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n188_), .B(ori_ori_n43_), .Y(ori_ori_n473_));
  NO3        o451(.A(ori_ori_n473_), .B(ori_ori_n228_), .C(ori_ori_n190_), .Y(ori_ori_n474_));
  NO2        o452(.A(ori_ori_n110_), .B(ori_ori_n37_), .Y(ori_ori_n475_));
  NO2        o453(.A(ori_ori_n475_), .B(i_6_), .Y(ori_ori_n476_));
  NO2        o454(.A(ori_ori_n81_), .B(i_9_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n477_), .B(ori_ori_n58_), .Y(ori_ori_n478_));
  NO2        o456(.A(ori_ori_n478_), .B(ori_ori_n440_), .Y(ori_ori_n479_));
  NO4        o457(.A(ori_ori_n479_), .B(ori_ori_n476_), .C(ori_ori_n474_), .D(i_4_), .Y(ori_ori_n480_));
  NA2        o458(.A(i_1_), .B(i_3_), .Y(ori_ori_n481_));
  NO2        o459(.A(ori_ori_n323_), .B(ori_ori_n90_), .Y(ori_ori_n482_));
  AOI210     o460(.A0(ori_ori_n473_), .A1(ori_ori_n388_), .B0(ori_ori_n482_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n483_), .B(ori_ori_n481_), .Y(ori_ori_n484_));
  NO3        o462(.A(ori_ori_n484_), .B(ori_ori_n480_), .C(ori_ori_n472_), .Y(ori_ori_n485_));
  NA3        o463(.A(ori_ori_n485_), .B(ori_ori_n467_), .C(ori_ori_n444_), .Y(ori_ori_n486_));
  NA2        o464(.A(ori_ori_n263_), .B(ori_ori_n262_), .Y(ori_ori_n487_));
  NA3        o465(.A(ori_ori_n340_), .B(ori_ori_n362_), .C(ori_ori_n45_), .Y(ori_ori_n488_));
  NA3        o466(.A(ori_ori_n142_), .B(ori_ori_n79_), .C(ori_ori_n81_), .Y(ori_ori_n489_));
  NA3        o467(.A(ori_ori_n489_), .B(ori_ori_n488_), .C(ori_ori_n487_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n490_), .B(i_1_), .Y(ori_ori_n491_));
  AOI210     o469(.A0(ori_ori_n211_), .A1(ori_ori_n95_), .B0(i_1_), .Y(ori_ori_n492_));
  NO2        o470(.A(ori_ori_n261_), .B(i_2_), .Y(ori_ori_n493_));
  NA2        o471(.A(ori_ori_n493_), .B(ori_ori_n492_), .Y(ori_ori_n494_));
  OAI210     o472(.A0(ori_ori_n457_), .A1(ori_ori_n314_), .B0(ori_ori_n494_), .Y(ori_ori_n495_));
  INV        o473(.A(ori_ori_n495_), .Y(ori_ori_n496_));
  AOI210     o474(.A0(ori_ori_n496_), .A1(ori_ori_n491_), .B0(i_13_), .Y(ori_ori_n497_));
  OR2        o475(.A(i_11_), .B(i_7_), .Y(ori_ori_n498_));
  NA3        o476(.A(ori_ori_n498_), .B(ori_ori_n102_), .C(ori_ori_n129_), .Y(ori_ori_n499_));
  AOI220     o477(.A0(ori_ori_n334_), .A1(ori_ori_n142_), .B0(ori_ori_n316_), .B1(ori_ori_n129_), .Y(ori_ori_n500_));
  OAI210     o478(.A0(ori_ori_n500_), .A1(ori_ori_n43_), .B0(ori_ori_n499_), .Y(ori_ori_n501_));
  NO2        o479(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n502_));
  INV        o480(.A(ori_ori_n502_), .Y(ori_ori_n503_));
  NA2        o481(.A(i_7_), .B(ori_ori_n469_), .Y(ori_ori_n504_));
  OAI220     o482(.A0(ori_ori_n504_), .A1(ori_ori_n40_), .B0(ori_ori_n503_), .B1(ori_ori_n90_), .Y(ori_ori_n505_));
  AOI210     o483(.A0(ori_ori_n501_), .A1(ori_ori_n241_), .B0(ori_ori_n505_), .Y(ori_ori_n506_));
  INV        o484(.A(ori_ori_n109_), .Y(ori_ori_n507_));
  AOI220     o485(.A0(ori_ori_n507_), .A1(ori_ori_n67_), .B0(ori_ori_n278_), .B1(ori_ori_n455_), .Y(ori_ori_n508_));
  NO2        o486(.A(ori_ori_n508_), .B(ori_ori_n194_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n118_), .B(i_13_), .Y(ori_ori_n510_));
  NO2        o488(.A(ori_ori_n510_), .B(ori_ori_n492_), .Y(ori_ori_n511_));
  NO3        o489(.A(ori_ori_n66_), .B(ori_ori_n32_), .C(ori_ori_n97_), .Y(ori_ori_n512_));
  AOI220     o490(.A0(ori_ori_n278_), .A1(ori_ori_n455_), .B0(ori_ori_n89_), .B1(ori_ori_n98_), .Y(ori_ori_n513_));
  OAI220     o491(.A0(ori_ori_n513_), .A1(ori_ori_n416_), .B0(ori_ori_n765_), .B1(ori_ori_n425_), .Y(ori_ori_n514_));
  NO3        o492(.A(ori_ori_n514_), .B(ori_ori_n511_), .C(ori_ori_n509_), .Y(ori_ori_n515_));
  NA3        o493(.A(ori_ori_n300_), .B(ori_ori_n419_), .C(ori_ori_n95_), .Y(ori_ori_n516_));
  NA2        o494(.A(ori_ori_n447_), .B(i_13_), .Y(ori_ori_n517_));
  NAi21      o495(.An(i_11_), .B(i_12_), .Y(ori_ori_n518_));
  NOi41      o496(.An(ori_ori_n107_), .B(ori_ori_n518_), .C(i_13_), .D(ori_ori_n81_), .Y(ori_ori_n519_));
  INV        o497(.A(ori_ori_n519_), .Y(ori_ori_n520_));
  NA3        o498(.A(ori_ori_n520_), .B(ori_ori_n517_), .C(ori_ori_n516_), .Y(ori_ori_n521_));
  NA2        o499(.A(ori_ori_n521_), .B(ori_ori_n58_), .Y(ori_ori_n522_));
  NO2        o500(.A(i_2_), .B(i_12_), .Y(ori_ori_n523_));
  NA2        o501(.A(ori_ori_n260_), .B(ori_ori_n523_), .Y(ori_ori_n524_));
  NA2        o502(.A(i_8_), .B(ori_ori_n25_), .Y(ori_ori_n525_));
  NO2        o503(.A(ori_ori_n525_), .B(ori_ori_n276_), .Y(ori_ori_n526_));
  OAI210     o504(.A0(ori_ori_n526_), .A1(ori_ori_n262_), .B0(ori_ori_n260_), .Y(ori_ori_n527_));
  NA2        o505(.A(ori_ori_n527_), .B(ori_ori_n524_), .Y(ori_ori_n528_));
  NA3        o506(.A(ori_ori_n528_), .B(ori_ori_n44_), .C(ori_ori_n182_), .Y(ori_ori_n529_));
  NA4        o507(.A(ori_ori_n529_), .B(ori_ori_n522_), .C(ori_ori_n515_), .D(ori_ori_n506_), .Y(ori_ori_n530_));
  OR4        o508(.A(ori_ori_n530_), .B(ori_ori_n497_), .C(ori_ori_n486_), .D(ori_ori_n427_), .Y(ori5));
  NA2        o509(.A(ori_ori_n468_), .B(ori_ori_n214_), .Y(ori_ori_n532_));
  AN2        o510(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n533_));
  NA3        o511(.A(ori_ori_n533_), .B(ori_ori_n523_), .C(ori_ori_n104_), .Y(ori_ori_n534_));
  NO2        o512(.A(ori_ori_n416_), .B(i_11_), .Y(ori_ori_n535_));
  NA2        o513(.A(ori_ori_n84_), .B(ori_ori_n535_), .Y(ori_ori_n536_));
  NA3        o514(.A(ori_ori_n536_), .B(ori_ori_n534_), .C(ori_ori_n532_), .Y(ori_ori_n537_));
  NO3        o515(.A(i_11_), .B(ori_ori_n189_), .C(i_13_), .Y(ori_ori_n538_));
  NO2        o516(.A(ori_ori_n115_), .B(ori_ori_n23_), .Y(ori_ori_n539_));
  NA2        o517(.A(i_12_), .B(i_8_), .Y(ori_ori_n540_));
  INV        o518(.A(ori_ori_n313_), .Y(ori_ori_n541_));
  AOI220     o519(.A0(ori_ori_n231_), .A1(ori_ori_n392_), .B0(i_12_), .B1(ori_ori_n539_), .Y(ori_ori_n542_));
  INV        o520(.A(ori_ori_n542_), .Y(ori_ori_n543_));
  NO2        o521(.A(ori_ori_n543_), .B(ori_ori_n537_), .Y(ori_ori_n544_));
  INV        o522(.A(ori_ori_n145_), .Y(ori_ori_n545_));
  INV        o523(.A(ori_ori_n196_), .Y(ori_ori_n546_));
  OAI210     o524(.A0(ori_ori_n493_), .A1(ori_ori_n315_), .B0(ori_ori_n107_), .Y(ori_ori_n547_));
  AOI210     o525(.A0(ori_ori_n547_), .A1(ori_ori_n546_), .B0(ori_ori_n545_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n323_), .B(ori_ori_n26_), .Y(ori_ori_n549_));
  NO2        o527(.A(ori_ori_n549_), .B(ori_ori_n304_), .Y(ori_ori_n550_));
  NA2        o528(.A(ori_ori_n550_), .B(i_2_), .Y(ori_ori_n551_));
  INV        o529(.A(ori_ori_n551_), .Y(ori_ori_n552_));
  AOI210     o530(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n302_), .Y(ori_ori_n553_));
  AOI210     o531(.A0(ori_ori_n553_), .A1(ori_ori_n552_), .B0(ori_ori_n548_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n156_), .B(ori_ori_n116_), .Y(ori_ori_n555_));
  OAI210     o533(.A0(ori_ori_n555_), .A1(ori_ori_n539_), .B0(i_2_), .Y(ori_ori_n556_));
  INV        o534(.A(ori_ori_n146_), .Y(ori_ori_n557_));
  NA2        o535(.A(ori_ori_n557_), .B(ori_ori_n84_), .Y(ori_ori_n558_));
  AOI210     o536(.A0(ori_ori_n558_), .A1(ori_ori_n556_), .B0(ori_ori_n157_), .Y(ori_ori_n559_));
  OA210      o537(.A0(ori_ori_n430_), .A1(ori_ori_n117_), .B0(i_13_), .Y(ori_ori_n560_));
  NA2        o538(.A(ori_ori_n161_), .B(ori_ori_n164_), .Y(ori_ori_n561_));
  NO2        o539(.A(ori_ori_n561_), .B(ori_ori_n265_), .Y(ori_ori_n562_));
  AOI210     o540(.A0(ori_ori_n169_), .A1(ori_ori_n136_), .B0(ori_ori_n362_), .Y(ori_ori_n563_));
  NA2        o541(.A(ori_ori_n563_), .B(ori_ori_n304_), .Y(ori_ori_n564_));
  NO2        o542(.A(ori_ori_n98_), .B(ori_ori_n43_), .Y(ori_ori_n565_));
  INV        o543(.A(ori_ori_n225_), .Y(ori_ori_n566_));
  NA4        o544(.A(ori_ori_n566_), .B(ori_ori_n226_), .C(ori_ori_n115_), .D(ori_ori_n41_), .Y(ori_ori_n567_));
  OAI210     o545(.A0(ori_ori_n567_), .A1(ori_ori_n565_), .B0(ori_ori_n564_), .Y(ori_ori_n568_));
  NO4        o546(.A(ori_ori_n568_), .B(ori_ori_n562_), .C(ori_ori_n560_), .D(ori_ori_n559_), .Y(ori_ori_n569_));
  NO2        o547(.A(ori_ori_n57_), .B(i_12_), .Y(ori_ori_n570_));
  NO2        o548(.A(ori_ori_n570_), .B(ori_ori_n117_), .Y(ori_ori_n571_));
  NO2        o549(.A(ori_ori_n571_), .B(ori_ori_n412_), .Y(ori_ori_n572_));
  NA2        o550(.A(ori_ori_n572_), .B(ori_ori_n36_), .Y(ori_ori_n573_));
  NA4        o551(.A(ori_ori_n573_), .B(ori_ori_n569_), .C(ori_ori_n554_), .D(ori_ori_n544_), .Y(ori6));
  NA4        o552(.A(ori_ori_n281_), .B(ori_ori_n339_), .C(ori_ori_n66_), .D(ori_ori_n97_), .Y(ori_ori_n575_));
  INV        o553(.A(ori_ori_n575_), .Y(ori_ori_n576_));
  NO2        o554(.A(i_11_), .B(i_9_), .Y(ori_ori_n577_));
  NO2        o555(.A(ori_ori_n576_), .B(ori_ori_n236_), .Y(ori_ori_n578_));
  OR2        o556(.A(ori_ori_n578_), .B(i_12_), .Y(ori_ori_n579_));
  NA2        o557(.A(ori_ori_n266_), .B(ori_ori_n242_), .Y(ori_ori_n580_));
  NA2        o558(.A(ori_ori_n398_), .B(ori_ori_n58_), .Y(ori_ori_n581_));
  BUFFER     o559(.A(ori_ori_n435_), .Y(ori_ori_n582_));
  NA3        o560(.A(ori_ori_n582_), .B(ori_ori_n581_), .C(ori_ori_n580_), .Y(ori_ori_n583_));
  INV        o561(.A(ori_ori_n159_), .Y(ori_ori_n584_));
  AOI220     o562(.A0(ori_ori_n584_), .A1(ori_ori_n577_), .B0(ori_ori_n583_), .B1(ori_ori_n68_), .Y(ori_ori_n585_));
  INV        o563(.A(ori_ori_n235_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n70_), .B(ori_ori_n122_), .Y(ori_ori_n587_));
  INV        o565(.A(ori_ori_n115_), .Y(ori_ori_n588_));
  NA2        o566(.A(ori_ori_n588_), .B(ori_ori_n45_), .Y(ori_ori_n589_));
  AOI210     o567(.A0(ori_ori_n589_), .A1(ori_ori_n587_), .B0(ori_ori_n586_), .Y(ori_ori_n590_));
  NO2        o568(.A(ori_ori_n198_), .B(i_9_), .Y(ori_ori_n591_));
  NA2        o569(.A(ori_ori_n591_), .B(ori_ori_n570_), .Y(ori_ori_n592_));
  AOI210     o570(.A0(ori_ori_n592_), .A1(ori_ori_n360_), .B0(ori_ori_n151_), .Y(ori_ori_n593_));
  NO2        o571(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n594_));
  NA3        o572(.A(ori_ori_n594_), .B(ori_ori_n337_), .C(ori_ori_n281_), .Y(ori_ori_n595_));
  INV        o573(.A(ori_ori_n595_), .Y(ori_ori_n596_));
  OR3        o574(.A(ori_ori_n596_), .B(ori_ori_n593_), .C(ori_ori_n590_), .Y(ori_ori_n597_));
  OR2        o575(.A(ori_ori_n430_), .B(ori_ori_n315_), .Y(ori_ori_n598_));
  NA3        o576(.A(ori_ori_n598_), .B(ori_ori_n135_), .C(ori_ori_n64_), .Y(ori_ori_n599_));
  AO210      o577(.A0(ori_ori_n346_), .A1(ori_ori_n541_), .B0(ori_ori_n36_), .Y(ori_ori_n600_));
  NA2        o578(.A(ori_ori_n600_), .B(ori_ori_n599_), .Y(ori_ori_n601_));
  OAI210     o579(.A0(i_6_), .A1(i_11_), .B0(ori_ori_n82_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n602_), .B(ori_ori_n387_), .Y(ori_ori_n603_));
  NA3        o581(.A(ori_ori_n265_), .B(ori_ori_n191_), .C(ori_ori_n135_), .Y(ori_ori_n604_));
  NA3        o582(.A(ori_ori_n604_), .B(ori_ori_n603_), .C(ori_ori_n418_), .Y(ori_ori_n605_));
  AO210      o583(.A0(ori_ori_n362_), .A1(ori_ori_n45_), .B0(ori_ori_n83_), .Y(ori_ori_n606_));
  NA3        o584(.A(ori_ori_n606_), .B(ori_ori_n340_), .C(ori_ori_n176_), .Y(ori_ori_n607_));
  AOI210     o585(.A0(ori_ori_n315_), .A1(ori_ori_n313_), .B0(ori_ori_n386_), .Y(ori_ori_n608_));
  NO2        o586(.A(ori_ori_n424_), .B(ori_ori_n98_), .Y(ori_ori_n609_));
  OAI210     o587(.A0(ori_ori_n609_), .A1(ori_ori_n108_), .B0(ori_ori_n299_), .Y(ori_ori_n610_));
  NA3        o588(.A(ori_ori_n610_), .B(ori_ori_n608_), .C(ori_ori_n607_), .Y(ori_ori_n611_));
  NO4        o589(.A(ori_ori_n611_), .B(ori_ori_n605_), .C(ori_ori_n601_), .D(ori_ori_n597_), .Y(ori_ori_n612_));
  NA4        o590(.A(ori_ori_n612_), .B(ori_ori_n585_), .C(ori_ori_n579_), .D(ori_ori_n272_), .Y(ori3));
  NA2        o591(.A(i_12_), .B(i_10_), .Y(ori_ori_n614_));
  NO2        o592(.A(i_11_), .B(ori_ori_n189_), .Y(ori_ori_n615_));
  NA3        o593(.A(ori_ori_n604_), .B(ori_ori_n418_), .C(ori_ori_n264_), .Y(ori_ori_n616_));
  NA2        o594(.A(ori_ori_n616_), .B(ori_ori_n39_), .Y(ori_ori_n617_));
  NOi21      o595(.An(ori_ori_n94_), .B(ori_ori_n550_), .Y(ori_ori_n618_));
  NA2        o596(.A(ori_ori_n300_), .B(ori_ori_n44_), .Y(ori_ori_n619_));
  AN2        o597(.A(ori_ori_n321_), .B(ori_ori_n53_), .Y(ori_ori_n620_));
  NO2        o598(.A(ori_ori_n620_), .B(ori_ori_n618_), .Y(ori_ori_n621_));
  AOI210     o599(.A0(ori_ori_n621_), .A1(ori_ori_n617_), .B0(ori_ori_n47_), .Y(ori_ori_n622_));
  NO4        o600(.A(ori_ori_n268_), .B(ori_ori_n275_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n623_));
  NA2        o601(.A(ori_ori_n151_), .B(ori_ori_n388_), .Y(ori_ori_n624_));
  NOi21      o602(.An(ori_ori_n624_), .B(ori_ori_n623_), .Y(ori_ori_n625_));
  NO2        o603(.A(ori_ori_n625_), .B(ori_ori_n58_), .Y(ori_ori_n626_));
  NO2        o604(.A(ori_ori_n626_), .B(ori_ori_n622_), .Y(ori_ori_n627_));
  NA2        o605(.A(ori_ori_n151_), .B(ori_ori_n24_), .Y(ori_ori_n628_));
  NO2        o606(.A(ori_ori_n475_), .B(ori_ori_n409_), .Y(ori_ori_n629_));
  NO2        o607(.A(ori_ori_n629_), .B(ori_ori_n628_), .Y(ori_ori_n630_));
  NA2        o608(.A(ori_ori_n230_), .B(ori_ori_n120_), .Y(ori_ori_n631_));
  NO2        o609(.A(ori_ori_n631_), .B(ori_ori_n293_), .Y(ori_ori_n632_));
  NO2        o610(.A(ori_ori_n632_), .B(ori_ori_n630_), .Y(ori_ori_n633_));
  NA2        o611(.A(ori_ori_n389_), .B(i_0_), .Y(ori_ori_n634_));
  NO3        o612(.A(ori_ori_n634_), .B(ori_ori_n277_), .C(ori_ori_n84_), .Y(ori_ori_n635_));
  NO3        o613(.A(ori_ori_n402_), .B(ori_ori_n173_), .C(ori_ori_n302_), .Y(ori_ori_n636_));
  AOI210     o614(.A0(ori_ori_n636_), .A1(i_11_), .B0(ori_ori_n635_), .Y(ori_ori_n637_));
  NA2        o615(.A(ori_ori_n538_), .B(ori_ori_n236_), .Y(ori_ori_n638_));
  AOI210     o616(.A0(ori_ori_n340_), .A1(ori_ori_n84_), .B0(ori_ori_n55_), .Y(ori_ori_n639_));
  NO2        o617(.A(ori_ori_n639_), .B(ori_ori_n638_), .Y(ori_ori_n640_));
  NO2        o618(.A(ori_ori_n200_), .B(ori_ori_n139_), .Y(ori_ori_n641_));
  NA2        o619(.A(i_0_), .B(i_10_), .Y(ori_ori_n642_));
  INV        o620(.A(ori_ori_n370_), .Y(ori_ori_n643_));
  NO3        o621(.A(ori_ori_n109_), .B(ori_ori_n470_), .C(i_5_), .Y(ori_ori_n644_));
  AO220      o622(.A0(ori_ori_n644_), .A1(ori_ori_n643_), .B0(ori_ori_n641_), .B1(i_6_), .Y(ori_ori_n645_));
  NO2        o623(.A(ori_ori_n645_), .B(ori_ori_n640_), .Y(ori_ori_n646_));
  NA3        o624(.A(ori_ori_n646_), .B(ori_ori_n637_), .C(ori_ori_n633_), .Y(ori_ori_n647_));
  NO2        o625(.A(ori_ori_n99_), .B(ori_ori_n37_), .Y(ori_ori_n648_));
  NA2        o626(.A(i_11_), .B(i_9_), .Y(ori_ori_n649_));
  NO3        o627(.A(i_12_), .B(ori_ori_n649_), .C(ori_ori_n417_), .Y(ori_ori_n650_));
  AN2        o628(.A(ori_ori_n650_), .B(ori_ori_n648_), .Y(ori_ori_n651_));
  NA2        o629(.A(ori_ori_n286_), .B(ori_ori_n150_), .Y(ori_ori_n652_));
  INV        o630(.A(ori_ori_n652_), .Y(ori_ori_n653_));
  NO2        o631(.A(ori_ori_n649_), .B(ori_ori_n68_), .Y(ori_ori_n654_));
  NO2        o632(.A(ori_ori_n148_), .B(i_0_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n653_), .B(ori_ori_n651_), .Y(ori_ori_n656_));
  NA2        o634(.A(ori_ori_n463_), .B(ori_ori_n112_), .Y(ori_ori_n657_));
  NO2        o635(.A(i_6_), .B(ori_ori_n657_), .Y(ori_ori_n658_));
  NA2        o636(.A(ori_ori_n145_), .B(ori_ori_n99_), .Y(ori_ori_n659_));
  NO2        o637(.A(ori_ori_n767_), .B(ori_ori_n619_), .Y(ori_ori_n660_));
  NO2        o638(.A(ori_ori_n660_), .B(ori_ori_n658_), .Y(ori_ori_n661_));
  NOi21      o639(.An(i_7_), .B(i_5_), .Y(ori_ori_n662_));
  NOi31      o640(.An(ori_ori_n662_), .B(i_0_), .C(ori_ori_n518_), .Y(ori_ori_n663_));
  NA3        o641(.A(ori_ori_n663_), .B(ori_ori_n276_), .C(i_6_), .Y(ori_ori_n664_));
  BUFFER     o642(.A(ori_ori_n664_), .Y(ori_ori_n665_));
  INV        o643(.A(ori_ori_n232_), .Y(ori_ori_n666_));
  NA3        o644(.A(ori_ori_n665_), .B(ori_ori_n661_), .C(ori_ori_n656_), .Y(ori_ori_n667_));
  NO2        o645(.A(ori_ori_n614_), .B(ori_ori_n231_), .Y(ori_ori_n668_));
  OA210      o646(.A0(ori_ori_n337_), .A1(ori_ori_n180_), .B0(ori_ori_n336_), .Y(ori_ori_n669_));
  NA2        o647(.A(ori_ori_n668_), .B(ori_ori_n654_), .Y(ori_ori_n670_));
  NA2        o648(.A(ori_ori_n654_), .B(ori_ori_n226_), .Y(ori_ori_n671_));
  OAI210     o649(.A0(i_3_), .A1(ori_ori_n153_), .B0(ori_ori_n671_), .Y(ori_ori_n672_));
  NA2        o650(.A(ori_ori_n672_), .B(ori_ori_n337_), .Y(ori_ori_n673_));
  NA3        o651(.A(i_5_), .B(ori_ori_n274_), .C(i_6_), .Y(ori_ori_n674_));
  NA2        o652(.A(ori_ori_n90_), .B(ori_ori_n43_), .Y(ori_ori_n675_));
  NO2        o653(.A(ori_ori_n70_), .B(ori_ori_n540_), .Y(ori_ori_n676_));
  AOI220     o654(.A0(ori_ori_n676_), .A1(ori_ori_n675_), .B0(ori_ori_n147_), .B1(ori_ori_n409_), .Y(ori_ori_n677_));
  AOI210     o655(.A0(ori_ori_n677_), .A1(ori_ori_n674_), .B0(ori_ori_n46_), .Y(ori_ori_n678_));
  NO3        o656(.A(ori_ori_n402_), .B(i_0_), .C(ori_ori_n24_), .Y(ori_ori_n679_));
  AOI210     o657(.A0(i_7_), .A1(ori_ori_n376_), .B0(ori_ori_n679_), .Y(ori_ori_n680_));
  NAi21      o658(.An(i_9_), .B(i_5_), .Y(ori_ori_n681_));
  NO2        o659(.A(ori_ori_n681_), .B(ori_ori_n294_), .Y(ori_ori_n682_));
  NA2        o660(.A(ori_ori_n682_), .B(ori_ori_n430_), .Y(ori_ori_n683_));
  OAI220     o661(.A0(ori_ori_n683_), .A1(ori_ori_n81_), .B0(ori_ori_n680_), .B1(ori_ori_n146_), .Y(ori_ori_n684_));
  NO3        o662(.A(ori_ori_n684_), .B(ori_ori_n678_), .C(ori_ori_n363_), .Y(ori_ori_n685_));
  NA3        o663(.A(ori_ori_n685_), .B(ori_ori_n673_), .C(ori_ori_n670_), .Y(ori_ori_n686_));
  NO3        o664(.A(ori_ori_n686_), .B(ori_ori_n667_), .C(ori_ori_n647_), .Y(ori_ori_n687_));
  NO2        o665(.A(i_0_), .B(ori_ori_n518_), .Y(ori_ori_n688_));
  AOI210     o666(.A0(ori_ori_n581_), .A1(ori_ori_n487_), .B0(ori_ori_n659_), .Y(ori_ori_n689_));
  INV        o667(.A(ori_ori_n689_), .Y(ori_ori_n690_));
  NA2        o668(.A(ori_ori_n195_), .B(ori_ori_n187_), .Y(ori_ori_n691_));
  AOI210     o669(.A0(ori_ori_n691_), .A1(ori_ori_n634_), .B0(ori_ori_n139_), .Y(ori_ori_n692_));
  INV        o670(.A(ori_ori_n692_), .Y(ori_ori_n693_));
  NA2        o671(.A(ori_ori_n693_), .B(ori_ori_n690_), .Y(ori_ori_n694_));
  NO3        o672(.A(ori_ori_n642_), .B(i_5_), .C(ori_ori_n156_), .Y(ori_ori_n695_));
  NA2        o673(.A(ori_ori_n695_), .B(i_11_), .Y(ori_ori_n696_));
  NO3        o674(.A(ori_ori_n170_), .B(ori_ori_n275_), .C(i_0_), .Y(ori_ori_n697_));
  OAI210     o675(.A0(ori_ori_n697_), .A1(ori_ori_n71_), .B0(i_13_), .Y(ori_ori_n698_));
  NA2        o676(.A(ori_ori_n698_), .B(ori_ori_n696_), .Y(ori_ori_n699_));
  NO2        o677(.A(ori_ori_n194_), .B(ori_ori_n90_), .Y(ori_ori_n700_));
  AOI210     o678(.A0(ori_ori_n700_), .A1(ori_ori_n688_), .B0(ori_ori_n105_), .Y(ori_ori_n701_));
  OR2        o679(.A(ori_ori_n701_), .B(i_5_), .Y(ori_ori_n702_));
  AOI210     o680(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n148_), .Y(ori_ori_n703_));
  NA2        o681(.A(ori_ori_n703_), .B(ori_ori_n669_), .Y(ori_ori_n704_));
  NA2        o682(.A(ori_ori_n345_), .B(ori_ori_n341_), .Y(ori_ori_n705_));
  INV        o683(.A(ori_ori_n705_), .Y(ori_ori_n706_));
  NA3        o684(.A(ori_ori_n281_), .B(ori_ori_n145_), .C(ori_ori_n144_), .Y(ori_ori_n707_));
  NA3        o685(.A(i_5_), .B(ori_ori_n223_), .C(ori_ori_n187_), .Y(ori_ori_n708_));
  NA2        o686(.A(ori_ori_n708_), .B(ori_ori_n707_), .Y(ori_ori_n709_));
  NO3        o687(.A(ori_ori_n649_), .B(ori_ori_n176_), .C(ori_ori_n156_), .Y(ori_ori_n710_));
  NO2        o688(.A(ori_ori_n710_), .B(ori_ori_n709_), .Y(ori_ori_n711_));
  NA4        o689(.A(ori_ori_n711_), .B(ori_ori_n706_), .C(ori_ori_n704_), .D(ori_ori_n702_), .Y(ori_ori_n712_));
  NO2        o690(.A(ori_ori_n81_), .B(i_5_), .Y(ori_ori_n713_));
  NA3        o691(.A(ori_ori_n615_), .B(ori_ori_n106_), .C(ori_ori_n115_), .Y(ori_ori_n714_));
  INV        o692(.A(ori_ori_n714_), .Y(ori_ori_n715_));
  NA2        o693(.A(ori_ori_n715_), .B(ori_ori_n713_), .Y(ori_ori_n716_));
  NA2        o694(.A(ori_ori_n226_), .B(i_5_), .Y(ori_ori_n717_));
  NAi31      o695(.An(ori_ori_n193_), .B(ori_ori_n717_), .C(ori_ori_n194_), .Y(ori_ori_n718_));
  NO4        o696(.A(ori_ori_n192_), .B(ori_ori_n170_), .C(i_0_), .D(i_12_), .Y(ori_ori_n719_));
  AOI220     o697(.A0(ori_ori_n719_), .A1(ori_ori_n718_), .B0(ori_ori_n576_), .B1(ori_ori_n149_), .Y(ori_ori_n720_));
  AN2        o698(.A(ori_ori_n642_), .B(ori_ori_n139_), .Y(ori_ori_n721_));
  NO3        o699(.A(ori_ori_n721_), .B(i_12_), .C(ori_ori_n452_), .Y(ori_ori_n722_));
  NA2        o700(.A(ori_ori_n722_), .B(ori_ori_n176_), .Y(ori_ori_n723_));
  NA2        o701(.A(ori_ori_n662_), .B(ori_ori_n334_), .Y(ori_ori_n724_));
  NA2        o702(.A(ori_ori_n59_), .B(ori_ori_n97_), .Y(ori_ori_n725_));
  OAI220     o703(.A0(ori_ori_n725_), .A1(ori_ori_n717_), .B0(ori_ori_n724_), .B1(ori_ori_n478_), .Y(ori_ori_n726_));
  NA2        o704(.A(ori_ori_n726_), .B(ori_ori_n655_), .Y(ori_ori_n727_));
  NA4        o705(.A(ori_ori_n727_), .B(ori_ori_n723_), .C(ori_ori_n720_), .D(ori_ori_n716_), .Y(ori_ori_n728_));
  NO4        o706(.A(ori_ori_n728_), .B(ori_ori_n712_), .C(ori_ori_n699_), .D(ori_ori_n694_), .Y(ori_ori_n729_));
  NA2        o707(.A(ori_ori_n594_), .B(ori_ori_n37_), .Y(ori_ori_n730_));
  NA2        o708(.A(ori_ori_n730_), .B(ori_ori_n423_), .Y(ori_ori_n731_));
  NA2        o709(.A(ori_ori_n731_), .B(ori_ori_n168_), .Y(ori_ori_n732_));
  BUFFER     o710(.A(ori_ori_n498_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n152_), .B(ori_ori_n154_), .Y(ori_ori_n734_));
  AO210      o712(.A0(ori_ori_n733_), .A1(ori_ori_n33_), .B0(ori_ori_n734_), .Y(ori_ori_n735_));
  NAi31      o713(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n736_));
  NO2        o714(.A(ori_ori_n65_), .B(ori_ori_n736_), .Y(ori_ori_n737_));
  NO2        o715(.A(ori_ori_n737_), .B(ori_ori_n449_), .Y(ori_ori_n738_));
  NA2        o716(.A(ori_ori_n738_), .B(ori_ori_n735_), .Y(ori_ori_n739_));
  AOI210     o717(.A0(ori_ori_n739_), .A1(ori_ori_n47_), .B0(ori_ori_n636_), .Y(ori_ori_n740_));
  AOI210     o718(.A0(ori_ori_n740_), .A1(ori_ori_n732_), .B0(ori_ori_n68_), .Y(ori_ori_n741_));
  INV        o719(.A(ori_ori_n271_), .Y(ori_ori_n742_));
  NO2        o720(.A(ori_ori_n742_), .B(ori_ori_n545_), .Y(ori_ori_n743_));
  INV        o721(.A(ori_ori_n71_), .Y(ori_ori_n744_));
  AOI210     o722(.A0(ori_ori_n703_), .A1(i_5_), .B0(ori_ori_n663_), .Y(ori_ori_n745_));
  AOI210     o723(.A0(ori_ori_n745_), .A1(ori_ori_n744_), .B0(ori_ori_n481_), .Y(ori_ori_n746_));
  INV        o724(.A(ori_ori_n746_), .Y(ori_ori_n747_));
  NA2        o725(.A(ori_ori_n213_), .B(ori_ori_n84_), .Y(ori_ori_n748_));
  NA3        o726(.A(ori_ori_n549_), .B(ori_ori_n223_), .C(ori_ori_n75_), .Y(ori_ori_n749_));
  AOI210     o727(.A0(ori_ori_n749_), .A1(ori_ori_n748_), .B0(i_11_), .Y(ori_ori_n750_));
  NO3        o728(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(i_4_), .Y(ori_ori_n751_));
  OAI210     o729(.A0(ori_ori_n666_), .A1(ori_ori_n227_), .B0(ori_ori_n751_), .Y(ori_ori_n752_));
  NO2        o730(.A(ori_ori_n752_), .B(ori_ori_n518_), .Y(ori_ori_n753_));
  NO4        o731(.A(ori_ori_n681_), .B(i_11_), .C(ori_ori_n199_), .D(ori_ori_n198_), .Y(ori_ori_n754_));
  NO2        o732(.A(ori_ori_n754_), .B(ori_ori_n386_), .Y(ori_ori_n755_));
  INV        o733(.A(ori_ori_n253_), .Y(ori_ori_n756_));
  AOI210     o734(.A0(ori_ori_n756_), .A1(ori_ori_n755_), .B0(ori_ori_n40_), .Y(ori_ori_n757_));
  NO3        o735(.A(ori_ori_n757_), .B(ori_ori_n753_), .C(ori_ori_n750_), .Y(ori_ori_n758_));
  OAI210     o736(.A0(ori_ori_n747_), .A1(i_4_), .B0(ori_ori_n758_), .Y(ori_ori_n759_));
  NO3        o737(.A(ori_ori_n759_), .B(ori_ori_n743_), .C(ori_ori_n741_), .Y(ori_ori_n760_));
  NA4        o738(.A(ori_ori_n760_), .B(ori_ori_n729_), .C(ori_ori_n687_), .D(ori_ori_n627_), .Y(ori4));
  INV        o739(.A(i_6_), .Y(ori_ori_n764_));
  INV        o740(.A(ori_ori_n512_), .Y(ori_ori_n765_));
  INV        o741(.A(i_8_), .Y(ori_ori_n766_));
  INV        o742(.A(ori_ori_n236_), .Y(ori_ori_n767_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m021(.A(mai_mai_n35_), .Y(mai1));
  INV        m022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m024(.A(i_2_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_0_), .B(i_2_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_7_), .B(i_9_), .Y(mai_mai_n52_));
  NA3        m030(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n53_));
  NO2        m031(.A(i_1_), .B(i_6_), .Y(mai_mai_n54_));
  NA2        m032(.A(i_8_), .B(i_7_), .Y(mai_mai_n55_));
  OAI210     m033(.A0(mai_mai_n55_), .A1(mai_mai_n54_), .B0(mai_mai_n53_), .Y(mai_mai_n56_));
  NA2        m034(.A(mai_mai_n56_), .B(i_12_), .Y(mai_mai_n57_));
  NAi21      m035(.An(i_2_), .B(i_7_), .Y(mai_mai_n58_));
  INV        m036(.A(i_1_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(i_6_), .Y(mai_mai_n60_));
  NA3        m038(.A(mai_mai_n60_), .B(mai_mai_n58_), .C(mai_mai_n31_), .Y(mai_mai_n61_));
  NA2        m039(.A(i_1_), .B(i_10_), .Y(mai_mai_n62_));
  NO2        m040(.A(mai_mai_n62_), .B(i_6_), .Y(mai_mai_n63_));
  NAi31      m041(.An(mai_mai_n63_), .B(mai_mai_n61_), .C(mai_mai_n57_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n65_));
  AOI210     m043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_1_), .B(i_6_), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n67_), .B(mai_mai_n25_), .Y(mai_mai_n68_));
  INV        m046(.A(i_0_), .Y(mai_mai_n69_));
  NAi21      m047(.An(i_5_), .B(i_10_), .Y(mai_mai_n70_));
  NA2        m048(.A(i_5_), .B(i_9_), .Y(mai_mai_n71_));
  AOI210     m049(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n69_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n72_), .B(mai_mai_n68_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n66_), .A1(mai_mai_n65_), .B0(mai_mai_n73_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n74_), .A1(mai_mai_n64_), .B0(i_0_), .Y(mai_mai_n75_));
  NA2        m053(.A(i_12_), .B(i_5_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_2_), .B(i_8_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n54_), .Y(mai_mai_n78_));
  NO2        m056(.A(i_3_), .B(i_9_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_3_), .B(i_7_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n80_), .B(mai_mai_n79_), .C(mai_mai_n59_), .Y(mai_mai_n81_));
  INV        m059(.A(i_6_), .Y(mai_mai_n82_));
  OR4        m060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n83_));
  INV        m061(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  NO2        m062(.A(i_2_), .B(i_7_), .Y(mai_mai_n85_));
  OAI210     m063(.A0(mai_mai_n81_), .A1(mai_mai_n78_), .B0(i_2_), .Y(mai_mai_n86_));
  NAi21      m064(.An(i_6_), .B(i_10_), .Y(mai_mai_n87_));
  NA2        m065(.A(i_6_), .B(i_9_), .Y(mai_mai_n88_));
  AOI210     m066(.A0(mai_mai_n88_), .A1(mai_mai_n87_), .B0(mai_mai_n59_), .Y(mai_mai_n89_));
  NA2        m067(.A(i_2_), .B(i_6_), .Y(mai_mai_n90_));
  INV        m068(.A(mai_mai_n89_), .Y(mai_mai_n91_));
  AOI210     m069(.A0(mai_mai_n91_), .A1(mai_mai_n86_), .B0(mai_mai_n76_), .Y(mai_mai_n92_));
  AN3        m070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n93_));
  NAi21      m071(.An(i_6_), .B(i_11_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_5_), .B(i_8_), .Y(mai_mai_n95_));
  NOi21      m073(.An(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  AOI220     m074(.A0(mai_mai_n96_), .A1(mai_mai_n58_), .B0(mai_mai_n93_), .B1(mai_mai_n32_), .Y(mai_mai_n97_));
  INV        m075(.A(i_7_), .Y(mai_mai_n98_));
  NA2        m076(.A(mai_mai_n47_), .B(mai_mai_n98_), .Y(mai_mai_n99_));
  NO2        m077(.A(i_0_), .B(i_5_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n82_), .Y(mai_mai_n101_));
  NA2        m079(.A(i_12_), .B(i_3_), .Y(mai_mai_n102_));
  INV        m080(.A(mai_mai_n102_), .Y(mai_mai_n103_));
  NA3        m081(.A(mai_mai_n103_), .B(mai_mai_n101_), .C(mai_mai_n99_), .Y(mai_mai_n104_));
  NAi21      m082(.An(i_7_), .B(i_11_), .Y(mai_mai_n105_));
  AN2        m083(.A(i_2_), .B(i_10_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(i_7_), .Y(mai_mai_n107_));
  OR2        m085(.A(mai_mai_n76_), .B(mai_mai_n54_), .Y(mai_mai_n108_));
  NO2        m086(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n109_));
  NO3        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n110_));
  NA2        m088(.A(i_12_), .B(i_7_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n59_), .B(mai_mai_n26_), .Y(mai_mai_n112_));
  NA2        m090(.A(mai_mai_n112_), .B(i_0_), .Y(mai_mai_n113_));
  NA2        m091(.A(i_11_), .B(i_12_), .Y(mai_mai_n114_));
  OAI210     m092(.A0(mai_mai_n113_), .A1(mai_mai_n111_), .B0(mai_mai_n114_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n110_), .Y(mai_mai_n116_));
  NA3        m094(.A(mai_mai_n116_), .B(mai_mai_n104_), .C(mai_mai_n97_), .Y(mai_mai_n117_));
  NOi21      m095(.An(i_1_), .B(i_5_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n118_), .B(i_11_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n98_), .B(mai_mai_n37_), .Y(mai_mai_n120_));
  NA2        m098(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(mai_mai_n120_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n122_), .B(mai_mai_n47_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n124_));
  INV        m102(.A(mai_mai_n124_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_1_), .B(mai_mai_n82_), .Y(mai_mai_n126_));
  NO2        m104(.A(i_6_), .B(i_5_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(i_3_), .Y(mai_mai_n128_));
  OAI220     m106(.A0(mai_mai_n128_), .A1(mai_mai_n105_), .B0(mai_mai_n125_), .B1(mai_mai_n119_), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n117_), .C(mai_mai_n92_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n75_), .Y(mai2));
  NO2        m109(.A(mai_mai_n59_), .B(mai_mai_n37_), .Y(mai_mai_n132_));
  NA2        m110(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NA4        m112(.A(mai_mai_n134_), .B(mai_mai_n73_), .C(mai_mai_n65_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m113(.A(i_8_), .B(i_7_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n136_), .B(i_6_), .Y(mai_mai_n137_));
  NO2        m115(.A(i_12_), .B(i_13_), .Y(mai_mai_n138_));
  NAi21      m116(.An(i_5_), .B(i_11_), .Y(mai_mai_n139_));
  NOi21      m117(.An(mai_mai_n138_), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m118(.A(i_0_), .B(i_1_), .Y(mai_mai_n141_));
  NA2        m119(.A(i_2_), .B(i_3_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n142_), .B(i_4_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(mai_mai_n140_), .Y(mai_mai_n144_));
  AN2        m122(.A(mai_mai_n138_), .B(mai_mai_n79_), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n145_), .B(mai_mai_n27_), .Y(mai_mai_n146_));
  NA2        m124(.A(i_1_), .B(i_5_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n69_), .B(mai_mai_n47_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n150_));
  OR2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n76_), .C(i_13_), .Y(mai_mai_n152_));
  NAi32      m130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n153_));
  NAi21      m131(.An(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m132(.An(i_4_), .B(i_10_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NO2        m134(.A(i_3_), .B(i_5_), .Y(mai_mai_n157_));
  NO3        m135(.A(mai_mai_n69_), .B(i_2_), .C(i_1_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n154_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(mai_mai_n150_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(mai_mai_n161_), .A1(mai_mai_n144_), .B0(mai_mai_n137_), .Y(mai_mai_n162_));
  NA3        m140(.A(mai_mai_n69_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n163_));
  NOi21      m141(.An(i_4_), .B(i_9_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_11_), .B(i_13_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  NO2        m144(.A(i_4_), .B(i_5_), .Y(mai_mai_n167_));
  NAi21      m145(.An(i_12_), .B(i_11_), .Y(mai_mai_n168_));
  NO2        m146(.A(mai_mai_n168_), .B(i_13_), .Y(mai_mai_n169_));
  NA3        m147(.A(mai_mai_n169_), .B(mai_mai_n167_), .C(mai_mai_n79_), .Y(mai_mai_n170_));
  AOI210     m148(.A0(mai_mai_n170_), .A1(mai_mai_n166_), .B0(mai_mai_n163_), .Y(mai_mai_n171_));
  NO2        m149(.A(mai_mai_n69_), .B(mai_mai_n59_), .Y(mai_mai_n172_));
  INV        m150(.A(mai_mai_n172_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n174_));
  NAi31      m152(.An(mai_mai_n174_), .B(mai_mai_n145_), .C(i_11_), .Y(mai_mai_n175_));
  NA2        m153(.A(i_3_), .B(i_5_), .Y(mai_mai_n176_));
  OR2        m154(.A(mai_mai_n176_), .B(mai_mai_n166_), .Y(mai_mai_n177_));
  AOI210     m155(.A0(mai_mai_n177_), .A1(mai_mai_n175_), .B0(mai_mai_n173_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n69_), .B(i_5_), .Y(mai_mai_n179_));
  NO2        m157(.A(i_13_), .B(i_10_), .Y(mai_mai_n180_));
  NA3        m158(.A(mai_mai_n180_), .B(mai_mai_n179_), .C(mai_mai_n45_), .Y(mai_mai_n181_));
  NO2        m159(.A(i_2_), .B(i_1_), .Y(mai_mai_n182_));
  NAi21      m160(.An(i_4_), .B(i_12_), .Y(mai_mai_n183_));
  NO3        m161(.A(mai_mai_n183_), .B(i_2_), .C(mai_mai_n181_), .Y(mai_mai_n184_));
  NO3        m162(.A(mai_mai_n184_), .B(mai_mai_n178_), .C(mai_mai_n171_), .Y(mai_mai_n185_));
  INV        m163(.A(i_8_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n186_), .B(i_7_), .Y(mai_mai_n187_));
  NA2        m165(.A(mai_mai_n187_), .B(i_6_), .Y(mai_mai_n188_));
  NO3        m166(.A(i_3_), .B(mai_mai_n82_), .C(mai_mai_n48_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n109_), .Y(mai_mai_n190_));
  NO3        m168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n191_));
  NA3        m169(.A(mai_mai_n191_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n192_));
  NO3        m170(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n193_));
  OAI210     m171(.A0(mai_mai_n93_), .A1(i_12_), .B0(mai_mai_n193_), .Y(mai_mai_n194_));
  AOI210     m172(.A0(mai_mai_n194_), .A1(mai_mai_n192_), .B0(mai_mai_n190_), .Y(mai_mai_n195_));
  NO2        m173(.A(i_3_), .B(i_8_), .Y(mai_mai_n196_));
  NO3        m174(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n197_));
  NA3        m175(.A(mai_mai_n197_), .B(mai_mai_n196_), .C(mai_mai_n40_), .Y(mai_mai_n198_));
  NO2        m176(.A(mai_mai_n100_), .B(mai_mai_n54_), .Y(mai_mai_n199_));
  NO2        m177(.A(i_13_), .B(i_9_), .Y(mai_mai_n200_));
  NA3        m178(.A(mai_mai_n200_), .B(i_6_), .C(mai_mai_n186_), .Y(mai_mai_n201_));
  NAi21      m179(.An(i_12_), .B(i_3_), .Y(mai_mai_n202_));
  BUFFER     m180(.A(mai_mai_n201_), .Y(mai_mai_n203_));
  NO2        m181(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n204_));
  NO3        m182(.A(i_0_), .B(i_2_), .C(mai_mai_n59_), .Y(mai_mai_n205_));
  NA3        m183(.A(mai_mai_n205_), .B(mai_mai_n204_), .C(i_10_), .Y(mai_mai_n206_));
  OAI220     m184(.A0(mai_mai_n206_), .A1(mai_mai_n203_), .B0(mai_mai_n100_), .B1(mai_mai_n198_), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n207_), .A1(i_7_), .B0(mai_mai_n195_), .Y(mai_mai_n208_));
  OAI220     m186(.A0(mai_mai_n208_), .A1(i_4_), .B0(mai_mai_n188_), .B1(mai_mai_n185_), .Y(mai_mai_n209_));
  NAi21      m187(.An(i_12_), .B(i_7_), .Y(mai_mai_n210_));
  NA3        m188(.A(i_13_), .B(mai_mai_n186_), .C(i_10_), .Y(mai_mai_n211_));
  NA2        m189(.A(i_0_), .B(i_5_), .Y(mai_mai_n212_));
  NAi31      m190(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n69_), .B(mai_mai_n26_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n47_), .B(mai_mai_n59_), .Y(mai_mai_n216_));
  INV        m194(.A(i_13_), .Y(mai_mai_n217_));
  NO2        m195(.A(i_12_), .B(mai_mai_n217_), .Y(mai_mai_n218_));
  NO2        m196(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n176_), .B(i_4_), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n220_), .B(mai_mai_n219_), .Y(mai_mai_n221_));
  OR2        m199(.A(i_8_), .B(i_7_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n222_), .B(mai_mai_n82_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n51_), .B(i_1_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n225_));
  INV        m203(.A(i_12_), .Y(mai_mai_n226_));
  NO3        m204(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n227_));
  NA2        m205(.A(i_2_), .B(i_1_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n225_), .B(mai_mai_n221_), .Y(mai_mai_n229_));
  NAi21      m207(.An(i_4_), .B(i_3_), .Y(mai_mai_n230_));
  INV        m208(.A(mai_mai_n71_), .Y(mai_mai_n231_));
  NO2        m209(.A(i_0_), .B(i_6_), .Y(mai_mai_n232_));
  NOi41      m210(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n233_), .B(mai_mai_n232_), .Y(mai_mai_n234_));
  NAi21      m212(.An(mai_mai_n234_), .B(i_5_), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n235_), .Y(mai_mai_n236_));
  AOI210     m214(.A0(mai_mai_n236_), .A1(mai_mai_n40_), .B0(mai_mai_n229_), .Y(mai_mai_n237_));
  NO2        m215(.A(i_11_), .B(mai_mai_n217_), .Y(mai_mai_n238_));
  NOi21      m216(.An(i_1_), .B(i_6_), .Y(mai_mai_n239_));
  NAi21      m217(.An(i_3_), .B(i_7_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n226_), .B(i_9_), .Y(mai_mai_n241_));
  OR4        m219(.A(mai_mai_n241_), .B(mai_mai_n240_), .C(mai_mai_n239_), .D(mai_mai_n179_), .Y(mai_mai_n242_));
  NO2        m220(.A(i_12_), .B(i_3_), .Y(mai_mai_n243_));
  NA2        m221(.A(mai_mai_n69_), .B(i_5_), .Y(mai_mai_n244_));
  NA2        m222(.A(i_3_), .B(i_9_), .Y(mai_mai_n245_));
  NAi21      m223(.An(i_7_), .B(i_10_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n246_), .B(mai_mai_n245_), .Y(mai_mai_n247_));
  NA3        m225(.A(mai_mai_n247_), .B(mai_mai_n244_), .C(mai_mai_n60_), .Y(mai_mai_n248_));
  NA2        m226(.A(mai_mai_n248_), .B(mai_mai_n242_), .Y(mai_mai_n249_));
  NA3        m227(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n250_));
  INV        m228(.A(mai_mai_n137_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n226_), .B(i_13_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n252_), .B(mai_mai_n71_), .Y(mai_mai_n253_));
  AOI220     m231(.A0(mai_mai_n253_), .A1(mai_mai_n251_), .B0(mai_mai_n249_), .B1(mai_mai_n238_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n222_), .B(mai_mai_n37_), .Y(mai_mai_n255_));
  NA2        m233(.A(i_12_), .B(i_6_), .Y(mai_mai_n256_));
  OR2        m234(.A(i_13_), .B(i_9_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n230_), .B(i_2_), .Y(mai_mai_n258_));
  NA2        m236(.A(mai_mai_n238_), .B(i_9_), .Y(mai_mai_n259_));
  NA2        m237(.A(mai_mai_n148_), .B(mai_mai_n59_), .Y(mai_mai_n260_));
  NO3        m238(.A(i_11_), .B(mai_mai_n217_), .C(mai_mai_n25_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n240_), .B(i_8_), .Y(mai_mai_n262_));
  NA3        m240(.A(i_5_), .B(mai_mai_n262_), .C(mai_mai_n261_), .Y(mai_mai_n263_));
  NA3        m241(.A(i_6_), .B(mai_mai_n255_), .C(mai_mai_n218_), .Y(mai_mai_n264_));
  AOI210     m242(.A0(mai_mai_n264_), .A1(mai_mai_n263_), .B0(mai_mai_n260_), .Y(mai_mai_n265_));
  INV        m243(.A(mai_mai_n265_), .Y(mai_mai_n266_));
  NA3        m244(.A(mai_mai_n266_), .B(mai_mai_n254_), .C(mai_mai_n237_), .Y(mai_mai_n267_));
  NO3        m245(.A(i_12_), .B(mai_mai_n217_), .C(mai_mai_n37_), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n268_), .Y(mai_mai_n269_));
  NA2        m247(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n270_));
  NOi21      m248(.An(mai_mai_n157_), .B(mai_mai_n82_), .Y(mai_mai_n271_));
  NO3        m249(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n272_));
  AOI220     m250(.A0(mai_mai_n272_), .A1(mai_mai_n189_), .B0(mai_mai_n271_), .B1(mai_mai_n224_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n273_), .B(mai_mai_n270_), .Y(mai_mai_n274_));
  NO3        m252(.A(i_0_), .B(i_2_), .C(mai_mai_n59_), .Y(mai_mai_n275_));
  NO2        m253(.A(mai_mai_n228_), .B(i_0_), .Y(mai_mai_n276_));
  AOI220     m254(.A0(mai_mai_n276_), .A1(mai_mai_n187_), .B0(mai_mai_n275_), .B1(mai_mai_n136_), .Y(mai_mai_n277_));
  NA2        m255(.A(i_5_), .B(mai_mai_n26_), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n278_), .B(mai_mai_n277_), .Y(mai_mai_n279_));
  NA2        m257(.A(i_0_), .B(i_1_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n280_), .B(i_2_), .Y(mai_mai_n281_));
  NO2        m259(.A(mai_mai_n55_), .B(i_6_), .Y(mai_mai_n282_));
  NA3        m260(.A(mai_mai_n282_), .B(mai_mai_n281_), .C(mai_mai_n157_), .Y(mai_mai_n283_));
  OAI210     m261(.A0(mai_mai_n159_), .A1(mai_mai_n137_), .B0(mai_mai_n283_), .Y(mai_mai_n284_));
  NO3        m262(.A(mai_mai_n284_), .B(mai_mai_n279_), .C(mai_mai_n274_), .Y(mai_mai_n285_));
  NO2        m263(.A(i_3_), .B(i_10_), .Y(mai_mai_n286_));
  NA3        m264(.A(mai_mai_n286_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n287_));
  NO2        m265(.A(i_2_), .B(mai_mai_n98_), .Y(mai_mai_n288_));
  NO2        m266(.A(i_4_), .B(i_8_), .Y(mai_mai_n289_));
  NOi21      m267(.An(mai_mai_n212_), .B(mai_mai_n100_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n290_), .B(mai_mai_n289_), .C(mai_mai_n288_), .Y(mai_mai_n291_));
  AN2        m269(.A(i_3_), .B(i_10_), .Y(mai_mai_n292_));
  NA4        m270(.A(mai_mai_n292_), .B(mai_mai_n191_), .C(mai_mai_n169_), .D(mai_mai_n167_), .Y(mai_mai_n293_));
  NO2        m271(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n295_));
  OR2        m273(.A(mai_mai_n291_), .B(mai_mai_n287_), .Y(mai_mai_n296_));
  OAI220     m274(.A0(mai_mai_n296_), .A1(i_6_), .B0(mai_mai_n285_), .B1(mai_mai_n269_), .Y(mai_mai_n297_));
  NO4        m275(.A(mai_mai_n297_), .B(mai_mai_n267_), .C(mai_mai_n209_), .D(mai_mai_n162_), .Y(mai_mai_n298_));
  NO3        m276(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n55_), .B(mai_mai_n82_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n276_), .B(mai_mai_n300_), .Y(mai_mai_n301_));
  NO3        m279(.A(i_6_), .B(mai_mai_n186_), .C(i_7_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n302_), .B(mai_mai_n191_), .Y(mai_mai_n303_));
  AOI210     m281(.A0(mai_mai_n303_), .A1(mai_mai_n301_), .B0(i_5_), .Y(mai_mai_n304_));
  NO2        m282(.A(i_2_), .B(i_3_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n223_), .B(mai_mai_n305_), .C(i_1_), .Y(mai_mai_n306_));
  NA3        m284(.A(mai_mai_n276_), .B(mai_mai_n271_), .C(mai_mai_n109_), .Y(mai_mai_n307_));
  NO2        m285(.A(i_8_), .B(i_6_), .Y(mai_mai_n308_));
  NO2        m286(.A(mai_mai_n151_), .B(mai_mai_n47_), .Y(mai_mai_n309_));
  NA3        m287(.A(mai_mai_n309_), .B(mai_mai_n308_), .C(mai_mai_n157_), .Y(mai_mai_n310_));
  NA3        m288(.A(mai_mai_n310_), .B(mai_mai_n307_), .C(mai_mai_n306_), .Y(mai_mai_n311_));
  OAI210     m289(.A0(mai_mai_n311_), .A1(mai_mai_n304_), .B0(i_4_), .Y(mai_mai_n312_));
  NO2        m290(.A(i_12_), .B(i_10_), .Y(mai_mai_n313_));
  NOi21      m291(.An(i_5_), .B(i_0_), .Y(mai_mai_n314_));
  NA4        m292(.A(mai_mai_n80_), .B(mai_mai_n36_), .C(mai_mai_n82_), .D(i_8_), .Y(mai_mai_n315_));
  NO2        m293(.A(i_6_), .B(i_8_), .Y(mai_mai_n316_));
  AN2        m294(.A(i_0_), .B(mai_mai_n316_), .Y(mai_mai_n317_));
  NO2        m295(.A(i_1_), .B(i_7_), .Y(mai_mai_n318_));
  NA3        m296(.A(mai_mai_n316_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n319_));
  NA2        m297(.A(mai_mai_n319_), .B(mai_mai_n312_), .Y(mai_mai_n320_));
  NO3        m298(.A(mai_mai_n222_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n321_));
  NO3        m299(.A(i_8_), .B(i_2_), .C(i_1_), .Y(mai_mai_n322_));
  OAI210     m300(.A0(mai_mai_n322_), .A1(mai_mai_n321_), .B0(i_6_), .Y(mai_mai_n323_));
  INV        m301(.A(mai_mai_n323_), .Y(mai_mai_n324_));
  NOi21      m302(.An(mai_mai_n147_), .B(mai_mai_n101_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n325_), .B(mai_mai_n121_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n326_), .A1(mai_mai_n324_), .B0(i_3_), .Y(mai_mai_n327_));
  NO2        m305(.A(mai_mai_n280_), .B(mai_mai_n77_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n328_), .B(mai_mai_n127_), .Y(mai_mai_n329_));
  NO2        m307(.A(mai_mai_n90_), .B(mai_mai_n186_), .Y(mai_mai_n330_));
  NA3        m308(.A(mai_mai_n290_), .B(mai_mai_n330_), .C(mai_mai_n59_), .Y(mai_mai_n331_));
  AOI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n329_), .B0(i_7_), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n186_), .B(i_9_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n333_), .B(mai_mai_n199_), .Y(mai_mai_n334_));
  NO2        m312(.A(mai_mai_n334_), .B(mai_mai_n47_), .Y(mai_mai_n335_));
  NO3        m313(.A(mai_mai_n335_), .B(mai_mai_n332_), .C(mai_mai_n279_), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n327_), .B0(mai_mai_n156_), .Y(mai_mai_n337_));
  AOI210     m315(.A0(mai_mai_n320_), .A1(mai_mai_n299_), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  NOi32      m316(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n339_));
  INV        m317(.A(mai_mai_n339_), .Y(mai_mai_n340_));
  NAi21      m318(.An(i_1_), .B(i_5_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n341_), .B(i_0_), .Y(mai_mai_n342_));
  NA2        m320(.A(mai_mai_n342_), .B(mai_mai_n25_), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n153_), .B0(mai_mai_n234_), .Y(mai_mai_n344_));
  NAi41      m322(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n345_));
  OAI220     m323(.A0(mai_mai_n345_), .A1(mai_mai_n341_), .B0(mai_mai_n213_), .B1(mai_mai_n153_), .Y(mai_mai_n346_));
  NO2        m324(.A(mai_mai_n153_), .B(mai_mai_n151_), .Y(mai_mai_n347_));
  NOi32      m325(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n348_));
  NAi21      m326(.An(i_6_), .B(i_1_), .Y(mai_mai_n349_));
  NA3        m327(.A(mai_mai_n349_), .B(mai_mai_n348_), .C(mai_mai_n47_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n350_), .B(i_0_), .Y(mai_mai_n351_));
  OR3        m329(.A(mai_mai_n351_), .B(mai_mai_n347_), .C(mai_mai_n346_), .Y(mai_mai_n352_));
  NO2        m330(.A(i_1_), .B(mai_mai_n98_), .Y(mai_mai_n353_));
  NAi21      m331(.An(i_3_), .B(i_4_), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n354_), .B(i_9_), .Y(mai_mai_n355_));
  AN2        m333(.A(i_6_), .B(i_7_), .Y(mai_mai_n356_));
  NA2        m334(.A(i_2_), .B(i_7_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n354_), .B(i_10_), .Y(mai_mai_n358_));
  NA3        m336(.A(mai_mai_n358_), .B(mai_mai_n357_), .C(mai_mai_n232_), .Y(mai_mai_n359_));
  INV        m337(.A(mai_mai_n359_), .Y(mai_mai_n360_));
  AOI220     m338(.A0(mai_mai_n358_), .A1(mai_mai_n318_), .B0(mai_mai_n227_), .B1(mai_mai_n182_), .Y(mai_mai_n361_));
  NO3        m339(.A(mai_mai_n360_), .B(mai_mai_n352_), .C(mai_mai_n344_), .Y(mai_mai_n362_));
  NO2        m340(.A(mai_mai_n362_), .B(mai_mai_n340_), .Y(mai_mai_n363_));
  AN2        m341(.A(i_12_), .B(i_5_), .Y(mai_mai_n364_));
  NO2        m342(.A(i_11_), .B(i_6_), .Y(mai_mai_n365_));
  NO2        m343(.A(mai_mai_n230_), .B(i_5_), .Y(mai_mai_n366_));
  NO2        m344(.A(i_5_), .B(i_10_), .Y(mai_mai_n367_));
  AOI220     m345(.A0(mai_mai_n367_), .A1(mai_mai_n258_), .B0(mai_mai_n366_), .B1(mai_mai_n191_), .Y(mai_mai_n368_));
  NA2        m346(.A(mai_mai_n138_), .B(mai_mai_n46_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n369_), .B(mai_mai_n368_), .Y(mai_mai_n370_));
  NA2        m348(.A(mai_mai_n370_), .B(i_7_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n372_));
  NO3        m350(.A(mai_mai_n82_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n373_));
  INV        m351(.A(i_3_), .Y(mai_mai_n374_));
  NA3        m352(.A(mai_mai_n286_), .B(mai_mai_n88_), .C(mai_mai_n52_), .Y(mai_mai_n375_));
  NO2        m353(.A(i_11_), .B(i_12_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n376_), .B(mai_mai_n36_), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n375_), .B(mai_mai_n377_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n42_), .B(i_11_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(mai_mai_n213_), .Y(mai_mai_n380_));
  NAi21      m358(.An(i_13_), .B(i_0_), .Y(mai_mai_n381_));
  NO2        m359(.A(mai_mai_n381_), .B(mai_mai_n228_), .Y(mai_mai_n382_));
  OAI210     m360(.A0(mai_mai_n380_), .A1(mai_mai_n378_), .B0(mai_mai_n382_), .Y(mai_mai_n383_));
  NA2        m361(.A(mai_mai_n383_), .B(mai_mai_n371_), .Y(mai_mai_n384_));
  NO3        m362(.A(i_1_), .B(i_12_), .C(mai_mai_n82_), .Y(mai_mai_n385_));
  NO2        m363(.A(i_0_), .B(i_11_), .Y(mai_mai_n386_));
  AN2        m364(.A(i_1_), .B(i_6_), .Y(mai_mai_n387_));
  NOi21      m365(.An(i_2_), .B(i_12_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n388_), .B(mai_mai_n387_), .Y(mai_mai_n389_));
  INV        m367(.A(mai_mai_n389_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n391_));
  NO2        m369(.A(mai_mai_n391_), .B(i_4_), .Y(mai_mai_n392_));
  NA2        m370(.A(mai_mai_n390_), .B(mai_mai_n392_), .Y(mai_mai_n393_));
  NAi21      m371(.An(i_9_), .B(i_4_), .Y(mai_mai_n394_));
  OR2        m372(.A(i_13_), .B(i_10_), .Y(mai_mai_n395_));
  NO3        m373(.A(mai_mai_n395_), .B(mai_mai_n114_), .C(mai_mai_n394_), .Y(mai_mai_n396_));
  OR2        m374(.A(mai_mai_n211_), .B(mai_mai_n210_), .Y(mai_mai_n397_));
  NO2        m375(.A(mai_mai_n98_), .B(mai_mai_n25_), .Y(mai_mai_n398_));
  NA2        m376(.A(mai_mai_n268_), .B(mai_mai_n398_), .Y(mai_mai_n399_));
  NA2        m377(.A(i_5_), .B(mai_mai_n205_), .Y(mai_mai_n400_));
  OAI220     m378(.A0(mai_mai_n400_), .A1(mai_mai_n397_), .B0(mai_mai_n399_), .B1(mai_mai_n325_), .Y(mai_mai_n401_));
  INV        m379(.A(mai_mai_n401_), .Y(mai_mai_n402_));
  AOI210     m380(.A0(mai_mai_n402_), .A1(mai_mai_n393_), .B0(mai_mai_n26_), .Y(mai_mai_n403_));
  NA2        m381(.A(mai_mai_n307_), .B(mai_mai_n306_), .Y(mai_mai_n404_));
  AOI220     m382(.A0(mai_mai_n282_), .A1(mai_mai_n272_), .B0(mai_mai_n276_), .B1(mai_mai_n300_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n405_), .B(i_5_), .Y(mai_mai_n406_));
  AOI220     m384(.A0(i_3_), .A1(mai_mai_n281_), .B0(i_6_), .B1(mai_mai_n205_), .Y(mai_mai_n407_));
  NO2        m385(.A(mai_mai_n407_), .B(mai_mai_n270_), .Y(mai_mai_n408_));
  NO3        m386(.A(mai_mai_n408_), .B(mai_mai_n406_), .C(mai_mai_n404_), .Y(mai_mai_n409_));
  NA2        m387(.A(mai_mai_n189_), .B(mai_mai_n93_), .Y(mai_mai_n410_));
  NA3        m388(.A(mai_mai_n309_), .B(mai_mai_n157_), .C(mai_mai_n82_), .Y(mai_mai_n411_));
  AOI210     m389(.A0(mai_mai_n411_), .A1(mai_mai_n410_), .B0(i_8_), .Y(mai_mai_n412_));
  NA2        m390(.A(mai_mai_n186_), .B(i_10_), .Y(mai_mai_n413_));
  NA3        m391(.A(mai_mai_n244_), .B(mai_mai_n60_), .C(i_2_), .Y(mai_mai_n414_));
  NA2        m392(.A(mai_mai_n282_), .B(mai_mai_n224_), .Y(mai_mai_n415_));
  OAI220     m393(.A0(mai_mai_n415_), .A1(mai_mai_n176_), .B0(mai_mai_n414_), .B1(mai_mai_n413_), .Y(mai_mai_n416_));
  NO2        m394(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n417_));
  NA3        m395(.A(mai_mai_n318_), .B(mai_mai_n317_), .C(mai_mai_n417_), .Y(mai_mai_n418_));
  INV        m396(.A(mai_mai_n418_), .Y(mai_mai_n419_));
  NO3        m397(.A(mai_mai_n419_), .B(mai_mai_n416_), .C(mai_mai_n412_), .Y(mai_mai_n420_));
  AOI210     m398(.A0(mai_mai_n420_), .A1(mai_mai_n409_), .B0(mai_mai_n259_), .Y(mai_mai_n421_));
  NO4        m399(.A(mai_mai_n421_), .B(mai_mai_n403_), .C(mai_mai_n384_), .D(mai_mai_n363_), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n69_), .B(i_13_), .Y(mai_mai_n423_));
  NO2        m401(.A(i_10_), .B(i_9_), .Y(mai_mai_n424_));
  NAi21      m402(.An(i_12_), .B(i_8_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n425_), .B(i_3_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n295_), .B(i_0_), .Y(mai_mai_n427_));
  NO3        m405(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n428_));
  NA2        m406(.A(mai_mai_n256_), .B(mai_mai_n94_), .Y(mai_mai_n429_));
  NA2        m407(.A(mai_mai_n429_), .B(mai_mai_n428_), .Y(mai_mai_n430_));
  NA2        m408(.A(i_8_), .B(i_9_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n268_), .B(mai_mai_n199_), .Y(mai_mai_n432_));
  OAI220     m410(.A0(mai_mai_n432_), .A1(mai_mai_n431_), .B0(mai_mai_n430_), .B1(mai_mai_n427_), .Y(mai_mai_n433_));
  NA2        m411(.A(mai_mai_n238_), .B(mai_mai_n294_), .Y(mai_mai_n434_));
  NO3        m412(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n435_));
  INV        m413(.A(mai_mai_n435_), .Y(mai_mai_n436_));
  NA3        m414(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n437_));
  NA4        m415(.A(mai_mai_n139_), .B(mai_mai_n112_), .C(mai_mai_n76_), .D(mai_mai_n23_), .Y(mai_mai_n438_));
  OAI220     m416(.A0(mai_mai_n438_), .A1(mai_mai_n437_), .B0(mai_mai_n436_), .B1(mai_mai_n434_), .Y(mai_mai_n439_));
  NO2        m417(.A(mai_mai_n439_), .B(mai_mai_n433_), .Y(mai_mai_n440_));
  NA2        m418(.A(mai_mai_n281_), .B(mai_mai_n105_), .Y(mai_mai_n441_));
  OR2        m419(.A(mai_mai_n441_), .B(mai_mai_n201_), .Y(mai_mai_n442_));
  BUFFER     m420(.A(mai_mai_n283_), .Y(mai_mai_n443_));
  OA220      m421(.A0(mai_mai_n443_), .A1(mai_mai_n156_), .B0(mai_mai_n442_), .B1(mai_mai_n221_), .Y(mai_mai_n444_));
  NA2        m422(.A(mai_mai_n93_), .B(i_13_), .Y(mai_mai_n445_));
  NO3        m423(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n446_));
  NO2        m424(.A(i_6_), .B(i_7_), .Y(mai_mai_n447_));
  NA2        m425(.A(mai_mai_n447_), .B(mai_mai_n446_), .Y(mai_mai_n448_));
  NO2        m426(.A(i_11_), .B(i_1_), .Y(mai_mai_n449_));
  OR2        m427(.A(i_11_), .B(i_8_), .Y(mai_mai_n450_));
  NOi21      m428(.An(i_2_), .B(i_7_), .Y(mai_mai_n451_));
  NAi31      m429(.An(mai_mai_n450_), .B(mai_mai_n451_), .C(i_0_), .Y(mai_mai_n452_));
  NO2        m430(.A(mai_mai_n395_), .B(i_6_), .Y(mai_mai_n453_));
  NA2        m431(.A(mai_mai_n453_), .B(i_1_), .Y(mai_mai_n454_));
  NO2        m432(.A(mai_mai_n454_), .B(mai_mai_n452_), .Y(mai_mai_n455_));
  NO2        m433(.A(i_3_), .B(mai_mai_n186_), .Y(mai_mai_n456_));
  NO2        m434(.A(i_6_), .B(i_10_), .Y(mai_mai_n457_));
  NA4        m435(.A(mai_mai_n457_), .B(mai_mai_n299_), .C(mai_mai_n456_), .D(mai_mai_n226_), .Y(mai_mai_n458_));
  NO2        m436(.A(mai_mai_n458_), .B(mai_mai_n149_), .Y(mai_mai_n459_));
  NA2        m437(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n460_));
  NO2        m438(.A(mai_mai_n151_), .B(i_3_), .Y(mai_mai_n461_));
  NAi31      m439(.An(mai_mai_n460_), .B(mai_mai_n461_), .C(mai_mai_n218_), .Y(mai_mai_n462_));
  INV        m440(.A(mai_mai_n462_), .Y(mai_mai_n463_));
  NO3        m441(.A(mai_mai_n463_), .B(mai_mai_n459_), .C(mai_mai_n455_), .Y(mai_mai_n464_));
  NA2        m442(.A(mai_mai_n428_), .B(mai_mai_n364_), .Y(mai_mai_n465_));
  NAi21      m443(.An(mai_mai_n211_), .B(mai_mai_n376_), .Y(mai_mai_n466_));
  NO2        m444(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n467_));
  NA3        m445(.A(i_6_), .B(mai_mai_n467_), .C(mai_mai_n136_), .Y(mai_mai_n468_));
  OR3        m446(.A(i_4_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n469_));
  NO2        m447(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  NA2        m448(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n471_));
  NA2        m449(.A(mai_mai_n299_), .B(mai_mai_n227_), .Y(mai_mai_n472_));
  OAI220     m450(.A0(mai_mai_n472_), .A1(mai_mai_n414_), .B0(mai_mai_n471_), .B1(mai_mai_n445_), .Y(mai_mai_n473_));
  NA4        m451(.A(mai_mai_n292_), .B(mai_mai_n216_), .C(mai_mai_n69_), .D(mai_mai_n226_), .Y(mai_mai_n474_));
  NO2        m452(.A(mai_mai_n474_), .B(mai_mai_n448_), .Y(mai_mai_n475_));
  NO3        m453(.A(mai_mai_n475_), .B(mai_mai_n473_), .C(mai_mai_n470_), .Y(mai_mai_n476_));
  NA4        m454(.A(mai_mai_n476_), .B(mai_mai_n464_), .C(mai_mai_n444_), .D(mai_mai_n440_), .Y(mai_mai_n477_));
  NA3        m455(.A(mai_mai_n292_), .B(mai_mai_n169_), .C(mai_mai_n167_), .Y(mai_mai_n478_));
  OAI210     m456(.A0(mai_mai_n287_), .A1(mai_mai_n174_), .B0(mai_mai_n478_), .Y(mai_mai_n479_));
  AN2        m457(.A(mai_mai_n272_), .B(mai_mai_n223_), .Y(mai_mai_n480_));
  NA2        m458(.A(mai_mai_n480_), .B(mai_mai_n479_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n299_), .B(mai_mai_n158_), .Y(mai_mai_n482_));
  OAI210     m460(.A0(mai_mai_n482_), .A1(mai_mai_n221_), .B0(mai_mai_n293_), .Y(mai_mai_n483_));
  NA2        m461(.A(mai_mai_n483_), .B(mai_mai_n308_), .Y(mai_mai_n484_));
  NA2        m462(.A(mai_mai_n364_), .B(mai_mai_n217_), .Y(mai_mai_n485_));
  NA2        m463(.A(mai_mai_n339_), .B(mai_mai_n69_), .Y(mai_mai_n486_));
  NA2        m464(.A(mai_mai_n356_), .B(mai_mai_n348_), .Y(mai_mai_n487_));
  OR2        m465(.A(mai_mai_n485_), .B(mai_mai_n487_), .Y(mai_mai_n488_));
  NO2        m466(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n489_));
  NAi41      m467(.An(mai_mai_n486_), .B(mai_mai_n457_), .C(mai_mai_n489_), .D(mai_mai_n47_), .Y(mai_mai_n490_));
  AOI210     m468(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n396_), .Y(mai_mai_n491_));
  NA3        m469(.A(mai_mai_n491_), .B(mai_mai_n490_), .C(mai_mai_n488_), .Y(mai_mai_n492_));
  INV        m470(.A(mai_mai_n492_), .Y(mai_mai_n493_));
  AOI210     m471(.A0(mai_mai_n187_), .A1(i_9_), .B0(mai_mai_n255_), .Y(mai_mai_n494_));
  NO2        m472(.A(mai_mai_n494_), .B(mai_mai_n192_), .Y(mai_mai_n495_));
  NO2        m473(.A(mai_mai_n176_), .B(mai_mai_n82_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n496_), .B(mai_mai_n495_), .Y(mai_mai_n497_));
  NA4        m475(.A(mai_mai_n497_), .B(mai_mai_n493_), .C(mai_mai_n484_), .D(mai_mai_n481_), .Y(mai_mai_n498_));
  NA2        m476(.A(mai_mai_n366_), .B(mai_mai_n281_), .Y(mai_mai_n499_));
  NA2        m477(.A(mai_mai_n163_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NO2        m478(.A(i_12_), .B(mai_mai_n186_), .Y(mai_mai_n501_));
  NO3        m479(.A(i_10_), .B(mai_mai_n186_), .C(mai_mai_n441_), .Y(mai_mai_n502_));
  NOi31      m480(.An(mai_mai_n302_), .B(mai_mai_n395_), .C(mai_mai_n38_), .Y(mai_mai_n503_));
  OAI210     m481(.A0(mai_mai_n503_), .A1(mai_mai_n502_), .B0(mai_mai_n500_), .Y(mai_mai_n504_));
  NO2        m482(.A(i_8_), .B(i_7_), .Y(mai_mai_n505_));
  OAI210     m483(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n506_));
  NA2        m484(.A(mai_mai_n506_), .B(mai_mai_n216_), .Y(mai_mai_n507_));
  AOI220     m485(.A0(mai_mai_n309_), .A1(mai_mai_n40_), .B0(mai_mai_n224_), .B1(mai_mai_n200_), .Y(mai_mai_n508_));
  OAI220     m486(.A0(mai_mai_n508_), .A1(mai_mai_n176_), .B0(mai_mai_n507_), .B1(mai_mai_n230_), .Y(mai_mai_n509_));
  NA2        m487(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n510_));
  NO2        m488(.A(mai_mai_n510_), .B(i_6_), .Y(mai_mai_n511_));
  NA3        m489(.A(mai_mai_n511_), .B(mai_mai_n509_), .C(mai_mai_n505_), .Y(mai_mai_n512_));
  NO2        m490(.A(mai_mai_n445_), .B(mai_mai_n128_), .Y(mai_mai_n513_));
  NA2        m491(.A(mai_mai_n513_), .B(mai_mai_n255_), .Y(mai_mai_n514_));
  NO2        m492(.A(mai_mai_n287_), .B(mai_mai_n174_), .Y(mai_mai_n515_));
  NA2        m493(.A(mai_mai_n515_), .B(mai_mai_n435_), .Y(mai_mai_n516_));
  NA4        m494(.A(mai_mai_n516_), .B(mai_mai_n514_), .C(mai_mai_n512_), .D(mai_mai_n504_), .Y(mai_mai_n517_));
  NA3        m495(.A(mai_mai_n212_), .B(mai_mai_n67_), .C(mai_mai_n45_), .Y(mai_mai_n518_));
  NA2        m496(.A(mai_mai_n268_), .B(mai_mai_n80_), .Y(mai_mai_n519_));
  AOI210     m497(.A0(mai_mai_n518_), .A1(mai_mai_n329_), .B0(mai_mai_n519_), .Y(mai_mai_n520_));
  NA2        m498(.A(mai_mai_n282_), .B(mai_mai_n272_), .Y(mai_mai_n521_));
  NO2        m499(.A(mai_mai_n521_), .B(mai_mai_n166_), .Y(mai_mai_n522_));
  NA2        m500(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n523_));
  NA2        m501(.A(mai_mai_n424_), .B(mai_mai_n214_), .Y(mai_mai_n524_));
  NO2        m502(.A(mai_mai_n523_), .B(mai_mai_n524_), .Y(mai_mai_n525_));
  NA2        m503(.A(i_0_), .B(mai_mai_n48_), .Y(mai_mai_n526_));
  NA3        m504(.A(mai_mai_n501_), .B(mai_mai_n261_), .C(mai_mai_n526_), .Y(mai_mai_n527_));
  NO2        m505(.A(i_2_), .B(mai_mai_n527_), .Y(mai_mai_n528_));
  NO4        m506(.A(mai_mai_n528_), .B(mai_mai_n525_), .C(mai_mai_n522_), .D(mai_mai_n520_), .Y(mai_mai_n529_));
  NO4        m507(.A(mai_mai_n239_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n530_));
  NO3        m508(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n222_), .B(mai_mai_n36_), .Y(mai_mai_n532_));
  AN2        m510(.A(mai_mai_n532_), .B(mai_mai_n531_), .Y(mai_mai_n533_));
  AN2        m511(.A(mai_mai_n530_), .B(mai_mai_n339_), .Y(mai_mai_n534_));
  NO2        m512(.A(mai_mai_n395_), .B(i_1_), .Y(mai_mai_n535_));
  NOi31      m513(.An(mai_mai_n535_), .B(mai_mai_n429_), .C(mai_mai_n69_), .Y(mai_mai_n536_));
  AN4        m514(.A(mai_mai_n536_), .B(mai_mai_n392_), .C(mai_mai_n467_), .D(i_2_), .Y(mai_mai_n537_));
  NO2        m515(.A(mai_mai_n405_), .B(mai_mai_n170_), .Y(mai_mai_n538_));
  NO3        m516(.A(mai_mai_n538_), .B(mai_mai_n537_), .C(mai_mai_n534_), .Y(mai_mai_n539_));
  NOi21      m517(.An(i_10_), .B(i_6_), .Y(mai_mai_n540_));
  NO2        m518(.A(mai_mai_n111_), .B(mai_mai_n23_), .Y(mai_mai_n541_));
  NA2        m519(.A(mai_mai_n302_), .B(mai_mai_n158_), .Y(mai_mai_n542_));
  AOI220     m520(.A0(mai_mai_n542_), .A1(mai_mai_n415_), .B0(mai_mai_n177_), .B1(mai_mai_n175_), .Y(mai_mai_n543_));
  NOi21      m521(.An(mai_mai_n140_), .B(mai_mai_n315_), .Y(mai_mai_n544_));
  NO2        m522(.A(mai_mai_n544_), .B(mai_mai_n543_), .Y(mai_mai_n545_));
  INV        m523(.A(mai_mai_n305_), .Y(mai_mai_n546_));
  NO2        m524(.A(i_12_), .B(mai_mai_n82_), .Y(mai_mai_n547_));
  NA2        m525(.A(mai_mai_n167_), .B(i_0_), .Y(mai_mai_n548_));
  NO3        m526(.A(mai_mai_n548_), .B(mai_mai_n323_), .C(mai_mai_n287_), .Y(mai_mai_n549_));
  OR2        m527(.A(i_2_), .B(i_5_), .Y(mai_mai_n550_));
  OR2        m528(.A(mai_mai_n550_), .B(mai_mai_n387_), .Y(mai_mai_n551_));
  AOI210     m529(.A0(mai_mai_n357_), .A1(mai_mai_n232_), .B0(mai_mai_n191_), .Y(mai_mai_n552_));
  AOI210     m530(.A0(mai_mai_n552_), .A1(mai_mai_n551_), .B0(mai_mai_n466_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n553_), .B(mai_mai_n549_), .Y(mai_mai_n554_));
  NA4        m532(.A(mai_mai_n554_), .B(mai_mai_n545_), .C(mai_mai_n539_), .D(mai_mai_n529_), .Y(mai_mai_n555_));
  NO4        m533(.A(mai_mai_n555_), .B(mai_mai_n517_), .C(mai_mai_n498_), .D(mai_mai_n477_), .Y(mai_mai_n556_));
  NA4        m534(.A(mai_mai_n556_), .B(mai_mai_n422_), .C(mai_mai_n338_), .D(mai_mai_n298_), .Y(mai7));
  NO2        m535(.A(mai_mai_n90_), .B(mai_mai_n52_), .Y(mai_mai_n558_));
  NA2        m536(.A(mai_mai_n457_), .B(mai_mai_n80_), .Y(mai_mai_n559_));
  NA2        m537(.A(i_11_), .B(mai_mai_n186_), .Y(mai_mai_n560_));
  NA3        m538(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n561_));
  NO2        m539(.A(mai_mai_n226_), .B(i_4_), .Y(mai_mai_n562_));
  NO2        m540(.A(mai_mai_n102_), .B(mai_mai_n561_), .Y(mai_mai_n563_));
  NA2        m541(.A(i_2_), .B(mai_mai_n82_), .Y(mai_mai_n564_));
  OAI210     m542(.A0(mai_mai_n85_), .A1(mai_mai_n196_), .B0(mai_mai_n197_), .Y(mai_mai_n565_));
  NO2        m543(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n566_));
  NA2        m544(.A(i_4_), .B(i_8_), .Y(mai_mai_n567_));
  AOI210     m545(.A0(mai_mai_n567_), .A1(mai_mai_n292_), .B0(mai_mai_n566_), .Y(mai_mai_n568_));
  NO2        m546(.A(mai_mai_n568_), .B(mai_mai_n564_), .Y(mai_mai_n569_));
  NO3        m547(.A(mai_mai_n569_), .B(mai_mai_n563_), .C(mai_mai_n558_), .Y(mai_mai_n570_));
  AOI210     m548(.A0(i_3_), .A1(mai_mai_n58_), .B0(i_10_), .Y(mai_mai_n571_));
  AOI210     m549(.A0(mai_mai_n571_), .A1(mai_mai_n226_), .B0(mai_mai_n155_), .Y(mai_mai_n572_));
  OR2        m550(.A(i_6_), .B(i_10_), .Y(mai_mai_n573_));
  NO2        m551(.A(mai_mai_n573_), .B(mai_mai_n23_), .Y(mai_mai_n574_));
  OR3        m552(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n575_));
  NO3        m553(.A(mai_mai_n575_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n576_));
  INV        m554(.A(mai_mai_n193_), .Y(mai_mai_n577_));
  NO2        m555(.A(mai_mai_n576_), .B(mai_mai_n574_), .Y(mai_mai_n578_));
  OA220      m556(.A0(mai_mai_n578_), .A1(mai_mai_n546_), .B0(mai_mai_n572_), .B1(mai_mai_n257_), .Y(mai_mai_n579_));
  AOI210     m557(.A0(mai_mai_n579_), .A1(mai_mai_n570_), .B0(mai_mai_n59_), .Y(mai_mai_n580_));
  NOi21      m558(.An(i_11_), .B(i_7_), .Y(mai_mai_n581_));
  AO210      m559(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n582_), .B(mai_mai_n581_), .Y(mai_mai_n583_));
  NA2        m561(.A(mai_mai_n84_), .B(mai_mai_n59_), .Y(mai_mai_n584_));
  AO210      m562(.A0(mai_mai_n584_), .A1(mai_mai_n361_), .B0(mai_mai_n41_), .Y(mai_mai_n585_));
  NA2        m563(.A(mai_mai_n218_), .B(mai_mai_n59_), .Y(mai_mai_n586_));
  NA2        m564(.A(mai_mai_n388_), .B(mai_mai_n31_), .Y(mai_mai_n587_));
  OR2        m565(.A(mai_mai_n202_), .B(mai_mai_n105_), .Y(mai_mai_n588_));
  NA2        m566(.A(mai_mai_n588_), .B(mai_mai_n587_), .Y(mai_mai_n589_));
  NO2        m567(.A(mai_mai_n59_), .B(i_9_), .Y(mai_mai_n590_));
  NO2        m568(.A(mai_mai_n590_), .B(i_4_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n591_), .B(mai_mai_n589_), .Y(mai_mai_n592_));
  NO2        m570(.A(i_1_), .B(i_12_), .Y(mai_mai_n593_));
  NA3        m571(.A(mai_mai_n593_), .B(mai_mai_n106_), .C(mai_mai_n24_), .Y(mai_mai_n594_));
  BUFFER     m572(.A(mai_mai_n594_), .Y(mai_mai_n595_));
  NA4        m573(.A(mai_mai_n595_), .B(mai_mai_n592_), .C(mai_mai_n586_), .D(mai_mai_n585_), .Y(mai_mai_n596_));
  NA2        m574(.A(mai_mai_n596_), .B(i_6_), .Y(mai_mai_n597_));
  NO2        m575(.A(i_6_), .B(i_11_), .Y(mai_mai_n598_));
  INV        m576(.A(mai_mai_n430_), .Y(mai_mai_n599_));
  NO4        m577(.A(mai_mai_n210_), .B(i_3_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n600_));
  NA2        m578(.A(mai_mai_n600_), .B(mai_mai_n590_), .Y(mai_mai_n601_));
  NA2        m579(.A(i_1_), .B(mai_mai_n247_), .Y(mai_mai_n602_));
  OAI210     m580(.A0(mai_mai_n602_), .A1(mai_mai_n45_), .B0(mai_mai_n601_), .Y(mai_mai_n603_));
  INV        m581(.A(i_2_), .Y(mai_mai_n604_));
  NA2        m582(.A(mai_mai_n132_), .B(i_9_), .Y(mai_mai_n605_));
  NA3        m583(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n606_));
  NO2        m584(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n607_));
  NA3        m585(.A(mai_mai_n607_), .B(mai_mai_n256_), .C(mai_mai_n45_), .Y(mai_mai_n608_));
  OAI220     m586(.A0(mai_mai_n608_), .A1(mai_mai_n606_), .B0(mai_mai_n605_), .B1(mai_mai_n604_), .Y(mai_mai_n609_));
  NO2        m587(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n610_));
  NA2        m588(.A(mai_mai_n610_), .B(mai_mai_n24_), .Y(mai_mai_n611_));
  NO3        m589(.A(mai_mai_n609_), .B(mai_mai_n603_), .C(mai_mai_n599_), .Y(mai_mai_n612_));
  NO2        m590(.A(mai_mai_n226_), .B(mai_mai_n98_), .Y(mai_mai_n613_));
  NO2        m591(.A(mai_mai_n613_), .B(mai_mai_n581_), .Y(mai_mai_n614_));
  NA2        m592(.A(mai_mai_n614_), .B(i_1_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n615_), .B(mai_mai_n575_), .Y(mai_mai_n616_));
  NA2        m594(.A(mai_mai_n616_), .B(mai_mai_n47_), .Y(mai_mai_n617_));
  NA2        m595(.A(i_3_), .B(mai_mai_n186_), .Y(mai_mai_n618_));
  NO2        m596(.A(mai_mai_n618_), .B(mai_mai_n111_), .Y(mai_mai_n619_));
  AN2        m597(.A(mai_mai_n619_), .B(mai_mai_n511_), .Y(mai_mai_n620_));
  NO2        m598(.A(mai_mai_n222_), .B(mai_mai_n45_), .Y(mai_mai_n621_));
  NO3        m599(.A(mai_mai_n621_), .B(mai_mai_n295_), .C(i_12_), .Y(mai_mai_n622_));
  NO2        m600(.A(mai_mai_n114_), .B(mai_mai_n37_), .Y(mai_mai_n623_));
  NO2        m601(.A(mai_mai_n623_), .B(i_6_), .Y(mai_mai_n624_));
  NO2        m602(.A(mai_mai_n82_), .B(i_9_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n625_), .B(mai_mai_n59_), .Y(mai_mai_n626_));
  NO2        m604(.A(mai_mai_n626_), .B(mai_mai_n593_), .Y(mai_mai_n627_));
  NO4        m605(.A(mai_mai_n627_), .B(mai_mai_n624_), .C(mai_mai_n622_), .D(i_4_), .Y(mai_mai_n628_));
  NA2        m606(.A(i_1_), .B(i_3_), .Y(mai_mai_n629_));
  NO2        m607(.A(mai_mai_n431_), .B(mai_mai_n90_), .Y(mai_mai_n630_));
  AOI210     m608(.A0(mai_mai_n621_), .A1(mai_mai_n540_), .B0(mai_mai_n630_), .Y(mai_mai_n631_));
  NO2        m609(.A(mai_mai_n631_), .B(mai_mai_n629_), .Y(mai_mai_n632_));
  NO3        m610(.A(mai_mai_n632_), .B(mai_mai_n628_), .C(mai_mai_n620_), .Y(mai_mai_n633_));
  NA4        m611(.A(mai_mai_n633_), .B(mai_mai_n617_), .C(mai_mai_n612_), .D(mai_mai_n597_), .Y(mai_mai_n634_));
  NO3        m612(.A(mai_mai_n450_), .B(i_3_), .C(i_7_), .Y(mai_mai_n635_));
  NOi21      m613(.An(mai_mai_n635_), .B(i_10_), .Y(mai_mai_n636_));
  OA210      m614(.A0(mai_mai_n636_), .A1(mai_mai_n233_), .B0(mai_mai_n82_), .Y(mai_mai_n637_));
  NA2        m615(.A(mai_mai_n356_), .B(mai_mai_n355_), .Y(mai_mai_n638_));
  NA3        m616(.A(mai_mai_n457_), .B(mai_mai_n489_), .C(mai_mai_n47_), .Y(mai_mai_n639_));
  NO3        m617(.A(mai_mai_n451_), .B(mai_mai_n567_), .C(mai_mai_n82_), .Y(mai_mai_n640_));
  NA2        m618(.A(mai_mai_n640_), .B(mai_mai_n25_), .Y(mai_mai_n641_));
  NA3        m619(.A(mai_mai_n155_), .B(mai_mai_n80_), .C(mai_mai_n82_), .Y(mai_mai_n642_));
  NA3        m620(.A(mai_mai_n642_), .B(mai_mai_n641_), .C(mai_mai_n639_), .Y(mai_mai_n643_));
  OAI210     m621(.A0(mai_mai_n643_), .A1(mai_mai_n637_), .B0(i_1_), .Y(mai_mai_n644_));
  AOI210     m622(.A0(mai_mai_n256_), .A1(mai_mai_n94_), .B0(i_1_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n354_), .B(i_2_), .Y(mai_mai_n646_));
  NA2        m624(.A(mai_mai_n646_), .B(mai_mai_n645_), .Y(mai_mai_n647_));
  AOI210     m625(.A0(mai_mai_n647_), .A1(mai_mai_n644_), .B0(i_13_), .Y(mai_mai_n648_));
  OR2        m626(.A(i_11_), .B(i_7_), .Y(mai_mai_n649_));
  NO2        m627(.A(mai_mai_n52_), .B(i_12_), .Y(mai_mai_n650_));
  INV        m628(.A(mai_mai_n650_), .Y(mai_mai_n651_));
  NA2        m629(.A(mai_mai_n233_), .B(mai_mai_n126_), .Y(mai_mai_n652_));
  OAI220     m630(.A0(mai_mai_n652_), .A1(mai_mai_n41_), .B0(mai_mai_n651_), .B1(mai_mai_n90_), .Y(mai_mai_n653_));
  INV        m631(.A(mai_mai_n653_), .Y(mai_mai_n654_));
  NA2        m632(.A(mai_mai_n365_), .B(mai_mai_n607_), .Y(mai_mai_n655_));
  NO2        m633(.A(mai_mai_n655_), .B(mai_mai_n230_), .Y(mai_mai_n656_));
  AOI210     m634(.A0(mai_mai_n425_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n657_));
  NOi31      m635(.An(mai_mai_n657_), .B(mai_mai_n559_), .C(mai_mai_n45_), .Y(mai_mai_n658_));
  NA2        m636(.A(mai_mai_n124_), .B(i_13_), .Y(mai_mai_n659_));
  NO2        m637(.A(mai_mai_n606_), .B(mai_mai_n111_), .Y(mai_mai_n660_));
  INV        m638(.A(mai_mai_n660_), .Y(mai_mai_n661_));
  OAI220     m639(.A0(mai_mai_n661_), .A1(mai_mai_n67_), .B0(mai_mai_n659_), .B1(mai_mai_n645_), .Y(mai_mai_n662_));
  NA2        m640(.A(mai_mai_n26_), .B(mai_mai_n186_), .Y(mai_mai_n663_));
  NA2        m641(.A(mai_mai_n663_), .B(i_7_), .Y(mai_mai_n664_));
  NO3        m642(.A(mai_mai_n451_), .B(mai_mai_n226_), .C(mai_mai_n82_), .Y(mai_mai_n665_));
  NA2        m643(.A(mai_mai_n665_), .B(mai_mai_n664_), .Y(mai_mai_n666_));
  NO2        m644(.A(mai_mai_n666_), .B(mai_mai_n577_), .Y(mai_mai_n667_));
  NO4        m645(.A(mai_mai_n667_), .B(mai_mai_n662_), .C(mai_mai_n658_), .D(mai_mai_n656_), .Y(mai_mai_n668_));
  OR2        m646(.A(i_11_), .B(i_6_), .Y(mai_mai_n669_));
  NA2        m647(.A(mai_mai_n562_), .B(i_7_), .Y(mai_mai_n670_));
  AOI210     m648(.A0(mai_mai_n670_), .A1(mai_mai_n661_), .B0(mai_mai_n669_), .Y(mai_mai_n671_));
  NA3        m649(.A(mai_mai_n388_), .B(mai_mai_n566_), .C(mai_mai_n94_), .Y(mai_mai_n672_));
  NA2        m650(.A(mai_mai_n598_), .B(i_13_), .Y(mai_mai_n673_));
  NA2        m651(.A(mai_mai_n99_), .B(mai_mai_n663_), .Y(mai_mai_n674_));
  NAi21      m652(.An(i_11_), .B(i_12_), .Y(mai_mai_n675_));
  NOi41      m653(.An(mai_mai_n107_), .B(mai_mai_n675_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n676_));
  NO3        m654(.A(mai_mai_n451_), .B(mai_mai_n547_), .C(mai_mai_n567_), .Y(mai_mai_n677_));
  AOI220     m655(.A0(mai_mai_n677_), .A1(mai_mai_n299_), .B0(mai_mai_n676_), .B1(mai_mai_n674_), .Y(mai_mai_n678_));
  NA3        m656(.A(mai_mai_n678_), .B(mai_mai_n673_), .C(mai_mai_n672_), .Y(mai_mai_n679_));
  OAI210     m657(.A0(mai_mai_n679_), .A1(mai_mai_n671_), .B0(mai_mai_n59_), .Y(mai_mai_n680_));
  NO3        m658(.A(i_9_), .B(i_3_), .C(mai_mai_n562_), .Y(mai_mai_n681_));
  NA2        m659(.A(mai_mai_n681_), .B(mai_mai_n353_), .Y(mai_mai_n682_));
  NO2        m660(.A(i_3_), .B(i_2_), .Y(mai_mai_n683_));
  NA2        m661(.A(mai_mai_n683_), .B(mai_mai_n593_), .Y(mai_mai_n684_));
  NA2        m662(.A(mai_mai_n684_), .B(mai_mai_n682_), .Y(mai_mai_n685_));
  NA3        m663(.A(mai_mai_n685_), .B(mai_mai_n46_), .C(mai_mai_n217_), .Y(mai_mai_n686_));
  NA4        m664(.A(mai_mai_n686_), .B(mai_mai_n680_), .C(mai_mai_n668_), .D(mai_mai_n654_), .Y(mai_mai_n687_));
  OR4        m665(.A(mai_mai_n687_), .B(mai_mai_n648_), .C(mai_mai_n634_), .D(mai_mai_n580_), .Y(mai5));
  NA2        m666(.A(mai_mai_n614_), .B(mai_mai_n258_), .Y(mai_mai_n689_));
  INV        m667(.A(mai_mai_n689_), .Y(mai_mai_n690_));
  NO3        m668(.A(i_11_), .B(mai_mai_n226_), .C(i_13_), .Y(mai_mai_n691_));
  NO2        m669(.A(mai_mai_n121_), .B(mai_mai_n23_), .Y(mai_mai_n692_));
  INV        m670(.A(mai_mai_n424_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n305_), .B(mai_mai_n541_), .Y(mai_mai_n694_));
  INV        m672(.A(mai_mai_n694_), .Y(mai_mai_n695_));
  NO2        m673(.A(mai_mai_n695_), .B(mai_mai_n690_), .Y(mai_mai_n696_));
  INV        m674(.A(mai_mai_n165_), .Y(mai_mai_n697_));
  INV        m675(.A(mai_mai_n233_), .Y(mai_mai_n698_));
  OAI210     m676(.A0(mai_mai_n646_), .A1(mai_mai_n426_), .B0(mai_mai_n107_), .Y(mai_mai_n699_));
  AOI210     m677(.A0(mai_mai_n699_), .A1(mai_mai_n698_), .B0(mai_mai_n697_), .Y(mai_mai_n700_));
  NO2        m678(.A(mai_mai_n431_), .B(mai_mai_n26_), .Y(mai_mai_n701_));
  NO2        m679(.A(mai_mai_n701_), .B(mai_mai_n398_), .Y(mai_mai_n702_));
  NA2        m680(.A(mai_mai_n702_), .B(i_2_), .Y(mai_mai_n703_));
  INV        m681(.A(mai_mai_n703_), .Y(mai_mai_n704_));
  AOI210     m682(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n395_), .Y(mai_mai_n705_));
  AOI210     m683(.A0(mai_mai_n705_), .A1(mai_mai_n704_), .B0(mai_mai_n700_), .Y(mai_mai_n706_));
  NO2        m684(.A(mai_mai_n183_), .B(mai_mai_n122_), .Y(mai_mai_n707_));
  OAI210     m685(.A0(mai_mai_n707_), .A1(mai_mai_n692_), .B0(i_2_), .Y(mai_mai_n708_));
  INV        m686(.A(mai_mai_n166_), .Y(mai_mai_n709_));
  NO3        m687(.A(mai_mai_n582_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n710_));
  AOI210     m688(.A0(mai_mai_n709_), .A1(mai_mai_n85_), .B0(mai_mai_n710_), .Y(mai_mai_n711_));
  AOI210     m689(.A0(mai_mai_n711_), .A1(mai_mai_n708_), .B0(mai_mai_n186_), .Y(mai_mai_n712_));
  OA210      m690(.A0(mai_mai_n583_), .A1(mai_mai_n123_), .B0(i_13_), .Y(mai_mai_n713_));
  NA2        m691(.A(mai_mai_n193_), .B(mai_mai_n196_), .Y(mai_mai_n714_));
  INV        m692(.A(mai_mai_n145_), .Y(mai_mai_n715_));
  AOI210     m693(.A0(mai_mai_n715_), .A1(mai_mai_n714_), .B0(mai_mai_n357_), .Y(mai_mai_n716_));
  AOI210     m694(.A0(mai_mai_n202_), .A1(mai_mai_n142_), .B0(mai_mai_n489_), .Y(mai_mai_n717_));
  NA2        m695(.A(mai_mai_n717_), .B(mai_mai_n398_), .Y(mai_mai_n718_));
  NO2        m696(.A(mai_mai_n99_), .B(mai_mai_n45_), .Y(mai_mai_n719_));
  INV        m697(.A(mai_mai_n288_), .Y(mai_mai_n720_));
  NA4        m698(.A(mai_mai_n720_), .B(mai_mai_n292_), .C(mai_mai_n121_), .D(mai_mai_n43_), .Y(mai_mai_n721_));
  OAI210     m699(.A0(mai_mai_n721_), .A1(mai_mai_n719_), .B0(mai_mai_n718_), .Y(mai_mai_n722_));
  NO4        m700(.A(mai_mai_n722_), .B(mai_mai_n716_), .C(mai_mai_n713_), .D(mai_mai_n712_), .Y(mai_mai_n723_));
  NA2        m701(.A(mai_mai_n541_), .B(mai_mai_n28_), .Y(mai_mai_n724_));
  NA2        m702(.A(mai_mai_n691_), .B(mai_mai_n262_), .Y(mai_mai_n725_));
  NA2        m703(.A(mai_mai_n725_), .B(mai_mai_n724_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n58_), .B(i_12_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n727_), .B(mai_mai_n123_), .Y(mai_mai_n728_));
  NO2        m706(.A(mai_mai_n728_), .B(mai_mai_n560_), .Y(mai_mai_n729_));
  AOI220     m707(.A0(mai_mai_n729_), .A1(mai_mai_n36_), .B0(mai_mai_n726_), .B1(mai_mai_n47_), .Y(mai_mai_n730_));
  NA4        m708(.A(mai_mai_n730_), .B(mai_mai_n723_), .C(mai_mai_n706_), .D(mai_mai_n696_), .Y(mai6));
  NO3        m709(.A(i_9_), .B(mai_mai_n294_), .C(i_1_), .Y(mai_mai_n732_));
  NO2        m710(.A(mai_mai_n179_), .B(mai_mai_n133_), .Y(mai_mai_n733_));
  OAI210     m711(.A0(mai_mai_n733_), .A1(mai_mai_n732_), .B0(mai_mai_n683_), .Y(mai_mai_n734_));
  NA4        m712(.A(mai_mai_n367_), .B(mai_mai_n456_), .C(mai_mai_n67_), .D(mai_mai_n98_), .Y(mai_mai_n735_));
  INV        m713(.A(mai_mai_n735_), .Y(mai_mai_n736_));
  NO2        m714(.A(mai_mai_n213_), .B(mai_mai_n460_), .Y(mai_mai_n737_));
  NO2        m715(.A(i_11_), .B(i_9_), .Y(mai_mai_n738_));
  NO2        m716(.A(mai_mai_n736_), .B(mai_mai_n314_), .Y(mai_mai_n739_));
  AO210      m717(.A0(mai_mai_n739_), .A1(mai_mai_n734_), .B0(i_12_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n358_), .B(mai_mai_n318_), .Y(mai_mai_n741_));
  NA2        m719(.A(mai_mai_n547_), .B(mai_mai_n59_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n636_), .B(mai_mai_n67_), .Y(mai_mai_n743_));
  BUFFER     m721(.A(mai_mai_n584_), .Y(mai_mai_n744_));
  NA4        m722(.A(mai_mai_n744_), .B(mai_mai_n743_), .C(mai_mai_n742_), .D(mai_mai_n741_), .Y(mai_mai_n745_));
  INV        m723(.A(mai_mai_n190_), .Y(mai_mai_n746_));
  AOI220     m724(.A0(mai_mai_n746_), .A1(mai_mai_n738_), .B0(mai_mai_n745_), .B1(mai_mai_n69_), .Y(mai_mai_n747_));
  INV        m725(.A(mai_mai_n313_), .Y(mai_mai_n748_));
  NA2        m726(.A(mai_mai_n71_), .B(mai_mai_n126_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n749_), .B(mai_mai_n748_), .Y(mai_mai_n750_));
  NO2        m728(.A(mai_mai_n239_), .B(i_9_), .Y(mai_mai_n751_));
  NA2        m729(.A(mai_mai_n751_), .B(mai_mai_n727_), .Y(mai_mai_n752_));
  AOI210     m730(.A0(mai_mai_n752_), .A1(mai_mai_n487_), .B0(mai_mai_n179_), .Y(mai_mai_n753_));
  NAi32      m731(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n754_));
  NO2        m732(.A(mai_mai_n669_), .B(mai_mai_n754_), .Y(mai_mai_n755_));
  OAI210     m733(.A0(mai_mai_n635_), .A1(mai_mai_n532_), .B0(mai_mai_n531_), .Y(mai_mai_n756_));
  NAi21      m734(.An(mai_mai_n755_), .B(mai_mai_n756_), .Y(mai_mai_n757_));
  OR3        m735(.A(mai_mai_n757_), .B(mai_mai_n753_), .C(mai_mai_n750_), .Y(mai_mai_n758_));
  NO2        m736(.A(mai_mai_n649_), .B(i_2_), .Y(mai_mai_n759_));
  NA2        m737(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n760_));
  NO2        m738(.A(mai_mai_n760_), .B(mai_mai_n387_), .Y(mai_mai_n761_));
  NA2        m739(.A(mai_mai_n761_), .B(mai_mai_n759_), .Y(mai_mai_n762_));
  AO220      m740(.A0(mai_mai_n342_), .A1(mai_mai_n333_), .B0(mai_mai_n373_), .B1(mai_mai_n560_), .Y(mai_mai_n763_));
  NA3        m741(.A(mai_mai_n763_), .B(mai_mai_n243_), .C(i_7_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n426_), .B(mai_mai_n141_), .Y(mai_mai_n765_));
  OR2        m743(.A(mai_mai_n693_), .B(mai_mai_n36_), .Y(mai_mai_n766_));
  NA4        m744(.A(mai_mai_n766_), .B(mai_mai_n765_), .C(mai_mai_n764_), .D(mai_mai_n762_), .Y(mai_mai_n767_));
  OAI210     m745(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n83_), .Y(mai_mai_n768_));
  AOI220     m746(.A0(mai_mai_n768_), .A1(mai_mai_n531_), .B0(mai_mai_n737_), .B1(mai_mai_n664_), .Y(mai_mai_n769_));
  NA2        m747(.A(mai_mai_n373_), .B(mai_mai_n66_), .Y(mai_mai_n770_));
  NA3        m748(.A(mai_mai_n770_), .B(mai_mai_n769_), .C(mai_mai_n565_), .Y(mai_mai_n771_));
  AO210      m749(.A0(mai_mai_n489_), .A1(mai_mai_n47_), .B0(mai_mai_n84_), .Y(mai_mai_n772_));
  NA3        m750(.A(mai_mai_n772_), .B(mai_mai_n457_), .C(mai_mai_n212_), .Y(mai_mai_n773_));
  AOI210     m751(.A0(mai_mai_n426_), .A1(mai_mai_n424_), .B0(mai_mai_n530_), .Y(mai_mai_n774_));
  NA2        m752(.A(mai_mai_n108_), .B(mai_mai_n386_), .Y(mai_mai_n775_));
  INV        m753(.A(mai_mai_n551_), .Y(mai_mai_n776_));
  NA3        m754(.A(mai_mai_n776_), .B(mai_mai_n313_), .C(i_7_), .Y(mai_mai_n777_));
  NA4        m755(.A(mai_mai_n777_), .B(mai_mai_n775_), .C(mai_mai_n774_), .D(mai_mai_n773_), .Y(mai_mai_n778_));
  NO4        m756(.A(mai_mai_n778_), .B(mai_mai_n771_), .C(mai_mai_n767_), .D(mai_mai_n758_), .Y(mai_mai_n779_));
  NA4        m757(.A(mai_mai_n779_), .B(mai_mai_n747_), .C(mai_mai_n740_), .D(mai_mai_n362_), .Y(mai3));
  NA2        m758(.A(i_12_), .B(i_10_), .Y(mai_mai_n781_));
  NA2        m759(.A(i_6_), .B(i_7_), .Y(mai_mai_n782_));
  NO2        m760(.A(mai_mai_n782_), .B(i_0_), .Y(mai_mai_n783_));
  NO2        m761(.A(i_11_), .B(mai_mai_n226_), .Y(mai_mai_n784_));
  NA2        m762(.A(mai_mai_n276_), .B(mai_mai_n784_), .Y(mai_mai_n785_));
  NO2        m763(.A(mai_mai_n785_), .B(mai_mai_n186_), .Y(mai_mai_n786_));
  NO3        m764(.A(mai_mai_n427_), .B(mai_mai_n87_), .C(mai_mai_n45_), .Y(mai_mai_n787_));
  OA210      m765(.A0(mai_mai_n787_), .A1(mai_mai_n786_), .B0(mai_mai_n167_), .Y(mai_mai_n788_));
  NO2        m766(.A(mai_mai_n588_), .B(mai_mai_n431_), .Y(mai_mai_n789_));
  NA2        m767(.A(mai_mai_n388_), .B(mai_mai_n46_), .Y(mai_mai_n790_));
  NO2        m768(.A(mai_mai_n962_), .B(mai_mai_n48_), .Y(mai_mai_n791_));
  NA2        m769(.A(mai_mai_n657_), .B(mai_mai_n625_), .Y(mai_mai_n792_));
  NA2        m770(.A(i_0_), .B(mai_mai_n417_), .Y(mai_mai_n793_));
  NO2        m771(.A(mai_mai_n793_), .B(mai_mai_n792_), .Y(mai_mai_n794_));
  NOi21      m772(.An(i_5_), .B(i_9_), .Y(mai_mai_n795_));
  NA2        m773(.A(mai_mai_n795_), .B(mai_mai_n423_), .Y(mai_mai_n796_));
  BUFFER     m774(.A(mai_mai_n256_), .Y(mai_mai_n797_));
  AOI210     m775(.A0(mai_mai_n797_), .A1(mai_mai_n449_), .B0(mai_mai_n640_), .Y(mai_mai_n798_));
  NO3        m776(.A(mai_mai_n391_), .B(mai_mai_n256_), .C(mai_mai_n69_), .Y(mai_mai_n799_));
  NO2        m777(.A(mai_mai_n168_), .B(mai_mai_n142_), .Y(mai_mai_n800_));
  AOI210     m778(.A0(mai_mai_n800_), .A1(mai_mai_n232_), .B0(mai_mai_n799_), .Y(mai_mai_n801_));
  OAI220     m779(.A0(mai_mai_n801_), .A1(mai_mai_n174_), .B0(mai_mai_n798_), .B1(mai_mai_n796_), .Y(mai_mai_n802_));
  NO4        m780(.A(mai_mai_n802_), .B(mai_mai_n794_), .C(mai_mai_n791_), .D(mai_mai_n788_), .Y(mai_mai_n803_));
  NA2        m781(.A(mai_mai_n179_), .B(mai_mai_n24_), .Y(mai_mai_n804_));
  NAi21      m782(.An(mai_mai_n156_), .B(mai_mai_n417_), .Y(mai_mai_n805_));
  NO2        m783(.A(mai_mai_n805_), .B(i_2_), .Y(mai_mai_n806_));
  INV        m784(.A(mai_mai_n806_), .Y(mai_mai_n807_));
  INV        m785(.A(mai_mai_n280_), .Y(mai_mai_n808_));
  NA2        m786(.A(mai_mai_n808_), .B(mai_mai_n660_), .Y(mai_mai_n809_));
  NO4        m787(.A(mai_mai_n550_), .B(mai_mai_n210_), .C(mai_mai_n395_), .D(mai_mai_n387_), .Y(mai_mai_n810_));
  NA2        m788(.A(mai_mai_n810_), .B(i_11_), .Y(mai_mai_n811_));
  AN2        m789(.A(mai_mai_n93_), .B(mai_mai_n231_), .Y(mai_mai_n812_));
  NA2        m790(.A(mai_mai_n691_), .B(mai_mai_n314_), .Y(mai_mai_n813_));
  INV        m791(.A(mai_mai_n54_), .Y(mai_mai_n814_));
  OAI220     m792(.A0(mai_mai_n814_), .A1(mai_mai_n813_), .B0(mai_mai_n611_), .B1(mai_mai_n507_), .Y(mai_mai_n815_));
  NO2        m793(.A(mai_mai_n241_), .B(mai_mai_n147_), .Y(mai_mai_n816_));
  INV        m794(.A(mai_mai_n510_), .Y(mai_mai_n817_));
  NO4        m795(.A(mai_mai_n111_), .B(mai_mai_n54_), .C(mai_mai_n618_), .D(i_5_), .Y(mai_mai_n818_));
  AO220      m796(.A0(mai_mai_n818_), .A1(mai_mai_n817_), .B0(mai_mai_n816_), .B1(i_6_), .Y(mai_mai_n819_));
  NA2        m797(.A(mai_mai_n179_), .B(mai_mai_n80_), .Y(mai_mai_n820_));
  NA2        m798(.A(mai_mai_n535_), .B(i_4_), .Y(mai_mai_n821_));
  NA2        m799(.A(mai_mai_n182_), .B(mai_mai_n196_), .Y(mai_mai_n822_));
  OAI220     m800(.A0(mai_mai_n822_), .A1(mai_mai_n813_), .B0(mai_mai_n821_), .B1(mai_mai_n820_), .Y(mai_mai_n823_));
  NO4        m801(.A(mai_mai_n823_), .B(mai_mai_n819_), .C(mai_mai_n815_), .D(mai_mai_n812_), .Y(mai_mai_n824_));
  NA4        m802(.A(mai_mai_n824_), .B(mai_mai_n811_), .C(mai_mai_n809_), .D(mai_mai_n807_), .Y(mai_mai_n825_));
  NA2        m803(.A(i_11_), .B(i_9_), .Y(mai_mai_n826_));
  NO2        m804(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n372_), .B(mai_mai_n172_), .Y(mai_mai_n828_));
  NA2        m806(.A(mai_mai_n828_), .B(mai_mai_n154_), .Y(mai_mai_n829_));
  NO2        m807(.A(mai_mai_n826_), .B(mai_mai_n69_), .Y(mai_mai_n830_));
  NA2        m808(.A(mai_mai_n447_), .B(mai_mai_n220_), .Y(mai_mai_n831_));
  AOI210     m809(.A0(mai_mai_n356_), .A1(mai_mai_n42_), .B0(mai_mai_n385_), .Y(mai_mai_n832_));
  OAI220     m810(.A0(mai_mai_n832_), .A1(mai_mai_n796_), .B0(mai_mai_n831_), .B1(mai_mai_n168_), .Y(mai_mai_n833_));
  NO2        m811(.A(mai_mai_n833_), .B(mai_mai_n829_), .Y(mai_mai_n834_));
  NA2        m812(.A(mai_mai_n610_), .B(mai_mai_n118_), .Y(mai_mai_n835_));
  NO2        m813(.A(i_6_), .B(mai_mai_n835_), .Y(mai_mai_n836_));
  AOI210     m814(.A0(mai_mai_n425_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n837_));
  NA2        m815(.A(mai_mai_n165_), .B(mai_mai_n100_), .Y(mai_mai_n838_));
  NOi32      m816(.An(mai_mai_n837_), .Bn(mai_mai_n182_), .C(mai_mai_n838_), .Y(mai_mai_n839_));
  NA2        m817(.A(mai_mai_n566_), .B(mai_mai_n314_), .Y(mai_mai_n840_));
  NO2        m818(.A(mai_mai_n840_), .B(mai_mai_n790_), .Y(mai_mai_n841_));
  NO3        m819(.A(mai_mai_n841_), .B(mai_mai_n839_), .C(mai_mai_n836_), .Y(mai_mai_n842_));
  INV        m820(.A(i_5_), .Y(mai_mai_n843_));
  OR2        m821(.A(mai_mai_n838_), .B(mai_mai_n487_), .Y(mai_mai_n844_));
  NO3        m822(.A(mai_mai_n381_), .B(mai_mai_n345_), .C(mai_mai_n341_), .Y(mai_mai_n845_));
  NO2        m823(.A(mai_mai_n250_), .B(i_5_), .Y(mai_mai_n846_));
  NO2        m824(.A(mai_mai_n675_), .B(mai_mai_n245_), .Y(mai_mai_n847_));
  AOI210     m825(.A0(mai_mai_n847_), .A1(mai_mai_n846_), .B0(mai_mai_n845_), .Y(mai_mai_n848_));
  NA4        m826(.A(mai_mai_n848_), .B(mai_mai_n844_), .C(mai_mai_n842_), .D(mai_mai_n834_), .Y(mai_mai_n849_));
  NO2        m827(.A(mai_mai_n804_), .B(mai_mai_n228_), .Y(mai_mai_n850_));
  AN2        m828(.A(mai_mai_n316_), .B(mai_mai_n314_), .Y(mai_mai_n851_));
  AN2        m829(.A(mai_mai_n851_), .B(mai_mai_n800_), .Y(mai_mai_n852_));
  OAI210     m830(.A0(mai_mai_n852_), .A1(mai_mai_n850_), .B0(i_10_), .Y(mai_mai_n853_));
  INV        m831(.A(mai_mai_n781_), .Y(mai_mai_n854_));
  NA2        m832(.A(mai_mai_n854_), .B(mai_mai_n830_), .Y(mai_mai_n855_));
  NA3        m833(.A(mai_mai_n446_), .B(mai_mai_n388_), .C(mai_mai_n46_), .Y(mai_mai_n856_));
  OAI210     m834(.A0(mai_mai_n805_), .A1(i_7_), .B0(mai_mai_n856_), .Y(mai_mai_n857_));
  NA2        m835(.A(mai_mai_n830_), .B(mai_mai_n292_), .Y(mai_mai_n858_));
  OAI210     m836(.A0(i_2_), .A1(mai_mai_n181_), .B0(mai_mai_n858_), .Y(mai_mai_n859_));
  AOI220     m837(.A0(mai_mai_n859_), .A1(mai_mai_n447_), .B0(mai_mai_n857_), .B1(mai_mai_n69_), .Y(mai_mai_n860_));
  NAi21      m838(.An(i_9_), .B(i_5_), .Y(mai_mai_n861_));
  NO2        m839(.A(mai_mai_n861_), .B(mai_mai_n381_), .Y(mai_mai_n862_));
  NO2        m840(.A(mai_mai_n561_), .B(mai_mai_n102_), .Y(mai_mai_n863_));
  AOI220     m841(.A0(mai_mai_n863_), .A1(i_0_), .B0(mai_mai_n862_), .B1(mai_mai_n583_), .Y(mai_mai_n864_));
  NO2        m842(.A(mai_mai_n864_), .B(mai_mai_n82_), .Y(mai_mai_n865_));
  NO2        m843(.A(mai_mai_n865_), .B(mai_mai_n492_), .Y(mai_mai_n866_));
  NA4        m844(.A(mai_mai_n866_), .B(mai_mai_n860_), .C(mai_mai_n855_), .D(mai_mai_n853_), .Y(mai_mai_n867_));
  NO3        m845(.A(mai_mai_n867_), .B(mai_mai_n849_), .C(mai_mai_n825_), .Y(mai_mai_n868_));
  NO2        m846(.A(i_0_), .B(mai_mai_n675_), .Y(mai_mai_n869_));
  NA2        m847(.A(mai_mai_n69_), .B(mai_mai_n45_), .Y(mai_mai_n870_));
  NO3        m848(.A(mai_mai_n102_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n871_));
  AO220      m849(.A0(mai_mai_n871_), .A1(mai_mai_n45_), .B0(mai_mai_n869_), .B1(mai_mai_n167_), .Y(mai_mai_n872_));
  AOI210     m850(.A0(mai_mai_n742_), .A1(mai_mai_n638_), .B0(mai_mai_n838_), .Y(mai_mai_n873_));
  AOI210     m851(.A0(mai_mai_n872_), .A1(mai_mai_n330_), .B0(mai_mai_n873_), .Y(mai_mai_n874_));
  NA3        m852(.A(mai_mai_n140_), .B(mai_mai_n625_), .C(mai_mai_n69_), .Y(mai_mai_n875_));
  NO2        m853(.A(mai_mai_n756_), .B(mai_mai_n381_), .Y(mai_mai_n876_));
  NA3        m854(.A(mai_mai_n783_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n877_));
  NA2        m855(.A(mai_mai_n784_), .B(i_9_), .Y(mai_mai_n878_));
  AOI210     m856(.A0(mai_mai_n877_), .A1(mai_mai_n468_), .B0(mai_mai_n878_), .Y(mai_mai_n879_));
  NA2        m857(.A(mai_mai_n232_), .B(mai_mai_n219_), .Y(mai_mai_n880_));
  NO2        m858(.A(mai_mai_n880_), .B(mai_mai_n147_), .Y(mai_mai_n881_));
  NO3        m859(.A(mai_mai_n881_), .B(mai_mai_n879_), .C(mai_mai_n876_), .Y(mai_mai_n882_));
  NA3        m860(.A(mai_mai_n882_), .B(mai_mai_n875_), .C(mai_mai_n874_), .Y(mai_mai_n883_));
  NA2        m861(.A(mai_mai_n851_), .B(mai_mai_n357_), .Y(mai_mai_n884_));
  AOI210     m862(.A0(mai_mai_n287_), .A1(mai_mai_n156_), .B0(mai_mai_n884_), .Y(mai_mai_n885_));
  NA3        m863(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n886_));
  NA2        m864(.A(mai_mai_n827_), .B(mai_mai_n461_), .Y(mai_mai_n887_));
  AOI210     m865(.A0(mai_mai_n886_), .A1(mai_mai_n156_), .B0(mai_mai_n887_), .Y(mai_mai_n888_));
  NO2        m866(.A(mai_mai_n888_), .B(mai_mai_n885_), .Y(mai_mai_n889_));
  NA2        m867(.A(mai_mai_n536_), .B(mai_mai_n71_), .Y(mai_mai_n890_));
  NO3        m868(.A(mai_mai_n204_), .B(mai_mai_n364_), .C(i_0_), .Y(mai_mai_n891_));
  OAI210     m869(.A0(mai_mai_n891_), .A1(mai_mai_n72_), .B0(i_13_), .Y(mai_mai_n892_));
  INV        m870(.A(mai_mai_n212_), .Y(mai_mai_n893_));
  NO2        m871(.A(i_12_), .B(mai_mai_n577_), .Y(mai_mai_n894_));
  NA3        m872(.A(mai_mai_n894_), .B(mai_mai_n374_), .C(mai_mai_n893_), .Y(mai_mai_n895_));
  NA4        m873(.A(mai_mai_n895_), .B(mai_mai_n892_), .C(mai_mai_n890_), .D(mai_mai_n889_), .Y(mai_mai_n896_));
  NA2        m874(.A(mai_mai_n843_), .B(mai_mai_n461_), .Y(mai_mai_n897_));
  NA2        m875(.A(mai_mai_n333_), .B(mai_mai_n169_), .Y(mai_mai_n898_));
  OR2        m876(.A(mai_mai_n898_), .B(mai_mai_n897_), .Y(mai_mai_n899_));
  NA3        m877(.A(mai_mai_n574_), .B(mai_mai_n179_), .C(mai_mai_n80_), .Y(mai_mai_n900_));
  INV        m878(.A(mai_mai_n900_), .Y(mai_mai_n901_));
  NO3        m879(.A(mai_mai_n790_), .B(mai_mai_n52_), .C(mai_mai_n48_), .Y(mai_mai_n902_));
  INV        m880(.A(mai_mai_n465_), .Y(mai_mai_n903_));
  NO3        m881(.A(mai_mai_n903_), .B(mai_mai_n902_), .C(mai_mai_n901_), .Y(mai_mai_n904_));
  NA3        m882(.A(mai_mai_n367_), .B(mai_mai_n165_), .C(mai_mai_n164_), .Y(mai_mai_n905_));
  NA3        m883(.A(mai_mai_n827_), .B(mai_mai_n276_), .C(mai_mai_n219_), .Y(mai_mai_n906_));
  NA2        m884(.A(mai_mai_n906_), .B(mai_mai_n905_), .Y(mai_mai_n907_));
  NA3        m885(.A(mai_mai_n367_), .B(mai_mai_n317_), .C(mai_mai_n214_), .Y(mai_mai_n908_));
  INV        m886(.A(mai_mai_n908_), .Y(mai_mai_n909_));
  NOi31      m887(.An(mai_mai_n366_), .B(mai_mai_n870_), .C(mai_mai_n228_), .Y(mai_mai_n910_));
  NO3        m888(.A(mai_mai_n826_), .B(mai_mai_n212_), .C(mai_mai_n183_), .Y(mai_mai_n911_));
  NO4        m889(.A(mai_mai_n911_), .B(mai_mai_n910_), .C(mai_mai_n909_), .D(mai_mai_n907_), .Y(mai_mai_n912_));
  NA3        m890(.A(mai_mai_n912_), .B(mai_mai_n904_), .C(mai_mai_n899_), .Y(mai_mai_n913_));
  INV        m891(.A(mai_mai_n576_), .Y(mai_mai_n914_));
  NO3        m892(.A(mai_mai_n914_), .B(mai_mai_n526_), .C(i_7_), .Y(mai_mai_n915_));
  INV        m893(.A(mai_mai_n915_), .Y(mai_mai_n916_));
  NA2        m894(.A(mai_mai_n736_), .B(mai_mai_n169_), .Y(mai_mai_n917_));
  NA3        m895(.A(mai_mai_n95_), .B(mai_mai_n540_), .C(i_11_), .Y(mai_mai_n918_));
  NO2        m896(.A(mai_mai_n918_), .B(mai_mai_n149_), .Y(mai_mai_n919_));
  INV        m897(.A(mai_mai_n919_), .Y(mai_mai_n920_));
  NA3        m898(.A(mai_mai_n920_), .B(mai_mai_n917_), .C(mai_mai_n916_), .Y(mai_mai_n921_));
  NO4        m899(.A(mai_mai_n921_), .B(mai_mai_n913_), .C(mai_mai_n896_), .D(mai_mai_n883_), .Y(mai_mai_n922_));
  NA2        m900(.A(mai_mai_n759_), .B(mai_mai_n37_), .Y(mai_mai_n923_));
  NA3        m901(.A(mai_mai_n837_), .B(mai_mai_n353_), .C(i_5_), .Y(mai_mai_n924_));
  NA3        m902(.A(mai_mai_n924_), .B(mai_mai_n923_), .C(mai_mai_n572_), .Y(mai_mai_n925_));
  NA2        m903(.A(mai_mai_n925_), .B(mai_mai_n200_), .Y(mai_mai_n926_));
  NA2        m904(.A(mai_mai_n180_), .B(mai_mai_n182_), .Y(mai_mai_n927_));
  OAI210     m905(.A0(mai_mai_n576_), .A1(mai_mai_n574_), .B0(mai_mai_n305_), .Y(mai_mai_n928_));
  NAi31      m906(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n929_));
  NO2        m907(.A(mai_mai_n66_), .B(mai_mai_n929_), .Y(mai_mai_n930_));
  INV        m908(.A(mai_mai_n930_), .Y(mai_mai_n931_));
  NA3        m909(.A(mai_mai_n931_), .B(mai_mai_n928_), .C(mai_mai_n927_), .Y(mai_mai_n932_));
  NO2        m910(.A(mai_mai_n437_), .B(mai_mai_n256_), .Y(mai_mai_n933_));
  NO4        m911(.A(mai_mai_n222_), .B(mai_mai_n139_), .C(mai_mai_n629_), .D(mai_mai_n37_), .Y(mai_mai_n934_));
  NO3        m912(.A(mai_mai_n934_), .B(mai_mai_n933_), .C(mai_mai_n810_), .Y(mai_mai_n935_));
  NA2        m913(.A(mai_mai_n918_), .B(mai_mai_n935_), .Y(mai_mai_n936_));
  AOI210     m914(.A0(mai_mai_n932_), .A1(mai_mai_n48_), .B0(mai_mai_n936_), .Y(mai_mai_n937_));
  AOI210     m915(.A0(mai_mai_n937_), .A1(mai_mai_n926_), .B0(mai_mai_n69_), .Y(mai_mai_n938_));
  INV        m916(.A(mai_mai_n533_), .Y(mai_mai_n939_));
  NO2        m917(.A(mai_mai_n939_), .B(mai_mai_n697_), .Y(mai_mai_n940_));
  NA2        m918(.A(mai_mai_n250_), .B(mai_mai_n53_), .Y(mai_mai_n941_));
  NA2        m919(.A(mai_mai_n941_), .B(mai_mai_n72_), .Y(mai_mai_n942_));
  NO2        m920(.A(mai_mai_n942_), .B(mai_mai_n226_), .Y(mai_mai_n943_));
  NA3        m921(.A(mai_mai_n93_), .B(mai_mai_n294_), .C(mai_mai_n31_), .Y(mai_mai_n944_));
  INV        m922(.A(mai_mai_n944_), .Y(mai_mai_n945_));
  NO2        m923(.A(mai_mai_n945_), .B(mai_mai_n943_), .Y(mai_mai_n946_));
  NA2        m924(.A(mai_mai_n152_), .B(mai_mai_n85_), .Y(mai_mai_n947_));
  NO2        m925(.A(mai_mai_n947_), .B(i_11_), .Y(mai_mai_n948_));
  OAI210     m926(.A0(mai_mai_n963_), .A1(mai_mai_n837_), .B0(mai_mai_n200_), .Y(mai_mai_n949_));
  NA2        m927(.A(mai_mai_n158_), .B(i_5_), .Y(mai_mai_n950_));
  NO2        m928(.A(mai_mai_n949_), .B(mai_mai_n950_), .Y(mai_mai_n951_));
  NO4        m929(.A(mai_mai_n861_), .B(mai_mai_n450_), .C(mai_mai_n240_), .D(mai_mai_n239_), .Y(mai_mai_n952_));
  NO2        m930(.A(mai_mai_n952_), .B(mai_mai_n530_), .Y(mai_mai_n953_));
  INV        m931(.A(mai_mai_n346_), .Y(mai_mai_n954_));
  AOI210     m932(.A0(mai_mai_n954_), .A1(mai_mai_n953_), .B0(mai_mai_n41_), .Y(mai_mai_n955_));
  NO3        m933(.A(mai_mai_n955_), .B(mai_mai_n951_), .C(mai_mai_n948_), .Y(mai_mai_n956_));
  OAI210     m934(.A0(mai_mai_n946_), .A1(i_4_), .B0(mai_mai_n956_), .Y(mai_mai_n957_));
  NO3        m935(.A(mai_mai_n957_), .B(mai_mai_n940_), .C(mai_mai_n938_), .Y(mai_mai_n958_));
  NA4        m936(.A(mai_mai_n958_), .B(mai_mai_n922_), .C(mai_mai_n868_), .D(mai_mai_n803_), .Y(mai4));
  INV        m937(.A(mai_mai_n789_), .Y(mai_mai_n962_));
  INV        m938(.A(i_12_), .Y(mai_mai_n963_));
  NAi21      u000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u002(.A(i_9_), .Y(men_men_n25_));
  INV        u003(.A(i_3_), .Y(men_men_n26_));
  NO2        u004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u013(.A(i_4_), .Y(men_men_n36_));
  INV        u014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u021(.A(men_men_n35_), .Y(men1));
  INV        u022(.A(i_11_), .Y(men_men_n45_));
  NO2        u023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u024(.A(i_2_), .Y(men_men_n47_));
  NA2        u025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u026(.A(i_5_), .Y(men_men_n49_));
  NO2        u027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  NA2        u034(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n57_));
  NA3        u035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n58_));
  NO2        u036(.A(i_1_), .B(i_6_), .Y(men_men_n59_));
  NA2        u037(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  OAI210     u038(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n58_), .Y(men_men_n61_));
  NA2        u039(.A(men_men_n61_), .B(i_12_), .Y(men_men_n62_));
  NAi21      u040(.An(i_2_), .B(i_7_), .Y(men_men_n63_));
  INV        u041(.A(i_1_), .Y(men_men_n64_));
  INV        u042(.A(men_men_n62_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n51_), .B(i_2_), .Y(men_men_n66_));
  AOI210     u044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n67_));
  NA2        u045(.A(i_1_), .B(i_6_), .Y(men_men_n68_));
  NO2        u046(.A(men_men_n68_), .B(men_men_n25_), .Y(men_men_n69_));
  INV        u047(.A(i_0_), .Y(men_men_n70_));
  NAi21      u048(.An(i_5_), .B(i_10_), .Y(men_men_n71_));
  NA2        u049(.A(i_5_), .B(i_9_), .Y(men_men_n72_));
  AOI210     u050(.A0(men_men_n72_), .A1(men_men_n71_), .B0(men_men_n70_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n73_), .B(men_men_n69_), .Y(men_men_n74_));
  OAI210     u052(.A0(men_men_n67_), .A1(men_men_n66_), .B0(men_men_n74_), .Y(men_men_n75_));
  OAI210     u053(.A0(men_men_n75_), .A1(men_men_n65_), .B0(i_0_), .Y(men_men_n76_));
  NA2        u054(.A(i_12_), .B(i_5_), .Y(men_men_n77_));
  NA2        u055(.A(i_2_), .B(i_8_), .Y(men_men_n78_));
  NO2        u056(.A(i_3_), .B(i_9_), .Y(men_men_n79_));
  NO2        u057(.A(i_3_), .B(i_7_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n79_), .B(men_men_n64_), .Y(men_men_n81_));
  INV        u059(.A(i_6_), .Y(men_men_n82_));
  NO2        u060(.A(i_2_), .B(i_7_), .Y(men_men_n83_));
  NA2        u061(.A(men_men_n81_), .B(i_7_), .Y(men_men_n84_));
  NAi21      u062(.An(i_6_), .B(i_10_), .Y(men_men_n85_));
  NA2        u063(.A(i_6_), .B(i_9_), .Y(men_men_n86_));
  AOI210     u064(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n64_), .Y(men_men_n87_));
  NA2        u065(.A(i_2_), .B(i_6_), .Y(men_men_n88_));
  NO3        u066(.A(men_men_n88_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n89_));
  NO2        u067(.A(men_men_n89_), .B(men_men_n87_), .Y(men_men_n90_));
  AOI210     u068(.A0(men_men_n90_), .A1(men_men_n84_), .B0(men_men_n77_), .Y(men_men_n91_));
  AN3        u069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n92_));
  NAi21      u070(.An(i_6_), .B(i_11_), .Y(men_men_n93_));
  NO2        u071(.A(i_5_), .B(i_8_), .Y(men_men_n94_));
  NOi21      u072(.An(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  AOI220     u073(.A0(men_men_n95_), .A1(men_men_n63_), .B0(men_men_n92_), .B1(men_men_n32_), .Y(men_men_n96_));
  INV        u074(.A(i_7_), .Y(men_men_n97_));
  NA2        u075(.A(men_men_n47_), .B(men_men_n97_), .Y(men_men_n98_));
  NO2        u076(.A(i_0_), .B(i_5_), .Y(men_men_n99_));
  NO2        u077(.A(men_men_n99_), .B(men_men_n82_), .Y(men_men_n100_));
  NA2        u078(.A(i_12_), .B(i_3_), .Y(men_men_n101_));
  INV        u079(.A(men_men_n101_), .Y(men_men_n102_));
  NA3        u080(.A(men_men_n102_), .B(men_men_n100_), .C(men_men_n98_), .Y(men_men_n103_));
  NAi21      u081(.An(i_7_), .B(i_11_), .Y(men_men_n104_));
  NO3        u082(.A(men_men_n104_), .B(men_men_n85_), .C(men_men_n54_), .Y(men_men_n105_));
  AN2        u083(.A(i_2_), .B(i_10_), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(i_7_), .Y(men_men_n107_));
  OR2        u085(.A(men_men_n77_), .B(men_men_n59_), .Y(men_men_n108_));
  NO2        u086(.A(i_8_), .B(men_men_n97_), .Y(men_men_n109_));
  NO3        u087(.A(men_men_n109_), .B(men_men_n108_), .C(men_men_n107_), .Y(men_men_n110_));
  NA2        u088(.A(i_12_), .B(i_7_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n64_), .B(men_men_n26_), .Y(men_men_n112_));
  NA2        u090(.A(men_men_n112_), .B(i_0_), .Y(men_men_n113_));
  NA2        u091(.A(i_11_), .B(i_12_), .Y(men_men_n114_));
  OAI210     u092(.A0(men_men_n113_), .A1(men_men_n111_), .B0(men_men_n114_), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n115_), .B(men_men_n110_), .Y(men_men_n116_));
  NAi41      u094(.An(men_men_n105_), .B(men_men_n116_), .C(men_men_n103_), .D(men_men_n96_), .Y(men_men_n117_));
  NOi21      u095(.An(i_1_), .B(i_5_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n118_), .B(i_11_), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n97_), .B(men_men_n37_), .Y(men_men_n120_));
  NA2        u098(.A(i_7_), .B(men_men_n25_), .Y(men_men_n121_));
  NA2        u099(.A(men_men_n121_), .B(men_men_n120_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(men_men_n47_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n86_), .B(men_men_n85_), .Y(men_men_n124_));
  NAi21      u102(.An(i_3_), .B(i_8_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n125_), .B(men_men_n63_), .Y(men_men_n126_));
  NOi31      u104(.An(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .Y(men_men_n127_));
  NO2        u105(.A(i_1_), .B(men_men_n82_), .Y(men_men_n128_));
  NO2        u106(.A(i_6_), .B(i_5_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n129_), .B(i_3_), .Y(men_men_n130_));
  AO210      u108(.A0(men_men_n130_), .A1(men_men_n48_), .B0(men_men_n128_), .Y(men_men_n131_));
  OAI220     u109(.A0(men_men_n131_), .A1(men_men_n104_), .B0(men_men_n127_), .B1(men_men_n119_), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n132_), .B(men_men_n117_), .C(men_men_n91_), .Y(men_men_n133_));
  NA3        u111(.A(men_men_n133_), .B(men_men_n76_), .C(men_men_n57_), .Y(men2));
  NO2        u112(.A(men_men_n64_), .B(men_men_n37_), .Y(men_men_n135_));
  NA2        u113(.A(i_6_), .B(men_men_n25_), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n136_), .B(men_men_n135_), .Y(men_men_n137_));
  NA4        u115(.A(men_men_n137_), .B(men_men_n74_), .C(men_men_n66_), .D(men_men_n30_), .Y(men0));
  AN2        u116(.A(i_8_), .B(i_7_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(i_6_), .Y(men_men_n140_));
  NO2        u118(.A(i_12_), .B(i_13_), .Y(men_men_n141_));
  NAi21      u119(.An(i_5_), .B(i_11_), .Y(men_men_n142_));
  NOi21      u120(.An(men_men_n141_), .B(men_men_n142_), .Y(men_men_n143_));
  NO2        u121(.A(i_0_), .B(i_1_), .Y(men_men_n144_));
  NA2        u122(.A(i_2_), .B(i_3_), .Y(men_men_n145_));
  NO2        u123(.A(men_men_n145_), .B(i_4_), .Y(men_men_n146_));
  NA3        u124(.A(men_men_n146_), .B(men_men_n144_), .C(men_men_n143_), .Y(men_men_n147_));
  OR2        u125(.A(men_men_n147_), .B(men_men_n25_), .Y(men_men_n148_));
  AN2        u126(.A(men_men_n141_), .B(men_men_n79_), .Y(men_men_n149_));
  NA2        u127(.A(i_1_), .B(i_5_), .Y(men_men_n150_));
  NO2        u128(.A(men_men_n70_), .B(men_men_n47_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n151_), .B(men_men_n36_), .Y(men_men_n152_));
  NO3        u130(.A(men_men_n152_), .B(men_men_n150_), .C(i_13_), .Y(men_men_n153_));
  OR2        u131(.A(i_0_), .B(i_1_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n154_), .B(men_men_n77_), .C(i_13_), .Y(men_men_n155_));
  NAi32      u133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n156_));
  NAi21      u134(.An(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  NOi21      u135(.An(i_4_), .B(i_10_), .Y(men_men_n158_));
  NA2        u136(.A(men_men_n158_), .B(men_men_n40_), .Y(men_men_n159_));
  NO2        u137(.A(i_3_), .B(i_5_), .Y(men_men_n160_));
  NO3        u138(.A(men_men_n70_), .B(i_2_), .C(i_1_), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n162_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n163_));
  NO2        u141(.A(men_men_n163_), .B(men_men_n153_), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n148_), .B0(men_men_n140_), .Y(men_men_n165_));
  NA2        u143(.A(i_3_), .B(men_men_n49_), .Y(men_men_n166_));
  NOi21      u144(.An(i_4_), .B(i_9_), .Y(men_men_n167_));
  NOi21      u145(.An(i_11_), .B(i_13_), .Y(men_men_n168_));
  NA2        u146(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NO2        u147(.A(i_4_), .B(i_5_), .Y(men_men_n170_));
  NAi21      u148(.An(i_12_), .B(i_11_), .Y(men_men_n171_));
  NO2        u149(.A(men_men_n171_), .B(i_13_), .Y(men_men_n172_));
  NA3        u150(.A(men_men_n172_), .B(men_men_n170_), .C(men_men_n79_), .Y(men_men_n173_));
  NO2        u151(.A(men_men_n173_), .B(men_men_n989_), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n70_), .B(men_men_n64_), .Y(men_men_n175_));
  NA2        u153(.A(men_men_n175_), .B(men_men_n47_), .Y(men_men_n176_));
  NA2        u154(.A(men_men_n36_), .B(i_5_), .Y(men_men_n177_));
  NAi31      u155(.An(men_men_n177_), .B(men_men_n149_), .C(i_11_), .Y(men_men_n178_));
  NA2        u156(.A(i_3_), .B(i_5_), .Y(men_men_n179_));
  AOI210     u157(.A0(men_men_n169_), .A1(men_men_n178_), .B0(men_men_n176_), .Y(men_men_n180_));
  NO2        u158(.A(men_men_n70_), .B(i_5_), .Y(men_men_n181_));
  NO2        u159(.A(i_13_), .B(i_10_), .Y(men_men_n182_));
  NA3        u160(.A(men_men_n182_), .B(men_men_n181_), .C(men_men_n45_), .Y(men_men_n183_));
  NO2        u161(.A(i_2_), .B(i_1_), .Y(men_men_n184_));
  NA2        u162(.A(men_men_n184_), .B(i_3_), .Y(men_men_n185_));
  NAi21      u163(.An(i_4_), .B(i_12_), .Y(men_men_n186_));
  NO4        u164(.A(men_men_n186_), .B(men_men_n185_), .C(men_men_n183_), .D(men_men_n25_), .Y(men_men_n187_));
  NO3        u165(.A(men_men_n187_), .B(men_men_n180_), .C(men_men_n174_), .Y(men_men_n188_));
  INV        u166(.A(i_8_), .Y(men_men_n189_));
  NA2        u167(.A(i_8_), .B(i_6_), .Y(men_men_n190_));
  NO3        u168(.A(i_3_), .B(men_men_n82_), .C(men_men_n49_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n191_), .B(men_men_n109_), .Y(men_men_n192_));
  NO3        u170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n193_));
  NA3        u171(.A(men_men_n193_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n194_));
  NO3        u172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n195_));
  NA2        u173(.A(men_men_n92_), .B(men_men_n195_), .Y(men_men_n196_));
  AOI210     u174(.A0(men_men_n196_), .A1(men_men_n194_), .B0(men_men_n192_), .Y(men_men_n197_));
  NO2        u175(.A(i_3_), .B(i_8_), .Y(men_men_n198_));
  NO3        u176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n199_));
  NA3        u177(.A(men_men_n199_), .B(men_men_n198_), .C(men_men_n40_), .Y(men_men_n200_));
  NO2        u178(.A(i_13_), .B(i_9_), .Y(men_men_n201_));
  NA3        u179(.A(men_men_n201_), .B(i_6_), .C(men_men_n189_), .Y(men_men_n202_));
  NAi21      u180(.An(i_12_), .B(i_3_), .Y(men_men_n203_));
  OR2        u181(.A(men_men_n203_), .B(men_men_n202_), .Y(men_men_n204_));
  NO2        u182(.A(men_men_n45_), .B(i_5_), .Y(men_men_n205_));
  NO3        u183(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n206_));
  INV        u184(.A(men_men_n206_), .Y(men_men_n207_));
  OAI220     u185(.A0(men_men_n207_), .A1(men_men_n204_), .B0(men_men_n59_), .B1(men_men_n200_), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n208_), .A1(i_7_), .B0(men_men_n197_), .Y(men_men_n209_));
  OAI220     u187(.A0(men_men_n209_), .A1(i_4_), .B0(men_men_n190_), .B1(men_men_n188_), .Y(men_men_n210_));
  NAi21      u188(.An(i_12_), .B(i_7_), .Y(men_men_n211_));
  NA3        u189(.A(i_13_), .B(men_men_n189_), .C(i_10_), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  NA2        u191(.A(i_0_), .B(i_5_), .Y(men_men_n214_));
  NA2        u192(.A(men_men_n214_), .B(men_men_n100_), .Y(men_men_n215_));
  OAI220     u193(.A0(men_men_n215_), .A1(men_men_n185_), .B0(men_men_n176_), .B1(men_men_n130_), .Y(men_men_n216_));
  NAi31      u194(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n36_), .B(i_13_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n70_), .B(men_men_n26_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n47_), .B(men_men_n64_), .Y(men_men_n220_));
  NA3        u198(.A(men_men_n220_), .B(men_men_n219_), .C(men_men_n218_), .Y(men_men_n221_));
  INV        u199(.A(i_13_), .Y(men_men_n222_));
  NO2        u200(.A(i_12_), .B(men_men_n222_), .Y(men_men_n223_));
  NA3        u201(.A(men_men_n223_), .B(men_men_n193_), .C(men_men_n191_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n221_), .A1(men_men_n217_), .B0(men_men_n224_), .Y(men_men_n225_));
  AOI220     u203(.A0(men_men_n225_), .A1(men_men_n139_), .B0(men_men_n216_), .B1(men_men_n213_), .Y(men_men_n226_));
  NO2        u204(.A(i_12_), .B(men_men_n37_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n179_), .B(i_4_), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n228_), .B(men_men_n227_), .Y(men_men_n229_));
  OR2        u207(.A(i_8_), .B(i_7_), .Y(men_men_n230_));
  NO2        u208(.A(men_men_n230_), .B(men_men_n82_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n54_), .B(i_1_), .Y(men_men_n232_));
  INV        u210(.A(i_12_), .Y(men_men_n233_));
  NO3        u211(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n234_));
  NA2        u212(.A(i_2_), .B(i_1_), .Y(men_men_n235_));
  NO3        u213(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n236_));
  NAi21      u214(.An(i_4_), .B(i_3_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n237_), .B(men_men_n72_), .Y(men_men_n238_));
  NO2        u216(.A(i_0_), .B(i_6_), .Y(men_men_n239_));
  NOi41      u217(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n240_));
  NA2        u218(.A(men_men_n240_), .B(men_men_n239_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n235_), .B(men_men_n179_), .Y(men_men_n242_));
  NAi21      u220(.An(men_men_n241_), .B(men_men_n242_), .Y(men_men_n243_));
  NO2        u221(.A(i_11_), .B(men_men_n222_), .Y(men_men_n244_));
  NAi21      u222(.An(i_3_), .B(i_7_), .Y(men_men_n245_));
  NO2        u223(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n246_));
  NO2        u224(.A(i_12_), .B(i_3_), .Y(men_men_n247_));
  NA2        u225(.A(men_men_n70_), .B(i_5_), .Y(men_men_n248_));
  NA3        u226(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n249_));
  INV        u227(.A(men_men_n140_), .Y(men_men_n250_));
  NA2        u228(.A(men_men_n233_), .B(i_13_), .Y(men_men_n251_));
  NO2        u229(.A(men_men_n251_), .B(men_men_n72_), .Y(men_men_n252_));
  NA2        u230(.A(men_men_n252_), .B(men_men_n250_), .Y(men_men_n253_));
  NO2        u231(.A(men_men_n230_), .B(men_men_n37_), .Y(men_men_n254_));
  NA2        u232(.A(i_12_), .B(i_6_), .Y(men_men_n255_));
  OR2        u233(.A(i_13_), .B(i_9_), .Y(men_men_n256_));
  NO3        u234(.A(men_men_n256_), .B(men_men_n255_), .C(men_men_n49_), .Y(men_men_n257_));
  NO2        u235(.A(men_men_n237_), .B(i_2_), .Y(men_men_n258_));
  NA3        u236(.A(men_men_n258_), .B(men_men_n257_), .C(men_men_n45_), .Y(men_men_n259_));
  NA2        u237(.A(men_men_n244_), .B(i_9_), .Y(men_men_n260_));
  OAI210     u238(.A0(men_men_n70_), .A1(men_men_n260_), .B0(men_men_n259_), .Y(men_men_n261_));
  NO3        u239(.A(i_11_), .B(men_men_n222_), .C(men_men_n25_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n245_), .B(i_8_), .Y(men_men_n263_));
  NO2        u241(.A(i_6_), .B(men_men_n49_), .Y(men_men_n264_));
  NA3        u242(.A(men_men_n264_), .B(men_men_n263_), .C(men_men_n262_), .Y(men_men_n265_));
  NO3        u243(.A(men_men_n26_), .B(men_men_n82_), .C(i_5_), .Y(men_men_n266_));
  NA3        u244(.A(men_men_n266_), .B(men_men_n254_), .C(men_men_n223_), .Y(men_men_n267_));
  AOI210     u245(.A0(men_men_n267_), .A1(men_men_n265_), .B0(i_1_), .Y(men_men_n268_));
  AOI210     u246(.A0(men_men_n261_), .A1(men_men_n254_), .B0(men_men_n268_), .Y(men_men_n269_));
  NA4        u247(.A(men_men_n269_), .B(men_men_n253_), .C(men_men_n243_), .D(men_men_n226_), .Y(men_men_n270_));
  NO3        u248(.A(i_12_), .B(men_men_n222_), .C(men_men_n37_), .Y(men_men_n271_));
  INV        u249(.A(men_men_n271_), .Y(men_men_n272_));
  NA2        u250(.A(i_8_), .B(men_men_n97_), .Y(men_men_n273_));
  NO3        u251(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n274_));
  AOI220     u252(.A0(men_men_n274_), .A1(men_men_n191_), .B0(men_men_n160_), .B1(men_men_n232_), .Y(men_men_n275_));
  NO2        u253(.A(men_men_n275_), .B(men_men_n273_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n235_), .B(i_0_), .Y(men_men_n277_));
  AOI220     u255(.A0(men_men_n277_), .A1(i_8_), .B0(i_1_), .B1(men_men_n139_), .Y(men_men_n278_));
  NA2        u256(.A(men_men_n264_), .B(men_men_n26_), .Y(men_men_n279_));
  NO2        u257(.A(men_men_n279_), .B(men_men_n278_), .Y(men_men_n280_));
  NA2        u258(.A(i_0_), .B(i_1_), .Y(men_men_n281_));
  NO2        u259(.A(men_men_n281_), .B(i_2_), .Y(men_men_n282_));
  NO2        u260(.A(men_men_n60_), .B(i_6_), .Y(men_men_n283_));
  NA3        u261(.A(men_men_n283_), .B(men_men_n282_), .C(men_men_n160_), .Y(men_men_n284_));
  OAI210     u262(.A0(men_men_n162_), .A1(men_men_n140_), .B0(men_men_n284_), .Y(men_men_n285_));
  NO3        u263(.A(men_men_n285_), .B(men_men_n280_), .C(men_men_n276_), .Y(men_men_n286_));
  NO2        u264(.A(i_3_), .B(i_10_), .Y(men_men_n287_));
  NA3        u265(.A(men_men_n287_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n288_));
  NO2        u266(.A(i_2_), .B(men_men_n97_), .Y(men_men_n289_));
  NA2        u267(.A(i_1_), .B(men_men_n36_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n290_), .B(i_8_), .Y(men_men_n291_));
  NA2        u269(.A(men_men_n291_), .B(men_men_n289_), .Y(men_men_n292_));
  AN2        u270(.A(i_3_), .B(i_10_), .Y(men_men_n293_));
  NA3        u271(.A(men_men_n293_), .B(men_men_n172_), .C(men_men_n170_), .Y(men_men_n294_));
  NO2        u272(.A(i_5_), .B(men_men_n37_), .Y(men_men_n295_));
  NO2        u273(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n296_));
  OR2        u274(.A(men_men_n292_), .B(men_men_n288_), .Y(men_men_n297_));
  OAI220     u275(.A0(men_men_n297_), .A1(i_6_), .B0(men_men_n286_), .B1(men_men_n272_), .Y(men_men_n298_));
  NO4        u276(.A(men_men_n298_), .B(men_men_n270_), .C(men_men_n210_), .D(men_men_n165_), .Y(men_men_n299_));
  NO3        u277(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n300_));
  NO3        u278(.A(i_6_), .B(men_men_n189_), .C(i_7_), .Y(men_men_n301_));
  NO2        u279(.A(men_men_n189_), .B(men_men_n166_), .Y(men_men_n302_));
  NO2        u280(.A(i_2_), .B(i_3_), .Y(men_men_n303_));
  OR2        u281(.A(i_0_), .B(i_5_), .Y(men_men_n304_));
  NA2        u282(.A(men_men_n214_), .B(men_men_n304_), .Y(men_men_n305_));
  NA4        u283(.A(men_men_n305_), .B(men_men_n231_), .C(men_men_n303_), .D(i_1_), .Y(men_men_n306_));
  NA3        u284(.A(men_men_n277_), .B(men_men_n160_), .C(men_men_n109_), .Y(men_men_n307_));
  NAi21      u285(.An(i_8_), .B(i_7_), .Y(men_men_n308_));
  NO2        u286(.A(men_men_n308_), .B(i_6_), .Y(men_men_n309_));
  NO2        u287(.A(men_men_n154_), .B(men_men_n47_), .Y(men_men_n310_));
  NA3        u288(.A(men_men_n310_), .B(men_men_n309_), .C(men_men_n160_), .Y(men_men_n311_));
  NA3        u289(.A(men_men_n311_), .B(men_men_n307_), .C(men_men_n306_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n312_), .A1(men_men_n302_), .B0(i_4_), .Y(men_men_n313_));
  NO2        u291(.A(i_12_), .B(i_10_), .Y(men_men_n314_));
  NOi21      u292(.An(i_5_), .B(i_0_), .Y(men_men_n315_));
  NO2        u293(.A(men_men_n290_), .B(men_men_n125_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n316_), .B(men_men_n314_), .Y(men_men_n317_));
  NO2        u295(.A(i_6_), .B(i_8_), .Y(men_men_n318_));
  NOi21      u296(.An(i_0_), .B(i_2_), .Y(men_men_n319_));
  AN2        u297(.A(men_men_n319_), .B(men_men_n318_), .Y(men_men_n320_));
  NO2        u298(.A(i_1_), .B(i_7_), .Y(men_men_n321_));
  AO220      u299(.A0(men_men_n321_), .A1(men_men_n320_), .B0(men_men_n309_), .B1(men_men_n232_), .Y(men_men_n322_));
  NA2        u300(.A(men_men_n322_), .B(men_men_n42_), .Y(men_men_n323_));
  NA3        u301(.A(men_men_n323_), .B(men_men_n317_), .C(men_men_n313_), .Y(men_men_n324_));
  NO3        u302(.A(men_men_n230_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n325_));
  NO3        u303(.A(men_men_n308_), .B(i_2_), .C(i_1_), .Y(men_men_n326_));
  OAI210     u304(.A0(men_men_n326_), .A1(men_men_n325_), .B0(i_6_), .Y(men_men_n327_));
  NA2        u305(.A(i_1_), .B(men_men_n289_), .Y(men_men_n328_));
  AOI210     u306(.A0(men_men_n328_), .A1(men_men_n327_), .B0(men_men_n305_), .Y(men_men_n329_));
  NOi21      u307(.An(men_men_n150_), .B(men_men_n100_), .Y(men_men_n330_));
  NO2        u308(.A(men_men_n330_), .B(men_men_n121_), .Y(men_men_n331_));
  OAI210     u309(.A0(men_men_n331_), .A1(men_men_n329_), .B0(i_3_), .Y(men_men_n332_));
  INV        u310(.A(men_men_n80_), .Y(men_men_n333_));
  NO2        u311(.A(men_men_n281_), .B(men_men_n78_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n334_), .B(men_men_n129_), .Y(men_men_n335_));
  NO2        u313(.A(men_men_n88_), .B(men_men_n189_), .Y(men_men_n336_));
  NA2        u314(.A(men_men_n336_), .B(men_men_n64_), .Y(men_men_n337_));
  AOI210     u315(.A0(men_men_n337_), .A1(men_men_n335_), .B0(men_men_n333_), .Y(men_men_n338_));
  NO2        u316(.A(men_men_n189_), .B(i_9_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n339_), .B(i_6_), .Y(men_men_n340_));
  NO2        u318(.A(men_men_n338_), .B(men_men_n280_), .Y(men_men_n341_));
  AOI210     u319(.A0(men_men_n341_), .A1(men_men_n332_), .B0(men_men_n159_), .Y(men_men_n342_));
  AOI210     u320(.A0(men_men_n324_), .A1(men_men_n300_), .B0(men_men_n342_), .Y(men_men_n343_));
  NOi32      u321(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n344_));
  INV        u322(.A(men_men_n344_), .Y(men_men_n345_));
  NAi21      u323(.An(i_0_), .B(i_6_), .Y(men_men_n346_));
  NAi21      u324(.An(i_1_), .B(i_5_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n348_), .B(men_men_n25_), .Y(men_men_n349_));
  OAI210     u327(.A0(men_men_n349_), .A1(men_men_n156_), .B0(men_men_n241_), .Y(men_men_n350_));
  NAi41      u328(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n351_));
  AOI210     u329(.A0(men_men_n351_), .A1(men_men_n156_), .B0(men_men_n154_), .Y(men_men_n352_));
  NOi32      u330(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n353_));
  NO2        u331(.A(i_1_), .B(men_men_n97_), .Y(men_men_n354_));
  NAi21      u332(.An(i_3_), .B(i_4_), .Y(men_men_n355_));
  NO2        u333(.A(men_men_n355_), .B(i_9_), .Y(men_men_n356_));
  AN2        u334(.A(i_6_), .B(i_7_), .Y(men_men_n357_));
  OAI210     u335(.A0(men_men_n357_), .A1(men_men_n354_), .B0(men_men_n356_), .Y(men_men_n358_));
  NA2        u336(.A(i_2_), .B(i_7_), .Y(men_men_n359_));
  NO2        u337(.A(men_men_n355_), .B(i_10_), .Y(men_men_n360_));
  NA3        u338(.A(men_men_n360_), .B(men_men_n359_), .C(men_men_n239_), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n361_), .A1(men_men_n358_), .B0(men_men_n181_), .Y(men_men_n362_));
  AOI210     u340(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n363_));
  OAI210     u341(.A0(men_men_n363_), .A1(men_men_n184_), .B0(men_men_n360_), .Y(men_men_n364_));
  AOI220     u342(.A0(men_men_n360_), .A1(men_men_n321_), .B0(men_men_n234_), .B1(men_men_n184_), .Y(men_men_n365_));
  AOI210     u343(.A0(men_men_n365_), .A1(men_men_n364_), .B0(i_5_), .Y(men_men_n366_));
  NO4        u344(.A(men_men_n366_), .B(men_men_n362_), .C(men_men_n352_), .D(men_men_n350_), .Y(men_men_n367_));
  NO2        u345(.A(men_men_n367_), .B(men_men_n345_), .Y(men_men_n368_));
  NO2        u346(.A(men_men_n60_), .B(men_men_n25_), .Y(men_men_n369_));
  AN2        u347(.A(i_12_), .B(i_5_), .Y(men_men_n370_));
  NO2        u348(.A(i_4_), .B(men_men_n26_), .Y(men_men_n371_));
  NA2        u349(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  NO2        u350(.A(i_11_), .B(i_6_), .Y(men_men_n373_));
  NA3        u351(.A(men_men_n373_), .B(men_men_n310_), .C(men_men_n222_), .Y(men_men_n374_));
  NO2        u352(.A(men_men_n374_), .B(men_men_n372_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n237_), .B(i_5_), .Y(men_men_n376_));
  NO2        u354(.A(i_5_), .B(i_10_), .Y(men_men_n377_));
  NA2        u355(.A(men_men_n376_), .B(men_men_n193_), .Y(men_men_n378_));
  NO2        u356(.A(i_12_), .B(men_men_n378_), .Y(men_men_n379_));
  OAI210     u357(.A0(men_men_n379_), .A1(men_men_n375_), .B0(men_men_n369_), .Y(men_men_n380_));
  NO2        u358(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n381_));
  INV        u359(.A(men_men_n147_), .Y(men_men_n382_));
  OAI210     u360(.A0(men_men_n382_), .A1(men_men_n375_), .B0(men_men_n381_), .Y(men_men_n383_));
  NO3        u361(.A(men_men_n82_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n384_));
  NO2        u362(.A(i_11_), .B(i_12_), .Y(men_men_n385_));
  NA2        u363(.A(men_men_n377_), .B(men_men_n233_), .Y(men_men_n386_));
  NA2        u364(.A(men_men_n109_), .B(men_men_n42_), .Y(men_men_n387_));
  NO2        u365(.A(men_men_n387_), .B(men_men_n217_), .Y(men_men_n388_));
  NAi21      u366(.An(i_13_), .B(i_0_), .Y(men_men_n389_));
  NO2        u367(.A(men_men_n389_), .B(men_men_n235_), .Y(men_men_n390_));
  NA2        u368(.A(men_men_n388_), .B(men_men_n390_), .Y(men_men_n391_));
  NA3        u369(.A(men_men_n391_), .B(men_men_n383_), .C(men_men_n380_), .Y(men_men_n392_));
  NO3        u370(.A(i_1_), .B(i_12_), .C(men_men_n82_), .Y(men_men_n393_));
  NO2        u371(.A(i_0_), .B(i_11_), .Y(men_men_n394_));
  INV        u372(.A(i_5_), .Y(men_men_n395_));
  AN2        u373(.A(i_1_), .B(i_6_), .Y(men_men_n396_));
  NOi21      u374(.An(i_2_), .B(i_12_), .Y(men_men_n397_));
  NA2        u375(.A(men_men_n397_), .B(men_men_n396_), .Y(men_men_n398_));
  NO2        u376(.A(men_men_n398_), .B(men_men_n395_), .Y(men_men_n399_));
  NA2        u377(.A(men_men_n139_), .B(i_9_), .Y(men_men_n400_));
  NO2        u378(.A(men_men_n400_), .B(i_4_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n399_), .B(men_men_n401_), .Y(men_men_n402_));
  NAi21      u380(.An(i_9_), .B(i_4_), .Y(men_men_n403_));
  OR2        u381(.A(i_13_), .B(i_10_), .Y(men_men_n404_));
  NO3        u382(.A(men_men_n404_), .B(men_men_n114_), .C(men_men_n403_), .Y(men_men_n405_));
  NO2        u383(.A(men_men_n169_), .B(men_men_n120_), .Y(men_men_n406_));
  BUFFER     u384(.A(men_men_n212_), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n97_), .B(men_men_n25_), .Y(men_men_n408_));
  NA2        u386(.A(men_men_n271_), .B(men_men_n408_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n264_), .B(men_men_n206_), .Y(men_men_n410_));
  OAI220     u388(.A0(men_men_n410_), .A1(men_men_n407_), .B0(men_men_n409_), .B1(men_men_n330_), .Y(men_men_n411_));
  INV        u389(.A(men_men_n411_), .Y(men_men_n412_));
  AOI210     u390(.A0(men_men_n412_), .A1(men_men_n402_), .B0(men_men_n26_), .Y(men_men_n413_));
  NA2        u391(.A(men_men_n307_), .B(men_men_n306_), .Y(men_men_n414_));
  AOI220     u392(.A0(men_men_n283_), .A1(men_men_n274_), .B0(men_men_n277_), .B1(i_6_), .Y(men_men_n415_));
  NO2        u393(.A(men_men_n415_), .B(men_men_n166_), .Y(men_men_n416_));
  NO2        u394(.A(men_men_n179_), .B(men_men_n82_), .Y(men_men_n417_));
  AOI220     u395(.A0(men_men_n417_), .A1(men_men_n282_), .B0(men_men_n266_), .B1(men_men_n206_), .Y(men_men_n418_));
  NO2        u396(.A(men_men_n418_), .B(men_men_n273_), .Y(men_men_n419_));
  NO3        u397(.A(men_men_n419_), .B(men_men_n416_), .C(men_men_n414_), .Y(men_men_n420_));
  NA2        u398(.A(men_men_n191_), .B(men_men_n92_), .Y(men_men_n421_));
  NA3        u399(.A(men_men_n310_), .B(men_men_n160_), .C(men_men_n82_), .Y(men_men_n422_));
  AOI210     u400(.A0(men_men_n422_), .A1(men_men_n421_), .B0(men_men_n308_), .Y(men_men_n423_));
  NA2        u401(.A(men_men_n283_), .B(men_men_n232_), .Y(men_men_n424_));
  NO2        u402(.A(men_men_n424_), .B(men_men_n179_), .Y(men_men_n425_));
  NA3        u403(.A(men_men_n321_), .B(men_men_n320_), .C(i_5_), .Y(men_men_n426_));
  INV        u404(.A(men_men_n301_), .Y(men_men_n427_));
  OAI210     u405(.A0(men_men_n427_), .A1(men_men_n185_), .B0(men_men_n426_), .Y(men_men_n428_));
  NO3        u406(.A(men_men_n428_), .B(men_men_n425_), .C(men_men_n423_), .Y(men_men_n429_));
  AOI210     u407(.A0(men_men_n429_), .A1(men_men_n420_), .B0(men_men_n260_), .Y(men_men_n430_));
  NO4        u408(.A(men_men_n430_), .B(men_men_n413_), .C(men_men_n392_), .D(men_men_n368_), .Y(men_men_n431_));
  NO2        u409(.A(men_men_n64_), .B(i_4_), .Y(men_men_n432_));
  NO2        u410(.A(men_men_n70_), .B(i_13_), .Y(men_men_n433_));
  NO2        u411(.A(i_10_), .B(i_9_), .Y(men_men_n434_));
  NAi21      u412(.An(i_12_), .B(i_8_), .Y(men_men_n435_));
  NA2        u413(.A(men_men_n296_), .B(i_0_), .Y(men_men_n436_));
  NO3        u414(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n437_));
  NA2        u415(.A(men_men_n255_), .B(men_men_n93_), .Y(men_men_n438_));
  NA2        u416(.A(i_8_), .B(i_9_), .Y(men_men_n439_));
  NA2        u417(.A(men_men_n244_), .B(men_men_n295_), .Y(men_men_n440_));
  NO3        u418(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n441_));
  INV        u419(.A(men_men_n441_), .Y(men_men_n442_));
  NA3        u420(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n443_));
  NA4        u421(.A(men_men_n142_), .B(men_men_n112_), .C(men_men_n77_), .D(men_men_n23_), .Y(men_men_n444_));
  OAI220     u422(.A0(men_men_n444_), .A1(men_men_n443_), .B0(men_men_n442_), .B1(men_men_n440_), .Y(men_men_n445_));
  INV        u423(.A(men_men_n445_), .Y(men_men_n446_));
  OA210      u424(.A0(men_men_n340_), .A1(men_men_n97_), .B0(men_men_n284_), .Y(men_men_n447_));
  OA220      u425(.A0(men_men_n447_), .A1(men_men_n159_), .B0(men_men_n202_), .B1(men_men_n229_), .Y(men_men_n448_));
  NA2        u426(.A(men_men_n92_), .B(i_13_), .Y(men_men_n449_));
  NA2        u427(.A(men_men_n417_), .B(men_men_n369_), .Y(men_men_n450_));
  NO2        u428(.A(i_2_), .B(i_13_), .Y(men_men_n451_));
  NO2        u429(.A(men_men_n450_), .B(men_men_n449_), .Y(men_men_n452_));
  NO3        u430(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n453_));
  NO2        u431(.A(i_6_), .B(i_7_), .Y(men_men_n454_));
  NA2        u432(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  NO2        u433(.A(i_11_), .B(i_1_), .Y(men_men_n456_));
  NOi21      u434(.An(i_2_), .B(i_7_), .Y(men_men_n457_));
  NAi31      u435(.An(i_11_), .B(men_men_n457_), .C(men_men_n993_), .Y(men_men_n458_));
  INV        u436(.A(men_men_n404_), .Y(men_men_n459_));
  NA3        u437(.A(men_men_n459_), .B(men_men_n432_), .C(men_men_n72_), .Y(men_men_n460_));
  NO2        u438(.A(men_men_n460_), .B(men_men_n458_), .Y(men_men_n461_));
  NO2        u439(.A(i_6_), .B(i_10_), .Y(men_men_n462_));
  NA4        u440(.A(men_men_n462_), .B(men_men_n300_), .C(i_8_), .D(men_men_n233_), .Y(men_men_n463_));
  NO2        u441(.A(men_men_n463_), .B(men_men_n152_), .Y(men_men_n464_));
  NA3        u442(.A(men_men_n240_), .B(men_men_n168_), .C(men_men_n129_), .Y(men_men_n465_));
  NA2        u443(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n466_));
  NO2        u444(.A(men_men_n154_), .B(i_3_), .Y(men_men_n467_));
  NAi31      u445(.An(men_men_n466_), .B(men_men_n467_), .C(men_men_n223_), .Y(men_men_n468_));
  NA3        u446(.A(men_men_n381_), .B(men_men_n175_), .C(men_men_n146_), .Y(men_men_n469_));
  NA3        u447(.A(men_men_n469_), .B(men_men_n468_), .C(men_men_n465_), .Y(men_men_n470_));
  NO4        u448(.A(men_men_n470_), .B(men_men_n464_), .C(men_men_n461_), .D(men_men_n452_), .Y(men_men_n471_));
  NA2        u449(.A(men_men_n441_), .B(men_men_n377_), .Y(men_men_n472_));
  NO2        u450(.A(men_men_n472_), .B(men_men_n221_), .Y(men_men_n473_));
  NAi21      u451(.An(men_men_n212_), .B(men_men_n385_), .Y(men_men_n474_));
  NA3        u452(.A(men_men_n992_), .B(i_3_), .C(men_men_n139_), .Y(men_men_n475_));
  OR3        u453(.A(men_men_n290_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n476_));
  NO2        u454(.A(men_men_n476_), .B(men_men_n475_), .Y(men_men_n477_));
  NA2        u455(.A(men_men_n27_), .B(i_10_), .Y(men_men_n478_));
  NO2        u456(.A(men_men_n478_), .B(men_men_n449_), .Y(men_men_n479_));
  NA3        u457(.A(men_men_n293_), .B(men_men_n220_), .C(men_men_n70_), .Y(men_men_n480_));
  NO2        u458(.A(men_men_n480_), .B(men_men_n455_), .Y(men_men_n481_));
  NO4        u459(.A(men_men_n481_), .B(men_men_n479_), .C(men_men_n477_), .D(men_men_n473_), .Y(men_men_n482_));
  NA4        u460(.A(men_men_n482_), .B(men_men_n471_), .C(men_men_n448_), .D(men_men_n446_), .Y(men_men_n483_));
  AN2        u461(.A(men_men_n274_), .B(men_men_n231_), .Y(men_men_n484_));
  NA2        u462(.A(men_men_n484_), .B(men_men_n172_), .Y(men_men_n485_));
  NA2        u463(.A(men_men_n119_), .B(men_men_n108_), .Y(men_men_n486_));
  AN2        u464(.A(men_men_n486_), .B(men_men_n437_), .Y(men_men_n487_));
  OAI210     u465(.A0(i_2_), .A1(men_men_n229_), .B0(men_men_n294_), .Y(men_men_n488_));
  AOI220     u466(.A0(men_men_n488_), .A1(men_men_n309_), .B0(men_men_n487_), .B1(men_men_n296_), .Y(men_men_n489_));
  NA2        u467(.A(men_men_n344_), .B(men_men_n70_), .Y(men_men_n490_));
  NA2        u468(.A(men_men_n357_), .B(men_men_n353_), .Y(men_men_n491_));
  NO2        u469(.A(men_men_n36_), .B(i_8_), .Y(men_men_n492_));
  NAi41      u470(.An(men_men_n490_), .B(men_men_n462_), .C(men_men_n492_), .D(men_men_n47_), .Y(men_men_n493_));
  AOI210     u471(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n405_), .Y(men_men_n494_));
  NA2        u472(.A(men_men_n494_), .B(men_men_n493_), .Y(men_men_n495_));
  INV        u473(.A(men_men_n495_), .Y(men_men_n496_));
  INV        u474(.A(men_men_n248_), .Y(men_men_n497_));
  OAI210     u475(.A0(i_8_), .A1(men_men_n497_), .B0(men_men_n131_), .Y(men_men_n498_));
  NO2        u476(.A(i_7_), .B(men_men_n194_), .Y(men_men_n499_));
  OR2        u477(.A(men_men_n179_), .B(i_4_), .Y(men_men_n500_));
  INV        u478(.A(men_men_n500_), .Y(men_men_n501_));
  AOI220     u479(.A0(men_men_n501_), .A1(men_men_n499_), .B0(men_men_n498_), .B1(men_men_n406_), .Y(men_men_n502_));
  NA4        u480(.A(men_men_n502_), .B(men_men_n496_), .C(men_men_n489_), .D(men_men_n485_), .Y(men_men_n503_));
  NA2        u481(.A(men_men_n376_), .B(men_men_n282_), .Y(men_men_n504_));
  NA2        u482(.A(men_men_n372_), .B(men_men_n504_), .Y(men_men_n505_));
  NO2        u483(.A(i_12_), .B(men_men_n189_), .Y(men_men_n506_));
  NA2        u484(.A(men_men_n506_), .B(men_men_n222_), .Y(men_men_n507_));
  NA2        u485(.A(men_men_n462_), .B(men_men_n27_), .Y(men_men_n508_));
  NO2        u486(.A(men_men_n508_), .B(men_men_n507_), .Y(men_men_n509_));
  NOi31      u487(.An(men_men_n301_), .B(men_men_n404_), .C(men_men_n38_), .Y(men_men_n510_));
  OAI210     u488(.A0(men_men_n510_), .A1(men_men_n509_), .B0(men_men_n505_), .Y(men_men_n511_));
  NO2        u489(.A(i_8_), .B(i_7_), .Y(men_men_n512_));
  INV        u490(.A(men_men_n220_), .Y(men_men_n513_));
  OAI220     u491(.A0(men_men_n47_), .A1(men_men_n500_), .B0(men_men_n513_), .B1(men_men_n237_), .Y(men_men_n514_));
  NA2        u492(.A(men_men_n45_), .B(i_10_), .Y(men_men_n515_));
  NO2        u493(.A(men_men_n515_), .B(i_6_), .Y(men_men_n516_));
  NA3        u494(.A(men_men_n516_), .B(men_men_n514_), .C(men_men_n512_), .Y(men_men_n517_));
  AOI210     u495(.A0(men_men_n417_), .A1(men_men_n310_), .B0(men_men_n242_), .Y(men_men_n518_));
  NO2        u496(.A(men_men_n518_), .B(men_men_n251_), .Y(men_men_n519_));
  NA2        u497(.A(men_men_n519_), .B(men_men_n254_), .Y(men_men_n520_));
  NOi31      u498(.An(men_men_n277_), .B(men_men_n288_), .C(men_men_n177_), .Y(men_men_n521_));
  NA3        u499(.A(men_men_n293_), .B(men_men_n170_), .C(men_men_n92_), .Y(men_men_n522_));
  NO2        u500(.A(men_men_n218_), .B(men_men_n45_), .Y(men_men_n523_));
  NO2        u501(.A(men_men_n154_), .B(i_5_), .Y(men_men_n524_));
  NA2        u502(.A(men_men_n524_), .B(men_men_n303_), .Y(men_men_n525_));
  OAI210     u503(.A0(men_men_n525_), .A1(men_men_n523_), .B0(men_men_n522_), .Y(men_men_n526_));
  OAI210     u504(.A0(men_men_n526_), .A1(men_men_n521_), .B0(men_men_n441_), .Y(men_men_n527_));
  NA4        u505(.A(men_men_n527_), .B(men_men_n520_), .C(men_men_n517_), .D(men_men_n511_), .Y(men_men_n528_));
  NA3        u506(.A(men_men_n214_), .B(men_men_n68_), .C(men_men_n45_), .Y(men_men_n529_));
  NA2        u507(.A(men_men_n271_), .B(men_men_n80_), .Y(men_men_n530_));
  AOI210     u508(.A0(men_men_n529_), .A1(men_men_n335_), .B0(men_men_n530_), .Y(men_men_n531_));
  NA2        u509(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n532_));
  NA2        u510(.A(men_men_n434_), .B(men_men_n218_), .Y(men_men_n533_));
  NO2        u511(.A(men_men_n532_), .B(men_men_n533_), .Y(men_men_n534_));
  NA2        u512(.A(i_0_), .B(men_men_n49_), .Y(men_men_n535_));
  NA3        u513(.A(men_men_n506_), .B(men_men_n262_), .C(men_men_n535_), .Y(men_men_n536_));
  NO2        u514(.A(i_1_), .B(men_men_n536_), .Y(men_men_n537_));
  NO3        u515(.A(men_men_n537_), .B(men_men_n534_), .C(men_men_n531_), .Y(men_men_n538_));
  NO4        u516(.A(i_1_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n539_));
  NO3        u517(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n540_));
  NO2        u518(.A(men_men_n230_), .B(men_men_n36_), .Y(men_men_n541_));
  AN2        u519(.A(men_men_n541_), .B(men_men_n540_), .Y(men_men_n542_));
  OA210      u520(.A0(men_men_n542_), .A1(men_men_n539_), .B0(men_men_n344_), .Y(men_men_n543_));
  NO2        u521(.A(men_men_n404_), .B(i_1_), .Y(men_men_n544_));
  NOi31      u522(.An(men_men_n544_), .B(men_men_n438_), .C(men_men_n70_), .Y(men_men_n545_));
  AN3        u523(.A(men_men_n545_), .B(men_men_n401_), .C(i_3_), .Y(men_men_n546_));
  NO2        u524(.A(men_men_n415_), .B(men_men_n173_), .Y(men_men_n547_));
  NO3        u525(.A(men_men_n547_), .B(men_men_n546_), .C(men_men_n543_), .Y(men_men_n548_));
  NOi21      u526(.An(i_10_), .B(i_6_), .Y(men_men_n549_));
  NO2        u527(.A(men_men_n82_), .B(men_men_n25_), .Y(men_men_n550_));
  AOI220     u528(.A0(men_men_n271_), .A1(men_men_n550_), .B0(men_men_n262_), .B1(men_men_n549_), .Y(men_men_n551_));
  NO2        u529(.A(men_men_n551_), .B(men_men_n436_), .Y(men_men_n552_));
  NO2        u530(.A(men_men_n111_), .B(men_men_n23_), .Y(men_men_n553_));
  NA2        u531(.A(men_men_n301_), .B(men_men_n161_), .Y(men_men_n554_));
  AOI220     u532(.A0(men_men_n554_), .A1(men_men_n424_), .B0(men_men_n169_), .B1(men_men_n178_), .Y(men_men_n555_));
  NO2        u533(.A(men_men_n555_), .B(men_men_n552_), .Y(men_men_n556_));
  NO2        u534(.A(men_men_n490_), .B(men_men_n365_), .Y(men_men_n557_));
  INV        u535(.A(men_men_n303_), .Y(men_men_n558_));
  NO2        u536(.A(i_12_), .B(men_men_n82_), .Y(men_men_n559_));
  NA3        u537(.A(men_men_n559_), .B(men_men_n262_), .C(men_men_n535_), .Y(men_men_n560_));
  NA3        u538(.A(men_men_n373_), .B(men_men_n271_), .C(men_men_n214_), .Y(men_men_n561_));
  AOI210     u539(.A0(men_men_n561_), .A1(men_men_n560_), .B0(men_men_n558_), .Y(men_men_n562_));
  NO3        u540(.A(i_4_), .B(men_men_n327_), .C(men_men_n288_), .Y(men_men_n563_));
  OR2        u541(.A(i_2_), .B(i_5_), .Y(men_men_n564_));
  OR2        u542(.A(men_men_n564_), .B(men_men_n396_), .Y(men_men_n565_));
  NO2        u543(.A(men_men_n565_), .B(men_men_n474_), .Y(men_men_n566_));
  NO4        u544(.A(men_men_n566_), .B(men_men_n563_), .C(men_men_n562_), .D(men_men_n557_), .Y(men_men_n567_));
  NA4        u545(.A(men_men_n567_), .B(men_men_n556_), .C(men_men_n548_), .D(men_men_n538_), .Y(men_men_n568_));
  NO4        u546(.A(men_men_n568_), .B(men_men_n528_), .C(men_men_n503_), .D(men_men_n483_), .Y(men_men_n569_));
  NA4        u547(.A(men_men_n569_), .B(men_men_n431_), .C(men_men_n343_), .D(men_men_n299_), .Y(men7));
  NO2        u548(.A(men_men_n88_), .B(men_men_n55_), .Y(men_men_n571_));
  NO2        u549(.A(men_men_n104_), .B(men_men_n85_), .Y(men_men_n572_));
  NA2        u550(.A(men_men_n462_), .B(men_men_n80_), .Y(men_men_n573_));
  NA2        u551(.A(i_11_), .B(men_men_n189_), .Y(men_men_n574_));
  NA3        u552(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n575_));
  NO2        u553(.A(men_men_n233_), .B(i_4_), .Y(men_men_n576_));
  NA2        u554(.A(men_men_n576_), .B(i_8_), .Y(men_men_n577_));
  NO2        u555(.A(men_men_n101_), .B(men_men_n575_), .Y(men_men_n578_));
  NA2        u556(.A(i_2_), .B(men_men_n82_), .Y(men_men_n579_));
  OAI210     u557(.A0(men_men_n83_), .A1(men_men_n198_), .B0(men_men_n199_), .Y(men_men_n580_));
  NA2        u558(.A(i_4_), .B(i_8_), .Y(men_men_n581_));
  OAI220     u559(.A0(men_men_n991_), .A1(men_men_n579_), .B0(men_men_n580_), .B1(i_13_), .Y(men_men_n582_));
  NO4        u560(.A(men_men_n582_), .B(men_men_n578_), .C(men_men_n572_), .D(men_men_n571_), .Y(men_men_n583_));
  INV        u561(.A(men_men_n158_), .Y(men_men_n584_));
  OR2        u562(.A(i_6_), .B(i_10_), .Y(men_men_n585_));
  NO2        u563(.A(men_men_n585_), .B(men_men_n23_), .Y(men_men_n586_));
  OR3        u564(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n587_));
  NO3        u565(.A(men_men_n587_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n588_));
  INV        u566(.A(men_men_n195_), .Y(men_men_n589_));
  NO2        u567(.A(men_men_n588_), .B(men_men_n586_), .Y(men_men_n590_));
  OA220      u568(.A0(men_men_n590_), .A1(men_men_n558_), .B0(men_men_n584_), .B1(men_men_n256_), .Y(men_men_n591_));
  AOI210     u569(.A0(men_men_n591_), .A1(men_men_n583_), .B0(men_men_n64_), .Y(men_men_n592_));
  NOi21      u570(.An(i_11_), .B(i_7_), .Y(men_men_n593_));
  AO210      u571(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n594_));
  NO2        u572(.A(men_men_n594_), .B(men_men_n593_), .Y(men_men_n595_));
  NA2        u573(.A(men_men_n595_), .B(men_men_n201_), .Y(men_men_n596_));
  NA3        u574(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n597_));
  NAi31      u575(.An(men_men_n597_), .B(men_men_n211_), .C(i_11_), .Y(men_men_n598_));
  AOI210     u576(.A0(men_men_n598_), .A1(men_men_n596_), .B0(men_men_n64_), .Y(men_men_n599_));
  NA2        u577(.A(men_men_n223_), .B(men_men_n64_), .Y(men_men_n600_));
  NA2        u578(.A(men_men_n397_), .B(men_men_n31_), .Y(men_men_n601_));
  OR2        u579(.A(men_men_n203_), .B(men_men_n104_), .Y(men_men_n602_));
  NA2        u580(.A(men_men_n602_), .B(men_men_n601_), .Y(men_men_n603_));
  NO2        u581(.A(men_men_n64_), .B(i_9_), .Y(men_men_n604_));
  NA2        u582(.A(men_men_n64_), .B(men_men_n603_), .Y(men_men_n605_));
  NO2        u583(.A(i_1_), .B(i_12_), .Y(men_men_n606_));
  NA2        u584(.A(men_men_n605_), .B(men_men_n600_), .Y(men_men_n607_));
  OAI210     u585(.A0(men_men_n607_), .A1(men_men_n599_), .B0(i_6_), .Y(men_men_n608_));
  NO2        u586(.A(men_men_n233_), .B(men_men_n82_), .Y(men_men_n609_));
  NO2        u587(.A(men_men_n609_), .B(i_11_), .Y(men_men_n610_));
  NO4        u588(.A(men_men_n211_), .B(men_men_n125_), .C(i_13_), .D(men_men_n82_), .Y(men_men_n611_));
  NA2        u589(.A(men_men_n611_), .B(men_men_n604_), .Y(men_men_n612_));
  NA2        u590(.A(men_men_n233_), .B(i_6_), .Y(men_men_n613_));
  NO3        u591(.A(men_men_n585_), .B(men_men_n230_), .C(men_men_n23_), .Y(men_men_n614_));
  INV        u592(.A(men_men_n614_), .Y(men_men_n615_));
  OAI210     u593(.A0(men_men_n615_), .A1(men_men_n45_), .B0(men_men_n612_), .Y(men_men_n616_));
  NA3        u594(.A(men_men_n512_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n617_));
  NA2        u595(.A(men_men_n135_), .B(i_9_), .Y(men_men_n618_));
  NA3        u596(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n619_));
  NO2        u597(.A(men_men_n47_), .B(i_1_), .Y(men_men_n620_));
  NA3        u598(.A(men_men_n620_), .B(men_men_n255_), .C(men_men_n45_), .Y(men_men_n621_));
  OAI220     u599(.A0(men_men_n621_), .A1(men_men_n619_), .B0(men_men_n618_), .B1(men_men_n987_), .Y(men_men_n622_));
  NA3        u600(.A(men_men_n604_), .B(men_men_n303_), .C(i_6_), .Y(men_men_n623_));
  NO2        u601(.A(men_men_n623_), .B(men_men_n23_), .Y(men_men_n624_));
  AOI210     u602(.A0(men_men_n456_), .A1(men_men_n408_), .B0(men_men_n236_), .Y(men_men_n625_));
  NO2        u603(.A(men_men_n625_), .B(men_men_n579_), .Y(men_men_n626_));
  NA2        u604(.A(men_men_n620_), .B(men_men_n255_), .Y(men_men_n627_));
  NO2        u605(.A(i_11_), .B(men_men_n37_), .Y(men_men_n628_));
  NA2        u606(.A(men_men_n628_), .B(men_men_n24_), .Y(men_men_n629_));
  NO2        u607(.A(men_men_n629_), .B(men_men_n627_), .Y(men_men_n630_));
  OR4        u608(.A(men_men_n630_), .B(men_men_n626_), .C(men_men_n624_), .D(men_men_n622_), .Y(men_men_n631_));
  NO2        u609(.A(men_men_n631_), .B(men_men_n616_), .Y(men_men_n632_));
  NO2        u610(.A(men_men_n233_), .B(men_men_n97_), .Y(men_men_n633_));
  NO2        u611(.A(men_men_n633_), .B(men_men_n593_), .Y(men_men_n634_));
  NA2        u612(.A(men_men_n634_), .B(i_1_), .Y(men_men_n635_));
  NO2        u613(.A(men_men_n635_), .B(men_men_n587_), .Y(men_men_n636_));
  NO2        u614(.A(men_men_n403_), .B(men_men_n82_), .Y(men_men_n637_));
  NA2        u615(.A(men_men_n636_), .B(men_men_n47_), .Y(men_men_n638_));
  NO2        u616(.A(men_men_n114_), .B(men_men_n37_), .Y(men_men_n639_));
  NO2        u617(.A(men_men_n82_), .B(i_9_), .Y(men_men_n640_));
  NO2        u618(.A(men_men_n640_), .B(men_men_n64_), .Y(men_men_n641_));
  NA2        u619(.A(i_1_), .B(i_3_), .Y(men_men_n642_));
  NA3        u620(.A(men_men_n638_), .B(men_men_n632_), .C(men_men_n608_), .Y(men_men_n643_));
  NO3        u621(.A(i_11_), .B(i_3_), .C(i_7_), .Y(men_men_n644_));
  NOi21      u622(.An(men_men_n644_), .B(i_10_), .Y(men_men_n645_));
  OA210      u623(.A0(men_men_n645_), .A1(men_men_n240_), .B0(men_men_n82_), .Y(men_men_n646_));
  NO3        u624(.A(men_men_n457_), .B(men_men_n581_), .C(men_men_n82_), .Y(men_men_n647_));
  NA2        u625(.A(men_men_n647_), .B(men_men_n25_), .Y(men_men_n648_));
  INV        u626(.A(men_men_n648_), .Y(men_men_n649_));
  OAI210     u627(.A0(men_men_n649_), .A1(men_men_n646_), .B0(i_1_), .Y(men_men_n650_));
  AOI210     u628(.A0(men_men_n255_), .A1(men_men_n93_), .B0(i_1_), .Y(men_men_n651_));
  NO2        u629(.A(men_men_n355_), .B(i_2_), .Y(men_men_n652_));
  NA2        u630(.A(men_men_n652_), .B(men_men_n651_), .Y(men_men_n653_));
  OAI210     u631(.A0(men_men_n623_), .A1(men_men_n435_), .B0(men_men_n653_), .Y(men_men_n654_));
  INV        u632(.A(men_men_n654_), .Y(men_men_n655_));
  AOI210     u633(.A0(men_men_n655_), .A1(men_men_n650_), .B0(i_13_), .Y(men_men_n656_));
  OR2        u634(.A(i_11_), .B(i_7_), .Y(men_men_n657_));
  NA3        u635(.A(men_men_n657_), .B(men_men_n102_), .C(men_men_n135_), .Y(men_men_n658_));
  AOI220     u636(.A0(men_men_n451_), .A1(men_men_n158_), .B0(i_2_), .B1(men_men_n135_), .Y(men_men_n659_));
  OAI210     u637(.A0(men_men_n659_), .A1(men_men_n45_), .B0(men_men_n658_), .Y(men_men_n660_));
  NO2        u638(.A(men_men_n457_), .B(men_men_n24_), .Y(men_men_n661_));
  AOI220     u639(.A0(men_men_n661_), .A1(men_men_n637_), .B0(men_men_n240_), .B1(men_men_n128_), .Y(men_men_n662_));
  NO2        u640(.A(men_men_n662_), .B(men_men_n41_), .Y(men_men_n663_));
  AOI210     u641(.A0(men_men_n660_), .A1(men_men_n318_), .B0(men_men_n663_), .Y(men_men_n664_));
  AOI210     u642(.A0(men_men_n435_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n665_));
  NOi31      u643(.An(men_men_n665_), .B(men_men_n573_), .C(men_men_n45_), .Y(men_men_n666_));
  NA2        u644(.A(men_men_n124_), .B(i_13_), .Y(men_men_n667_));
  NO2        u645(.A(men_men_n619_), .B(men_men_n111_), .Y(men_men_n668_));
  INV        u646(.A(men_men_n668_), .Y(men_men_n669_));
  OAI220     u647(.A0(men_men_n669_), .A1(men_men_n68_), .B0(men_men_n667_), .B1(men_men_n651_), .Y(men_men_n670_));
  NO3        u648(.A(men_men_n68_), .B(men_men_n32_), .C(men_men_n97_), .Y(men_men_n671_));
  NA2        u649(.A(men_men_n26_), .B(men_men_n189_), .Y(men_men_n672_));
  NA2        u650(.A(men_men_n672_), .B(i_7_), .Y(men_men_n673_));
  NO3        u651(.A(men_men_n457_), .B(men_men_n233_), .C(men_men_n82_), .Y(men_men_n674_));
  AOI210     u652(.A0(men_men_n674_), .A1(men_men_n673_), .B0(men_men_n671_), .Y(men_men_n675_));
  AOI220     u653(.A0(men_men_n373_), .A1(men_men_n620_), .B0(men_men_n87_), .B1(men_men_n98_), .Y(men_men_n676_));
  OAI220     u654(.A0(men_men_n676_), .A1(men_men_n577_), .B0(men_men_n675_), .B1(men_men_n589_), .Y(men_men_n677_));
  NO3        u655(.A(men_men_n677_), .B(men_men_n670_), .C(men_men_n666_), .Y(men_men_n678_));
  OR2        u656(.A(i_11_), .B(i_6_), .Y(men_men_n679_));
  NA3        u657(.A(men_men_n576_), .B(men_men_n672_), .C(i_7_), .Y(men_men_n680_));
  AOI210     u658(.A0(men_men_n680_), .A1(men_men_n669_), .B0(men_men_n679_), .Y(men_men_n681_));
  NA2        u659(.A(men_men_n610_), .B(i_13_), .Y(men_men_n682_));
  NAi21      u660(.An(i_11_), .B(i_12_), .Y(men_men_n683_));
  NO2        u661(.A(men_men_n559_), .B(men_men_n581_), .Y(men_men_n684_));
  NA2        u662(.A(men_men_n684_), .B(men_men_n300_), .Y(men_men_n685_));
  NA2        u663(.A(men_men_n685_), .B(men_men_n682_), .Y(men_men_n686_));
  OAI210     u664(.A0(men_men_n686_), .A1(men_men_n681_), .B0(men_men_n64_), .Y(men_men_n687_));
  NO2        u665(.A(i_2_), .B(i_12_), .Y(men_men_n688_));
  NA2        u666(.A(men_men_n354_), .B(men_men_n688_), .Y(men_men_n689_));
  NO2        u667(.A(men_men_n125_), .B(i_2_), .Y(men_men_n690_));
  NA2        u668(.A(men_men_n690_), .B(men_men_n606_), .Y(men_men_n691_));
  NA2        u669(.A(men_men_n691_), .B(men_men_n689_), .Y(men_men_n692_));
  NA3        u670(.A(men_men_n692_), .B(men_men_n46_), .C(men_men_n222_), .Y(men_men_n693_));
  NA4        u671(.A(men_men_n693_), .B(men_men_n687_), .C(men_men_n678_), .D(men_men_n664_), .Y(men_men_n694_));
  OR4        u672(.A(men_men_n694_), .B(men_men_n656_), .C(men_men_n643_), .D(men_men_n592_), .Y(men5));
  AOI210     u673(.A0(men_men_n634_), .A1(men_men_n258_), .B0(men_men_n406_), .Y(men_men_n696_));
  AN2        u674(.A(men_men_n24_), .B(i_10_), .Y(men_men_n697_));
  NA3        u675(.A(men_men_n697_), .B(men_men_n688_), .C(men_men_n104_), .Y(men_men_n698_));
  NO2        u676(.A(men_men_n577_), .B(i_11_), .Y(men_men_n699_));
  NA2        u677(.A(men_men_n83_), .B(men_men_n699_), .Y(men_men_n700_));
  NA3        u678(.A(men_men_n700_), .B(men_men_n698_), .C(men_men_n696_), .Y(men_men_n701_));
  NO3        u679(.A(i_11_), .B(men_men_n233_), .C(i_13_), .Y(men_men_n702_));
  NO2        u680(.A(men_men_n121_), .B(men_men_n23_), .Y(men_men_n703_));
  NA2        u681(.A(i_12_), .B(i_8_), .Y(men_men_n704_));
  OAI210     u682(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n704_), .Y(men_men_n705_));
  INV        u683(.A(men_men_n434_), .Y(men_men_n706_));
  AOI220     u684(.A0(men_men_n303_), .A1(men_men_n553_), .B0(men_men_n705_), .B1(men_men_n703_), .Y(men_men_n707_));
  INV        u685(.A(men_men_n707_), .Y(men_men_n708_));
  NO2        u686(.A(men_men_n708_), .B(men_men_n701_), .Y(men_men_n709_));
  INV        u687(.A(men_men_n168_), .Y(men_men_n710_));
  NA2        u688(.A(men_men_n652_), .B(men_men_n107_), .Y(men_men_n711_));
  NO2        u689(.A(men_men_n711_), .B(men_men_n710_), .Y(men_men_n712_));
  NO2        u690(.A(men_men_n439_), .B(men_men_n26_), .Y(men_men_n713_));
  NO2        u691(.A(men_men_n713_), .B(men_men_n408_), .Y(men_men_n714_));
  NA2        u692(.A(men_men_n714_), .B(i_2_), .Y(men_men_n715_));
  INV        u693(.A(men_men_n715_), .Y(men_men_n716_));
  AOI210     u694(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n404_), .Y(men_men_n717_));
  AOI210     u695(.A0(men_men_n717_), .A1(men_men_n716_), .B0(men_men_n712_), .Y(men_men_n718_));
  NO2        u696(.A(men_men_n186_), .B(men_men_n122_), .Y(men_men_n719_));
  OAI210     u697(.A0(men_men_n719_), .A1(men_men_n703_), .B0(i_2_), .Y(men_men_n720_));
  NO3        u698(.A(men_men_n594_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n721_));
  AOI210     u699(.A0(men_men_n990_), .A1(men_men_n720_), .B0(men_men_n189_), .Y(men_men_n722_));
  OA210      u700(.A0(men_men_n595_), .A1(men_men_n123_), .B0(i_13_), .Y(men_men_n723_));
  NA2        u701(.A(men_men_n149_), .B(men_men_n574_), .Y(men_men_n724_));
  NO2        u702(.A(men_men_n724_), .B(men_men_n359_), .Y(men_men_n725_));
  AOI210     u703(.A0(men_men_n203_), .A1(men_men_n145_), .B0(men_men_n492_), .Y(men_men_n726_));
  NA2        u704(.A(men_men_n726_), .B(men_men_n408_), .Y(men_men_n727_));
  NO2        u705(.A(men_men_n98_), .B(men_men_n45_), .Y(men_men_n728_));
  INV        u706(.A(men_men_n289_), .Y(men_men_n729_));
  NA4        u707(.A(men_men_n729_), .B(men_men_n293_), .C(men_men_n121_), .D(men_men_n43_), .Y(men_men_n730_));
  OAI210     u708(.A0(men_men_n730_), .A1(men_men_n728_), .B0(men_men_n727_), .Y(men_men_n731_));
  NO4        u709(.A(men_men_n731_), .B(men_men_n725_), .C(men_men_n723_), .D(men_men_n722_), .Y(men_men_n732_));
  NA2        u710(.A(men_men_n553_), .B(men_men_n28_), .Y(men_men_n733_));
  NA2        u711(.A(men_men_n702_), .B(men_men_n263_), .Y(men_men_n734_));
  NA2        u712(.A(men_men_n734_), .B(men_men_n733_), .Y(men_men_n735_));
  NO2        u713(.A(men_men_n63_), .B(i_12_), .Y(men_men_n736_));
  NO2        u714(.A(men_men_n736_), .B(men_men_n123_), .Y(men_men_n737_));
  NO2        u715(.A(men_men_n737_), .B(men_men_n574_), .Y(men_men_n738_));
  AOI220     u716(.A0(men_men_n738_), .A1(men_men_n36_), .B0(men_men_n735_), .B1(men_men_n47_), .Y(men_men_n739_));
  NA4        u717(.A(men_men_n739_), .B(men_men_n732_), .C(men_men_n718_), .D(men_men_n709_), .Y(men6));
  NO3        u718(.A(men_men_n246_), .B(men_men_n295_), .C(i_1_), .Y(men_men_n741_));
  NO2        u719(.A(men_men_n181_), .B(men_men_n136_), .Y(men_men_n742_));
  OAI210     u720(.A0(men_men_n742_), .A1(men_men_n741_), .B0(men_men_n690_), .Y(men_men_n743_));
  NO2        u721(.A(men_men_n217_), .B(men_men_n466_), .Y(men_men_n744_));
  AO210      u722(.A0(men_men_n988_), .A1(men_men_n743_), .B0(i_12_), .Y(men_men_n745_));
  NA2        u723(.A(men_men_n645_), .B(men_men_n70_), .Y(men_men_n746_));
  INV        u724(.A(men_men_n314_), .Y(men_men_n747_));
  NA2        u725(.A(men_men_n72_), .B(men_men_n128_), .Y(men_men_n748_));
  INV        u726(.A(men_men_n121_), .Y(men_men_n749_));
  NA2        u727(.A(men_men_n749_), .B(men_men_n47_), .Y(men_men_n750_));
  AOI210     u728(.A0(men_men_n750_), .A1(men_men_n748_), .B0(men_men_n747_), .Y(men_men_n751_));
  NO2        u729(.A(men_men_n32_), .B(i_11_), .Y(men_men_n752_));
  NA3        u730(.A(men_men_n752_), .B(men_men_n454_), .C(men_men_n377_), .Y(men_men_n753_));
  NAi32      u731(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n754_));
  NO2        u732(.A(men_men_n679_), .B(men_men_n754_), .Y(men_men_n755_));
  OAI210     u733(.A0(men_men_n644_), .A1(men_men_n541_), .B0(men_men_n540_), .Y(men_men_n756_));
  NAi31      u734(.An(men_men_n755_), .B(men_men_n756_), .C(men_men_n753_), .Y(men_men_n757_));
  OR2        u735(.A(men_men_n757_), .B(men_men_n751_), .Y(men_men_n758_));
  NO2        u736(.A(men_men_n657_), .B(i_2_), .Y(men_men_n759_));
  NA2        u737(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n760_));
  NO2        u738(.A(men_men_n760_), .B(men_men_n396_), .Y(men_men_n761_));
  NA2        u739(.A(men_men_n761_), .B(men_men_n759_), .Y(men_men_n762_));
  AO210      u740(.A0(men_men_n348_), .A1(men_men_n339_), .B0(men_men_n384_), .Y(men_men_n763_));
  NA3        u741(.A(men_men_n763_), .B(men_men_n247_), .C(i_7_), .Y(men_men_n764_));
  BUFFER     u742(.A(men_men_n595_), .Y(men_men_n765_));
  NA2        u743(.A(men_men_n765_), .B(men_men_n144_), .Y(men_men_n766_));
  AO210      u744(.A0(men_men_n472_), .A1(men_men_n706_), .B0(men_men_n36_), .Y(men_men_n767_));
  NA4        u745(.A(men_men_n767_), .B(men_men_n766_), .C(men_men_n764_), .D(men_men_n762_), .Y(men_men_n768_));
  NO2        u746(.A(men_men_n609_), .B(i_11_), .Y(men_men_n769_));
  AOI220     u747(.A0(men_men_n769_), .A1(men_men_n540_), .B0(men_men_n744_), .B1(men_men_n673_), .Y(men_men_n770_));
  NA3        u748(.A(men_men_n359_), .B(men_men_n234_), .C(men_men_n144_), .Y(men_men_n771_));
  NA2        u749(.A(men_men_n384_), .B(men_men_n67_), .Y(men_men_n772_));
  NA4        u750(.A(men_men_n772_), .B(men_men_n771_), .C(men_men_n770_), .D(men_men_n580_), .Y(men_men_n773_));
  NO2        u751(.A(men_men_n585_), .B(men_men_n98_), .Y(men_men_n774_));
  OAI210     u752(.A0(men_men_n774_), .A1(men_men_n108_), .B0(men_men_n394_), .Y(men_men_n775_));
  INV        u753(.A(men_men_n565_), .Y(men_men_n776_));
  NA3        u754(.A(men_men_n776_), .B(men_men_n314_), .C(i_7_), .Y(men_men_n777_));
  NA2        u755(.A(men_men_n777_), .B(men_men_n775_), .Y(men_men_n778_));
  NO4        u756(.A(men_men_n778_), .B(men_men_n773_), .C(men_men_n768_), .D(men_men_n758_), .Y(men_men_n779_));
  NA4        u757(.A(men_men_n779_), .B(men_men_n746_), .C(men_men_n745_), .D(men_men_n367_), .Y(men3));
  NA2        u758(.A(i_6_), .B(i_7_), .Y(men_men_n781_));
  NO2        u759(.A(men_men_n781_), .B(i_0_), .Y(men_men_n782_));
  NO2        u760(.A(i_11_), .B(men_men_n233_), .Y(men_men_n783_));
  OAI210     u761(.A0(men_men_n782_), .A1(men_men_n277_), .B0(men_men_n783_), .Y(men_men_n784_));
  INV        u762(.A(men_men_n784_), .Y(men_men_n785_));
  NO3        u763(.A(men_men_n436_), .B(men_men_n85_), .C(men_men_n45_), .Y(men_men_n786_));
  OA210      u764(.A0(men_men_n786_), .A1(men_men_n785_), .B0(men_men_n170_), .Y(men_men_n787_));
  NA3        u765(.A(men_men_n771_), .B(men_men_n580_), .C(men_men_n358_), .Y(men_men_n788_));
  NA2        u766(.A(men_men_n788_), .B(men_men_n40_), .Y(men_men_n789_));
  NO3        u767(.A(men_men_n602_), .B(men_men_n439_), .C(men_men_n128_), .Y(men_men_n790_));
  AN2        u768(.A(men_men_n438_), .B(men_men_n56_), .Y(men_men_n791_));
  NO2        u769(.A(men_men_n791_), .B(men_men_n790_), .Y(men_men_n792_));
  AOI210     u770(.A0(men_men_n792_), .A1(men_men_n789_), .B0(men_men_n49_), .Y(men_men_n793_));
  NO4        u771(.A(men_men_n363_), .B(men_men_n370_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n794_));
  NA2        u772(.A(men_men_n181_), .B(men_men_n549_), .Y(men_men_n795_));
  NOi21      u773(.An(men_men_n795_), .B(men_men_n794_), .Y(men_men_n796_));
  NA2        u774(.A(men_men_n665_), .B(men_men_n640_), .Y(men_men_n797_));
  NA2        u775(.A(men_men_n319_), .B(i_5_), .Y(men_men_n798_));
  OAI220     u776(.A0(men_men_n798_), .A1(men_men_n797_), .B0(men_men_n796_), .B1(men_men_n64_), .Y(men_men_n799_));
  NOi21      u777(.An(i_5_), .B(i_9_), .Y(men_men_n800_));
  NA2        u778(.A(men_men_n800_), .B(men_men_n433_), .Y(men_men_n801_));
  AOI210     u779(.A0(men_men_n255_), .A1(men_men_n456_), .B0(men_men_n647_), .Y(men_men_n802_));
  NO3        u780(.A(men_men_n400_), .B(men_men_n255_), .C(men_men_n70_), .Y(men_men_n803_));
  NO2        u781(.A(men_men_n171_), .B(men_men_n145_), .Y(men_men_n804_));
  INV        u782(.A(men_men_n803_), .Y(men_men_n805_));
  OAI220     u783(.A0(men_men_n805_), .A1(men_men_n177_), .B0(men_men_n802_), .B1(men_men_n801_), .Y(men_men_n806_));
  NO4        u784(.A(men_men_n806_), .B(men_men_n799_), .C(men_men_n793_), .D(men_men_n787_), .Y(men_men_n807_));
  NA2        u785(.A(men_men_n181_), .B(men_men_n24_), .Y(men_men_n808_));
  NO2        u786(.A(men_men_n639_), .B(men_men_n572_), .Y(men_men_n809_));
  NO2        u787(.A(men_men_n809_), .B(men_men_n808_), .Y(men_men_n810_));
  NA2        u788(.A(men_men_n300_), .B(men_men_n126_), .Y(men_men_n811_));
  NAi21      u789(.An(men_men_n159_), .B(i_5_), .Y(men_men_n812_));
  NO2        u790(.A(men_men_n811_), .B(men_men_n386_), .Y(men_men_n813_));
  NO2        u791(.A(men_men_n813_), .B(men_men_n810_), .Y(men_men_n814_));
  NO2        u792(.A(men_men_n377_), .B(men_men_n281_), .Y(men_men_n815_));
  NA2        u793(.A(men_men_n815_), .B(men_men_n668_), .Y(men_men_n816_));
  NA2        u794(.A(men_men_n550_), .B(i_0_), .Y(men_men_n817_));
  NO2        u795(.A(men_men_n817_), .B(men_men_n372_), .Y(men_men_n818_));
  INV        u796(.A(men_men_n818_), .Y(men_men_n819_));
  AN2        u797(.A(men_men_n92_), .B(men_men_n238_), .Y(men_men_n820_));
  NA2        u798(.A(men_men_n702_), .B(men_men_n315_), .Y(men_men_n821_));
  AOI210     u799(.A0(men_men_n462_), .A1(men_men_n83_), .B0(men_men_n59_), .Y(men_men_n822_));
  OAI220     u800(.A0(men_men_n822_), .A1(men_men_n821_), .B0(men_men_n629_), .B1(men_men_n513_), .Y(men_men_n823_));
  NA2        u801(.A(i_0_), .B(i_10_), .Y(men_men_n824_));
  NA2        u802(.A(men_men_n319_), .B(men_men_n94_), .Y(men_men_n825_));
  NA2        u803(.A(men_men_n544_), .B(i_4_), .Y(men_men_n826_));
  NA2        u804(.A(men_men_n184_), .B(men_men_n198_), .Y(men_men_n827_));
  OAI220     u805(.A0(men_men_n827_), .A1(men_men_n821_), .B0(men_men_n826_), .B1(men_men_n825_), .Y(men_men_n828_));
  NO3        u806(.A(men_men_n828_), .B(men_men_n823_), .C(men_men_n820_), .Y(men_men_n829_));
  NA4        u807(.A(men_men_n829_), .B(men_men_n819_), .C(men_men_n816_), .D(men_men_n814_), .Y(men_men_n830_));
  NO2        u808(.A(men_men_n99_), .B(men_men_n37_), .Y(men_men_n831_));
  NA2        u809(.A(i_11_), .B(i_9_), .Y(men_men_n832_));
  NO3        u810(.A(i_12_), .B(men_men_n832_), .C(men_men_n579_), .Y(men_men_n833_));
  AN2        u811(.A(men_men_n833_), .B(men_men_n831_), .Y(men_men_n834_));
  NO2        u812(.A(men_men_n49_), .B(i_7_), .Y(men_men_n835_));
  NA2        u813(.A(men_men_n381_), .B(men_men_n175_), .Y(men_men_n836_));
  NA2        u814(.A(men_men_n836_), .B(men_men_n157_), .Y(men_men_n837_));
  NO2        u815(.A(men_men_n171_), .B(i_0_), .Y(men_men_n838_));
  INV        u816(.A(men_men_n838_), .Y(men_men_n839_));
  NA2        u817(.A(men_men_n454_), .B(men_men_n228_), .Y(men_men_n840_));
  AOI210     u818(.A0(men_men_n357_), .A1(men_men_n42_), .B0(men_men_n393_), .Y(men_men_n841_));
  OAI220     u819(.A0(men_men_n841_), .A1(men_men_n801_), .B0(men_men_n840_), .B1(men_men_n839_), .Y(men_men_n842_));
  NO3        u820(.A(men_men_n842_), .B(men_men_n837_), .C(men_men_n834_), .Y(men_men_n843_));
  NA2        u821(.A(men_men_n628_), .B(men_men_n118_), .Y(men_men_n844_));
  NO2        u822(.A(i_6_), .B(men_men_n844_), .Y(men_men_n845_));
  AOI210     u823(.A0(men_men_n435_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n846_));
  NA2        u824(.A(men_men_n168_), .B(men_men_n99_), .Y(men_men_n847_));
  NOi32      u825(.An(men_men_n846_), .Bn(men_men_n184_), .C(men_men_n847_), .Y(men_men_n848_));
  NO2        u826(.A(men_men_n848_), .B(men_men_n845_), .Y(men_men_n849_));
  NOi21      u827(.An(i_7_), .B(i_5_), .Y(men_men_n850_));
  NOi31      u828(.An(men_men_n850_), .B(i_0_), .C(men_men_n683_), .Y(men_men_n851_));
  OR2        u829(.A(men_men_n847_), .B(men_men_n491_), .Y(men_men_n852_));
  NO3        u830(.A(men_men_n389_), .B(men_men_n351_), .C(men_men_n347_), .Y(men_men_n853_));
  NO2        u831(.A(men_men_n249_), .B(men_men_n304_), .Y(men_men_n854_));
  INV        u832(.A(men_men_n683_), .Y(men_men_n855_));
  AOI210     u833(.A0(men_men_n855_), .A1(men_men_n854_), .B0(men_men_n853_), .Y(men_men_n856_));
  NA4        u834(.A(men_men_n856_), .B(men_men_n852_), .C(men_men_n849_), .D(men_men_n843_), .Y(men_men_n857_));
  NO2        u835(.A(men_men_n808_), .B(men_men_n235_), .Y(men_men_n858_));
  AN2        u836(.A(men_men_n318_), .B(men_men_n315_), .Y(men_men_n859_));
  AN2        u837(.A(men_men_n859_), .B(men_men_n804_), .Y(men_men_n860_));
  OAI210     u838(.A0(men_men_n860_), .A1(men_men_n858_), .B0(i_10_), .Y(men_men_n861_));
  OA210      u839(.A0(men_men_n454_), .A1(men_men_n220_), .B0(men_men_n453_), .Y(men_men_n862_));
  NA3        u840(.A(men_men_n453_), .B(men_men_n397_), .C(men_men_n46_), .Y(men_men_n863_));
  OAI210     u841(.A0(men_men_n812_), .A1(i_6_), .B0(men_men_n863_), .Y(men_men_n864_));
  NO2        u842(.A(men_men_n247_), .B(men_men_n47_), .Y(men_men_n865_));
  NO2        u843(.A(men_men_n865_), .B(men_men_n183_), .Y(men_men_n866_));
  AOI220     u844(.A0(men_men_n866_), .A1(men_men_n454_), .B0(men_men_n864_), .B1(men_men_n70_), .Y(men_men_n867_));
  NA3        u845(.A(men_men_n760_), .B(men_men_n369_), .C(men_men_n609_), .Y(men_men_n868_));
  NA2        u846(.A(men_men_n88_), .B(men_men_n45_), .Y(men_men_n869_));
  NO2        u847(.A(men_men_n72_), .B(men_men_n704_), .Y(men_men_n870_));
  AOI220     u848(.A0(men_men_n870_), .A1(men_men_n869_), .B0(men_men_n170_), .B1(men_men_n572_), .Y(men_men_n871_));
  AOI210     u849(.A0(men_men_n871_), .A1(men_men_n868_), .B0(men_men_n48_), .Y(men_men_n872_));
  NO3        u850(.A(men_men_n564_), .B(men_men_n346_), .C(men_men_n24_), .Y(men_men_n873_));
  AOI210     u851(.A0(men_men_n661_), .A1(men_men_n524_), .B0(men_men_n873_), .Y(men_men_n874_));
  NO2        u852(.A(men_men_n575_), .B(men_men_n101_), .Y(men_men_n875_));
  NA2        u853(.A(men_men_n875_), .B(i_0_), .Y(men_men_n876_));
  OAI220     u854(.A0(men_men_n876_), .A1(men_men_n82_), .B0(men_men_n874_), .B1(men_men_n169_), .Y(men_men_n877_));
  NO3        u855(.A(men_men_n877_), .B(men_men_n872_), .C(men_men_n495_), .Y(men_men_n878_));
  NA3        u856(.A(men_men_n878_), .B(men_men_n867_), .C(men_men_n861_), .Y(men_men_n879_));
  NO3        u857(.A(men_men_n879_), .B(men_men_n857_), .C(men_men_n830_), .Y(men_men_n880_));
  NO2        u858(.A(i_0_), .B(men_men_n683_), .Y(men_men_n881_));
  NO3        u859(.A(men_men_n101_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n882_));
  AO220      u860(.A0(men_men_n882_), .A1(men_men_n70_), .B0(men_men_n881_), .B1(men_men_n170_), .Y(men_men_n883_));
  NA2        u861(.A(men_men_n883_), .B(men_men_n336_), .Y(men_men_n884_));
  NA2        u862(.A(men_men_n690_), .B(men_men_n143_), .Y(men_men_n885_));
  INV        u863(.A(men_men_n885_), .Y(men_men_n886_));
  NA2        u864(.A(men_men_n886_), .B(men_men_n640_), .Y(men_men_n887_));
  NO2        u865(.A(men_men_n756_), .B(men_men_n389_), .Y(men_men_n888_));
  NA2        u866(.A(men_men_n782_), .B(men_men_n49_), .Y(men_men_n889_));
  NA2        u867(.A(men_men_n783_), .B(i_9_), .Y(men_men_n890_));
  NO2        u868(.A(men_men_n889_), .B(men_men_n890_), .Y(men_men_n891_));
  NA2        u869(.A(men_men_n239_), .B(men_men_n227_), .Y(men_men_n892_));
  AOI210     u870(.A0(men_men_n892_), .A1(men_men_n817_), .B0(men_men_n150_), .Y(men_men_n893_));
  NO3        u871(.A(men_men_n893_), .B(men_men_n891_), .C(men_men_n888_), .Y(men_men_n894_));
  NA3        u872(.A(men_men_n894_), .B(men_men_n887_), .C(men_men_n884_), .Y(men_men_n895_));
  NA2        u873(.A(men_men_n859_), .B(men_men_n359_), .Y(men_men_n896_));
  AOI210     u874(.A0(men_men_n288_), .A1(men_men_n159_), .B0(men_men_n896_), .Y(men_men_n897_));
  NA2        u875(.A(men_men_n40_), .B(men_men_n45_), .Y(men_men_n898_));
  NA2        u876(.A(men_men_n835_), .B(men_men_n467_), .Y(men_men_n899_));
  AOI210     u877(.A0(men_men_n898_), .A1(men_men_n159_), .B0(men_men_n899_), .Y(men_men_n900_));
  NO2        u878(.A(men_men_n900_), .B(men_men_n897_), .Y(men_men_n901_));
  NO3        u879(.A(men_men_n824_), .B(men_men_n800_), .C(men_men_n186_), .Y(men_men_n902_));
  AOI220     u880(.A0(men_men_n902_), .A1(i_11_), .B0(men_men_n545_), .B1(men_men_n72_), .Y(men_men_n903_));
  NO3        u881(.A(men_men_n205_), .B(men_men_n370_), .C(i_0_), .Y(men_men_n904_));
  OAI210     u882(.A0(men_men_n904_), .A1(men_men_n73_), .B0(i_13_), .Y(men_men_n905_));
  INV        u883(.A(men_men_n214_), .Y(men_men_n906_));
  OAI220     u884(.A0(men_men_n507_), .A1(men_men_n136_), .B0(men_men_n613_), .B1(men_men_n589_), .Y(men_men_n907_));
  NA3        u885(.A(men_men_n907_), .B(i_7_), .C(men_men_n906_), .Y(men_men_n908_));
  NA4        u886(.A(men_men_n908_), .B(men_men_n905_), .C(men_men_n903_), .D(men_men_n901_), .Y(men_men_n909_));
  NO2        u887(.A(men_men_n237_), .B(men_men_n88_), .Y(men_men_n910_));
  AOI210     u888(.A0(men_men_n910_), .A1(men_men_n881_), .B0(men_men_n105_), .Y(men_men_n911_));
  AOI220     u889(.A0(men_men_n850_), .A1(men_men_n467_), .B0(men_men_n782_), .B1(men_men_n160_), .Y(men_men_n912_));
  NA2        u890(.A(men_men_n339_), .B(men_men_n172_), .Y(men_men_n913_));
  OA220      u891(.A0(men_men_n913_), .A1(men_men_n912_), .B0(men_men_n911_), .B1(i_5_), .Y(men_men_n914_));
  AOI210     u892(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n171_), .Y(men_men_n915_));
  NA2        u893(.A(men_men_n915_), .B(men_men_n862_), .Y(men_men_n916_));
  NA3        u894(.A(men_men_n586_), .B(men_men_n181_), .C(men_men_n80_), .Y(men_men_n917_));
  NA2        u895(.A(men_men_n917_), .B(men_men_n522_), .Y(men_men_n918_));
  INV        u896(.A(men_men_n465_), .Y(men_men_n919_));
  NO2        u897(.A(men_men_n919_), .B(men_men_n918_), .Y(men_men_n920_));
  NA3        u898(.A(men_men_n377_), .B(men_men_n320_), .C(men_men_n218_), .Y(men_men_n921_));
  NA4        u899(.A(men_men_n921_), .B(men_men_n920_), .C(men_men_n916_), .D(men_men_n914_), .Y(men_men_n922_));
  INV        u900(.A(men_men_n588_), .Y(men_men_n923_));
  NO3        u901(.A(men_men_n923_), .B(men_men_n535_), .C(men_men_n333_), .Y(men_men_n924_));
  NO2        u902(.A(men_men_n82_), .B(i_5_), .Y(men_men_n925_));
  NA3        u903(.A(men_men_n783_), .B(men_men_n106_), .C(men_men_n121_), .Y(men_men_n926_));
  INV        u904(.A(men_men_n926_), .Y(men_men_n927_));
  AOI210     u905(.A0(men_men_n927_), .A1(men_men_n925_), .B0(men_men_n924_), .Y(men_men_n928_));
  NA3        u906(.A(men_men_n293_), .B(i_5_), .C(men_men_n189_), .Y(men_men_n929_));
  NAi31      u907(.An(men_men_n236_), .B(men_men_n929_), .C(men_men_n237_), .Y(men_men_n930_));
  NO4        u908(.A(men_men_n235_), .B(men_men_n205_), .C(i_0_), .D(i_12_), .Y(men_men_n931_));
  NA2        u909(.A(men_men_n931_), .B(men_men_n930_), .Y(men_men_n932_));
  AN2        u910(.A(men_men_n824_), .B(men_men_n150_), .Y(men_men_n933_));
  NO4        u911(.A(men_men_n933_), .B(i_12_), .C(men_men_n617_), .D(men_men_n128_), .Y(men_men_n934_));
  NA2        u912(.A(men_men_n934_), .B(men_men_n214_), .Y(men_men_n935_));
  NA3        u913(.A(men_men_n94_), .B(men_men_n549_), .C(i_11_), .Y(men_men_n936_));
  NO2        u914(.A(men_men_n936_), .B(men_men_n152_), .Y(men_men_n937_));
  NA2        u915(.A(men_men_n850_), .B(men_men_n451_), .Y(men_men_n938_));
  OAI220     u916(.A0(i_7_), .A1(men_men_n929_), .B0(men_men_n938_), .B1(men_men_n641_), .Y(men_men_n939_));
  AOI210     u917(.A0(men_men_n939_), .A1(men_men_n838_), .B0(men_men_n937_), .Y(men_men_n940_));
  NA4        u918(.A(men_men_n940_), .B(men_men_n935_), .C(men_men_n932_), .D(men_men_n928_), .Y(men_men_n941_));
  NO4        u919(.A(men_men_n941_), .B(men_men_n922_), .C(men_men_n909_), .D(men_men_n895_), .Y(men_men_n942_));
  OAI210     u920(.A0(men_men_n759_), .A1(men_men_n752_), .B0(men_men_n37_), .Y(men_men_n943_));
  NA3        u921(.A(men_men_n846_), .B(men_men_n354_), .C(i_5_), .Y(men_men_n944_));
  NA3        u922(.A(men_men_n944_), .B(men_men_n943_), .C(men_men_n584_), .Y(men_men_n945_));
  NA2        u923(.A(men_men_n945_), .B(men_men_n201_), .Y(men_men_n946_));
  BUFFER     u924(.A(men_men_n355_), .Y(men_men_n947_));
  NA2        u925(.A(men_men_n182_), .B(men_men_n184_), .Y(men_men_n948_));
  AO210      u926(.A0(men_men_n947_), .A1(men_men_n33_), .B0(men_men_n948_), .Y(men_men_n949_));
  OAI210     u927(.A0(men_men_n588_), .A1(men_men_n586_), .B0(men_men_n303_), .Y(men_men_n950_));
  INV        u928(.A(men_men_n614_), .Y(men_men_n951_));
  NA3        u929(.A(men_men_n951_), .B(men_men_n950_), .C(men_men_n949_), .Y(men_men_n952_));
  NO2        u930(.A(men_men_n443_), .B(men_men_n255_), .Y(men_men_n953_));
  NO4        u931(.A(men_men_n230_), .B(men_men_n142_), .C(men_men_n642_), .D(men_men_n37_), .Y(men_men_n954_));
  NO2        u932(.A(men_men_n954_), .B(men_men_n953_), .Y(men_men_n955_));
  OAI210     u933(.A0(men_men_n936_), .A1(men_men_n145_), .B0(men_men_n955_), .Y(men_men_n956_));
  AOI210     u934(.A0(men_men_n952_), .A1(men_men_n49_), .B0(men_men_n956_), .Y(men_men_n957_));
  AOI210     u935(.A0(men_men_n957_), .A1(men_men_n946_), .B0(men_men_n70_), .Y(men_men_n958_));
  NO2        u936(.A(men_men_n542_), .B(men_men_n366_), .Y(men_men_n959_));
  NO2        u937(.A(men_men_n959_), .B(men_men_n710_), .Y(men_men_n960_));
  OAI210     u938(.A0(men_men_n77_), .A1(men_men_n55_), .B0(men_men_n104_), .Y(men_men_n961_));
  NA2        u939(.A(men_men_n961_), .B(men_men_n73_), .Y(men_men_n962_));
  AOI210     u940(.A0(men_men_n915_), .A1(men_men_n835_), .B0(men_men_n851_), .Y(men_men_n963_));
  AOI210     u941(.A0(men_men_n963_), .A1(men_men_n962_), .B0(men_men_n642_), .Y(men_men_n964_));
  NA2        u942(.A(men_men_n249_), .B(men_men_n58_), .Y(men_men_n965_));
  AOI220     u943(.A0(men_men_n965_), .A1(men_men_n73_), .B0(men_men_n334_), .B1(men_men_n246_), .Y(men_men_n966_));
  NO2        u944(.A(men_men_n966_), .B(men_men_n233_), .Y(men_men_n967_));
  NA3        u945(.A(men_men_n92_), .B(men_men_n295_), .C(men_men_n31_), .Y(men_men_n968_));
  INV        u946(.A(men_men_n968_), .Y(men_men_n969_));
  NO3        u947(.A(men_men_n969_), .B(men_men_n967_), .C(men_men_n964_), .Y(men_men_n970_));
  OAI210     u948(.A0(men_men_n257_), .A1(men_men_n155_), .B0(men_men_n83_), .Y(men_men_n971_));
  NA3        u949(.A(men_men_n713_), .B(men_men_n277_), .C(men_men_n77_), .Y(men_men_n972_));
  AOI210     u950(.A0(men_men_n972_), .A1(men_men_n971_), .B0(i_11_), .Y(men_men_n973_));
  NA2        u951(.A(men_men_n581_), .B(men_men_n211_), .Y(men_men_n974_));
  OAI210     u952(.A0(men_men_n974_), .A1(men_men_n846_), .B0(men_men_n201_), .Y(men_men_n975_));
  NA2        u953(.A(men_men_n161_), .B(i_5_), .Y(men_men_n976_));
  NO2        u954(.A(men_men_n975_), .B(men_men_n976_), .Y(men_men_n977_));
  NO3        u955(.A(men_men_n60_), .B(men_men_n59_), .C(i_4_), .Y(men_men_n978_));
  OAI210     u956(.A0(men_men_n854_), .A1(men_men_n295_), .B0(men_men_n978_), .Y(men_men_n979_));
  NO2        u957(.A(men_men_n979_), .B(men_men_n683_), .Y(men_men_n980_));
  NO3        u958(.A(men_men_n980_), .B(men_men_n977_), .C(men_men_n973_), .Y(men_men_n981_));
  OAI210     u959(.A0(men_men_n970_), .A1(i_4_), .B0(men_men_n981_), .Y(men_men_n982_));
  NO3        u960(.A(men_men_n982_), .B(men_men_n960_), .C(men_men_n958_), .Y(men_men_n983_));
  NA4        u961(.A(men_men_n983_), .B(men_men_n942_), .C(men_men_n880_), .D(men_men_n807_), .Y(men4));
  INV        u962(.A(i_2_), .Y(men_men_n987_));
  INV        u963(.A(men_men_n315_), .Y(men_men_n988_));
  INV        u964(.A(i_1_), .Y(men_men_n989_));
  INV        u965(.A(men_men_n721_), .Y(men_men_n990_));
  INV        u966(.A(men_men_n293_), .Y(men_men_n991_));
  INV        u967(.A(i_0_), .Y(men_men_n992_));
  INV        u968(.A(i_3_), .Y(men_men_n993_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule