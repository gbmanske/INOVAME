library verilog;
use verilog.vl_types.all;
entity shifter_vlg_vec_tst is
end shifter_vlg_vec_tst;
