//Benchmark atmr_alu4_1266_0.25

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n118_, ori_ori_n119_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  INV        o019(.A(ori_ori_n35_), .Y(ori1));
  INV        o020(.A(i_11_), .Y(ori_ori_n43_));
  NO2        o021(.A(ori_ori_n43_), .B(i_6_), .Y(ori_ori_n44_));
  INV        o022(.A(i_2_), .Y(ori_ori_n45_));
  NA2        o023(.A(i_0_), .B(i_3_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_5_), .A1(ori_ori_n46_), .B0(ori_ori_n45_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_0_), .B(i_2_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NA2        o031(.A(ori_ori_n50_), .B(ori_ori_n44_), .Y(ori_ori_n54_));
  NO2        o032(.A(i_1_), .B(i_6_), .Y(ori_ori_n55_));
  NA2        o033(.A(i_8_), .B(i_7_), .Y(ori_ori_n56_));
  INV        o034(.A(ori_ori_n56_), .Y(ori_ori_n57_));
  NA2        o035(.A(ori_ori_n57_), .B(i_12_), .Y(ori_ori_n58_));
  NAi21      o036(.An(i_2_), .B(i_7_), .Y(ori_ori_n59_));
  INV        o037(.A(i_1_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_6_), .Y(ori_ori_n61_));
  NA2        o039(.A(i_1_), .B(i_10_), .Y(ori_ori_n62_));
  NO2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NAi21      o041(.An(ori_ori_n63_), .B(ori_ori_n58_), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n65_));
  AOI210     o043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n66_));
  NA2        o044(.A(i_1_), .B(i_6_), .Y(ori_ori_n67_));
  NO2        o045(.A(ori_ori_n67_), .B(ori_ori_n25_), .Y(ori_ori_n68_));
  INV        o046(.A(i_0_), .Y(ori_ori_n69_));
  NAi21      o047(.An(i_5_), .B(i_10_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_5_), .B(i_9_), .Y(ori_ori_n71_));
  AOI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n70_), .B0(ori_ori_n69_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n72_), .B(ori_ori_n68_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n66_), .A1(ori_ori_n65_), .B0(ori_ori_n73_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n64_), .B0(i_0_), .Y(ori_ori_n75_));
  NA2        o053(.A(i_12_), .B(i_5_), .Y(ori_ori_n76_));
  NO2        o054(.A(i_3_), .B(i_9_), .Y(ori_ori_n77_));
  NO2        o055(.A(i_3_), .B(i_7_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n77_), .B(ori_ori_n60_), .Y(ori_ori_n79_));
  INV        o057(.A(i_6_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_2_), .B(i_7_), .Y(ori_ori_n81_));
  INV        o059(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  OAI210     o060(.A0(ori_ori_n79_), .A1(i_8_), .B0(ori_ori_n82_), .Y(ori_ori_n83_));
  NAi21      o061(.An(i_6_), .B(i_10_), .Y(ori_ori_n84_));
  NA2        o062(.A(i_6_), .B(i_9_), .Y(ori_ori_n85_));
  AOI210     o063(.A0(ori_ori_n85_), .A1(ori_ori_n84_), .B0(ori_ori_n60_), .Y(ori_ori_n86_));
  NA2        o064(.A(i_2_), .B(i_6_), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n87_), .B(ori_ori_n25_), .Y(ori_ori_n88_));
  NO2        o066(.A(ori_ori_n88_), .B(ori_ori_n86_), .Y(ori_ori_n89_));
  AOI210     o067(.A0(ori_ori_n89_), .A1(ori_ori_n83_), .B0(ori_ori_n76_), .Y(ori_ori_n90_));
  AN3        o068(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n91_));
  NAi21      o069(.An(i_6_), .B(i_11_), .Y(ori_ori_n92_));
  INV        o070(.A(i_7_), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n45_), .B(ori_ori_n93_), .Y(ori_ori_n94_));
  NO2        o072(.A(i_0_), .B(i_5_), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n95_), .B(ori_ori_n80_), .Y(ori_ori_n96_));
  NA2        o074(.A(i_12_), .B(i_3_), .Y(ori_ori_n97_));
  INV        o075(.A(ori_ori_n97_), .Y(ori_ori_n98_));
  NA3        o076(.A(ori_ori_n98_), .B(ori_ori_n96_), .C(ori_ori_n94_), .Y(ori_ori_n99_));
  NAi21      o077(.An(i_7_), .B(i_11_), .Y(ori_ori_n100_));
  AN2        o078(.A(i_2_), .B(i_10_), .Y(ori_ori_n101_));
  BUFFER     o079(.A(ori_ori_n76_), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n60_), .B(ori_ori_n26_), .Y(ori_ori_n103_));
  NA2        o081(.A(i_11_), .B(i_12_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n104_), .B(ori_ori_n99_), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n93_), .B(ori_ori_n37_), .Y(ori_ori_n106_));
  NA2        o084(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n107_), .B(ori_ori_n106_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n108_), .B(ori_ori_n45_), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n110_));
  NAi21      o088(.An(i_3_), .B(i_8_), .Y(ori_ori_n111_));
  NO2        o089(.A(i_1_), .B(ori_ori_n80_), .Y(ori_ori_n112_));
  NO2        o090(.A(i_6_), .B(i_5_), .Y(ori_ori_n113_));
  AO210      o091(.A0(i_5_), .A1(ori_ori_n46_), .B0(ori_ori_n112_), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n114_), .B(ori_ori_n100_), .Y(ori_ori_n115_));
  NO3        o093(.A(ori_ori_n115_), .B(ori_ori_n105_), .C(ori_ori_n90_), .Y(ori_ori_n116_));
  NA3        o094(.A(ori_ori_n116_), .B(ori_ori_n75_), .C(ori_ori_n54_), .Y(ori2));
  NO2        o095(.A(ori_ori_n60_), .B(ori_ori_n37_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n479_), .B(ori_ori_n118_), .Y(ori_ori_n119_));
  NA4        o097(.A(ori_ori_n119_), .B(ori_ori_n73_), .C(ori_ori_n65_), .D(ori_ori_n30_), .Y(ori0));
  NA2        o098(.A(i_7_), .B(i_6_), .Y(ori_ori_n121_));
  NO2        o099(.A(i_12_), .B(i_13_), .Y(ori_ori_n122_));
  NAi21      o100(.An(i_5_), .B(i_11_), .Y(ori_ori_n123_));
  NO2        o101(.A(i_0_), .B(i_1_), .Y(ori_ori_n124_));
  AN2        o102(.A(ori_ori_n122_), .B(ori_ori_n77_), .Y(ori_ori_n125_));
  NA2        o103(.A(i_1_), .B(i_5_), .Y(ori_ori_n126_));
  OR2        o104(.A(i_0_), .B(i_1_), .Y(ori_ori_n127_));
  NOi21      o105(.An(i_4_), .B(i_10_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n40_), .Y(ori_ori_n129_));
  NOi21      o107(.An(i_4_), .B(i_9_), .Y(ori_ori_n130_));
  NOi21      o108(.An(i_11_), .B(i_13_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n131_), .B(ori_ori_n130_), .Y(ori_ori_n132_));
  NO2        o110(.A(ori_ori_n69_), .B(ori_ori_n60_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n69_), .B(i_5_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_2_), .B(i_1_), .Y(ori_ori_n135_));
  NAi21      o113(.An(i_4_), .B(i_12_), .Y(ori_ori_n136_));
  INV        o114(.A(i_8_), .Y(ori_ori_n137_));
  NO2        o115(.A(i_3_), .B(i_8_), .Y(ori_ori_n138_));
  NO3        o116(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n95_), .B(ori_ori_n55_), .Y(ori_ori_n140_));
  NO2        o118(.A(i_13_), .B(i_9_), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n43_), .B(i_5_), .Y(ori_ori_n142_));
  NA2        o120(.A(i_0_), .B(i_5_), .Y(ori_ori_n143_));
  NAi31      o121(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n144_));
  INV        o122(.A(i_13_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_12_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  INV        o124(.A(i_12_), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n43_), .B(ori_ori_n147_), .Y(ori_ori_n148_));
  NO3        o126(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n149_));
  NA2        o127(.A(i_2_), .B(i_1_), .Y(ori_ori_n150_));
  NO3        o128(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n151_));
  NAi21      o129(.An(i_4_), .B(i_3_), .Y(ori_ori_n152_));
  NOi41      o130(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n153_));
  NO2        o131(.A(i_11_), .B(ori_ori_n145_), .Y(ori_ori_n154_));
  NOi21      o132(.An(i_1_), .B(i_6_), .Y(ori_ori_n155_));
  INV        o133(.A(i_7_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n147_), .B(i_9_), .Y(ori_ori_n157_));
  OR4        o135(.A(ori_ori_n157_), .B(ori_ori_n156_), .C(ori_ori_n155_), .D(ori_ori_n134_), .Y(ori_ori_n158_));
  NA2        o136(.A(ori_ori_n69_), .B(i_5_), .Y(ori_ori_n159_));
  NA2        o137(.A(i_3_), .B(i_9_), .Y(ori_ori_n160_));
  NAi21      o138(.An(i_7_), .B(i_10_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n161_), .B(ori_ori_n160_), .Y(ori_ori_n162_));
  NA3        o140(.A(ori_ori_n162_), .B(ori_ori_n159_), .C(ori_ori_n61_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n163_), .B(ori_ori_n158_), .Y(ori_ori_n164_));
  INV        o142(.A(ori_ori_n121_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n147_), .B(i_13_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n166_), .B(ori_ori_n71_), .Y(ori_ori_n167_));
  AOI220     o145(.A0(ori_ori_n167_), .A1(ori_ori_n165_), .B0(ori_ori_n164_), .B1(ori_ori_n154_), .Y(ori_ori_n168_));
  NA2        o146(.A(i_12_), .B(i_6_), .Y(ori_ori_n169_));
  OR2        o147(.A(i_13_), .B(i_9_), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n152_), .B(i_2_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n154_), .B(i_9_), .Y(ori_ori_n172_));
  NO3        o150(.A(i_12_), .B(ori_ori_n145_), .C(ori_ori_n37_), .Y(ori_ori_n173_));
  AN2        o151(.A(i_3_), .B(i_10_), .Y(ori_ori_n174_));
  NO2        o152(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n45_), .B(ori_ori_n26_), .Y(ori_ori_n176_));
  NO3        o154(.A(ori_ori_n43_), .B(i_13_), .C(i_9_), .Y(ori_ori_n177_));
  NO2        o155(.A(i_2_), .B(i_3_), .Y(ori_ori_n178_));
  NO2        o156(.A(i_12_), .B(i_10_), .Y(ori_ori_n179_));
  NOi21      o157(.An(i_5_), .B(i_0_), .Y(ori_ori_n180_));
  NOi21      o158(.An(ori_ori_n126_), .B(ori_ori_n96_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n181_), .B(ori_ori_n107_), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n182_), .B(i_3_), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n137_), .B(i_9_), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n184_), .B(ori_ori_n140_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n185_), .B(ori_ori_n45_), .Y(ori_ori_n186_));
  INV        o164(.A(ori_ori_n186_), .Y(ori_ori_n187_));
  AOI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n183_), .B0(ori_ori_n129_), .Y(ori_ori_n188_));
  INV        o166(.A(ori_ori_n188_), .Y(ori_ori_n189_));
  NOi32      o167(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n190_));
  INV        o168(.A(ori_ori_n190_), .Y(ori_ori_n191_));
  NOi32      o169(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n192_));
  NO2        o170(.A(i_1_), .B(ori_ori_n93_), .Y(ori_ori_n193_));
  NAi21      o171(.An(i_3_), .B(i_4_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n194_), .B(i_9_), .Y(ori_ori_n195_));
  AN2        o173(.A(i_6_), .B(i_7_), .Y(ori_ori_n196_));
  OAI210     o174(.A0(ori_ori_n196_), .A1(ori_ori_n193_), .B0(ori_ori_n195_), .Y(ori_ori_n197_));
  NA2        o175(.A(i_2_), .B(i_7_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n194_), .B(i_10_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n197_), .B(ori_ori_n134_), .Y(ori_ori_n200_));
  AOI210     o178(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n201_));
  OAI210     o179(.A0(ori_ori_n201_), .A1(ori_ori_n135_), .B0(ori_ori_n199_), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n202_), .B(i_5_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n203_), .B(ori_ori_n200_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(ori_ori_n191_), .Y(ori_ori_n205_));
  AN2        o183(.A(i_12_), .B(i_5_), .Y(ori_ori_n206_));
  NO2        o184(.A(i_11_), .B(i_6_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_5_), .B(i_10_), .Y(ori_ori_n208_));
  NO2        o186(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n209_));
  NO3        o187(.A(i_1_), .B(i_12_), .C(ori_ori_n80_), .Y(ori_ori_n210_));
  NO2        o188(.A(i_0_), .B(i_11_), .Y(ori_ori_n211_));
  BUFFER     o189(.A(i_6_), .Y(ori_ori_n212_));
  NAi21      o190(.An(i_9_), .B(i_4_), .Y(ori_ori_n213_));
  OR2        o191(.A(i_13_), .B(i_10_), .Y(ori_ori_n214_));
  NO3        o192(.A(ori_ori_n214_), .B(ori_ori_n104_), .C(ori_ori_n213_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n93_), .B(ori_ori_n25_), .Y(ori_ori_n216_));
  NA2        o194(.A(ori_ori_n173_), .B(ori_ori_n216_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n217_), .B(ori_ori_n181_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n137_), .B(i_10_), .Y(ori_ori_n219_));
  NA3        o197(.A(ori_ori_n159_), .B(ori_ori_n61_), .C(i_2_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n221_));
  INV        o199(.A(ori_ori_n221_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n222_), .B(ori_ori_n172_), .Y(ori_ori_n223_));
  NO3        o201(.A(ori_ori_n223_), .B(ori_ori_n218_), .C(ori_ori_n205_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n69_), .B(i_13_), .Y(ori_ori_n225_));
  NO2        o203(.A(i_10_), .B(i_9_), .Y(ori_ori_n226_));
  NO3        o204(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n169_), .B(ori_ori_n92_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n228_), .B(ori_ori_n227_), .Y(ori_ori_n229_));
  NA2        o207(.A(i_8_), .B(i_9_), .Y(ori_ori_n230_));
  NO2        o208(.A(i_7_), .B(i_2_), .Y(ori_ori_n231_));
  OR2        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n173_), .B(ori_ori_n140_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n233_), .B(ori_ori_n232_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n154_), .B(ori_ori_n175_), .Y(ori_ori_n235_));
  NO3        o213(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NA3        o215(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n238_));
  NA4        o216(.A(ori_ori_n123_), .B(ori_ori_n103_), .C(ori_ori_n76_), .D(ori_ori_n23_), .Y(ori_ori_n239_));
  OAI220     o217(.A0(ori_ori_n239_), .A1(ori_ori_n238_), .B0(ori_ori_n237_), .B1(ori_ori_n235_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n240_), .B(ori_ori_n234_), .Y(ori_ori_n241_));
  NA2        o219(.A(ori_ori_n91_), .B(i_13_), .Y(ori_ori_n242_));
  NO2        o220(.A(i_11_), .B(i_1_), .Y(ori_ori_n243_));
  NA3        o221(.A(ori_ori_n153_), .B(ori_ori_n131_), .C(ori_ori_n113_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n45_), .B(ori_ori_n43_), .Y(ori_ori_n245_));
  NO2        o223(.A(ori_ori_n127_), .B(i_3_), .Y(ori_ori_n246_));
  NAi31      o224(.An(ori_ori_n245_), .B(ori_ori_n246_), .C(ori_ori_n146_), .Y(ori_ori_n247_));
  NA2        o225(.A(ori_ori_n247_), .B(ori_ori_n244_), .Y(ori_ori_n248_));
  INV        o226(.A(ori_ori_n248_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n227_), .B(ori_ori_n206_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n236_), .B(ori_ori_n208_), .Y(ori_ori_n251_));
  NA2        o229(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n177_), .B(ori_ori_n149_), .Y(ori_ori_n253_));
  OAI220     o231(.A0(ori_ori_n253_), .A1(ori_ori_n220_), .B0(ori_ori_n252_), .B1(ori_ori_n242_), .Y(ori_ori_n254_));
  INV        o232(.A(ori_ori_n254_), .Y(ori_ori_n255_));
  NA3        o233(.A(ori_ori_n255_), .B(ori_ori_n249_), .C(ori_ori_n241_), .Y(ori_ori_n256_));
  NA2        o234(.A(ori_ori_n206_), .B(ori_ori_n145_), .Y(ori_ori_n257_));
  NA2        o235(.A(ori_ori_n196_), .B(ori_ori_n192_), .Y(ori_ori_n258_));
  OR2        o236(.A(ori_ori_n257_), .B(ori_ori_n258_), .Y(ori_ori_n259_));
  AOI210     o237(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n215_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n260_), .B(ori_ori_n259_), .Y(ori_ori_n261_));
  NA3        o239(.A(ori_ori_n143_), .B(ori_ori_n67_), .C(ori_ori_n43_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n173_), .B(ori_ori_n78_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n262_), .B(ori_ori_n263_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n214_), .B(i_1_), .Y(ori_ori_n265_));
  NOi31      o243(.An(ori_ori_n265_), .B(ori_ori_n228_), .C(ori_ori_n69_), .Y(ori_ori_n266_));
  NOi21      o244(.An(i_10_), .B(i_6_), .Y(ori_ori_n267_));
  OR2        o245(.A(i_2_), .B(i_5_), .Y(ori_ori_n268_));
  NO3        o246(.A(ori_ori_n264_), .B(ori_ori_n261_), .C(ori_ori_n256_), .Y(ori_ori_n269_));
  NA4        o247(.A(ori_ori_n269_), .B(ori_ori_n224_), .C(ori_ori_n189_), .D(ori_ori_n168_), .Y(ori7));
  NO2        o248(.A(ori_ori_n87_), .B(ori_ori_n52_), .Y(ori_ori_n271_));
  NA2        o249(.A(i_11_), .B(ori_ori_n137_), .Y(ori_ori_n272_));
  NA3        o250(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n273_));
  NO2        o251(.A(ori_ori_n147_), .B(i_4_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n274_), .B(i_8_), .Y(ori_ori_n275_));
  NO2        o253(.A(ori_ori_n97_), .B(ori_ori_n273_), .Y(ori_ori_n276_));
  NA2        o254(.A(i_2_), .B(ori_ori_n80_), .Y(ori_ori_n277_));
  OAI210     o255(.A0(ori_ori_n81_), .A1(ori_ori_n138_), .B0(ori_ori_n139_), .Y(ori_ori_n278_));
  NO2        o256(.A(ori_ori_n276_), .B(ori_ori_n271_), .Y(ori_ori_n279_));
  AOI210     o257(.A0(ori_ori_n111_), .A1(ori_ori_n59_), .B0(i_10_), .Y(ori_ori_n280_));
  AOI210     o258(.A0(ori_ori_n280_), .A1(ori_ori_n147_), .B0(ori_ori_n128_), .Y(ori_ori_n281_));
  OR2        o259(.A(i_6_), .B(i_10_), .Y(ori_ori_n282_));
  OR3        o260(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n283_));
  OR2        o261(.A(ori_ori_n281_), .B(ori_ori_n170_), .Y(ori_ori_n284_));
  AOI210     o262(.A0(ori_ori_n284_), .A1(ori_ori_n279_), .B0(ori_ori_n60_), .Y(ori_ori_n285_));
  NOi21      o263(.An(i_11_), .B(i_7_), .Y(ori_ori_n286_));
  AO210      o264(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n287_));
  NO2        o265(.A(ori_ori_n287_), .B(ori_ori_n286_), .Y(ori_ori_n288_));
  NA2        o266(.A(ori_ori_n288_), .B(ori_ori_n141_), .Y(ori_ori_n289_));
  NA3        o267(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n290_));
  NO2        o268(.A(ori_ori_n289_), .B(ori_ori_n60_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n146_), .B(ori_ori_n60_), .Y(ori_ori_n292_));
  NO2        o270(.A(i_1_), .B(i_12_), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n292_), .Y(ori_ori_n294_));
  OAI210     o272(.A0(ori_ori_n294_), .A1(ori_ori_n291_), .B0(i_6_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n290_), .B(ori_ori_n100_), .Y(ori_ori_n296_));
  NA2        o274(.A(ori_ori_n296_), .B(i_6_), .Y(ori_ori_n297_));
  NO2        o275(.A(i_6_), .B(i_11_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n297_), .B(ori_ori_n229_), .Y(ori_ori_n299_));
  NO3        o277(.A(ori_ori_n282_), .B(i_7_), .C(ori_ori_n23_), .Y(ori_ori_n300_));
  AOI210     o278(.A0(i_1_), .A1(ori_ori_n162_), .B0(ori_ori_n300_), .Y(ori_ori_n301_));
  NO2        o279(.A(ori_ori_n301_), .B(ori_ori_n43_), .Y(ori_ori_n302_));
  INV        o280(.A(i_2_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n118_), .B(i_9_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n304_), .B(ori_ori_n303_), .Y(ori_ori_n305_));
  AOI210     o283(.A0(ori_ori_n243_), .A1(ori_ori_n216_), .B0(ori_ori_n151_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n306_), .B(ori_ori_n277_), .Y(ori_ori_n307_));
  OR2        o285(.A(ori_ori_n307_), .B(ori_ori_n305_), .Y(ori_ori_n308_));
  NO3        o286(.A(ori_ori_n308_), .B(ori_ori_n302_), .C(ori_ori_n299_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n147_), .B(ori_ori_n93_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n310_), .B(ori_ori_n286_), .Y(ori_ori_n311_));
  NA2        o289(.A(ori_ori_n311_), .B(i_1_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n312_), .B(ori_ori_n283_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n213_), .B(ori_ori_n80_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n313_), .B(ori_ori_n45_), .Y(ori_ori_n315_));
  NO2        o293(.A(i_7_), .B(ori_ori_n43_), .Y(ori_ori_n316_));
  NO3        o294(.A(ori_ori_n316_), .B(ori_ori_n176_), .C(ori_ori_n148_), .Y(ori_ori_n317_));
  NO2        o295(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n318_));
  NO2        o296(.A(ori_ori_n318_), .B(i_6_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n80_), .B(i_9_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n320_), .B(ori_ori_n60_), .Y(ori_ori_n321_));
  NO2        o299(.A(ori_ori_n321_), .B(ori_ori_n293_), .Y(ori_ori_n322_));
  NO4        o300(.A(ori_ori_n322_), .B(ori_ori_n319_), .C(ori_ori_n317_), .D(i_4_), .Y(ori_ori_n323_));
  INV        o301(.A(ori_ori_n323_), .Y(ori_ori_n324_));
  NA4        o302(.A(ori_ori_n324_), .B(ori_ori_n315_), .C(ori_ori_n309_), .D(ori_ori_n295_), .Y(ori_ori_n325_));
  AOI210     o303(.A0(ori_ori_n169_), .A1(ori_ori_n92_), .B0(i_1_), .Y(ori_ori_n326_));
  NO2        o304(.A(ori_ori_n194_), .B(i_2_), .Y(ori_ori_n327_));
  NA2        o305(.A(ori_ori_n327_), .B(ori_ori_n326_), .Y(ori_ori_n328_));
  NO2        o306(.A(ori_ori_n328_), .B(i_13_), .Y(ori_ori_n329_));
  OR2        o307(.A(i_11_), .B(i_7_), .Y(ori_ori_n330_));
  NO2        o308(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n331_));
  INV        o309(.A(ori_ori_n331_), .Y(ori_ori_n332_));
  NA2        o310(.A(i_7_), .B(ori_ori_n314_), .Y(ori_ori_n333_));
  OAI220     o311(.A0(ori_ori_n333_), .A1(ori_ori_n41_), .B0(ori_ori_n332_), .B1(ori_ori_n87_), .Y(ori_ori_n334_));
  INV        o312(.A(ori_ori_n334_), .Y(ori_ori_n335_));
  NA2        o313(.A(ori_ori_n110_), .B(i_13_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n336_), .B(ori_ori_n326_), .Y(ori_ori_n337_));
  INV        o315(.A(i_7_), .Y(ori_ori_n338_));
  AOI220     o316(.A0(ori_ori_n207_), .A1(ori_ori_n481_), .B0(ori_ori_n86_), .B1(ori_ori_n94_), .Y(ori_ori_n339_));
  NO2        o317(.A(ori_ori_n339_), .B(ori_ori_n275_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n340_), .B(ori_ori_n337_), .Y(ori_ori_n341_));
  OR2        o319(.A(i_11_), .B(i_6_), .Y(ori_ori_n342_));
  NA2        o320(.A(ori_ori_n274_), .B(i_7_), .Y(ori_ori_n343_));
  NO2        o321(.A(ori_ori_n343_), .B(ori_ori_n342_), .Y(ori_ori_n344_));
  NA2        o322(.A(ori_ori_n298_), .B(i_13_), .Y(ori_ori_n345_));
  INV        o323(.A(ori_ori_n345_), .Y(ori_ori_n346_));
  OAI210     o324(.A0(ori_ori_n346_), .A1(ori_ori_n344_), .B0(ori_ori_n60_), .Y(ori_ori_n347_));
  NO2        o325(.A(i_2_), .B(i_12_), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n193_), .B(ori_ori_n348_), .Y(ori_ori_n349_));
  NA2        o327(.A(ori_ori_n195_), .B(ori_ori_n193_), .Y(ori_ori_n350_));
  NA2        o328(.A(ori_ori_n350_), .B(ori_ori_n349_), .Y(ori_ori_n351_));
  NA3        o329(.A(ori_ori_n351_), .B(ori_ori_n44_), .C(ori_ori_n145_), .Y(ori_ori_n352_));
  NA4        o330(.A(ori_ori_n352_), .B(ori_ori_n347_), .C(ori_ori_n341_), .D(ori_ori_n335_), .Y(ori_ori_n353_));
  OR4        o331(.A(ori_ori_n353_), .B(ori_ori_n329_), .C(ori_ori_n325_), .D(ori_ori_n285_), .Y(ori5));
  NA2        o332(.A(ori_ori_n311_), .B(ori_ori_n171_), .Y(ori_ori_n355_));
  NA3        o333(.A(ori_ori_n24_), .B(ori_ori_n348_), .C(ori_ori_n100_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(ori_ori_n355_), .Y(ori_ori_n357_));
  NO2        o335(.A(ori_ori_n107_), .B(ori_ori_n23_), .Y(ori_ori_n358_));
  INV        o336(.A(ori_ori_n226_), .Y(ori_ori_n359_));
  NO2        o337(.A(ori_ori_n358_), .B(ori_ori_n357_), .Y(ori_ori_n360_));
  INV        o338(.A(ori_ori_n153_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n361_), .B(i_13_), .Y(ori_ori_n362_));
  INV        o340(.A(ori_ori_n362_), .Y(ori_ori_n363_));
  NO2        o341(.A(ori_ori_n136_), .B(ori_ori_n108_), .Y(ori_ori_n364_));
  OAI210     o342(.A0(ori_ori_n364_), .A1(ori_ori_n358_), .B0(i_2_), .Y(ori_ori_n365_));
  INV        o343(.A(ori_ori_n132_), .Y(ori_ori_n366_));
  NO3        o344(.A(ori_ori_n287_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n367_));
  NO2        o345(.A(ori_ori_n366_), .B(ori_ori_n367_), .Y(ori_ori_n368_));
  AOI210     o346(.A0(ori_ori_n368_), .A1(ori_ori_n365_), .B0(ori_ori_n137_), .Y(ori_ori_n369_));
  OA210      o347(.A0(ori_ori_n288_), .A1(ori_ori_n109_), .B0(i_13_), .Y(ori_ori_n370_));
  INV        o348(.A(ori_ori_n125_), .Y(ori_ori_n371_));
  NO2        o349(.A(ori_ori_n371_), .B(ori_ori_n198_), .Y(ori_ori_n372_));
  NA3        o350(.A(i_2_), .B(ori_ori_n174_), .C(ori_ori_n107_), .Y(ori_ori_n373_));
  INV        o351(.A(ori_ori_n373_), .Y(ori_ori_n374_));
  NO4        o352(.A(ori_ori_n374_), .B(ori_ori_n372_), .C(ori_ori_n370_), .D(ori_ori_n369_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n376_), .B(ori_ori_n109_), .Y(ori_ori_n377_));
  NO2        o355(.A(ori_ori_n377_), .B(ori_ori_n272_), .Y(ori_ori_n378_));
  NA2        o356(.A(ori_ori_n378_), .B(ori_ori_n36_), .Y(ori_ori_n379_));
  NA4        o357(.A(ori_ori_n379_), .B(ori_ori_n375_), .C(ori_ori_n363_), .D(ori_ori_n360_), .Y(ori6));
  NO2        o358(.A(ori_ori_n144_), .B(ori_ori_n245_), .Y(ori_ori_n381_));
  INV        o359(.A(ori_ori_n180_), .Y(ori_ori_n382_));
  OR2        o360(.A(ori_ori_n382_), .B(i_12_), .Y(ori_ori_n383_));
  INV        o361(.A(ori_ori_n179_), .Y(ori_ori_n384_));
  NA2        o362(.A(ori_ori_n71_), .B(ori_ori_n112_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n155_), .B(i_9_), .Y(ori_ori_n387_));
  NA2        o365(.A(ori_ori_n387_), .B(ori_ori_n376_), .Y(ori_ori_n388_));
  AOI210     o366(.A0(ori_ori_n388_), .A1(ori_ori_n258_), .B0(ori_ori_n134_), .Y(ori_ori_n389_));
  NAi32      o367(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n342_), .B(ori_ori_n390_), .Y(ori_ori_n391_));
  OR3        o369(.A(ori_ori_n391_), .B(ori_ori_n389_), .C(ori_ori_n386_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n330_), .B(i_2_), .Y(ori_ori_n393_));
  BUFFER     o371(.A(ori_ori_n288_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n394_), .B(ori_ori_n124_), .Y(ori_ori_n395_));
  AO210      o373(.A0(ori_ori_n251_), .A1(ori_ori_n359_), .B0(ori_ori_n36_), .Y(ori_ori_n396_));
  NA2        o374(.A(ori_ori_n396_), .B(ori_ori_n395_), .Y(ori_ori_n397_));
  NA2        o375(.A(ori_ori_n381_), .B(ori_ori_n338_), .Y(ori_ori_n398_));
  NA2        o376(.A(ori_ori_n398_), .B(ori_ori_n278_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n282_), .B(ori_ori_n94_), .Y(ori_ori_n400_));
  OAI210     o378(.A0(ori_ori_n400_), .A1(ori_ori_n102_), .B0(ori_ori_n211_), .Y(ori_ori_n401_));
  NA3        o379(.A(ori_ori_n480_), .B(ori_ori_n179_), .C(i_7_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n402_), .B(ori_ori_n401_), .Y(ori_ori_n403_));
  NO4        o381(.A(ori_ori_n403_), .B(ori_ori_n399_), .C(ori_ori_n397_), .D(ori_ori_n392_), .Y(ori_ori_n404_));
  NA3        o382(.A(ori_ori_n404_), .B(ori_ori_n383_), .C(ori_ori_n204_), .Y(ori3));
  NA2        o383(.A(i_12_), .B(i_10_), .Y(ori_ori_n406_));
  NO2        o384(.A(i_11_), .B(ori_ori_n147_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n278_), .B(ori_ori_n197_), .Y(ori_ori_n408_));
  NA2        o386(.A(ori_ori_n408_), .B(ori_ori_n40_), .Y(ori_ori_n409_));
  NOi21      o387(.An(ori_ori_n91_), .B(ori_ori_n25_), .Y(ori_ori_n410_));
  AN2        o388(.A(ori_ori_n228_), .B(ori_ori_n53_), .Y(ori_ori_n411_));
  NO2        o389(.A(ori_ori_n411_), .B(ori_ori_n410_), .Y(ori_ori_n412_));
  AOI210     o390(.A0(ori_ori_n412_), .A1(ori_ori_n409_), .B0(ori_ori_n47_), .Y(ori_ori_n413_));
  NO3        o391(.A(ori_ori_n206_), .B(ori_ori_n38_), .C(i_0_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n134_), .B(ori_ori_n267_), .Y(ori_ori_n415_));
  NOi21      o393(.An(ori_ori_n415_), .B(ori_ori_n414_), .Y(ori_ori_n416_));
  NO2        o394(.A(ori_ori_n416_), .B(ori_ori_n60_), .Y(ori_ori_n417_));
  NOi21      o395(.An(i_5_), .B(i_9_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n418_), .B(ori_ori_n225_), .Y(ori_ori_n419_));
  BUFFER     o397(.A(ori_ori_n169_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n420_), .B(ori_ori_n243_), .Y(ori_ori_n421_));
  NO2        o399(.A(ori_ori_n421_), .B(ori_ori_n419_), .Y(ori_ori_n422_));
  NO3        o400(.A(ori_ori_n422_), .B(ori_ori_n417_), .C(ori_ori_n413_), .Y(ori_ori_n423_));
  NO4        o401(.A(ori_ori_n268_), .B(i_12_), .C(ori_ori_n214_), .D(ori_ori_n212_), .Y(ori_ori_n424_));
  NA2        o402(.A(ori_ori_n424_), .B(i_11_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n157_), .B(ori_ori_n126_), .Y(ori_ori_n426_));
  NA2        o404(.A(i_0_), .B(i_10_), .Y(ori_ori_n427_));
  AN2        o405(.A(ori_ori_n426_), .B(i_6_), .Y(ori_ori_n428_));
  INV        o406(.A(ori_ori_n428_), .Y(ori_ori_n429_));
  NA2        o407(.A(ori_ori_n429_), .B(ori_ori_n425_), .Y(ori_ori_n430_));
  NA2        o408(.A(i_11_), .B(i_9_), .Y(ori_ori_n431_));
  NO3        o409(.A(i_12_), .B(ori_ori_n431_), .C(ori_ori_n277_), .Y(ori_ori_n432_));
  AN2        o410(.A(ori_ori_n432_), .B(i_5_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n209_), .B(ori_ori_n133_), .Y(ori_ori_n434_));
  INV        o412(.A(ori_ori_n434_), .Y(ori_ori_n435_));
  NO2        o413(.A(ori_ori_n431_), .B(ori_ori_n69_), .Y(ori_ori_n436_));
  INV        o414(.A(ori_ori_n210_), .Y(ori_ori_n437_));
  NO2        o415(.A(ori_ori_n437_), .B(ori_ori_n419_), .Y(ori_ori_n438_));
  NO3        o416(.A(ori_ori_n438_), .B(ori_ori_n435_), .C(ori_ori_n433_), .Y(ori_ori_n439_));
  INV        o417(.A(ori_ori_n439_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n406_), .B(ori_ori_n178_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n441_), .B(ori_ori_n436_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n259_), .B(ori_ori_n442_), .Y(ori_ori_n443_));
  NO3        o421(.A(ori_ori_n443_), .B(ori_ori_n440_), .C(ori_ori_n430_), .Y(ori_ori_n444_));
  NO3        o422(.A(ori_ori_n427_), .B(ori_ori_n418_), .C(ori_ori_n136_), .Y(ori_ori_n445_));
  AOI220     o423(.A0(ori_ori_n445_), .A1(i_11_), .B0(ori_ori_n266_), .B1(ori_ori_n71_), .Y(ori_ori_n446_));
  NO3        o424(.A(ori_ori_n142_), .B(ori_ori_n206_), .C(i_0_), .Y(ori_ori_n447_));
  OAI210     o425(.A0(ori_ori_n447_), .A1(ori_ori_n72_), .B0(i_13_), .Y(ori_ori_n448_));
  NA2        o426(.A(ori_ori_n448_), .B(ori_ori_n446_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n250_), .B(ori_ori_n244_), .Y(ori_ori_n450_));
  INV        o428(.A(ori_ori_n450_), .Y(ori_ori_n451_));
  NA3        o429(.A(ori_ori_n208_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n452_));
  INV        o430(.A(ori_ori_n452_), .Y(ori_ori_n453_));
  NO3        o431(.A(ori_ori_n431_), .B(ori_ori_n143_), .C(ori_ori_n136_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n454_), .B(ori_ori_n453_), .Y(ori_ori_n455_));
  NA2        o433(.A(ori_ori_n455_), .B(ori_ori_n451_), .Y(ori_ori_n456_));
  NO2        o434(.A(ori_ori_n80_), .B(i_5_), .Y(ori_ori_n457_));
  NA2        o435(.A(ori_ori_n407_), .B(ori_ori_n101_), .Y(ori_ori_n458_));
  INV        o436(.A(ori_ori_n458_), .Y(ori_ori_n459_));
  NA2        o437(.A(ori_ori_n459_), .B(ori_ori_n457_), .Y(ori_ori_n460_));
  NAi21      o438(.An(ori_ori_n151_), .B(ori_ori_n152_), .Y(ori_ori_n461_));
  NO4        o439(.A(ori_ori_n150_), .B(ori_ori_n142_), .C(i_0_), .D(i_12_), .Y(ori_ori_n462_));
  NA2        o440(.A(ori_ori_n462_), .B(ori_ori_n461_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n463_), .B(ori_ori_n460_), .Y(ori_ori_n464_));
  NO3        o442(.A(ori_ori_n464_), .B(ori_ori_n456_), .C(ori_ori_n449_), .Y(ori_ori_n465_));
  NA2        o443(.A(ori_ori_n393_), .B(ori_ori_n37_), .Y(ori_ori_n466_));
  NA2        o444(.A(ori_ori_n466_), .B(ori_ori_n281_), .Y(ori_ori_n467_));
  NA2        o445(.A(ori_ori_n467_), .B(ori_ori_n141_), .Y(ori_ori_n468_));
  NA2        o446(.A(i_2_), .B(i_10_), .Y(ori_ori_n469_));
  NO2        o447(.A(ori_ori_n66_), .B(ori_ori_n469_), .Y(ori_ori_n470_));
  AOI210     o448(.A0(ori_ori_n470_), .A1(ori_ori_n47_), .B0(ori_ori_n424_), .Y(ori_ori_n471_));
  AOI210     o449(.A0(ori_ori_n471_), .A1(ori_ori_n468_), .B0(ori_ori_n69_), .Y(ori_ori_n472_));
  INV        o450(.A(ori_ori_n203_), .Y(ori_ori_n473_));
  NO2        o451(.A(ori_ori_n473_), .B(i_13_), .Y(ori_ori_n474_));
  NO2        o452(.A(ori_ori_n474_), .B(ori_ori_n472_), .Y(ori_ori_n475_));
  NA4        o453(.A(ori_ori_n475_), .B(ori_ori_n465_), .C(ori_ori_n444_), .D(ori_ori_n423_), .Y(ori4));
  INV        o454(.A(i_6_), .Y(ori_ori_n479_));
  INV        o455(.A(ori_ori_n268_), .Y(ori_ori_n480_));
  INV        o456(.A(i_1_), .Y(ori_ori_n481_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_0_), .B(i_2_), .Y(mai_mai_n51_));
  NA3        m029(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n52_));
  NO2        m030(.A(i_1_), .B(i_6_), .Y(mai_mai_n53_));
  NA2        m031(.A(i_8_), .B(i_7_), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n53_), .B0(mai_mai_n52_), .Y(mai_mai_n55_));
  NA2        m033(.A(mai_mai_n55_), .B(i_12_), .Y(mai_mai_n56_));
  INV        m034(.A(i_1_), .Y(mai_mai_n57_));
  NA2        m035(.A(i_1_), .B(i_10_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(i_6_), .Y(mai_mai_n59_));
  NAi31      m037(.An(mai_mai_n59_), .B(mai_mai_n946_), .C(mai_mai_n56_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n61_));
  AOI210     m039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_1_), .B(i_6_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(mai_mai_n25_), .Y(mai_mai_n64_));
  INV        m042(.A(i_0_), .Y(mai_mai_n65_));
  NAi21      m043(.An(i_5_), .B(i_10_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_5_), .B(i_9_), .Y(mai_mai_n67_));
  AOI210     m045(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n64_), .Y(mai_mai_n69_));
  INV        m047(.A(mai_mai_n69_), .Y(mai_mai_n70_));
  OAI210     m048(.A0(mai_mai_n70_), .A1(mai_mai_n60_), .B0(i_0_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_12_), .B(i_5_), .Y(mai_mai_n72_));
  NA2        m050(.A(i_2_), .B(i_8_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n53_), .Y(mai_mai_n74_));
  NO2        m052(.A(i_3_), .B(i_9_), .Y(mai_mai_n75_));
  NO2        m053(.A(i_3_), .B(i_7_), .Y(mai_mai_n76_));
  INV        m054(.A(i_6_), .Y(mai_mai_n77_));
  OR4        m055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n78_));
  INV        m056(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_2_), .B(i_7_), .Y(mai_mai_n80_));
  NAi21      m058(.An(i_6_), .B(i_10_), .Y(mai_mai_n81_));
  NA2        m059(.A(i_6_), .B(i_9_), .Y(mai_mai_n82_));
  AOI210     m060(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n57_), .Y(mai_mai_n83_));
  NA2        m061(.A(i_2_), .B(i_6_), .Y(mai_mai_n84_));
  INV        m062(.A(mai_mai_n83_), .Y(mai_mai_n85_));
  AOI210     m063(.A0(mai_mai_n85_), .A1(mai_mai_n936_), .B0(mai_mai_n72_), .Y(mai_mai_n86_));
  AN3        m064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n87_));
  NAi21      m065(.An(i_6_), .B(i_11_), .Y(mai_mai_n88_));
  NO2        m066(.A(i_5_), .B(i_8_), .Y(mai_mai_n89_));
  NOi21      m067(.An(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n90_));
  AOI210     m068(.A0(mai_mai_n87_), .A1(mai_mai_n32_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  INV        m069(.A(i_7_), .Y(mai_mai_n92_));
  NA2        m070(.A(mai_mai_n46_), .B(mai_mai_n92_), .Y(mai_mai_n93_));
  NO2        m071(.A(i_0_), .B(i_5_), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n94_), .B(mai_mai_n77_), .Y(mai_mai_n95_));
  NA2        m073(.A(i_12_), .B(i_3_), .Y(mai_mai_n96_));
  INV        m074(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NA3        m075(.A(mai_mai_n97_), .B(mai_mai_n95_), .C(mai_mai_n93_), .Y(mai_mai_n98_));
  NAi21      m076(.An(i_7_), .B(i_11_), .Y(mai_mai_n99_));
  NO3        m077(.A(mai_mai_n99_), .B(mai_mai_n81_), .C(mai_mai_n51_), .Y(mai_mai_n100_));
  AN2        m078(.A(i_2_), .B(i_10_), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n101_), .B(i_7_), .Y(mai_mai_n102_));
  OR2        m080(.A(mai_mai_n72_), .B(mai_mai_n53_), .Y(mai_mai_n103_));
  NO2        m081(.A(i_8_), .B(mai_mai_n92_), .Y(mai_mai_n104_));
  NO3        m082(.A(mai_mai_n104_), .B(mai_mai_n103_), .C(mai_mai_n102_), .Y(mai_mai_n105_));
  NA2        m083(.A(i_12_), .B(i_7_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n57_), .B(mai_mai_n26_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n107_), .B(i_0_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_11_), .B(i_12_), .Y(mai_mai_n109_));
  OAI210     m087(.A0(mai_mai_n108_), .A1(mai_mai_n106_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n110_), .B(mai_mai_n105_), .Y(mai_mai_n111_));
  NAi41      m089(.An(mai_mai_n100_), .B(mai_mai_n111_), .C(mai_mai_n98_), .D(mai_mai_n91_), .Y(mai_mai_n112_));
  NOi21      m090(.An(i_1_), .B(i_5_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n113_), .B(i_11_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n92_), .B(mai_mai_n37_), .Y(mai_mai_n115_));
  NA2        m093(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n117_), .B(mai_mai_n46_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n119_));
  NAi21      m097(.An(i_3_), .B(i_8_), .Y(mai_mai_n120_));
  INV        m098(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NOi21      m099(.An(mai_mai_n121_), .B(mai_mai_n119_), .Y(mai_mai_n122_));
  NO2        m100(.A(i_1_), .B(mai_mai_n77_), .Y(mai_mai_n123_));
  NO2        m101(.A(i_6_), .B(i_5_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(i_3_), .Y(mai_mai_n125_));
  AO210      m103(.A0(mai_mai_n125_), .A1(mai_mai_n47_), .B0(mai_mai_n123_), .Y(mai_mai_n126_));
  OAI220     m104(.A0(mai_mai_n126_), .A1(mai_mai_n99_), .B0(mai_mai_n122_), .B1(mai_mai_n114_), .Y(mai_mai_n127_));
  NO3        m105(.A(mai_mai_n127_), .B(mai_mai_n112_), .C(mai_mai_n86_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n71_), .Y(mai2));
  NO2        m107(.A(mai_mai_n57_), .B(mai_mai_n37_), .Y(mai_mai_n130_));
  NA2        m108(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(mai_mai_n130_), .Y(mai_mai_n132_));
  NA4        m110(.A(mai_mai_n132_), .B(mai_mai_n69_), .C(mai_mai_n61_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m111(.A(i_8_), .B(i_7_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n134_), .B(i_6_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_12_), .B(i_13_), .Y(mai_mai_n136_));
  NAi21      m114(.An(i_5_), .B(i_11_), .Y(mai_mai_n137_));
  NOi21      m115(.An(mai_mai_n136_), .B(mai_mai_n137_), .Y(mai_mai_n138_));
  NO2        m116(.A(i_0_), .B(i_1_), .Y(mai_mai_n139_));
  NA2        m117(.A(i_2_), .B(i_3_), .Y(mai_mai_n140_));
  NO2        m118(.A(mai_mai_n140_), .B(i_4_), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n141_), .B(mai_mai_n138_), .Y(mai_mai_n142_));
  AN2        m120(.A(mai_mai_n136_), .B(mai_mai_n75_), .Y(mai_mai_n143_));
  NA2        m121(.A(i_1_), .B(i_5_), .Y(mai_mai_n144_));
  NA2        m122(.A(i_0_), .B(mai_mai_n36_), .Y(mai_mai_n145_));
  NO3        m123(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(i_13_), .Y(mai_mai_n146_));
  OR2        m124(.A(i_0_), .B(i_1_), .Y(mai_mai_n147_));
  NO3        m125(.A(mai_mai_n147_), .B(mai_mai_n72_), .C(i_13_), .Y(mai_mai_n148_));
  NAi32      m126(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n149_));
  NAi21      m127(.An(mai_mai_n149_), .B(mai_mai_n148_), .Y(mai_mai_n150_));
  NOi21      m128(.An(i_4_), .B(i_10_), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n151_), .B(mai_mai_n40_), .Y(mai_mai_n152_));
  NO2        m130(.A(i_3_), .B(i_5_), .Y(mai_mai_n153_));
  NO3        m131(.A(mai_mai_n65_), .B(i_2_), .C(i_1_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  OAI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n152_), .B0(mai_mai_n150_), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n156_), .B(mai_mai_n146_), .Y(mai_mai_n157_));
  AOI210     m135(.A0(mai_mai_n157_), .A1(mai_mai_n142_), .B0(mai_mai_n135_), .Y(mai_mai_n158_));
  NA3        m136(.A(mai_mai_n65_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n159_));
  NA2        m137(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n160_));
  NOi21      m138(.An(i_4_), .B(i_9_), .Y(mai_mai_n161_));
  NOi21      m139(.An(i_11_), .B(i_13_), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  OR2        m141(.A(mai_mai_n163_), .B(mai_mai_n160_), .Y(mai_mai_n164_));
  NO2        m142(.A(i_4_), .B(i_5_), .Y(mai_mai_n165_));
  NAi21      m143(.An(i_12_), .B(i_11_), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n166_), .B(i_13_), .Y(mai_mai_n167_));
  NA3        m145(.A(mai_mai_n167_), .B(mai_mai_n165_), .C(mai_mai_n75_), .Y(mai_mai_n168_));
  AOI210     m146(.A0(mai_mai_n168_), .A1(mai_mai_n164_), .B0(mai_mai_n159_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n65_), .B(mai_mai_n57_), .Y(mai_mai_n170_));
  NA2        m148(.A(mai_mai_n170_), .B(mai_mai_n46_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n172_));
  NAi31      m150(.An(mai_mai_n172_), .B(mai_mai_n143_), .C(i_11_), .Y(mai_mai_n173_));
  NA2        m151(.A(i_3_), .B(i_5_), .Y(mai_mai_n174_));
  OR2        m152(.A(mai_mai_n174_), .B(mai_mai_n163_), .Y(mai_mai_n175_));
  AOI210     m153(.A0(mai_mai_n175_), .A1(mai_mai_n173_), .B0(mai_mai_n171_), .Y(mai_mai_n176_));
  NO2        m154(.A(mai_mai_n65_), .B(i_5_), .Y(mai_mai_n177_));
  NO2        m155(.A(i_13_), .B(i_10_), .Y(mai_mai_n178_));
  NA3        m156(.A(mai_mai_n178_), .B(mai_mai_n177_), .C(mai_mai_n44_), .Y(mai_mai_n179_));
  NO2        m157(.A(i_2_), .B(i_1_), .Y(mai_mai_n180_));
  NAi21      m158(.An(i_4_), .B(i_12_), .Y(mai_mai_n181_));
  NO3        m159(.A(mai_mai_n181_), .B(mai_mai_n944_), .C(mai_mai_n179_), .Y(mai_mai_n182_));
  NO3        m160(.A(mai_mai_n182_), .B(mai_mai_n176_), .C(mai_mai_n169_), .Y(mai_mai_n183_));
  INV        m161(.A(i_8_), .Y(mai_mai_n184_));
  INV        m162(.A(i_6_), .Y(mai_mai_n185_));
  NO3        m163(.A(i_3_), .B(mai_mai_n77_), .C(mai_mai_n48_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n186_), .B(mai_mai_n104_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n188_));
  NA3        m166(.A(mai_mai_n188_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n189_));
  NO3        m167(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n190_));
  NO2        m168(.A(i_13_), .B(mai_mai_n187_), .Y(mai_mai_n191_));
  NO2        m169(.A(i_3_), .B(i_8_), .Y(mai_mai_n192_));
  NO3        m170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n193_));
  NA3        m171(.A(mai_mai_n193_), .B(mai_mai_n192_), .C(mai_mai_n40_), .Y(mai_mai_n194_));
  NO2        m172(.A(i_13_), .B(i_9_), .Y(mai_mai_n195_));
  NAi21      m173(.An(i_12_), .B(i_3_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n197_));
  NO3        m175(.A(i_0_), .B(i_2_), .C(mai_mai_n57_), .Y(mai_mai_n198_));
  NA3        m176(.A(mai_mai_n198_), .B(mai_mai_n197_), .C(i_10_), .Y(mai_mai_n199_));
  OAI220     m177(.A0(mai_mai_n199_), .A1(i_13_), .B0(mai_mai_n53_), .B1(mai_mai_n194_), .Y(mai_mai_n200_));
  AOI210     m178(.A0(mai_mai_n200_), .A1(i_7_), .B0(mai_mai_n191_), .Y(mai_mai_n201_));
  OAI220     m179(.A0(mai_mai_n201_), .A1(i_4_), .B0(mai_mai_n185_), .B1(mai_mai_n183_), .Y(mai_mai_n202_));
  NA3        m180(.A(i_13_), .B(mai_mai_n184_), .C(i_10_), .Y(mai_mai_n203_));
  NO2        m181(.A(mai_mai_n203_), .B(i_12_), .Y(mai_mai_n204_));
  NA2        m182(.A(i_0_), .B(i_5_), .Y(mai_mai_n205_));
  NAi31      m183(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n206_));
  NO2        m184(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n46_), .B(mai_mai_n57_), .Y(mai_mai_n208_));
  NA3        m186(.A(mai_mai_n208_), .B(i_3_), .C(mai_mai_n207_), .Y(mai_mai_n209_));
  INV        m187(.A(i_13_), .Y(mai_mai_n210_));
  NO2        m188(.A(i_12_), .B(mai_mai_n210_), .Y(mai_mai_n211_));
  NA3        m189(.A(mai_mai_n211_), .B(mai_mai_n188_), .C(mai_mai_n186_), .Y(mai_mai_n212_));
  OAI210     m190(.A0(mai_mai_n209_), .A1(mai_mai_n206_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  AOI220     m191(.A0(mai_mai_n213_), .A1(mai_mai_n134_), .B0(i_3_), .B1(mai_mai_n204_), .Y(mai_mai_n214_));
  NO2        m192(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n174_), .B(i_4_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  OR2        m195(.A(i_8_), .B(i_7_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n218_), .B(mai_mai_n77_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n51_), .B(i_1_), .Y(mai_mai_n220_));
  INV        m198(.A(i_12_), .Y(mai_mai_n221_));
  NO3        m199(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n222_));
  NA2        m200(.A(i_2_), .B(i_1_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n51_), .B(mai_mai_n217_), .Y(mai_mai_n224_));
  NO3        m202(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n225_));
  NAi21      m203(.An(i_4_), .B(i_3_), .Y(mai_mai_n226_));
  NO2        m204(.A(i_0_), .B(i_6_), .Y(mai_mai_n227_));
  NOi41      m205(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n228_));
  NA2        m206(.A(mai_mai_n228_), .B(mai_mai_n227_), .Y(mai_mai_n229_));
  AOI210     m207(.A0(mai_mai_n940_), .A1(mai_mai_n40_), .B0(mai_mai_n224_), .Y(mai_mai_n230_));
  NO2        m208(.A(i_11_), .B(mai_mai_n210_), .Y(mai_mai_n231_));
  NOi21      m209(.An(i_1_), .B(i_6_), .Y(mai_mai_n232_));
  NAi21      m210(.An(i_3_), .B(i_7_), .Y(mai_mai_n233_));
  NO2        m211(.A(i_12_), .B(i_3_), .Y(mai_mai_n234_));
  NA3        m212(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n135_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n221_), .B(i_13_), .Y(mai_mai_n237_));
  NO2        m215(.A(mai_mai_n237_), .B(mai_mai_n67_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n238_), .B(mai_mai_n236_), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n218_), .B(mai_mai_n37_), .Y(mai_mai_n240_));
  NA2        m218(.A(i_12_), .B(i_6_), .Y(mai_mai_n241_));
  OR2        m219(.A(i_13_), .B(i_9_), .Y(mai_mai_n242_));
  NO3        m220(.A(mai_mai_n242_), .B(mai_mai_n241_), .C(mai_mai_n48_), .Y(mai_mai_n243_));
  NO2        m221(.A(mai_mai_n226_), .B(i_2_), .Y(mai_mai_n244_));
  NA3        m222(.A(mai_mai_n244_), .B(mai_mai_n243_), .C(mai_mai_n44_), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n231_), .B(i_9_), .Y(mai_mai_n246_));
  OAI210     m224(.A0(mai_mai_n57_), .A1(mai_mai_n246_), .B0(mai_mai_n245_), .Y(mai_mai_n247_));
  NO3        m225(.A(i_11_), .B(mai_mai_n210_), .C(mai_mai_n25_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n233_), .B(i_8_), .Y(mai_mai_n249_));
  NO2        m227(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n250_));
  NA2        m228(.A(mai_mai_n247_), .B(mai_mai_n240_), .Y(mai_mai_n251_));
  NA4        m229(.A(mai_mai_n251_), .B(mai_mai_n239_), .C(mai_mai_n230_), .D(mai_mai_n214_), .Y(mai_mai_n252_));
  NO3        m230(.A(i_12_), .B(mai_mai_n210_), .C(mai_mai_n37_), .Y(mai_mai_n253_));
  INV        m231(.A(mai_mai_n253_), .Y(mai_mai_n254_));
  NA2        m232(.A(i_8_), .B(mai_mai_n92_), .Y(mai_mai_n255_));
  NO3        m233(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n256_));
  NO2        m234(.A(mai_mai_n223_), .B(i_0_), .Y(mai_mai_n257_));
  NA2        m235(.A(mai_mai_n250_), .B(mai_mai_n26_), .Y(mai_mai_n258_));
  NO2        m236(.A(mai_mai_n258_), .B(mai_mai_n941_), .Y(mai_mai_n259_));
  NA2        m237(.A(i_0_), .B(i_1_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n260_), .B(i_2_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n54_), .B(i_6_), .Y(mai_mai_n262_));
  NA2        m240(.A(mai_mai_n262_), .B(mai_mai_n261_), .Y(mai_mai_n263_));
  OAI210     m241(.A0(mai_mai_n155_), .A1(mai_mai_n135_), .B0(mai_mai_n263_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n264_), .B(mai_mai_n259_), .Y(mai_mai_n265_));
  NO2        m243(.A(i_3_), .B(i_10_), .Y(mai_mai_n266_));
  NA3        m244(.A(mai_mai_n266_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n267_));
  NO2        m245(.A(i_2_), .B(mai_mai_n92_), .Y(mai_mai_n268_));
  NA2        m246(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n269_), .B(i_8_), .Y(mai_mai_n270_));
  NA2        m248(.A(mai_mai_n270_), .B(mai_mai_n268_), .Y(mai_mai_n271_));
  AN2        m249(.A(i_3_), .B(i_10_), .Y(mai_mai_n272_));
  NA3        m250(.A(mai_mai_n272_), .B(mai_mai_n167_), .C(mai_mai_n165_), .Y(mai_mai_n273_));
  NO2        m251(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n275_));
  OR2        m253(.A(mai_mai_n271_), .B(mai_mai_n267_), .Y(mai_mai_n276_));
  OAI220     m254(.A0(mai_mai_n276_), .A1(i_6_), .B0(mai_mai_n265_), .B1(mai_mai_n254_), .Y(mai_mai_n277_));
  NO4        m255(.A(mai_mai_n277_), .B(mai_mai_n252_), .C(mai_mai_n202_), .D(mai_mai_n158_), .Y(mai_mai_n278_));
  NO3        m256(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n279_));
  NO3        m257(.A(i_6_), .B(mai_mai_n184_), .C(i_7_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n280_), .B(mai_mai_n188_), .Y(mai_mai_n281_));
  AOI210     m259(.A0(mai_mai_n281_), .A1(mai_mai_n223_), .B0(mai_mai_n160_), .Y(mai_mai_n282_));
  NO2        m260(.A(i_2_), .B(i_3_), .Y(mai_mai_n283_));
  OR2        m261(.A(i_0_), .B(i_5_), .Y(mai_mai_n284_));
  NA3        m262(.A(mai_mai_n219_), .B(mai_mai_n283_), .C(i_1_), .Y(mai_mai_n285_));
  NA2        m263(.A(mai_mai_n257_), .B(mai_mai_n104_), .Y(mai_mai_n286_));
  NAi21      m264(.An(i_8_), .B(i_7_), .Y(mai_mai_n287_));
  NO2        m265(.A(mai_mai_n287_), .B(i_6_), .Y(mai_mai_n288_));
  NO2        m266(.A(mai_mai_n147_), .B(mai_mai_n46_), .Y(mai_mai_n289_));
  NA2        m267(.A(mai_mai_n289_), .B(mai_mai_n288_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n290_), .B(mai_mai_n286_), .C(mai_mai_n285_), .Y(mai_mai_n291_));
  OAI210     m269(.A0(mai_mai_n291_), .A1(mai_mai_n282_), .B0(i_4_), .Y(mai_mai_n292_));
  NO2        m270(.A(i_12_), .B(i_10_), .Y(mai_mai_n293_));
  NOi21      m271(.An(i_5_), .B(i_0_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n269_), .B(mai_mai_n120_), .Y(mai_mai_n295_));
  NA4        m273(.A(mai_mai_n76_), .B(mai_mai_n36_), .C(mai_mai_n77_), .D(i_8_), .Y(mai_mai_n296_));
  NA2        m274(.A(mai_mai_n295_), .B(mai_mai_n293_), .Y(mai_mai_n297_));
  NO2        m275(.A(i_6_), .B(i_8_), .Y(mai_mai_n298_));
  NOi21      m276(.An(i_0_), .B(i_2_), .Y(mai_mai_n299_));
  AN2        m277(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n300_));
  NO2        m278(.A(i_1_), .B(i_7_), .Y(mai_mai_n301_));
  AO220      m279(.A0(mai_mai_n301_), .A1(mai_mai_n300_), .B0(mai_mai_n288_), .B1(mai_mai_n220_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n302_), .B(i_4_), .Y(mai_mai_n303_));
  NA3        m281(.A(mai_mai_n303_), .B(mai_mai_n297_), .C(mai_mai_n292_), .Y(mai_mai_n304_));
  NO3        m282(.A(mai_mai_n218_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n305_));
  NO3        m283(.A(mai_mai_n287_), .B(i_2_), .C(i_1_), .Y(mai_mai_n306_));
  OAI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n305_), .B0(i_6_), .Y(mai_mai_n307_));
  NA2        m285(.A(mai_mai_n268_), .B(mai_mai_n184_), .Y(mai_mai_n308_));
  NA2        m286(.A(mai_mai_n308_), .B(mai_mai_n307_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n309_), .B(i_3_), .Y(mai_mai_n310_));
  INV        m288(.A(mai_mai_n76_), .Y(mai_mai_n311_));
  NO2        m289(.A(mai_mai_n84_), .B(mai_mai_n184_), .Y(mai_mai_n312_));
  NO2        m290(.A(mai_mai_n73_), .B(mai_mai_n311_), .Y(mai_mai_n313_));
  NO2        m291(.A(mai_mai_n184_), .B(i_9_), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n314_), .B(i_0_), .Y(mai_mai_n315_));
  NO2        m293(.A(mai_mai_n313_), .B(mai_mai_n259_), .Y(mai_mai_n316_));
  AOI210     m294(.A0(mai_mai_n316_), .A1(mai_mai_n310_), .B0(mai_mai_n152_), .Y(mai_mai_n317_));
  AOI210     m295(.A0(mai_mai_n304_), .A1(mai_mai_n279_), .B0(mai_mai_n317_), .Y(mai_mai_n318_));
  NOi32      m296(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n319_));
  INV        m297(.A(mai_mai_n319_), .Y(mai_mai_n320_));
  NAi21      m298(.An(i_0_), .B(i_6_), .Y(mai_mai_n321_));
  NAi21      m299(.An(i_1_), .B(i_5_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n322_), .B(mai_mai_n321_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n323_), .B(mai_mai_n25_), .Y(mai_mai_n324_));
  OAI210     m302(.A0(mai_mai_n324_), .A1(mai_mai_n149_), .B0(mai_mai_n229_), .Y(mai_mai_n325_));
  NAi41      m303(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n326_));
  OAI220     m304(.A0(mai_mai_n326_), .A1(mai_mai_n322_), .B0(mai_mai_n206_), .B1(mai_mai_n149_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n326_), .A1(mai_mai_n149_), .B0(mai_mai_n147_), .Y(mai_mai_n328_));
  NOi32      m306(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n329_));
  NAi21      m307(.An(i_6_), .B(i_1_), .Y(mai_mai_n330_));
  NA3        m308(.A(mai_mai_n330_), .B(mai_mai_n329_), .C(mai_mai_n46_), .Y(mai_mai_n331_));
  NO2        m309(.A(mai_mai_n331_), .B(i_0_), .Y(mai_mai_n332_));
  OR3        m310(.A(mai_mai_n332_), .B(mai_mai_n328_), .C(mai_mai_n327_), .Y(mai_mai_n333_));
  NO2        m311(.A(i_1_), .B(mai_mai_n92_), .Y(mai_mai_n334_));
  NAi21      m312(.An(i_3_), .B(i_4_), .Y(mai_mai_n335_));
  NO2        m313(.A(mai_mai_n335_), .B(i_9_), .Y(mai_mai_n336_));
  AN2        m314(.A(i_6_), .B(i_7_), .Y(mai_mai_n337_));
  NA2        m315(.A(i_2_), .B(i_7_), .Y(mai_mai_n338_));
  NO2        m316(.A(mai_mai_n335_), .B(i_10_), .Y(mai_mai_n339_));
  NA3        m317(.A(mai_mai_n339_), .B(mai_mai_n338_), .C(mai_mai_n227_), .Y(mai_mai_n340_));
  INV        m318(.A(mai_mai_n340_), .Y(mai_mai_n341_));
  AOI210     m319(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n342_));
  OAI210     m320(.A0(mai_mai_n342_), .A1(mai_mai_n180_), .B0(mai_mai_n339_), .Y(mai_mai_n343_));
  AOI220     m321(.A0(mai_mai_n339_), .A1(mai_mai_n301_), .B0(mai_mai_n222_), .B1(mai_mai_n180_), .Y(mai_mai_n344_));
  AOI210     m322(.A0(mai_mai_n344_), .A1(mai_mai_n343_), .B0(i_5_), .Y(mai_mai_n345_));
  NO4        m323(.A(mai_mai_n345_), .B(mai_mai_n341_), .C(mai_mai_n333_), .D(mai_mai_n325_), .Y(mai_mai_n346_));
  NO2        m324(.A(mai_mai_n346_), .B(mai_mai_n320_), .Y(mai_mai_n347_));
  NO2        m325(.A(mai_mai_n54_), .B(mai_mai_n25_), .Y(mai_mai_n348_));
  AN2        m326(.A(i_12_), .B(i_5_), .Y(mai_mai_n349_));
  NO2        m327(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n350_));
  NA2        m328(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n351_));
  NO2        m329(.A(i_11_), .B(i_6_), .Y(mai_mai_n352_));
  NA2        m330(.A(mai_mai_n352_), .B(mai_mai_n289_), .Y(mai_mai_n353_));
  NO2        m331(.A(mai_mai_n353_), .B(mai_mai_n351_), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n226_), .B(i_5_), .Y(mai_mai_n355_));
  NO2        m333(.A(i_5_), .B(i_10_), .Y(mai_mai_n356_));
  NA2        m334(.A(mai_mai_n136_), .B(mai_mai_n45_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n357_), .B(mai_mai_n226_), .Y(mai_mai_n358_));
  OAI210     m336(.A0(mai_mai_n358_), .A1(mai_mai_n354_), .B0(mai_mai_n348_), .Y(mai_mai_n359_));
  NO2        m337(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n360_));
  NA2        m338(.A(mai_mai_n354_), .B(mai_mai_n360_), .Y(mai_mai_n361_));
  NO3        m339(.A(mai_mai_n77_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n362_));
  NO2        m340(.A(i_11_), .B(i_12_), .Y(mai_mai_n363_));
  NA2        m341(.A(mai_mai_n356_), .B(mai_mai_n221_), .Y(mai_mai_n364_));
  NA2        m342(.A(mai_mai_n104_), .B(i_4_), .Y(mai_mai_n365_));
  OAI220     m343(.A0(mai_mai_n365_), .A1(mai_mai_n206_), .B0(mai_mai_n364_), .B1(mai_mai_n296_), .Y(mai_mai_n366_));
  NAi21      m344(.An(i_13_), .B(i_0_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n367_), .B(mai_mai_n223_), .Y(mai_mai_n368_));
  NA2        m346(.A(mai_mai_n366_), .B(mai_mai_n368_), .Y(mai_mai_n369_));
  NA3        m347(.A(mai_mai_n369_), .B(mai_mai_n361_), .C(mai_mai_n359_), .Y(mai_mai_n370_));
  NO2        m348(.A(i_0_), .B(i_11_), .Y(mai_mai_n371_));
  AN2        m349(.A(i_1_), .B(i_6_), .Y(mai_mai_n372_));
  NOi21      m350(.An(i_2_), .B(i_12_), .Y(mai_mai_n373_));
  NA2        m351(.A(mai_mai_n373_), .B(mai_mai_n372_), .Y(mai_mai_n374_));
  INV        m352(.A(mai_mai_n374_), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n134_), .B(i_9_), .Y(mai_mai_n376_));
  NO2        m354(.A(mai_mai_n376_), .B(i_4_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n375_), .B(mai_mai_n377_), .Y(mai_mai_n378_));
  OR2        m356(.A(i_13_), .B(i_10_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n163_), .B(mai_mai_n115_), .Y(mai_mai_n380_));
  NO2        m358(.A(mai_mai_n92_), .B(mai_mai_n25_), .Y(mai_mai_n381_));
  INV        m359(.A(mai_mai_n285_), .Y(mai_mai_n382_));
  AOI220     m360(.A0(mai_mai_n262_), .A1(mai_mai_n256_), .B0(mai_mai_n257_), .B1(i_8_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n383_), .B(mai_mai_n160_), .Y(mai_mai_n384_));
  NO2        m362(.A(i_2_), .B(mai_mai_n255_), .Y(mai_mai_n385_));
  NO3        m363(.A(mai_mai_n385_), .B(mai_mai_n384_), .C(mai_mai_n382_), .Y(mai_mai_n386_));
  NO2        m364(.A(i_3_), .B(mai_mai_n287_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n262_), .B(mai_mai_n220_), .Y(mai_mai_n388_));
  NO2        m366(.A(mai_mai_n388_), .B(mai_mai_n174_), .Y(mai_mai_n389_));
  NA3        m367(.A(mai_mai_n301_), .B(mai_mai_n300_), .C(i_5_), .Y(mai_mai_n390_));
  INV        m368(.A(mai_mai_n390_), .Y(mai_mai_n391_));
  NO3        m369(.A(mai_mai_n391_), .B(mai_mai_n389_), .C(mai_mai_n387_), .Y(mai_mai_n392_));
  AOI210     m370(.A0(mai_mai_n392_), .A1(mai_mai_n386_), .B0(mai_mai_n246_), .Y(mai_mai_n393_));
  NO4        m371(.A(mai_mai_n393_), .B(mai_mai_n943_), .C(mai_mai_n370_), .D(mai_mai_n347_), .Y(mai_mai_n394_));
  NO2        m372(.A(mai_mai_n57_), .B(i_4_), .Y(mai_mai_n395_));
  NO2        m373(.A(mai_mai_n65_), .B(i_13_), .Y(mai_mai_n396_));
  NA3        m374(.A(mai_mai_n396_), .B(mai_mai_n395_), .C(i_2_), .Y(mai_mai_n397_));
  NO2        m375(.A(i_10_), .B(i_9_), .Y(mai_mai_n398_));
  NAi21      m376(.An(i_12_), .B(i_8_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n399_), .B(i_3_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n400_), .B(mai_mai_n398_), .Y(mai_mai_n401_));
  NA2        m379(.A(i_2_), .B(mai_mai_n95_), .Y(mai_mai_n402_));
  OAI220     m380(.A0(mai_mai_n402_), .A1(mai_mai_n194_), .B0(mai_mai_n401_), .B1(mai_mai_n397_), .Y(mai_mai_n403_));
  NA2        m381(.A(mai_mai_n275_), .B(i_0_), .Y(mai_mai_n404_));
  NO3        m382(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n405_));
  NA2        m383(.A(mai_mai_n241_), .B(mai_mai_n88_), .Y(mai_mai_n406_));
  NA2        m384(.A(mai_mai_n406_), .B(mai_mai_n405_), .Y(mai_mai_n407_));
  NA2        m385(.A(i_8_), .B(i_9_), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n407_), .B(mai_mai_n404_), .Y(mai_mai_n409_));
  NA2        m387(.A(mai_mai_n231_), .B(mai_mai_n274_), .Y(mai_mai_n410_));
  NO3        m388(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n411_));
  INV        m389(.A(mai_mai_n411_), .Y(mai_mai_n412_));
  NA3        m390(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n413_));
  NA4        m391(.A(mai_mai_n137_), .B(mai_mai_n107_), .C(mai_mai_n72_), .D(mai_mai_n23_), .Y(mai_mai_n414_));
  OAI220     m392(.A0(mai_mai_n414_), .A1(mai_mai_n413_), .B0(mai_mai_n412_), .B1(mai_mai_n410_), .Y(mai_mai_n415_));
  NO3        m393(.A(mai_mai_n415_), .B(mai_mai_n409_), .C(mai_mai_n403_), .Y(mai_mai_n416_));
  OR2        m394(.A(mai_mai_n260_), .B(i_13_), .Y(mai_mai_n417_));
  OA210      m395(.A0(mai_mai_n315_), .A1(mai_mai_n92_), .B0(mai_mai_n263_), .Y(mai_mai_n418_));
  OA220      m396(.A0(mai_mai_n418_), .A1(mai_mai_n152_), .B0(mai_mai_n417_), .B1(mai_mai_n217_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n87_), .B(i_13_), .Y(mai_mai_n420_));
  NA2        m398(.A(i_3_), .B(mai_mai_n348_), .Y(mai_mai_n421_));
  NO2        m399(.A(i_2_), .B(i_13_), .Y(mai_mai_n422_));
  NA3        m400(.A(mai_mai_n422_), .B(mai_mai_n151_), .C(mai_mai_n90_), .Y(mai_mai_n423_));
  NO2        m401(.A(mai_mai_n421_), .B(mai_mai_n420_), .Y(mai_mai_n424_));
  NO3        m402(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n425_));
  NO2        m403(.A(i_6_), .B(i_7_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n426_), .B(mai_mai_n425_), .Y(mai_mai_n427_));
  NO2        m405(.A(i_11_), .B(i_1_), .Y(mai_mai_n428_));
  OR2        m406(.A(i_11_), .B(i_8_), .Y(mai_mai_n429_));
  NOi21      m407(.An(i_2_), .B(i_7_), .Y(mai_mai_n430_));
  NAi31      m408(.An(mai_mai_n429_), .B(mai_mai_n430_), .C(i_0_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n945_), .B(mai_mai_n395_), .Y(mai_mai_n432_));
  NO2        m410(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  NO2        m411(.A(i_3_), .B(mai_mai_n184_), .Y(mai_mai_n434_));
  NO2        m412(.A(i_6_), .B(i_10_), .Y(mai_mai_n435_));
  NA3        m413(.A(mai_mai_n435_), .B(mai_mai_n279_), .C(mai_mai_n434_), .Y(mai_mai_n436_));
  NO2        m414(.A(mai_mai_n436_), .B(mai_mai_n145_), .Y(mai_mai_n437_));
  NO2        m415(.A(mai_mai_n147_), .B(i_3_), .Y(mai_mai_n438_));
  NA3        m416(.A(mai_mai_n360_), .B(mai_mai_n170_), .C(mai_mai_n141_), .Y(mai_mai_n439_));
  INV        m417(.A(mai_mai_n439_), .Y(mai_mai_n440_));
  NO4        m418(.A(mai_mai_n440_), .B(mai_mai_n437_), .C(mai_mai_n433_), .D(mai_mai_n424_), .Y(mai_mai_n441_));
  NA2        m419(.A(mai_mai_n411_), .B(mai_mai_n356_), .Y(mai_mai_n442_));
  NO2        m420(.A(mai_mai_n442_), .B(mai_mai_n209_), .Y(mai_mai_n443_));
  NAi21      m421(.An(mai_mai_n203_), .B(mai_mai_n363_), .Y(mai_mai_n444_));
  NO2        m422(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n445_));
  NA3        m423(.A(mai_mai_n942_), .B(mai_mai_n445_), .C(mai_mai_n134_), .Y(mai_mai_n446_));
  OR3        m424(.A(mai_mai_n269_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n447_));
  NO2        m425(.A(mai_mai_n447_), .B(mai_mai_n446_), .Y(mai_mai_n448_));
  NA3        m426(.A(mai_mai_n272_), .B(mai_mai_n208_), .C(mai_mai_n65_), .Y(mai_mai_n449_));
  NO2        m427(.A(mai_mai_n449_), .B(mai_mai_n427_), .Y(mai_mai_n450_));
  NO3        m428(.A(mai_mai_n450_), .B(mai_mai_n448_), .C(mai_mai_n443_), .Y(mai_mai_n451_));
  NA4        m429(.A(mai_mai_n451_), .B(mai_mai_n441_), .C(mai_mai_n419_), .D(mai_mai_n416_), .Y(mai_mai_n452_));
  NA3        m430(.A(mai_mai_n272_), .B(mai_mai_n167_), .C(mai_mai_n165_), .Y(mai_mai_n453_));
  INV        m431(.A(mai_mai_n453_), .Y(mai_mai_n454_));
  BUFFER     m432(.A(mai_mai_n256_), .Y(mai_mai_n455_));
  NA2        m433(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n456_));
  AN2        m434(.A(i_12_), .B(mai_mai_n405_), .Y(mai_mai_n457_));
  OAI210     m435(.A0(mai_mai_n65_), .A1(mai_mai_n217_), .B0(mai_mai_n273_), .Y(mai_mai_n458_));
  AOI220     m436(.A0(mai_mai_n458_), .A1(mai_mai_n288_), .B0(mai_mai_n457_), .B1(mai_mai_n275_), .Y(mai_mai_n459_));
  NA4        m437(.A(mai_mai_n396_), .B(mai_mai_n395_), .C(mai_mai_n192_), .D(i_2_), .Y(mai_mai_n460_));
  INV        m438(.A(mai_mai_n460_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n319_), .B(mai_mai_n65_), .Y(mai_mai_n462_));
  INV        m440(.A(mai_mai_n329_), .Y(mai_mai_n463_));
  NO2        m441(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n464_));
  NA2        m442(.A(mai_mai_n39_), .B(i_13_), .Y(mai_mai_n465_));
  INV        m443(.A(mai_mai_n465_), .Y(mai_mai_n466_));
  AOI210     m444(.A0(mai_mai_n461_), .A1(mai_mai_n193_), .B0(mai_mai_n466_), .Y(mai_mai_n467_));
  OAI210     m445(.A0(i_8_), .A1(mai_mai_n57_), .B0(mai_mai_n126_), .Y(mai_mai_n468_));
  NO2        m446(.A(i_7_), .B(mai_mai_n189_), .Y(mai_mai_n469_));
  OR2        m447(.A(mai_mai_n174_), .B(i_4_), .Y(mai_mai_n470_));
  NO2        m448(.A(mai_mai_n470_), .B(mai_mai_n77_), .Y(mai_mai_n471_));
  AOI220     m449(.A0(mai_mai_n471_), .A1(mai_mai_n469_), .B0(mai_mai_n468_), .B1(mai_mai_n380_), .Y(mai_mai_n472_));
  NA4        m450(.A(mai_mai_n472_), .B(mai_mai_n467_), .C(mai_mai_n459_), .D(mai_mai_n456_), .Y(mai_mai_n473_));
  NA2        m451(.A(mai_mai_n355_), .B(mai_mai_n261_), .Y(mai_mai_n474_));
  OAI210     m452(.A0(mai_mai_n351_), .A1(mai_mai_n159_), .B0(mai_mai_n474_), .Y(mai_mai_n475_));
  NO2        m453(.A(i_12_), .B(mai_mai_n184_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n476_), .B(mai_mai_n210_), .Y(mai_mai_n477_));
  NO2        m455(.A(i_6_), .B(mai_mai_n477_), .Y(mai_mai_n478_));
  NOi21      m456(.An(mai_mai_n280_), .B(mai_mai_n38_), .Y(mai_mai_n479_));
  OAI210     m457(.A0(mai_mai_n479_), .A1(mai_mai_n478_), .B0(mai_mai_n475_), .Y(mai_mai_n480_));
  NO2        m458(.A(i_8_), .B(i_7_), .Y(mai_mai_n481_));
  INV        m459(.A(mai_mai_n208_), .Y(mai_mai_n482_));
  OAI220     m460(.A0(mai_mai_n46_), .A1(mai_mai_n470_), .B0(mai_mai_n482_), .B1(mai_mai_n226_), .Y(mai_mai_n483_));
  NA2        m461(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n484_));
  NO2        m462(.A(mai_mai_n484_), .B(i_6_), .Y(mai_mai_n485_));
  NA3        m463(.A(mai_mai_n485_), .B(mai_mai_n483_), .C(mai_mai_n481_), .Y(mai_mai_n486_));
  NO2        m464(.A(mai_mai_n420_), .B(mai_mai_n125_), .Y(mai_mai_n487_));
  NA2        m465(.A(mai_mai_n487_), .B(mai_mai_n240_), .Y(mai_mai_n488_));
  NO2        m466(.A(mai_mai_n267_), .B(mai_mai_n172_), .Y(mai_mai_n489_));
  NA3        m467(.A(mai_mai_n272_), .B(mai_mai_n165_), .C(mai_mai_n87_), .Y(mai_mai_n490_));
  NO2        m468(.A(mai_mai_n207_), .B(mai_mai_n44_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n147_), .B(i_5_), .Y(mai_mai_n492_));
  NA2        m470(.A(mai_mai_n492_), .B(mai_mai_n283_), .Y(mai_mai_n493_));
  OAI210     m471(.A0(mai_mai_n493_), .A1(mai_mai_n491_), .B0(mai_mai_n490_), .Y(mai_mai_n494_));
  OAI210     m472(.A0(mai_mai_n494_), .A1(mai_mai_n489_), .B0(mai_mai_n411_), .Y(mai_mai_n495_));
  NA4        m473(.A(mai_mai_n495_), .B(mai_mai_n488_), .C(mai_mai_n486_), .D(mai_mai_n480_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n253_), .B(mai_mai_n76_), .Y(mai_mai_n497_));
  NO2        m475(.A(mai_mai_n73_), .B(mai_mai_n497_), .Y(mai_mai_n498_));
  INV        m476(.A(mai_mai_n256_), .Y(mai_mai_n499_));
  NO2        m477(.A(mai_mai_n499_), .B(mai_mai_n164_), .Y(mai_mai_n500_));
  NA2        m478(.A(mai_mai_n208_), .B(i_3_), .Y(mai_mai_n501_));
  NA2        m479(.A(mai_mai_n398_), .B(mai_mai_n207_), .Y(mai_mai_n502_));
  NO2        m480(.A(mai_mai_n501_), .B(mai_mai_n502_), .Y(mai_mai_n503_));
  NA2        m481(.A(mai_mai_n476_), .B(mai_mai_n248_), .Y(mai_mai_n504_));
  NO2        m482(.A(mai_mai_n92_), .B(mai_mai_n504_), .Y(mai_mai_n505_));
  NO4        m483(.A(mai_mai_n505_), .B(mai_mai_n503_), .C(mai_mai_n500_), .D(mai_mai_n498_), .Y(mai_mai_n506_));
  NO4        m484(.A(mai_mai_n232_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n507_));
  NO3        m485(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n508_));
  NO2        m486(.A(mai_mai_n218_), .B(mai_mai_n36_), .Y(mai_mai_n509_));
  AN2        m487(.A(mai_mai_n509_), .B(mai_mai_n508_), .Y(mai_mai_n510_));
  OA210      m488(.A0(mai_mai_n510_), .A1(mai_mai_n507_), .B0(mai_mai_n319_), .Y(mai_mai_n511_));
  NO2        m489(.A(mai_mai_n379_), .B(i_1_), .Y(mai_mai_n512_));
  NOi31      m490(.An(mai_mai_n512_), .B(mai_mai_n406_), .C(mai_mai_n65_), .Y(mai_mai_n513_));
  AN3        m491(.A(mai_mai_n513_), .B(mai_mai_n377_), .C(mai_mai_n445_), .Y(mai_mai_n514_));
  NO2        m492(.A(mai_mai_n383_), .B(mai_mai_n168_), .Y(mai_mai_n515_));
  NO3        m493(.A(mai_mai_n515_), .B(mai_mai_n514_), .C(mai_mai_n511_), .Y(mai_mai_n516_));
  NOi21      m494(.An(i_10_), .B(i_6_), .Y(mai_mai_n517_));
  NO2        m495(.A(mai_mai_n77_), .B(mai_mai_n25_), .Y(mai_mai_n518_));
  NA2        m496(.A(mai_mai_n248_), .B(mai_mai_n517_), .Y(mai_mai_n519_));
  NO2        m497(.A(mai_mai_n519_), .B(mai_mai_n404_), .Y(mai_mai_n520_));
  NO2        m498(.A(mai_mai_n106_), .B(mai_mai_n23_), .Y(mai_mai_n521_));
  INV        m499(.A(mai_mai_n280_), .Y(mai_mai_n522_));
  AOI220     m500(.A0(mai_mai_n522_), .A1(mai_mai_n388_), .B0(mai_mai_n175_), .B1(mai_mai_n173_), .Y(mai_mai_n523_));
  NOi21      m501(.An(mai_mai_n138_), .B(mai_mai_n296_), .Y(mai_mai_n524_));
  NO3        m502(.A(mai_mai_n524_), .B(mai_mai_n523_), .C(mai_mai_n520_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n462_), .B(mai_mai_n344_), .Y(mai_mai_n526_));
  INV        m504(.A(mai_mai_n283_), .Y(mai_mai_n527_));
  NO2        m505(.A(i_12_), .B(mai_mai_n77_), .Y(mai_mai_n528_));
  NA2        m506(.A(mai_mai_n528_), .B(mai_mai_n248_), .Y(mai_mai_n529_));
  NA2        m507(.A(mai_mai_n352_), .B(mai_mai_n253_), .Y(mai_mai_n530_));
  AOI210     m508(.A0(mai_mai_n530_), .A1(mai_mai_n529_), .B0(mai_mai_n527_), .Y(mai_mai_n531_));
  NO3        m509(.A(i_4_), .B(mai_mai_n307_), .C(mai_mai_n267_), .Y(mai_mai_n532_));
  NO2        m510(.A(i_2_), .B(mai_mai_n444_), .Y(mai_mai_n533_));
  NO4        m511(.A(mai_mai_n533_), .B(mai_mai_n532_), .C(mai_mai_n531_), .D(mai_mai_n526_), .Y(mai_mai_n534_));
  NA4        m512(.A(mai_mai_n534_), .B(mai_mai_n525_), .C(mai_mai_n516_), .D(mai_mai_n506_), .Y(mai_mai_n535_));
  NO4        m513(.A(mai_mai_n535_), .B(mai_mai_n496_), .C(mai_mai_n473_), .D(mai_mai_n452_), .Y(mai_mai_n536_));
  NA4        m514(.A(mai_mai_n536_), .B(mai_mai_n394_), .C(mai_mai_n318_), .D(mai_mai_n278_), .Y(mai7));
  NA2        m515(.A(mai_mai_n435_), .B(mai_mai_n76_), .Y(mai_mai_n538_));
  NA2        m516(.A(mai_mai_n136_), .B(i_8_), .Y(mai_mai_n539_));
  NO2        m517(.A(mai_mai_n539_), .B(mai_mai_n538_), .Y(mai_mai_n540_));
  NA3        m518(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n541_));
  NO2        m519(.A(mai_mai_n221_), .B(i_4_), .Y(mai_mai_n542_));
  NA2        m520(.A(mai_mai_n542_), .B(i_8_), .Y(mai_mai_n543_));
  NA2        m521(.A(i_2_), .B(mai_mai_n77_), .Y(mai_mai_n544_));
  OAI210     m522(.A0(mai_mai_n80_), .A1(mai_mai_n192_), .B0(mai_mai_n193_), .Y(mai_mai_n545_));
  NA2        m523(.A(i_4_), .B(i_8_), .Y(mai_mai_n546_));
  OAI220     m524(.A0(mai_mai_n37_), .A1(mai_mai_n544_), .B0(mai_mai_n545_), .B1(i_13_), .Y(mai_mai_n547_));
  NO2        m525(.A(mai_mai_n547_), .B(mai_mai_n540_), .Y(mai_mai_n548_));
  OR2        m526(.A(i_6_), .B(i_10_), .Y(mai_mai_n549_));
  NO2        m527(.A(mai_mai_n549_), .B(mai_mai_n23_), .Y(mai_mai_n550_));
  OR3        m528(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n551_));
  NO3        m529(.A(mai_mai_n551_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n552_));
  INV        m530(.A(mai_mai_n190_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n552_), .B(mai_mai_n550_), .Y(mai_mai_n554_));
  OR2        m532(.A(mai_mai_n554_), .B(mai_mai_n527_), .Y(mai_mai_n555_));
  AOI210     m533(.A0(mai_mai_n555_), .A1(mai_mai_n548_), .B0(mai_mai_n57_), .Y(mai_mai_n556_));
  NOi21      m534(.An(i_11_), .B(i_7_), .Y(mai_mai_n557_));
  AO210      m535(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n558_));
  NO2        m536(.A(mai_mai_n558_), .B(mai_mai_n557_), .Y(mai_mai_n559_));
  NA3        m537(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n560_));
  NAi31      m538(.An(mai_mai_n560_), .B(i_12_), .C(i_11_), .Y(mai_mai_n561_));
  NO2        m539(.A(mai_mai_n561_), .B(mai_mai_n57_), .Y(mai_mai_n562_));
  NA2        m540(.A(mai_mai_n79_), .B(mai_mai_n57_), .Y(mai_mai_n563_));
  AO210      m541(.A0(mai_mai_n563_), .A1(mai_mai_n344_), .B0(mai_mai_n41_), .Y(mai_mai_n564_));
  NA2        m542(.A(mai_mai_n211_), .B(mai_mai_n57_), .Y(mai_mai_n565_));
  NA2        m543(.A(mai_mai_n373_), .B(mai_mai_n31_), .Y(mai_mai_n566_));
  OR2        m544(.A(mai_mai_n196_), .B(mai_mai_n99_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n567_), .B(mai_mai_n566_), .Y(mai_mai_n568_));
  NO2        m546(.A(mai_mai_n57_), .B(i_9_), .Y(mai_mai_n569_));
  NA2        m547(.A(mai_mai_n57_), .B(mai_mai_n568_), .Y(mai_mai_n570_));
  NO2        m548(.A(i_1_), .B(i_12_), .Y(mai_mai_n571_));
  NA3        m549(.A(mai_mai_n570_), .B(mai_mai_n565_), .C(mai_mai_n564_), .Y(mai_mai_n572_));
  OAI210     m550(.A0(mai_mai_n572_), .A1(mai_mai_n562_), .B0(i_6_), .Y(mai_mai_n573_));
  NO2        m551(.A(i_6_), .B(i_11_), .Y(mai_mai_n574_));
  INV        m552(.A(mai_mai_n407_), .Y(mai_mai_n575_));
  NO4        m553(.A(i_12_), .B(mai_mai_n120_), .C(i_13_), .D(mai_mai_n77_), .Y(mai_mai_n576_));
  NA2        m554(.A(mai_mai_n576_), .B(mai_mai_n569_), .Y(mai_mai_n577_));
  NA2        m555(.A(mai_mai_n221_), .B(i_6_), .Y(mai_mai_n578_));
  INV        m556(.A(mai_mai_n577_), .Y(mai_mai_n579_));
  NA3        m557(.A(mai_mai_n481_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n580_));
  NA2        m558(.A(mai_mai_n130_), .B(i_9_), .Y(mai_mai_n581_));
  NA3        m559(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n583_));
  NA3        m561(.A(mai_mai_n583_), .B(mai_mai_n241_), .C(mai_mai_n44_), .Y(mai_mai_n584_));
  OAI220     m562(.A0(mai_mai_n584_), .A1(mai_mai_n582_), .B0(mai_mai_n581_), .B1(mai_mai_n933_), .Y(mai_mai_n585_));
  NA3        m563(.A(mai_mai_n569_), .B(mai_mai_n283_), .C(i_6_), .Y(mai_mai_n586_));
  NO2        m564(.A(mai_mai_n586_), .B(mai_mai_n23_), .Y(mai_mai_n587_));
  AOI210     m565(.A0(mai_mai_n428_), .A1(mai_mai_n381_), .B0(mai_mai_n225_), .Y(mai_mai_n588_));
  NO2        m566(.A(mai_mai_n588_), .B(mai_mai_n544_), .Y(mai_mai_n589_));
  NAi21      m567(.An(mai_mai_n580_), .B(mai_mai_n83_), .Y(mai_mai_n590_));
  NO2        m568(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n591_), .B(mai_mai_n24_), .Y(mai_mai_n592_));
  INV        m570(.A(mai_mai_n590_), .Y(mai_mai_n593_));
  OR4        m571(.A(mai_mai_n593_), .B(mai_mai_n589_), .C(mai_mai_n587_), .D(mai_mai_n585_), .Y(mai_mai_n594_));
  NO3        m572(.A(mai_mai_n594_), .B(mai_mai_n579_), .C(mai_mai_n575_), .Y(mai_mai_n595_));
  NO2        m573(.A(mai_mai_n221_), .B(mai_mai_n92_), .Y(mai_mai_n596_));
  NO2        m574(.A(mai_mai_n596_), .B(mai_mai_n557_), .Y(mai_mai_n597_));
  NA2        m575(.A(mai_mai_n597_), .B(i_1_), .Y(mai_mai_n598_));
  NO2        m576(.A(mai_mai_n598_), .B(mai_mai_n551_), .Y(mai_mai_n599_));
  NA2        m577(.A(mai_mai_n599_), .B(mai_mai_n46_), .Y(mai_mai_n600_));
  NA2        m578(.A(i_3_), .B(mai_mai_n184_), .Y(mai_mai_n601_));
  NO2        m579(.A(mai_mai_n601_), .B(mai_mai_n106_), .Y(mai_mai_n602_));
  AN2        m580(.A(mai_mai_n602_), .B(mai_mai_n485_), .Y(mai_mai_n603_));
  NO2        m581(.A(mai_mai_n77_), .B(i_9_), .Y(mai_mai_n604_));
  NA2        m582(.A(i_1_), .B(i_3_), .Y(mai_mai_n605_));
  NO2        m583(.A(mai_mai_n408_), .B(mai_mai_n84_), .Y(mai_mai_n606_));
  AOI210     m584(.A0(i_11_), .A1(mai_mai_n517_), .B0(mai_mai_n606_), .Y(mai_mai_n607_));
  NO2        m585(.A(mai_mai_n607_), .B(mai_mai_n605_), .Y(mai_mai_n608_));
  NO2        m586(.A(mai_mai_n608_), .B(mai_mai_n603_), .Y(mai_mai_n609_));
  NA4        m587(.A(mai_mai_n609_), .B(mai_mai_n600_), .C(mai_mai_n595_), .D(mai_mai_n573_), .Y(mai_mai_n610_));
  NO3        m588(.A(mai_mai_n429_), .B(i_3_), .C(i_7_), .Y(mai_mai_n611_));
  NOi21      m589(.An(mai_mai_n611_), .B(i_10_), .Y(mai_mai_n612_));
  OA210      m590(.A0(mai_mai_n612_), .A1(mai_mai_n228_), .B0(mai_mai_n77_), .Y(mai_mai_n613_));
  NA2        m591(.A(mai_mai_n337_), .B(mai_mai_n336_), .Y(mai_mai_n614_));
  NA3        m592(.A(mai_mai_n435_), .B(mai_mai_n464_), .C(mai_mai_n46_), .Y(mai_mai_n615_));
  NO3        m593(.A(mai_mai_n430_), .B(mai_mai_n546_), .C(mai_mai_n77_), .Y(mai_mai_n616_));
  NA2        m594(.A(mai_mai_n616_), .B(mai_mai_n25_), .Y(mai_mai_n617_));
  NA3        m595(.A(mai_mai_n151_), .B(mai_mai_n76_), .C(mai_mai_n77_), .Y(mai_mai_n618_));
  NA4        m596(.A(mai_mai_n618_), .B(mai_mai_n617_), .C(mai_mai_n615_), .D(mai_mai_n614_), .Y(mai_mai_n619_));
  OAI210     m597(.A0(mai_mai_n619_), .A1(mai_mai_n613_), .B0(i_1_), .Y(mai_mai_n620_));
  AOI210     m598(.A0(mai_mai_n241_), .A1(mai_mai_n88_), .B0(i_1_), .Y(mai_mai_n621_));
  NO2        m599(.A(mai_mai_n335_), .B(i_2_), .Y(mai_mai_n622_));
  NA2        m600(.A(mai_mai_n622_), .B(mai_mai_n621_), .Y(mai_mai_n623_));
  AOI210     m601(.A0(mai_mai_n623_), .A1(mai_mai_n620_), .B0(i_13_), .Y(mai_mai_n624_));
  OR2        m602(.A(i_11_), .B(i_7_), .Y(mai_mai_n625_));
  AOI220     m603(.A0(mai_mai_n422_), .A1(mai_mai_n151_), .B0(i_2_), .B1(mai_mai_n130_), .Y(mai_mai_n626_));
  NO2        m604(.A(mai_mai_n626_), .B(mai_mai_n44_), .Y(mai_mai_n627_));
  NA2        m605(.A(mai_mai_n228_), .B(mai_mai_n123_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n628_), .B(mai_mai_n41_), .Y(mai_mai_n629_));
  AOI210     m607(.A0(mai_mai_n627_), .A1(mai_mai_n298_), .B0(mai_mai_n629_), .Y(mai_mai_n630_));
  INV        m608(.A(mai_mai_n106_), .Y(mai_mai_n631_));
  AOI220     m609(.A0(mai_mai_n631_), .A1(mai_mai_n64_), .B0(mai_mai_n352_), .B1(mai_mai_n583_), .Y(mai_mai_n632_));
  NO2        m610(.A(mai_mai_n632_), .B(mai_mai_n226_), .Y(mai_mai_n633_));
  AOI210     m611(.A0(mai_mai_n399_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n634_));
  NOi31      m612(.An(mai_mai_n634_), .B(mai_mai_n538_), .C(mai_mai_n44_), .Y(mai_mai_n635_));
  NA2        m613(.A(mai_mai_n119_), .B(i_13_), .Y(mai_mai_n636_));
  NO2        m614(.A(mai_mai_n582_), .B(mai_mai_n106_), .Y(mai_mai_n637_));
  INV        m615(.A(mai_mai_n637_), .Y(mai_mai_n638_));
  OAI220     m616(.A0(mai_mai_n638_), .A1(mai_mai_n63_), .B0(mai_mai_n636_), .B1(mai_mai_n621_), .Y(mai_mai_n639_));
  NO3        m617(.A(mai_mai_n63_), .B(mai_mai_n32_), .C(mai_mai_n92_), .Y(mai_mai_n640_));
  NA2        m618(.A(mai_mai_n26_), .B(mai_mai_n184_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n641_), .B(i_7_), .Y(mai_mai_n642_));
  NO3        m620(.A(mai_mai_n430_), .B(mai_mai_n221_), .C(mai_mai_n77_), .Y(mai_mai_n643_));
  AOI210     m621(.A0(mai_mai_n643_), .A1(mai_mai_n642_), .B0(mai_mai_n640_), .Y(mai_mai_n644_));
  NO2        m622(.A(mai_mai_n644_), .B(mai_mai_n553_), .Y(mai_mai_n645_));
  NO4        m623(.A(mai_mai_n645_), .B(mai_mai_n639_), .C(mai_mai_n635_), .D(mai_mai_n633_), .Y(mai_mai_n646_));
  OR2        m624(.A(i_11_), .B(i_6_), .Y(mai_mai_n647_));
  NA3        m625(.A(mai_mai_n542_), .B(mai_mai_n641_), .C(i_7_), .Y(mai_mai_n648_));
  AOI210     m626(.A0(mai_mai_n648_), .A1(mai_mai_n638_), .B0(mai_mai_n647_), .Y(mai_mai_n649_));
  NA3        m627(.A(mai_mai_n373_), .B(i_10_), .C(mai_mai_n88_), .Y(mai_mai_n650_));
  NA2        m628(.A(mai_mai_n574_), .B(i_13_), .Y(mai_mai_n651_));
  NA2        m629(.A(mai_mai_n93_), .B(mai_mai_n641_), .Y(mai_mai_n652_));
  NAi21      m630(.An(i_11_), .B(i_12_), .Y(mai_mai_n653_));
  NOi41      m631(.An(mai_mai_n102_), .B(mai_mai_n653_), .C(i_13_), .D(mai_mai_n77_), .Y(mai_mai_n654_));
  NO3        m632(.A(mai_mai_n430_), .B(mai_mai_n528_), .C(mai_mai_n546_), .Y(mai_mai_n655_));
  AOI220     m633(.A0(mai_mai_n655_), .A1(mai_mai_n279_), .B0(mai_mai_n654_), .B1(mai_mai_n652_), .Y(mai_mai_n656_));
  NA3        m634(.A(mai_mai_n656_), .B(mai_mai_n651_), .C(mai_mai_n650_), .Y(mai_mai_n657_));
  OAI210     m635(.A0(mai_mai_n657_), .A1(mai_mai_n649_), .B0(mai_mai_n57_), .Y(mai_mai_n658_));
  NO2        m636(.A(i_2_), .B(i_12_), .Y(mai_mai_n659_));
  NA2        m637(.A(mai_mai_n221_), .B(mai_mai_n334_), .Y(mai_mai_n660_));
  NO2        m638(.A(mai_mai_n120_), .B(i_2_), .Y(mai_mai_n661_));
  NA2        m639(.A(mai_mai_n661_), .B(mai_mai_n571_), .Y(mai_mai_n662_));
  NA2        m640(.A(mai_mai_n662_), .B(mai_mai_n660_), .Y(mai_mai_n663_));
  NA3        m641(.A(mai_mai_n663_), .B(mai_mai_n45_), .C(mai_mai_n210_), .Y(mai_mai_n664_));
  NA4        m642(.A(mai_mai_n664_), .B(mai_mai_n658_), .C(mai_mai_n646_), .D(mai_mai_n630_), .Y(mai_mai_n665_));
  OR4        m643(.A(mai_mai_n665_), .B(mai_mai_n624_), .C(mai_mai_n610_), .D(mai_mai_n556_), .Y(mai5));
  AOI210     m644(.A0(mai_mai_n597_), .A1(mai_mai_n244_), .B0(mai_mai_n380_), .Y(mai_mai_n667_));
  AN2        m645(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n668_));
  NA3        m646(.A(mai_mai_n668_), .B(mai_mai_n659_), .C(mai_mai_n99_), .Y(mai_mai_n669_));
  NO2        m647(.A(mai_mai_n543_), .B(i_11_), .Y(mai_mai_n670_));
  NA2        m648(.A(mai_mai_n80_), .B(mai_mai_n670_), .Y(mai_mai_n671_));
  NA3        m649(.A(mai_mai_n671_), .B(mai_mai_n669_), .C(mai_mai_n667_), .Y(mai_mai_n672_));
  NO3        m650(.A(i_11_), .B(mai_mai_n221_), .C(i_13_), .Y(mai_mai_n673_));
  NA2        m651(.A(i_12_), .B(i_8_), .Y(mai_mai_n674_));
  INV        m652(.A(mai_mai_n398_), .Y(mai_mai_n675_));
  NA2        m653(.A(mai_mai_n283_), .B(mai_mai_n521_), .Y(mai_mai_n676_));
  INV        m654(.A(mai_mai_n676_), .Y(mai_mai_n677_));
  NO2        m655(.A(mai_mai_n677_), .B(mai_mai_n672_), .Y(mai_mai_n678_));
  INV        m656(.A(mai_mai_n162_), .Y(mai_mai_n679_));
  OAI210     m657(.A0(mai_mai_n622_), .A1(mai_mai_n400_), .B0(mai_mai_n102_), .Y(mai_mai_n680_));
  NO2        m658(.A(mai_mai_n680_), .B(mai_mai_n679_), .Y(mai_mai_n681_));
  NO2        m659(.A(mai_mai_n408_), .B(mai_mai_n26_), .Y(mai_mai_n682_));
  AOI210     m660(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n379_), .Y(mai_mai_n683_));
  AOI210     m661(.A0(mai_mai_n683_), .A1(i_2_), .B0(mai_mai_n681_), .Y(mai_mai_n684_));
  INV        m662(.A(mai_mai_n163_), .Y(mai_mai_n685_));
  NO3        m663(.A(mai_mai_n558_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n686_));
  AOI210     m664(.A0(mai_mai_n685_), .A1(mai_mai_n80_), .B0(mai_mai_n686_), .Y(mai_mai_n687_));
  NO2        m665(.A(mai_mai_n687_), .B(mai_mai_n184_), .Y(mai_mai_n688_));
  OA210      m666(.A0(mai_mai_n559_), .A1(mai_mai_n118_), .B0(i_13_), .Y(mai_mai_n689_));
  NA2        m667(.A(mai_mai_n190_), .B(mai_mai_n192_), .Y(mai_mai_n690_));
  NA2        m668(.A(mai_mai_n143_), .B(i_8_), .Y(mai_mai_n691_));
  AOI210     m669(.A0(mai_mai_n691_), .A1(mai_mai_n690_), .B0(mai_mai_n338_), .Y(mai_mai_n692_));
  AOI210     m670(.A0(mai_mai_n196_), .A1(mai_mai_n140_), .B0(mai_mai_n464_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n693_), .B(mai_mai_n381_), .Y(mai_mai_n694_));
  NO2        m672(.A(mai_mai_n93_), .B(mai_mai_n44_), .Y(mai_mai_n695_));
  INV        m673(.A(mai_mai_n268_), .Y(mai_mai_n696_));
  NA4        m674(.A(mai_mai_n696_), .B(mai_mai_n272_), .C(mai_mai_n116_), .D(mai_mai_n42_), .Y(mai_mai_n697_));
  OAI210     m675(.A0(mai_mai_n697_), .A1(mai_mai_n695_), .B0(mai_mai_n694_), .Y(mai_mai_n698_));
  NO4        m676(.A(mai_mai_n698_), .B(mai_mai_n692_), .C(mai_mai_n689_), .D(mai_mai_n688_), .Y(mai_mai_n699_));
  NA2        m677(.A(mai_mai_n521_), .B(mai_mai_n28_), .Y(mai_mai_n700_));
  NA2        m678(.A(mai_mai_n673_), .B(mai_mai_n249_), .Y(mai_mai_n701_));
  NA2        m679(.A(mai_mai_n701_), .B(mai_mai_n700_), .Y(mai_mai_n702_));
  NA2        m680(.A(mai_mai_n702_), .B(mai_mai_n46_), .Y(mai_mai_n703_));
  NA4        m681(.A(mai_mai_n703_), .B(mai_mai_n699_), .C(mai_mai_n684_), .D(mai_mai_n678_), .Y(mai6));
  NO3        m682(.A(i_9_), .B(mai_mai_n274_), .C(i_1_), .Y(mai_mai_n705_));
  NO2        m683(.A(mai_mai_n177_), .B(mai_mai_n131_), .Y(mai_mai_n706_));
  OAI210     m684(.A0(mai_mai_n706_), .A1(mai_mai_n705_), .B0(mai_mai_n661_), .Y(mai_mai_n707_));
  NA4        m685(.A(mai_mai_n356_), .B(mai_mai_n434_), .C(mai_mai_n63_), .D(mai_mai_n92_), .Y(mai_mai_n708_));
  INV        m686(.A(mai_mai_n708_), .Y(mai_mai_n709_));
  NO2        m687(.A(i_11_), .B(i_9_), .Y(mai_mai_n710_));
  NO2        m688(.A(mai_mai_n709_), .B(mai_mai_n294_), .Y(mai_mai_n711_));
  AO210      m689(.A0(mai_mai_n711_), .A1(mai_mai_n707_), .B0(i_12_), .Y(mai_mai_n712_));
  NA2        m690(.A(mai_mai_n339_), .B(mai_mai_n301_), .Y(mai_mai_n713_));
  NA2        m691(.A(mai_mai_n528_), .B(mai_mai_n57_), .Y(mai_mai_n714_));
  NA2        m692(.A(mai_mai_n612_), .B(mai_mai_n63_), .Y(mai_mai_n715_));
  NA4        m693(.A(mai_mai_n563_), .B(mai_mai_n715_), .C(mai_mai_n714_), .D(mai_mai_n713_), .Y(mai_mai_n716_));
  INV        m694(.A(mai_mai_n187_), .Y(mai_mai_n717_));
  AOI220     m695(.A0(mai_mai_n717_), .A1(mai_mai_n710_), .B0(mai_mai_n716_), .B1(mai_mai_n65_), .Y(mai_mai_n718_));
  INV        m696(.A(mai_mai_n293_), .Y(mai_mai_n719_));
  NA2        m697(.A(mai_mai_n67_), .B(mai_mai_n123_), .Y(mai_mai_n720_));
  INV        m698(.A(mai_mai_n116_), .Y(mai_mai_n721_));
  NA2        m699(.A(mai_mai_n721_), .B(mai_mai_n46_), .Y(mai_mai_n722_));
  AOI210     m700(.A0(mai_mai_n722_), .A1(mai_mai_n720_), .B0(mai_mai_n719_), .Y(mai_mai_n723_));
  NO2        m701(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n724_));
  NA3        m702(.A(mai_mai_n724_), .B(mai_mai_n426_), .C(mai_mai_n356_), .Y(mai_mai_n725_));
  OAI210     m703(.A0(mai_mai_n611_), .A1(mai_mai_n509_), .B0(mai_mai_n508_), .Y(mai_mai_n726_));
  NA2        m704(.A(mai_mai_n726_), .B(mai_mai_n725_), .Y(mai_mai_n727_));
  OR2        m705(.A(mai_mai_n727_), .B(mai_mai_n723_), .Y(mai_mai_n728_));
  NO2        m706(.A(mai_mai_n625_), .B(i_2_), .Y(mai_mai_n729_));
  NA2        m707(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n730_));
  OAI210     m708(.A0(mai_mai_n730_), .A1(mai_mai_n372_), .B0(mai_mai_n324_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n731_), .B(mai_mai_n729_), .Y(mai_mai_n732_));
  AO220      m710(.A0(mai_mai_n323_), .A1(mai_mai_n314_), .B0(mai_mai_n362_), .B1(i_8_), .Y(mai_mai_n733_));
  NA3        m711(.A(mai_mai_n733_), .B(mai_mai_n234_), .C(i_7_), .Y(mai_mai_n734_));
  OR2        m712(.A(mai_mai_n559_), .B(mai_mai_n400_), .Y(mai_mai_n735_));
  NA2        m713(.A(mai_mai_n735_), .B(mai_mai_n139_), .Y(mai_mai_n736_));
  OR2        m714(.A(mai_mai_n675_), .B(mai_mai_n36_), .Y(mai_mai_n737_));
  NA4        m715(.A(mai_mai_n737_), .B(mai_mai_n736_), .C(mai_mai_n734_), .D(mai_mai_n732_), .Y(mai_mai_n738_));
  OAI210     m716(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n78_), .Y(mai_mai_n739_));
  NA2        m717(.A(mai_mai_n739_), .B(mai_mai_n508_), .Y(mai_mai_n740_));
  NA3        m718(.A(mai_mai_n338_), .B(mai_mai_n222_), .C(mai_mai_n139_), .Y(mai_mai_n741_));
  OAI210     m719(.A0(mai_mai_n362_), .A1(mai_mai_n193_), .B0(mai_mai_n62_), .Y(mai_mai_n742_));
  NA4        m720(.A(mai_mai_n742_), .B(mai_mai_n741_), .C(mai_mai_n740_), .D(mai_mai_n545_), .Y(mai_mai_n743_));
  AO210      m721(.A0(mai_mai_n464_), .A1(mai_mai_n46_), .B0(mai_mai_n79_), .Y(mai_mai_n744_));
  NA3        m722(.A(mai_mai_n744_), .B(mai_mai_n435_), .C(mai_mai_n205_), .Y(mai_mai_n745_));
  AOI210     m723(.A0(mai_mai_n400_), .A1(mai_mai_n398_), .B0(mai_mai_n507_), .Y(mai_mai_n746_));
  NA2        m724(.A(mai_mai_n103_), .B(mai_mai_n371_), .Y(mai_mai_n747_));
  NA3        m725(.A(mai_mai_n747_), .B(mai_mai_n746_), .C(mai_mai_n745_), .Y(mai_mai_n748_));
  NO4        m726(.A(mai_mai_n748_), .B(mai_mai_n743_), .C(mai_mai_n738_), .D(mai_mai_n728_), .Y(mai_mai_n749_));
  NA4        m727(.A(mai_mai_n749_), .B(mai_mai_n718_), .C(mai_mai_n712_), .D(mai_mai_n346_), .Y(mai3));
  NA2        m728(.A(i_6_), .B(i_7_), .Y(mai_mai_n751_));
  NO2        m729(.A(mai_mai_n751_), .B(i_0_), .Y(mai_mai_n752_));
  NO2        m730(.A(i_11_), .B(mai_mai_n221_), .Y(mai_mai_n753_));
  OAI210     m731(.A0(mai_mai_n752_), .A1(mai_mai_n257_), .B0(mai_mai_n753_), .Y(mai_mai_n754_));
  NO2        m732(.A(mai_mai_n754_), .B(mai_mai_n184_), .Y(mai_mai_n755_));
  NO3        m733(.A(mai_mai_n404_), .B(mai_mai_n81_), .C(mai_mai_n44_), .Y(mai_mai_n756_));
  OA210      m734(.A0(mai_mai_n756_), .A1(mai_mai_n755_), .B0(mai_mai_n165_), .Y(mai_mai_n757_));
  INV        m735(.A(mai_mai_n741_), .Y(mai_mai_n758_));
  NA2        m736(.A(mai_mai_n758_), .B(mai_mai_n40_), .Y(mai_mai_n759_));
  NO2        m737(.A(mai_mai_n567_), .B(mai_mai_n408_), .Y(mai_mai_n760_));
  NA2        m738(.A(mai_mai_n373_), .B(mai_mai_n45_), .Y(mai_mai_n761_));
  AOI210     m739(.A0(mai_mai_n934_), .A1(mai_mai_n759_), .B0(mai_mai_n48_), .Y(mai_mai_n762_));
  NO4        m740(.A(mai_mai_n342_), .B(mai_mai_n349_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n763_));
  NA2        m741(.A(mai_mai_n634_), .B(mai_mai_n604_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n299_), .B(i_5_), .Y(mai_mai_n765_));
  OAI220     m743(.A0(mai_mai_n765_), .A1(mai_mai_n764_), .B0(mai_mai_n938_), .B1(mai_mai_n57_), .Y(mai_mai_n766_));
  NOi21      m744(.An(i_5_), .B(i_9_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n767_), .B(mai_mai_n396_), .Y(mai_mai_n768_));
  NA2        m746(.A(mai_mai_n241_), .B(mai_mai_n428_), .Y(mai_mai_n769_));
  NO2        m747(.A(mai_mai_n166_), .B(mai_mai_n140_), .Y(mai_mai_n770_));
  INV        m748(.A(mai_mai_n770_), .Y(mai_mai_n771_));
  OAI220     m749(.A0(mai_mai_n771_), .A1(mai_mai_n172_), .B0(mai_mai_n769_), .B1(mai_mai_n768_), .Y(mai_mai_n772_));
  NO4        m750(.A(mai_mai_n772_), .B(mai_mai_n766_), .C(mai_mai_n762_), .D(mai_mai_n757_), .Y(mai_mai_n773_));
  NA2        m751(.A(mai_mai_n177_), .B(mai_mai_n24_), .Y(mai_mai_n774_));
  NO2        m752(.A(mai_mai_n37_), .B(mai_mai_n774_), .Y(mai_mai_n775_));
  NA2        m753(.A(mai_mai_n279_), .B(mai_mai_n121_), .Y(mai_mai_n776_));
  NAi21      m754(.An(mai_mai_n152_), .B(i_5_), .Y(mai_mai_n777_));
  NO2        m755(.A(mai_mai_n776_), .B(mai_mai_n364_), .Y(mai_mai_n778_));
  NO2        m756(.A(mai_mai_n778_), .B(mai_mai_n775_), .Y(mai_mai_n779_));
  NA2        m757(.A(mai_mai_n518_), .B(i_0_), .Y(mai_mai_n780_));
  NO3        m758(.A(mai_mai_n780_), .B(mai_mai_n351_), .C(mai_mai_n80_), .Y(mai_mai_n781_));
  INV        m759(.A(mai_mai_n781_), .Y(mai_mai_n782_));
  NA2        m760(.A(mai_mai_n673_), .B(mai_mai_n294_), .Y(mai_mai_n783_));
  OAI220     m761(.A0(i_6_), .A1(mai_mai_n783_), .B0(mai_mai_n592_), .B1(mai_mai_n482_), .Y(mai_mai_n784_));
  NA2        m762(.A(i_0_), .B(i_10_), .Y(mai_mai_n785_));
  NO4        m763(.A(mai_mai_n106_), .B(mai_mai_n53_), .C(mai_mai_n601_), .D(i_5_), .Y(mai_mai_n786_));
  AN2        m764(.A(mai_mai_n786_), .B(i_10_), .Y(mai_mai_n787_));
  NA2        m765(.A(mai_mai_n177_), .B(mai_mai_n76_), .Y(mai_mai_n788_));
  NA2        m766(.A(mai_mai_n512_), .B(i_4_), .Y(mai_mai_n789_));
  NA2        m767(.A(mai_mai_n180_), .B(mai_mai_n192_), .Y(mai_mai_n790_));
  OAI220     m768(.A0(mai_mai_n790_), .A1(mai_mai_n783_), .B0(mai_mai_n789_), .B1(mai_mai_n788_), .Y(mai_mai_n791_));
  NO3        m769(.A(mai_mai_n791_), .B(mai_mai_n787_), .C(mai_mai_n784_), .Y(mai_mai_n792_));
  NA3        m770(.A(mai_mai_n792_), .B(mai_mai_n782_), .C(mai_mai_n779_), .Y(mai_mai_n793_));
  NA2        m771(.A(i_11_), .B(i_9_), .Y(mai_mai_n794_));
  NO3        m772(.A(i_12_), .B(mai_mai_n794_), .C(mai_mai_n544_), .Y(mai_mai_n795_));
  AN2        m773(.A(mai_mai_n795_), .B(i_10_), .Y(mai_mai_n796_));
  NO2        m774(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n797_));
  NA2        m775(.A(mai_mai_n360_), .B(mai_mai_n170_), .Y(mai_mai_n798_));
  NA2        m776(.A(mai_mai_n798_), .B(mai_mai_n150_), .Y(mai_mai_n799_));
  NO2        m777(.A(mai_mai_n794_), .B(mai_mai_n65_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n166_), .B(i_0_), .Y(mai_mai_n801_));
  NA2        m779(.A(mai_mai_n426_), .B(mai_mai_n216_), .Y(mai_mai_n802_));
  NA2        m780(.A(mai_mai_n337_), .B(i_4_), .Y(mai_mai_n803_));
  OAI220     m781(.A0(mai_mai_n803_), .A1(mai_mai_n768_), .B0(mai_mai_n802_), .B1(mai_mai_n166_), .Y(mai_mai_n804_));
  NO3        m782(.A(mai_mai_n804_), .B(mai_mai_n799_), .C(mai_mai_n796_), .Y(mai_mai_n805_));
  NA2        m783(.A(mai_mai_n591_), .B(mai_mai_n113_), .Y(mai_mai_n806_));
  NO2        m784(.A(i_6_), .B(mai_mai_n806_), .Y(mai_mai_n807_));
  AOI210     m785(.A0(mai_mai_n399_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n808_));
  NA2        m786(.A(mai_mai_n162_), .B(mai_mai_n94_), .Y(mai_mai_n809_));
  NOi32      m787(.An(mai_mai_n808_), .Bn(mai_mai_n180_), .C(mai_mai_n809_), .Y(mai_mai_n810_));
  NA2        m788(.A(i_10_), .B(mai_mai_n294_), .Y(mai_mai_n811_));
  NO2        m789(.A(mai_mai_n811_), .B(mai_mai_n761_), .Y(mai_mai_n812_));
  NO3        m790(.A(mai_mai_n812_), .B(mai_mai_n810_), .C(mai_mai_n807_), .Y(mai_mai_n813_));
  NOi21      m791(.An(i_7_), .B(i_5_), .Y(mai_mai_n814_));
  NOi31      m792(.An(mai_mai_n814_), .B(i_0_), .C(mai_mai_n653_), .Y(mai_mai_n815_));
  NA3        m793(.A(mai_mai_n815_), .B(mai_mai_n350_), .C(i_6_), .Y(mai_mai_n816_));
  OA210      m794(.A0(mai_mai_n809_), .A1(mai_mai_n463_), .B0(mai_mai_n816_), .Y(mai_mai_n817_));
  NO3        m795(.A(mai_mai_n367_), .B(mai_mai_n326_), .C(mai_mai_n322_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n235_), .B(mai_mai_n284_), .Y(mai_mai_n819_));
  INV        m797(.A(mai_mai_n818_), .Y(mai_mai_n820_));
  NA4        m798(.A(mai_mai_n820_), .B(mai_mai_n817_), .C(mai_mai_n813_), .D(mai_mai_n805_), .Y(mai_mai_n821_));
  OA210      m799(.A0(mai_mai_n426_), .A1(mai_mai_n208_), .B0(mai_mai_n425_), .Y(mai_mai_n822_));
  NA3        m800(.A(mai_mai_n425_), .B(mai_mai_n373_), .C(mai_mai_n45_), .Y(mai_mai_n823_));
  OAI210     m801(.A0(mai_mai_n777_), .A1(i_6_), .B0(mai_mai_n823_), .Y(mai_mai_n824_));
  NA2        m802(.A(mai_mai_n800_), .B(mai_mai_n272_), .Y(mai_mai_n825_));
  NA2        m803(.A(mai_mai_n179_), .B(mai_mai_n825_), .Y(mai_mai_n826_));
  AOI220     m804(.A0(mai_mai_n826_), .A1(mai_mai_n426_), .B0(mai_mai_n824_), .B1(mai_mai_n65_), .Y(mai_mai_n827_));
  NO2        m805(.A(mai_mai_n67_), .B(mai_mai_n674_), .Y(mai_mai_n828_));
  AOI210     m806(.A0(mai_mai_n165_), .A1(i_10_), .B0(mai_mai_n828_), .Y(mai_mai_n829_));
  NO2        m807(.A(mai_mai_n829_), .B(mai_mai_n47_), .Y(mai_mai_n830_));
  NO3        m808(.A(i_5_), .B(mai_mai_n321_), .C(mai_mai_n24_), .Y(mai_mai_n831_));
  NO2        m809(.A(mai_mai_n492_), .B(mai_mai_n831_), .Y(mai_mai_n832_));
  NAi21      m810(.An(i_9_), .B(i_5_), .Y(mai_mai_n833_));
  NO2        m811(.A(mai_mai_n833_), .B(mai_mai_n367_), .Y(mai_mai_n834_));
  NO2        m812(.A(mai_mai_n541_), .B(mai_mai_n96_), .Y(mai_mai_n835_));
  AOI220     m813(.A0(mai_mai_n835_), .A1(i_0_), .B0(mai_mai_n834_), .B1(mai_mai_n559_), .Y(mai_mai_n836_));
  OAI220     m814(.A0(mai_mai_n836_), .A1(mai_mai_n77_), .B0(mai_mai_n832_), .B1(mai_mai_n163_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n837_), .B(mai_mai_n830_), .Y(mai_mai_n838_));
  NA2        m816(.A(mai_mai_n838_), .B(mai_mai_n827_), .Y(mai_mai_n839_));
  NO3        m817(.A(mai_mai_n839_), .B(mai_mai_n821_), .C(mai_mai_n793_), .Y(mai_mai_n840_));
  NO2        m818(.A(i_0_), .B(mai_mai_n653_), .Y(mai_mai_n841_));
  NA2        m819(.A(mai_mai_n65_), .B(mai_mai_n44_), .Y(mai_mai_n842_));
  NA2        m820(.A(mai_mai_n785_), .B(mai_mai_n842_), .Y(mai_mai_n843_));
  NO2        m821(.A(i_5_), .B(mai_mai_n25_), .Y(mai_mai_n844_));
  AO220      m822(.A0(mai_mai_n844_), .A1(mai_mai_n843_), .B0(mai_mai_n841_), .B1(mai_mai_n165_), .Y(mai_mai_n845_));
  NO2        m823(.A(mai_mai_n714_), .B(mai_mai_n809_), .Y(mai_mai_n846_));
  AOI210     m824(.A0(mai_mai_n845_), .A1(mai_mai_n312_), .B0(mai_mai_n846_), .Y(mai_mai_n847_));
  NA3        m825(.A(mai_mai_n138_), .B(mai_mai_n604_), .C(mai_mai_n65_), .Y(mai_mai_n848_));
  NO2        m826(.A(mai_mai_n726_), .B(mai_mai_n367_), .Y(mai_mai_n849_));
  NA3        m827(.A(mai_mai_n752_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n850_));
  NA2        m828(.A(mai_mai_n753_), .B(i_9_), .Y(mai_mai_n851_));
  AOI210     m829(.A0(mai_mai_n850_), .A1(mai_mai_n446_), .B0(mai_mai_n851_), .Y(mai_mai_n852_));
  NA2        m830(.A(mai_mai_n227_), .B(mai_mai_n215_), .Y(mai_mai_n853_));
  AOI210     m831(.A0(mai_mai_n853_), .A1(mai_mai_n780_), .B0(mai_mai_n144_), .Y(mai_mai_n854_));
  NO3        m832(.A(mai_mai_n854_), .B(mai_mai_n852_), .C(mai_mai_n849_), .Y(mai_mai_n855_));
  NA3        m833(.A(mai_mai_n855_), .B(mai_mai_n848_), .C(mai_mai_n847_), .Y(mai_mai_n856_));
  NA3        m834(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n857_));
  NA2        m835(.A(mai_mai_n797_), .B(mai_mai_n438_), .Y(mai_mai_n858_));
  AOI210     m836(.A0(mai_mai_n857_), .A1(mai_mai_n152_), .B0(mai_mai_n858_), .Y(mai_mai_n859_));
  INV        m837(.A(mai_mai_n859_), .Y(mai_mai_n860_));
  NA2        m838(.A(mai_mai_n513_), .B(mai_mai_n67_), .Y(mai_mai_n861_));
  NO3        m839(.A(mai_mai_n197_), .B(mai_mai_n349_), .C(i_0_), .Y(mai_mai_n862_));
  OAI210     m840(.A0(mai_mai_n862_), .A1(mai_mai_n68_), .B0(i_13_), .Y(mai_mai_n863_));
  INV        m841(.A(mai_mai_n205_), .Y(mai_mai_n864_));
  OAI220     m842(.A0(mai_mai_n477_), .A1(mai_mai_n131_), .B0(mai_mai_n578_), .B1(mai_mai_n553_), .Y(mai_mai_n865_));
  NA3        m843(.A(mai_mai_n865_), .B(i_7_), .C(mai_mai_n864_), .Y(mai_mai_n866_));
  NA4        m844(.A(mai_mai_n866_), .B(mai_mai_n863_), .C(mai_mai_n861_), .D(mai_mai_n860_), .Y(mai_mai_n867_));
  NO2        m845(.A(mai_mai_n226_), .B(mai_mai_n84_), .Y(mai_mai_n868_));
  AOI210     m846(.A0(mai_mai_n868_), .A1(mai_mai_n841_), .B0(mai_mai_n100_), .Y(mai_mai_n869_));
  NA2        m847(.A(mai_mai_n814_), .B(mai_mai_n438_), .Y(mai_mai_n870_));
  INV        m848(.A(mai_mai_n167_), .Y(mai_mai_n871_));
  OA220      m849(.A0(mai_mai_n871_), .A1(mai_mai_n870_), .B0(mai_mai_n869_), .B1(i_5_), .Y(mai_mai_n872_));
  AOI210     m850(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n166_), .Y(mai_mai_n873_));
  NA2        m851(.A(mai_mai_n873_), .B(mai_mai_n822_), .Y(mai_mai_n874_));
  NA3        m852(.A(mai_mai_n797_), .B(mai_mai_n257_), .C(mai_mai_n215_), .Y(mai_mai_n875_));
  INV        m853(.A(mai_mai_n875_), .Y(mai_mai_n876_));
  NA3        m854(.A(mai_mai_n356_), .B(mai_mai_n300_), .C(mai_mai_n207_), .Y(mai_mai_n877_));
  INV        m855(.A(mai_mai_n877_), .Y(mai_mai_n878_));
  NOi31      m856(.An(mai_mai_n355_), .B(mai_mai_n842_), .C(mai_mai_n223_), .Y(mai_mai_n879_));
  NO3        m857(.A(mai_mai_n794_), .B(mai_mai_n205_), .C(mai_mai_n181_), .Y(mai_mai_n880_));
  NO4        m858(.A(mai_mai_n880_), .B(mai_mai_n879_), .C(mai_mai_n878_), .D(mai_mai_n876_), .Y(mai_mai_n881_));
  NA4        m859(.A(mai_mai_n881_), .B(mai_mai_n423_), .C(mai_mai_n874_), .D(mai_mai_n872_), .Y(mai_mai_n882_));
  NA3        m860(.A(mai_mai_n272_), .B(i_5_), .C(mai_mai_n184_), .Y(mai_mai_n883_));
  NA2        m861(.A(mai_mai_n883_), .B(mai_mai_n226_), .Y(mai_mai_n884_));
  NO4        m862(.A(mai_mai_n223_), .B(mai_mai_n197_), .C(i_0_), .D(i_12_), .Y(mai_mai_n885_));
  AOI220     m863(.A0(mai_mai_n885_), .A1(mai_mai_n884_), .B0(mai_mai_n709_), .B1(mai_mai_n167_), .Y(mai_mai_n886_));
  AN2        m864(.A(mai_mai_n785_), .B(mai_mai_n144_), .Y(mai_mai_n887_));
  NO3        m865(.A(mai_mai_n887_), .B(i_12_), .C(mai_mai_n580_), .Y(mai_mai_n888_));
  INV        m866(.A(mai_mai_n888_), .Y(mai_mai_n889_));
  NA3        m867(.A(mai_mai_n89_), .B(mai_mai_n517_), .C(i_11_), .Y(mai_mai_n890_));
  NA2        m868(.A(mai_mai_n814_), .B(mai_mai_n422_), .Y(mai_mai_n891_));
  OAI220     m869(.A0(i_7_), .A1(mai_mai_n883_), .B0(mai_mai_n891_), .B1(i_1_), .Y(mai_mai_n892_));
  NA2        m870(.A(mai_mai_n892_), .B(mai_mai_n801_), .Y(mai_mai_n893_));
  NA3        m871(.A(mai_mai_n893_), .B(mai_mai_n889_), .C(mai_mai_n886_), .Y(mai_mai_n894_));
  NO4        m872(.A(mai_mai_n894_), .B(mai_mai_n882_), .C(mai_mai_n867_), .D(mai_mai_n856_), .Y(mai_mai_n895_));
  OAI210     m873(.A0(mai_mai_n729_), .A1(mai_mai_n724_), .B0(mai_mai_n37_), .Y(mai_mai_n896_));
  NA3        m874(.A(mai_mai_n808_), .B(mai_mai_n334_), .C(i_5_), .Y(mai_mai_n897_));
  NA3        m875(.A(mai_mai_n897_), .B(mai_mai_n896_), .C(mai_mai_n937_), .Y(mai_mai_n898_));
  NA2        m876(.A(mai_mai_n898_), .B(mai_mai_n195_), .Y(mai_mai_n899_));
  NA2        m877(.A(mai_mai_n178_), .B(mai_mai_n180_), .Y(mai_mai_n900_));
  AO210      m878(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n900_), .Y(mai_mai_n901_));
  OAI210     m879(.A0(mai_mai_n552_), .A1(mai_mai_n550_), .B0(mai_mai_n283_), .Y(mai_mai_n902_));
  NA2        m880(.A(mai_mai_n902_), .B(mai_mai_n901_), .Y(mai_mai_n903_));
  NA2        m881(.A(mai_mai_n890_), .B(mai_mai_n413_), .Y(mai_mai_n904_));
  AOI210     m882(.A0(mai_mai_n903_), .A1(mai_mai_n48_), .B0(mai_mai_n904_), .Y(mai_mai_n905_));
  AOI210     m883(.A0(mai_mai_n905_), .A1(mai_mai_n899_), .B0(mai_mai_n65_), .Y(mai_mai_n906_));
  NO2        m884(.A(mai_mai_n510_), .B(mai_mai_n345_), .Y(mai_mai_n907_));
  NO2        m885(.A(mai_mai_n907_), .B(mai_mai_n679_), .Y(mai_mai_n908_));
  INV        m886(.A(mai_mai_n68_), .Y(mai_mai_n909_));
  AOI210     m887(.A0(mai_mai_n873_), .A1(mai_mai_n797_), .B0(mai_mai_n815_), .Y(mai_mai_n910_));
  AOI210     m888(.A0(mai_mai_n910_), .A1(mai_mai_n909_), .B0(mai_mai_n605_), .Y(mai_mai_n911_));
  NA2        m889(.A(i_8_), .B(mai_mai_n68_), .Y(mai_mai_n912_));
  NO2        m890(.A(mai_mai_n912_), .B(mai_mai_n221_), .Y(mai_mai_n913_));
  NO2        m891(.A(mai_mai_n913_), .B(mai_mai_n911_), .Y(mai_mai_n914_));
  OAI210     m892(.A0(mai_mai_n243_), .A1(mai_mai_n148_), .B0(mai_mai_n80_), .Y(mai_mai_n915_));
  NA3        m893(.A(mai_mai_n682_), .B(mai_mai_n257_), .C(mai_mai_n72_), .Y(mai_mai_n916_));
  AOI210     m894(.A0(mai_mai_n916_), .A1(mai_mai_n915_), .B0(i_11_), .Y(mai_mai_n917_));
  OAI210     m895(.A0(mai_mai_n935_), .A1(mai_mai_n808_), .B0(mai_mai_n195_), .Y(mai_mai_n918_));
  NA2        m896(.A(mai_mai_n154_), .B(i_5_), .Y(mai_mai_n919_));
  AOI210     m897(.A0(mai_mai_n918_), .A1(mai_mai_n690_), .B0(mai_mai_n919_), .Y(mai_mai_n920_));
  NA2        m898(.A(mai_mai_n819_), .B(mai_mai_n939_), .Y(mai_mai_n921_));
  NO2        m899(.A(mai_mai_n921_), .B(mai_mai_n653_), .Y(mai_mai_n922_));
  NO3        m900(.A(mai_mai_n833_), .B(mai_mai_n429_), .C(mai_mai_n233_), .Y(mai_mai_n923_));
  NO2        m901(.A(mai_mai_n923_), .B(mai_mai_n507_), .Y(mai_mai_n924_));
  INV        m902(.A(mai_mai_n327_), .Y(mai_mai_n925_));
  AOI210     m903(.A0(mai_mai_n925_), .A1(mai_mai_n924_), .B0(mai_mai_n41_), .Y(mai_mai_n926_));
  NO4        m904(.A(mai_mai_n926_), .B(mai_mai_n922_), .C(mai_mai_n920_), .D(mai_mai_n917_), .Y(mai_mai_n927_));
  OAI210     m905(.A0(mai_mai_n914_), .A1(i_4_), .B0(mai_mai_n927_), .Y(mai_mai_n928_));
  NO3        m906(.A(mai_mai_n928_), .B(mai_mai_n908_), .C(mai_mai_n906_), .Y(mai_mai_n929_));
  NA4        m907(.A(mai_mai_n929_), .B(mai_mai_n895_), .C(mai_mai_n840_), .D(mai_mai_n773_), .Y(mai4));
  INV        m908(.A(i_2_), .Y(mai_mai_n933_));
  INV        m909(.A(mai_mai_n760_), .Y(mai_mai_n934_));
  INV        m910(.A(i_12_), .Y(mai_mai_n935_));
  INV        m911(.A(mai_mai_n74_), .Y(mai_mai_n936_));
  INV        m912(.A(mai_mai_n151_), .Y(mai_mai_n937_));
  INV        m913(.A(mai_mai_n763_), .Y(mai_mai_n938_));
  INV        m914(.A(i_4_), .Y(mai_mai_n939_));
  INV        m915(.A(mai_mai_n229_), .Y(mai_mai_n940_));
  INV        m916(.A(mai_mai_n134_), .Y(mai_mai_n941_));
  INV        m917(.A(i_0_), .Y(mai_mai_n942_));
  INV        m918(.A(mai_mai_n378_), .Y(mai_mai_n943_));
  INV        m919(.A(i_3_), .Y(mai_mai_n944_));
  INV        m920(.A(i_6_), .Y(mai_mai_n945_));
  INV        m921(.A(mai_mai_n31_), .Y(mai_mai_n946_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  OAI210     u0028(.A0(men_men_n50_), .A1(i_3_), .B0(men_men_n48_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  INV        u0037(.A(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(men_men_n65_), .B(men_men_n61_), .Y(men_men_n66_));
  NA2        u0044(.A(men_men_n50_), .B(i_2_), .Y(men_men_n67_));
  AOI210     u0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n68_));
  NA2        u0046(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO2        u0047(.A(men_men_n69_), .B(men_men_n25_), .Y(men_men_n70_));
  INV        u0048(.A(i_0_), .Y(men_men_n71_));
  NAi21      u0049(.An(i_5_), .B(i_10_), .Y(men_men_n72_));
  NA2        u0050(.A(i_5_), .B(i_9_), .Y(men_men_n73_));
  AOI210     u0051(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n71_), .Y(men_men_n74_));
  NO2        u0052(.A(men_men_n74_), .B(men_men_n70_), .Y(men_men_n75_));
  OAI210     u0053(.A0(men_men_n68_), .A1(men_men_n67_), .B0(men_men_n75_), .Y(men_men_n76_));
  OAI210     u0054(.A0(men_men_n76_), .A1(men_men_n66_), .B0(i_0_), .Y(men_men_n77_));
  NA2        u0055(.A(i_12_), .B(i_5_), .Y(men_men_n78_));
  NA2        u0056(.A(i_2_), .B(i_8_), .Y(men_men_n79_));
  NO2        u0057(.A(i_3_), .B(i_9_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_7_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n63_), .Y(men_men_n82_));
  INV        u0060(.A(i_6_), .Y(men_men_n83_));
  OR4        u0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n84_));
  NO2        u0062(.A(i_2_), .B(i_7_), .Y(men_men_n85_));
  NA2        u0063(.A(men_men_n82_), .B(men_men_n84_), .Y(men_men_n86_));
  NAi21      u0064(.An(i_6_), .B(i_10_), .Y(men_men_n87_));
  NA2        u0065(.A(i_6_), .B(i_9_), .Y(men_men_n88_));
  NO2        u0066(.A(men_men_n87_), .B(men_men_n63_), .Y(men_men_n89_));
  NA2        u0067(.A(i_2_), .B(i_6_), .Y(men_men_n90_));
  NO3        u0068(.A(men_men_n90_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n91_));
  INV        u0069(.A(men_men_n91_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n92_), .A1(men_men_n86_), .B0(men_men_n78_), .Y(men_men_n93_));
  AN3        u0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n94_));
  NAi21      u0072(.An(i_6_), .B(i_11_), .Y(men_men_n95_));
  NO2        u0073(.A(i_5_), .B(i_8_), .Y(men_men_n96_));
  NOi21      u0074(.An(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  NA2        u0075(.A(men_men_n94_), .B(men_men_n32_), .Y(men_men_n98_));
  INV        u0076(.A(i_7_), .Y(men_men_n99_));
  NO2        u0077(.A(i_0_), .B(i_5_), .Y(men_men_n100_));
  NO2        u0078(.A(men_men_n100_), .B(men_men_n83_), .Y(men_men_n101_));
  NA2        u0079(.A(i_12_), .B(i_3_), .Y(men_men_n102_));
  INV        u0080(.A(men_men_n102_), .Y(men_men_n103_));
  NAi21      u0081(.An(i_7_), .B(i_11_), .Y(men_men_n104_));
  NO3        u0082(.A(men_men_n104_), .B(men_men_n87_), .C(men_men_n53_), .Y(men_men_n105_));
  AN2        u0083(.A(i_2_), .B(i_10_), .Y(men_men_n106_));
  NO2        u0084(.A(men_men_n106_), .B(i_7_), .Y(men_men_n107_));
  OR2        u0085(.A(men_men_n78_), .B(men_men_n58_), .Y(men_men_n108_));
  NO2        u0086(.A(i_8_), .B(men_men_n99_), .Y(men_men_n109_));
  NO3        u0087(.A(men_men_n109_), .B(men_men_n108_), .C(men_men_n107_), .Y(men_men_n110_));
  NA2        u0088(.A(i_12_), .B(i_7_), .Y(men_men_n111_));
  NA2        u0089(.A(i_1_), .B(i_0_), .Y(men_men_n112_));
  NA2        u0090(.A(i_11_), .B(i_12_), .Y(men_men_n113_));
  OAI210     u0091(.A0(men_men_n112_), .A1(men_men_n111_), .B0(men_men_n113_), .Y(men_men_n114_));
  NO2        u0092(.A(men_men_n114_), .B(men_men_n110_), .Y(men_men_n115_));
  NAi31      u0093(.An(men_men_n105_), .B(men_men_n115_), .C(men_men_n98_), .Y(men_men_n116_));
  NOi21      u0094(.An(i_1_), .B(i_5_), .Y(men_men_n117_));
  NA2        u0095(.A(men_men_n117_), .B(i_11_), .Y(men_men_n118_));
  NA2        u0096(.A(men_men_n99_), .B(men_men_n37_), .Y(men_men_n119_));
  NA2        u0097(.A(i_7_), .B(men_men_n25_), .Y(men_men_n120_));
  NA2        u0098(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NO2        u0099(.A(men_men_n121_), .B(men_men_n46_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n88_), .B(men_men_n87_), .Y(men_men_n123_));
  NAi21      u0101(.An(i_3_), .B(i_8_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(men_men_n62_), .Y(men_men_n125_));
  NOi31      u0103(.An(men_men_n125_), .B(men_men_n123_), .C(men_men_n122_), .Y(men_men_n126_));
  NO2        u0104(.A(i_1_), .B(men_men_n83_), .Y(men_men_n127_));
  NO2        u0105(.A(i_6_), .B(i_5_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(i_3_), .Y(men_men_n129_));
  NO2        u0107(.A(men_men_n126_), .B(men_men_n118_), .Y(men_men_n130_));
  NO3        u0108(.A(men_men_n130_), .B(men_men_n116_), .C(men_men_n93_), .Y(men_men_n131_));
  NA3        u0109(.A(men_men_n131_), .B(men_men_n77_), .C(men_men_n56_), .Y(men2));
  NO2        u0110(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n133_));
  INV        u0111(.A(i_6_), .Y(men_men_n134_));
  NA2        u0112(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NA4        u0113(.A(men_men_n135_), .B(men_men_n75_), .C(men_men_n67_), .D(men_men_n30_), .Y(men0));
  AN2        u0114(.A(i_8_), .B(i_7_), .Y(men_men_n137_));
  NA2        u0115(.A(men_men_n137_), .B(i_6_), .Y(men_men_n138_));
  NO2        u0116(.A(i_12_), .B(i_13_), .Y(men_men_n139_));
  NAi21      u0117(.An(i_5_), .B(i_11_), .Y(men_men_n140_));
  NOi21      u0118(.An(men_men_n139_), .B(men_men_n140_), .Y(men_men_n141_));
  NO2        u0119(.A(i_0_), .B(i_1_), .Y(men_men_n142_));
  NA2        u0120(.A(i_2_), .B(i_3_), .Y(men_men_n143_));
  NO2        u0121(.A(men_men_n143_), .B(i_4_), .Y(men_men_n144_));
  NA3        u0122(.A(men_men_n144_), .B(men_men_n142_), .C(men_men_n141_), .Y(men_men_n145_));
  OR2        u0123(.A(men_men_n145_), .B(men_men_n25_), .Y(men_men_n146_));
  AN2        u0124(.A(men_men_n139_), .B(men_men_n80_), .Y(men_men_n147_));
  NO2        u0125(.A(men_men_n147_), .B(men_men_n27_), .Y(men_men_n148_));
  NA2        u0126(.A(i_1_), .B(i_5_), .Y(men_men_n149_));
  NO2        u0127(.A(men_men_n71_), .B(men_men_n46_), .Y(men_men_n150_));
  NA2        u0128(.A(men_men_n150_), .B(men_men_n36_), .Y(men_men_n151_));
  NO3        u0129(.A(men_men_n151_), .B(men_men_n149_), .C(men_men_n148_), .Y(men_men_n152_));
  OR2        u0130(.A(i_0_), .B(i_1_), .Y(men_men_n153_));
  NO3        u0131(.A(men_men_n153_), .B(men_men_n78_), .C(i_13_), .Y(men_men_n154_));
  NAi32      u0132(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n155_));
  NAi21      u0133(.An(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  NOi21      u0134(.An(i_4_), .B(i_10_), .Y(men_men_n157_));
  NA2        u0135(.A(men_men_n157_), .B(men_men_n39_), .Y(men_men_n158_));
  NO2        u0136(.A(i_3_), .B(i_5_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n71_), .B(i_2_), .C(i_1_), .Y(men_men_n160_));
  OAI210     u0138(.A0(i_2_), .A1(men_men_n158_), .B0(men_men_n156_), .Y(men_men_n161_));
  NO2        u0139(.A(men_men_n161_), .B(men_men_n152_), .Y(men_men_n162_));
  AOI210     u0140(.A0(men_men_n162_), .A1(men_men_n146_), .B0(men_men_n138_), .Y(men_men_n163_));
  NOi21      u0141(.An(i_4_), .B(i_9_), .Y(men_men_n164_));
  NOi21      u0142(.An(i_11_), .B(i_13_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  NO2        u0144(.A(i_4_), .B(i_5_), .Y(men_men_n167_));
  NAi21      u0145(.An(i_12_), .B(i_11_), .Y(men_men_n168_));
  NO2        u0146(.A(men_men_n168_), .B(i_13_), .Y(men_men_n169_));
  NA3        u0147(.A(men_men_n169_), .B(men_men_n167_), .C(men_men_n80_), .Y(men_men_n170_));
  AOI210     u0148(.A0(men_men_n170_), .A1(men_men_n166_), .B0(i_2_), .Y(men_men_n171_));
  NO2        u0149(.A(men_men_n71_), .B(men_men_n63_), .Y(men_men_n172_));
  NA2        u0150(.A(men_men_n172_), .B(men_men_n46_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n36_), .B(i_5_), .Y(men_men_n174_));
  NAi31      u0152(.An(men_men_n174_), .B(men_men_n147_), .C(i_11_), .Y(men_men_n175_));
  NA2        u0153(.A(i_3_), .B(i_5_), .Y(men_men_n176_));
  AOI210     u0154(.A0(men_men_n166_), .A1(men_men_n175_), .B0(men_men_n173_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n71_), .B(i_5_), .Y(men_men_n178_));
  NO2        u0156(.A(i_13_), .B(i_10_), .Y(men_men_n179_));
  NA3        u0157(.A(men_men_n179_), .B(men_men_n178_), .C(men_men_n44_), .Y(men_men_n180_));
  NO2        u0158(.A(i_2_), .B(i_1_), .Y(men_men_n181_));
  NA2        u0159(.A(men_men_n181_), .B(i_3_), .Y(men_men_n182_));
  NAi21      u0160(.An(i_4_), .B(i_12_), .Y(men_men_n183_));
  NO4        u0161(.A(men_men_n183_), .B(men_men_n182_), .C(men_men_n180_), .D(men_men_n25_), .Y(men_men_n184_));
  NO3        u0162(.A(men_men_n184_), .B(men_men_n177_), .C(men_men_n171_), .Y(men_men_n185_));
  INV        u0163(.A(i_8_), .Y(men_men_n186_));
  NO2        u0164(.A(men_men_n186_), .B(i_7_), .Y(men_men_n187_));
  NA2        u0165(.A(men_men_n187_), .B(i_6_), .Y(men_men_n188_));
  NO3        u0166(.A(i_3_), .B(men_men_n83_), .C(men_men_n48_), .Y(men_men_n189_));
  NA2        u0167(.A(men_men_n189_), .B(men_men_n109_), .Y(men_men_n190_));
  NO3        u0168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n191_));
  NA3        u0169(.A(men_men_n191_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n192_));
  NO3        u0170(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n193_));
  OAI210     u0171(.A0(men_men_n94_), .A1(i_12_), .B0(men_men_n193_), .Y(men_men_n194_));
  AOI210     u0172(.A0(men_men_n194_), .A1(men_men_n192_), .B0(men_men_n190_), .Y(men_men_n195_));
  NO2        u0173(.A(i_3_), .B(i_8_), .Y(men_men_n196_));
  NO3        u0174(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n197_));
  NA3        u0175(.A(men_men_n197_), .B(men_men_n196_), .C(men_men_n39_), .Y(men_men_n198_));
  NO2        u0176(.A(men_men_n100_), .B(men_men_n58_), .Y(men_men_n199_));
  NO2        u0177(.A(i_13_), .B(i_9_), .Y(men_men_n200_));
  NA3        u0178(.A(men_men_n200_), .B(i_6_), .C(men_men_n186_), .Y(men_men_n201_));
  NAi21      u0179(.An(i_12_), .B(i_3_), .Y(men_men_n202_));
  OR2        u0180(.A(men_men_n202_), .B(men_men_n201_), .Y(men_men_n203_));
  NO2        u0181(.A(men_men_n44_), .B(i_5_), .Y(men_men_n204_));
  NO3        u0182(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n205_));
  OAI220     u0183(.A0(i_2_), .A1(men_men_n203_), .B0(men_men_n100_), .B1(men_men_n198_), .Y(men_men_n206_));
  AOI210     u0184(.A0(men_men_n206_), .A1(i_7_), .B0(men_men_n195_), .Y(men_men_n207_));
  OAI220     u0185(.A0(men_men_n207_), .A1(i_4_), .B0(men_men_n188_), .B1(men_men_n185_), .Y(men_men_n208_));
  NAi21      u0186(.An(i_12_), .B(i_7_), .Y(men_men_n209_));
  NA3        u0187(.A(i_13_), .B(men_men_n186_), .C(i_10_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n210_), .B(men_men_n209_), .Y(men_men_n211_));
  NA2        u0189(.A(i_0_), .B(i_5_), .Y(men_men_n212_));
  NA2        u0190(.A(men_men_n212_), .B(men_men_n101_), .Y(men_men_n213_));
  OAI220     u0191(.A0(men_men_n213_), .A1(men_men_n182_), .B0(men_men_n173_), .B1(men_men_n129_), .Y(men_men_n214_));
  NAi31      u0192(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n215_));
  NO2        u0193(.A(men_men_n36_), .B(i_13_), .Y(men_men_n216_));
  NO2        u0194(.A(men_men_n71_), .B(men_men_n26_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n218_));
  NA3        u0196(.A(men_men_n218_), .B(men_men_n217_), .C(men_men_n216_), .Y(men_men_n219_));
  INV        u0197(.A(i_13_), .Y(men_men_n220_));
  NO2        u0198(.A(i_12_), .B(men_men_n220_), .Y(men_men_n221_));
  NA3        u0199(.A(men_men_n221_), .B(men_men_n191_), .C(men_men_n189_), .Y(men_men_n222_));
  OAI210     u0200(.A0(men_men_n219_), .A1(men_men_n215_), .B0(men_men_n222_), .Y(men_men_n223_));
  AOI220     u0201(.A0(men_men_n223_), .A1(men_men_n137_), .B0(men_men_n214_), .B1(men_men_n211_), .Y(men_men_n224_));
  NO2        u0202(.A(i_12_), .B(men_men_n37_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n176_), .B(i_4_), .Y(men_men_n226_));
  INV        u0204(.A(men_men_n226_), .Y(men_men_n227_));
  OR2        u0205(.A(i_8_), .B(i_7_), .Y(men_men_n228_));
  NO2        u0206(.A(men_men_n228_), .B(men_men_n83_), .Y(men_men_n229_));
  NO2        u0207(.A(men_men_n53_), .B(i_1_), .Y(men_men_n230_));
  NA2        u0208(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n231_));
  INV        u0209(.A(i_12_), .Y(men_men_n232_));
  NO3        u0210(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n233_));
  NA2        u0211(.A(i_2_), .B(i_1_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n231_), .B(men_men_n227_), .Y(men_men_n235_));
  NAi21      u0213(.An(i_4_), .B(i_3_), .Y(men_men_n236_));
  NO2        u0214(.A(men_men_n236_), .B(men_men_n73_), .Y(men_men_n237_));
  NO2        u0215(.A(i_0_), .B(i_6_), .Y(men_men_n238_));
  NOi41      u0216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n234_), .B(men_men_n176_), .Y(men_men_n241_));
  NAi21      u0219(.An(men_men_n240_), .B(men_men_n241_), .Y(men_men_n242_));
  INV        u0220(.A(men_men_n242_), .Y(men_men_n243_));
  AOI220     u0221(.A0(men_men_n243_), .A1(men_men_n39_), .B0(men_men_n235_), .B1(men_men_n200_), .Y(men_men_n244_));
  NO2        u0222(.A(i_11_), .B(men_men_n220_), .Y(men_men_n245_));
  NOi21      u0223(.An(i_1_), .B(i_6_), .Y(men_men_n246_));
  NAi21      u0224(.An(i_3_), .B(i_7_), .Y(men_men_n247_));
  NA2        u0225(.A(men_men_n232_), .B(i_9_), .Y(men_men_n248_));
  OR4        u0226(.A(men_men_n248_), .B(men_men_n247_), .C(men_men_n246_), .D(men_men_n178_), .Y(men_men_n249_));
  NO2        u0227(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n250_));
  NO2        u0228(.A(i_12_), .B(i_3_), .Y(men_men_n251_));
  NA2        u0229(.A(men_men_n71_), .B(i_5_), .Y(men_men_n252_));
  NA2        u0230(.A(i_3_), .B(i_9_), .Y(men_men_n253_));
  NAi21      u0231(.An(i_7_), .B(i_10_), .Y(men_men_n254_));
  NO2        u0232(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NA3        u0233(.A(men_men_n255_), .B(men_men_n252_), .C(men_men_n64_), .Y(men_men_n256_));
  NA2        u0234(.A(men_men_n256_), .B(men_men_n249_), .Y(men_men_n257_));
  NA3        u0235(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n258_));
  NA2        u0236(.A(men_men_n257_), .B(men_men_n245_), .Y(men_men_n259_));
  NO2        u0237(.A(men_men_n228_), .B(men_men_n37_), .Y(men_men_n260_));
  NA2        u0238(.A(i_12_), .B(i_6_), .Y(men_men_n261_));
  OR2        u0239(.A(i_13_), .B(i_9_), .Y(men_men_n262_));
  NO3        u0240(.A(men_men_n262_), .B(men_men_n261_), .C(men_men_n48_), .Y(men_men_n263_));
  NO2        u0241(.A(men_men_n236_), .B(i_2_), .Y(men_men_n264_));
  NA3        u0242(.A(men_men_n264_), .B(men_men_n263_), .C(men_men_n44_), .Y(men_men_n265_));
  NA2        u0243(.A(men_men_n245_), .B(i_9_), .Y(men_men_n266_));
  OAI210     u0244(.A0(men_men_n71_), .A1(men_men_n266_), .B0(men_men_n265_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n150_), .B(men_men_n63_), .Y(men_men_n268_));
  NO3        u0246(.A(i_11_), .B(men_men_n220_), .C(men_men_n25_), .Y(men_men_n269_));
  NO2        u0247(.A(men_men_n247_), .B(i_8_), .Y(men_men_n270_));
  NO2        u0248(.A(i_6_), .B(men_men_n48_), .Y(men_men_n271_));
  NA3        u0249(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n269_), .Y(men_men_n272_));
  NO3        u0250(.A(men_men_n26_), .B(men_men_n83_), .C(i_5_), .Y(men_men_n273_));
  NA3        u0251(.A(men_men_n273_), .B(men_men_n260_), .C(men_men_n221_), .Y(men_men_n274_));
  AOI210     u0252(.A0(men_men_n274_), .A1(men_men_n272_), .B0(men_men_n268_), .Y(men_men_n275_));
  AOI210     u0253(.A0(men_men_n267_), .A1(men_men_n260_), .B0(men_men_n275_), .Y(men_men_n276_));
  NA4        u0254(.A(men_men_n276_), .B(men_men_n259_), .C(men_men_n244_), .D(men_men_n224_), .Y(men_men_n277_));
  NO3        u0255(.A(i_12_), .B(men_men_n220_), .C(men_men_n37_), .Y(men_men_n278_));
  INV        u0256(.A(men_men_n278_), .Y(men_men_n279_));
  NOi21      u0257(.An(men_men_n159_), .B(men_men_n83_), .Y(men_men_n280_));
  NO3        u0258(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n281_));
  AOI220     u0259(.A0(men_men_n281_), .A1(men_men_n189_), .B0(men_men_n280_), .B1(men_men_n230_), .Y(men_men_n282_));
  NO2        u0260(.A(men_men_n282_), .B(i_7_), .Y(men_men_n283_));
  NO3        u0261(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n284_));
  NO2        u0262(.A(men_men_n234_), .B(i_0_), .Y(men_men_n285_));
  AOI220     u0263(.A0(men_men_n285_), .A1(men_men_n187_), .B0(men_men_n284_), .B1(men_men_n137_), .Y(men_men_n286_));
  NA2        u0264(.A(men_men_n271_), .B(men_men_n26_), .Y(men_men_n287_));
  NO2        u0265(.A(men_men_n287_), .B(men_men_n286_), .Y(men_men_n288_));
  NA2        u0266(.A(i_0_), .B(i_1_), .Y(men_men_n289_));
  NO2        u0267(.A(men_men_n289_), .B(i_2_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n59_), .B(i_6_), .Y(men_men_n291_));
  NA3        u0269(.A(men_men_n291_), .B(men_men_n290_), .C(men_men_n159_), .Y(men_men_n292_));
  OAI210     u0270(.A0(i_2_), .A1(men_men_n138_), .B0(men_men_n292_), .Y(men_men_n293_));
  NO3        u0271(.A(men_men_n293_), .B(men_men_n288_), .C(men_men_n283_), .Y(men_men_n294_));
  NO2        u0272(.A(i_3_), .B(i_10_), .Y(men_men_n295_));
  NA3        u0273(.A(men_men_n295_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n296_));
  NO2        u0274(.A(i_2_), .B(men_men_n99_), .Y(men_men_n297_));
  NOi21      u0275(.An(men_men_n212_), .B(men_men_n100_), .Y(men_men_n298_));
  NA3        u0276(.A(men_men_n298_), .B(i_1_), .C(men_men_n297_), .Y(men_men_n299_));
  AN2        u0277(.A(i_3_), .B(i_10_), .Y(men_men_n300_));
  NA4        u0278(.A(men_men_n300_), .B(men_men_n191_), .C(men_men_n169_), .D(men_men_n167_), .Y(men_men_n301_));
  NO2        u0279(.A(i_5_), .B(men_men_n37_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n303_));
  OR2        u0281(.A(men_men_n299_), .B(men_men_n296_), .Y(men_men_n304_));
  OAI220     u0282(.A0(men_men_n304_), .A1(i_6_), .B0(men_men_n294_), .B1(men_men_n279_), .Y(men_men_n305_));
  NO4        u0283(.A(men_men_n305_), .B(men_men_n277_), .C(men_men_n208_), .D(men_men_n163_), .Y(men_men_n306_));
  NO3        u0284(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n307_));
  NO2        u0285(.A(men_men_n59_), .B(men_men_n83_), .Y(men_men_n308_));
  NA2        u0286(.A(men_men_n285_), .B(men_men_n308_), .Y(men_men_n309_));
  NO3        u0287(.A(i_6_), .B(men_men_n186_), .C(i_7_), .Y(men_men_n310_));
  AOI210     u0288(.A0(men_men_n1030_), .A1(men_men_n309_), .B0(i_5_), .Y(men_men_n311_));
  NO2        u0289(.A(i_2_), .B(i_3_), .Y(men_men_n312_));
  OR2        u0290(.A(i_0_), .B(i_5_), .Y(men_men_n313_));
  NA2        u0291(.A(men_men_n212_), .B(men_men_n313_), .Y(men_men_n314_));
  NA4        u0292(.A(men_men_n314_), .B(men_men_n229_), .C(men_men_n312_), .D(i_1_), .Y(men_men_n315_));
  NA2        u0293(.A(men_men_n285_), .B(men_men_n280_), .Y(men_men_n316_));
  NO2        u0294(.A(men_men_n153_), .B(men_men_n46_), .Y(men_men_n317_));
  NA2        u0295(.A(men_men_n317_), .B(men_men_n159_), .Y(men_men_n318_));
  NA3        u0296(.A(men_men_n318_), .B(men_men_n316_), .C(men_men_n315_), .Y(men_men_n319_));
  OAI210     u0297(.A0(men_men_n319_), .A1(men_men_n311_), .B0(i_4_), .Y(men_men_n320_));
  NO2        u0298(.A(i_12_), .B(i_10_), .Y(men_men_n321_));
  NOi21      u0299(.An(i_5_), .B(i_0_), .Y(men_men_n322_));
  AOI210     u0300(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n99_), .Y(men_men_n323_));
  NO4        u0301(.A(men_men_n323_), .B(i_4_), .C(men_men_n322_), .D(men_men_n124_), .Y(men_men_n324_));
  NA4        u0302(.A(men_men_n81_), .B(men_men_n36_), .C(men_men_n83_), .D(i_8_), .Y(men_men_n325_));
  NA2        u0303(.A(men_men_n324_), .B(men_men_n321_), .Y(men_men_n326_));
  NO2        u0304(.A(i_6_), .B(i_8_), .Y(men_men_n327_));
  AN2        u0305(.A(i_0_), .B(men_men_n327_), .Y(men_men_n328_));
  NO2        u0306(.A(i_1_), .B(i_7_), .Y(men_men_n329_));
  NA3        u0307(.A(i_0_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n330_), .B(men_men_n326_), .C(men_men_n320_), .Y(men_men_n331_));
  NA2        u0309(.A(men_men_n1026_), .B(i_6_), .Y(men_men_n332_));
  NA3        u0310(.A(men_men_n246_), .B(men_men_n297_), .C(men_men_n186_), .Y(men_men_n333_));
  AOI210     u0311(.A0(men_men_n333_), .A1(men_men_n332_), .B0(men_men_n314_), .Y(men_men_n334_));
  NOi21      u0312(.An(men_men_n149_), .B(men_men_n101_), .Y(men_men_n335_));
  NO2        u0313(.A(men_men_n335_), .B(men_men_n120_), .Y(men_men_n336_));
  OAI210     u0314(.A0(men_men_n336_), .A1(men_men_n334_), .B0(i_3_), .Y(men_men_n337_));
  NO2        u0315(.A(men_men_n289_), .B(men_men_n79_), .Y(men_men_n338_));
  NA2        u0316(.A(men_men_n338_), .B(men_men_n128_), .Y(men_men_n339_));
  NO2        u0317(.A(men_men_n90_), .B(men_men_n186_), .Y(men_men_n340_));
  NA3        u0318(.A(men_men_n298_), .B(men_men_n340_), .C(men_men_n63_), .Y(men_men_n341_));
  AOI210     u0319(.A0(men_men_n341_), .A1(men_men_n339_), .B0(i_3_), .Y(men_men_n342_));
  NO2        u0320(.A(men_men_n186_), .B(i_9_), .Y(men_men_n343_));
  NA2        u0321(.A(men_men_n343_), .B(men_men_n199_), .Y(men_men_n344_));
  NO2        u0322(.A(men_men_n342_), .B(men_men_n288_), .Y(men_men_n345_));
  AOI210     u0323(.A0(men_men_n345_), .A1(men_men_n337_), .B0(men_men_n158_), .Y(men_men_n346_));
  AOI210     u0324(.A0(men_men_n331_), .A1(men_men_n307_), .B0(men_men_n346_), .Y(men_men_n347_));
  NOi32      u0325(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n348_));
  INV        u0326(.A(men_men_n348_), .Y(men_men_n349_));
  NAi21      u0327(.An(i_0_), .B(i_6_), .Y(men_men_n350_));
  INV        u0328(.A(men_men_n350_), .Y(men_men_n351_));
  NA2        u0329(.A(men_men_n351_), .B(men_men_n25_), .Y(men_men_n352_));
  OAI210     u0330(.A0(men_men_n352_), .A1(men_men_n155_), .B0(men_men_n240_), .Y(men_men_n353_));
  NAi41      u0331(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n354_));
  NO2        u0332(.A(men_men_n215_), .B(men_men_n155_), .Y(men_men_n355_));
  AOI210     u0333(.A0(men_men_n354_), .A1(men_men_n155_), .B0(men_men_n153_), .Y(men_men_n356_));
  NOi32      u0334(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n357_));
  NAi21      u0335(.An(i_6_), .B(i_1_), .Y(men_men_n358_));
  NA3        u0336(.A(men_men_n358_), .B(men_men_n357_), .C(men_men_n46_), .Y(men_men_n359_));
  NO2        u0337(.A(men_men_n359_), .B(i_0_), .Y(men_men_n360_));
  OR3        u0338(.A(men_men_n360_), .B(men_men_n356_), .C(men_men_n355_), .Y(men_men_n361_));
  NO2        u0339(.A(i_1_), .B(men_men_n99_), .Y(men_men_n362_));
  NAi21      u0340(.An(i_3_), .B(i_4_), .Y(men_men_n363_));
  NO2        u0341(.A(men_men_n363_), .B(i_9_), .Y(men_men_n364_));
  AN2        u0342(.A(i_6_), .B(i_7_), .Y(men_men_n365_));
  OAI210     u0343(.A0(men_men_n365_), .A1(men_men_n362_), .B0(men_men_n364_), .Y(men_men_n366_));
  NA2        u0344(.A(i_2_), .B(i_7_), .Y(men_men_n367_));
  NO2        u0345(.A(men_men_n363_), .B(i_10_), .Y(men_men_n368_));
  NA3        u0346(.A(men_men_n368_), .B(men_men_n367_), .C(men_men_n238_), .Y(men_men_n369_));
  AOI210     u0347(.A0(men_men_n369_), .A1(men_men_n366_), .B0(men_men_n178_), .Y(men_men_n370_));
  AOI220     u0348(.A0(men_men_n368_), .A1(men_men_n329_), .B0(men_men_n233_), .B1(men_men_n181_), .Y(men_men_n371_));
  NO2        u0349(.A(men_men_n371_), .B(i_5_), .Y(men_men_n372_));
  NO4        u0350(.A(men_men_n372_), .B(men_men_n370_), .C(men_men_n361_), .D(men_men_n353_), .Y(men_men_n373_));
  NO2        u0351(.A(men_men_n373_), .B(men_men_n349_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n375_));
  AN2        u0353(.A(i_12_), .B(i_5_), .Y(men_men_n376_));
  NO2        u0354(.A(i_4_), .B(men_men_n26_), .Y(men_men_n377_));
  NA2        u0355(.A(men_men_n377_), .B(men_men_n376_), .Y(men_men_n378_));
  NO2        u0356(.A(i_11_), .B(i_6_), .Y(men_men_n379_));
  NA3        u0357(.A(men_men_n379_), .B(men_men_n317_), .C(men_men_n220_), .Y(men_men_n380_));
  NO2        u0358(.A(men_men_n380_), .B(men_men_n378_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n236_), .B(i_5_), .Y(men_men_n382_));
  NO2        u0360(.A(i_5_), .B(i_10_), .Y(men_men_n383_));
  AOI220     u0361(.A0(men_men_n383_), .A1(men_men_n264_), .B0(men_men_n382_), .B1(men_men_n191_), .Y(men_men_n384_));
  INV        u0362(.A(men_men_n45_), .Y(men_men_n385_));
  NO2        u0363(.A(men_men_n385_), .B(men_men_n384_), .Y(men_men_n386_));
  OAI210     u0364(.A0(men_men_n386_), .A1(men_men_n381_), .B0(men_men_n375_), .Y(men_men_n387_));
  NO2        u0365(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n388_));
  NO2        u0366(.A(men_men_n145_), .B(men_men_n83_), .Y(men_men_n389_));
  OAI210     u0367(.A0(men_men_n389_), .A1(men_men_n381_), .B0(men_men_n388_), .Y(men_men_n390_));
  NO3        u0368(.A(men_men_n83_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n391_));
  INV        u0369(.A(i_3_), .Y(men_men_n392_));
  NO2        u0370(.A(i_11_), .B(i_12_), .Y(men_men_n393_));
  NAi21      u0371(.An(i_13_), .B(i_0_), .Y(men_men_n394_));
  NA2        u0372(.A(men_men_n390_), .B(men_men_n387_), .Y(men_men_n395_));
  NA2        u0373(.A(men_men_n44_), .B(men_men_n220_), .Y(men_men_n396_));
  NO3        u0374(.A(i_1_), .B(i_12_), .C(men_men_n83_), .Y(men_men_n397_));
  NO2        u0375(.A(i_0_), .B(i_11_), .Y(men_men_n398_));
  AN2        u0376(.A(i_1_), .B(i_6_), .Y(men_men_n399_));
  NOi21      u0377(.An(i_2_), .B(i_12_), .Y(men_men_n400_));
  NA2        u0378(.A(men_men_n400_), .B(men_men_n399_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n401_), .B(men_men_n1022_), .Y(men_men_n402_));
  NA2        u0380(.A(men_men_n137_), .B(i_9_), .Y(men_men_n403_));
  NO2        u0381(.A(men_men_n403_), .B(i_4_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n402_), .B(men_men_n404_), .Y(men_men_n405_));
  NAi21      u0383(.An(i_9_), .B(i_4_), .Y(men_men_n406_));
  OR2        u0384(.A(i_13_), .B(i_10_), .Y(men_men_n407_));
  NO3        u0385(.A(men_men_n407_), .B(men_men_n113_), .C(men_men_n406_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n166_), .B(men_men_n119_), .Y(men_men_n409_));
  OR2        u0387(.A(men_men_n210_), .B(men_men_n209_), .Y(men_men_n410_));
  NO2        u0388(.A(men_men_n99_), .B(men_men_n25_), .Y(men_men_n411_));
  NA2        u0389(.A(men_men_n278_), .B(men_men_n411_), .Y(men_men_n412_));
  NA2        u0390(.A(men_men_n271_), .B(men_men_n205_), .Y(men_men_n413_));
  OAI220     u0391(.A0(men_men_n413_), .A1(men_men_n410_), .B0(men_men_n412_), .B1(men_men_n335_), .Y(men_men_n414_));
  INV        u0392(.A(men_men_n414_), .Y(men_men_n415_));
  AOI210     u0393(.A0(men_men_n415_), .A1(men_men_n405_), .B0(men_men_n26_), .Y(men_men_n416_));
  NA2        u0394(.A(men_men_n316_), .B(men_men_n315_), .Y(men_men_n417_));
  AOI220     u0395(.A0(men_men_n291_), .A1(men_men_n281_), .B0(men_men_n285_), .B1(men_men_n308_), .Y(men_men_n418_));
  NO2        u0396(.A(men_men_n418_), .B(i_5_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n176_), .B(men_men_n83_), .Y(men_men_n420_));
  AOI220     u0398(.A0(men_men_n420_), .A1(men_men_n290_), .B0(men_men_n273_), .B1(men_men_n205_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n421_), .B(i_7_), .Y(men_men_n422_));
  NO3        u0400(.A(men_men_n422_), .B(men_men_n419_), .C(men_men_n417_), .Y(men_men_n423_));
  NA2        u0401(.A(men_men_n189_), .B(men_men_n94_), .Y(men_men_n424_));
  NA3        u0402(.A(men_men_n317_), .B(men_men_n159_), .C(men_men_n83_), .Y(men_men_n425_));
  AOI210     u0403(.A0(men_men_n425_), .A1(men_men_n424_), .B0(i_8_), .Y(men_men_n426_));
  NA3        u0404(.A(men_men_n252_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n291_), .B(men_men_n230_), .Y(men_men_n428_));
  OAI220     u0406(.A0(men_men_n428_), .A1(men_men_n176_), .B0(men_men_n427_), .B1(men_men_n1029_), .Y(men_men_n429_));
  NO2        u0407(.A(i_3_), .B(men_men_n48_), .Y(men_men_n430_));
  NA3        u0408(.A(men_men_n329_), .B(men_men_n328_), .C(men_men_n430_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n310_), .B(men_men_n314_), .Y(men_men_n432_));
  OAI210     u0410(.A0(men_men_n432_), .A1(men_men_n182_), .B0(men_men_n431_), .Y(men_men_n433_));
  NO3        u0411(.A(men_men_n433_), .B(men_men_n429_), .C(men_men_n426_), .Y(men_men_n434_));
  AOI210     u0412(.A0(men_men_n434_), .A1(men_men_n423_), .B0(men_men_n266_), .Y(men_men_n435_));
  NO4        u0413(.A(men_men_n435_), .B(men_men_n416_), .C(men_men_n395_), .D(men_men_n374_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n63_), .B(i_4_), .Y(men_men_n437_));
  NO2        u0415(.A(men_men_n71_), .B(i_13_), .Y(men_men_n438_));
  NA3        u0416(.A(men_men_n438_), .B(men_men_n437_), .C(i_2_), .Y(men_men_n439_));
  NO2        u0417(.A(i_10_), .B(i_9_), .Y(men_men_n440_));
  NAi21      u0418(.An(i_12_), .B(i_8_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n441_), .B(i_3_), .Y(men_men_n442_));
  NA2        u0420(.A(men_men_n442_), .B(men_men_n440_), .Y(men_men_n443_));
  NO2        u0421(.A(men_men_n46_), .B(i_4_), .Y(men_men_n444_));
  NA2        u0422(.A(men_men_n444_), .B(men_men_n101_), .Y(men_men_n445_));
  OAI220     u0423(.A0(men_men_n445_), .A1(men_men_n198_), .B0(men_men_n443_), .B1(men_men_n439_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n303_), .B(i_0_), .Y(men_men_n447_));
  NO3        u0425(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n448_));
  NA2        u0426(.A(men_men_n261_), .B(men_men_n95_), .Y(men_men_n449_));
  NA2        u0427(.A(i_8_), .B(i_9_), .Y(men_men_n450_));
  NA2        u0428(.A(men_men_n278_), .B(men_men_n199_), .Y(men_men_n451_));
  NO2        u0429(.A(men_men_n451_), .B(men_men_n450_), .Y(men_men_n452_));
  NO3        u0430(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n453_));
  NA3        u0431(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n452_), .B(men_men_n446_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n290_), .B(men_men_n104_), .Y(men_men_n456_));
  OR2        u0434(.A(men_men_n456_), .B(men_men_n201_), .Y(men_men_n457_));
  OA220      u0435(.A0(men_men_n344_), .A1(men_men_n158_), .B0(men_men_n457_), .B1(men_men_n227_), .Y(men_men_n458_));
  NA2        u0436(.A(men_men_n94_), .B(i_13_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n420_), .B(men_men_n375_), .Y(men_men_n460_));
  NO2        u0438(.A(i_2_), .B(i_13_), .Y(men_men_n461_));
  NA3        u0439(.A(men_men_n461_), .B(men_men_n157_), .C(men_men_n97_), .Y(men_men_n462_));
  OAI220     u0440(.A0(men_men_n462_), .A1(men_men_n232_), .B0(men_men_n460_), .B1(men_men_n459_), .Y(men_men_n463_));
  NO3        u0441(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n464_));
  NO2        u0442(.A(i_6_), .B(i_7_), .Y(men_men_n465_));
  NOi21      u0443(.An(i_2_), .B(i_7_), .Y(men_men_n466_));
  NAi31      u0444(.An(i_11_), .B(men_men_n466_), .C(men_men_n1023_), .Y(men_men_n467_));
  NO2        u0445(.A(men_men_n407_), .B(i_6_), .Y(men_men_n468_));
  NA3        u0446(.A(men_men_n468_), .B(men_men_n437_), .C(men_men_n73_), .Y(men_men_n469_));
  NO2        u0447(.A(men_men_n469_), .B(men_men_n467_), .Y(men_men_n470_));
  NO2        u0448(.A(i_3_), .B(men_men_n186_), .Y(men_men_n471_));
  NO2        u0449(.A(i_6_), .B(i_10_), .Y(men_men_n472_));
  NA3        u0450(.A(men_men_n239_), .B(men_men_n165_), .C(men_men_n128_), .Y(men_men_n473_));
  NA2        u0451(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n474_));
  NO2        u0452(.A(men_men_n153_), .B(i_3_), .Y(men_men_n475_));
  NAi31      u0453(.An(men_men_n474_), .B(men_men_n475_), .C(men_men_n221_), .Y(men_men_n476_));
  NA3        u0454(.A(men_men_n388_), .B(men_men_n172_), .C(men_men_n144_), .Y(men_men_n477_));
  NA3        u0455(.A(men_men_n477_), .B(men_men_n476_), .C(men_men_n473_), .Y(men_men_n478_));
  NO3        u0456(.A(men_men_n478_), .B(men_men_n470_), .C(men_men_n463_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n448_), .B(men_men_n376_), .Y(men_men_n480_));
  NA2        u0458(.A(men_men_n453_), .B(men_men_n383_), .Y(men_men_n481_));
  NO2        u0459(.A(men_men_n481_), .B(men_men_n219_), .Y(men_men_n482_));
  NAi21      u0460(.An(men_men_n210_), .B(men_men_n393_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n329_), .B(men_men_n212_), .Y(men_men_n484_));
  NO2        u0462(.A(i_0_), .B(men_men_n83_), .Y(men_men_n485_));
  NA3        u0463(.A(men_men_n485_), .B(i_3_), .C(men_men_n137_), .Y(men_men_n486_));
  OAI220     u0464(.A0(men_men_n38_), .A1(men_men_n486_), .B0(men_men_n484_), .B1(men_men_n483_), .Y(men_men_n487_));
  NA2        u0465(.A(men_men_n27_), .B(i_10_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n307_), .B(men_men_n233_), .Y(men_men_n489_));
  OAI220     u0467(.A0(men_men_n489_), .A1(men_men_n427_), .B0(men_men_n488_), .B1(men_men_n459_), .Y(men_men_n490_));
  NO3        u0468(.A(men_men_n490_), .B(men_men_n487_), .C(men_men_n482_), .Y(men_men_n491_));
  NA4        u0469(.A(men_men_n491_), .B(men_men_n479_), .C(men_men_n458_), .D(men_men_n455_), .Y(men_men_n492_));
  NA3        u0470(.A(men_men_n300_), .B(men_men_n169_), .C(men_men_n167_), .Y(men_men_n493_));
  OAI210     u0471(.A0(men_men_n296_), .A1(men_men_n174_), .B0(men_men_n493_), .Y(men_men_n494_));
  AN2        u0472(.A(men_men_n281_), .B(men_men_n229_), .Y(men_men_n495_));
  NA2        u0473(.A(men_men_n495_), .B(men_men_n494_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n118_), .B(men_men_n108_), .Y(men_men_n497_));
  AN2        u0475(.A(men_men_n497_), .B(men_men_n448_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n307_), .B(men_men_n160_), .Y(men_men_n499_));
  OAI210     u0477(.A0(men_men_n499_), .A1(men_men_n227_), .B0(men_men_n301_), .Y(men_men_n500_));
  AOI210     u0478(.A0(men_men_n498_), .A1(men_men_n303_), .B0(men_men_n500_), .Y(men_men_n501_));
  NA4        u0479(.A(men_men_n438_), .B(men_men_n437_), .C(men_men_n196_), .D(i_2_), .Y(men_men_n502_));
  INV        u0480(.A(men_men_n502_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n376_), .B(men_men_n220_), .Y(men_men_n504_));
  NA2        u0482(.A(men_men_n348_), .B(men_men_n71_), .Y(men_men_n505_));
  NA2        u0483(.A(men_men_n365_), .B(men_men_n357_), .Y(men_men_n506_));
  AO210      u0484(.A0(men_men_n505_), .A1(men_men_n504_), .B0(men_men_n506_), .Y(men_men_n507_));
  NO2        u0485(.A(men_men_n36_), .B(i_8_), .Y(men_men_n508_));
  INV        u0486(.A(men_men_n408_), .Y(men_men_n509_));
  NA2        u0487(.A(men_men_n509_), .B(men_men_n507_), .Y(men_men_n510_));
  AOI210     u0488(.A0(men_men_n503_), .A1(men_men_n197_), .B0(men_men_n510_), .Y(men_men_n511_));
  NA2        u0489(.A(men_men_n252_), .B(men_men_n64_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n512_), .B(men_men_n129_), .Y(men_men_n513_));
  AOI210     u0491(.A0(men_men_n187_), .A1(i_9_), .B0(men_men_n260_), .Y(men_men_n514_));
  NO2        u0492(.A(men_men_n514_), .B(men_men_n192_), .Y(men_men_n515_));
  AOI220     u0493(.A0(i_3_), .A1(men_men_n515_), .B0(men_men_n513_), .B1(men_men_n409_), .Y(men_men_n516_));
  NA4        u0494(.A(men_men_n516_), .B(men_men_n511_), .C(men_men_n501_), .D(men_men_n496_), .Y(men_men_n517_));
  NO2        u0495(.A(i_12_), .B(men_men_n186_), .Y(men_men_n518_));
  NA3        u0496(.A(men_men_n472_), .B(men_men_n167_), .C(men_men_n27_), .Y(men_men_n519_));
  NO3        u0497(.A(men_men_n519_), .B(i_13_), .C(men_men_n456_), .Y(men_men_n520_));
  NOi31      u0498(.An(men_men_n310_), .B(men_men_n407_), .C(men_men_n38_), .Y(men_men_n521_));
  OAI210     u0499(.A0(men_men_n521_), .A1(men_men_n520_), .B0(men_men_n377_), .Y(men_men_n522_));
  NO2        u0500(.A(i_8_), .B(i_7_), .Y(men_men_n523_));
  OAI210     u0501(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n524_), .B(men_men_n218_), .Y(men_men_n525_));
  AOI220     u0503(.A0(men_men_n317_), .A1(men_men_n39_), .B0(men_men_n230_), .B1(men_men_n200_), .Y(men_men_n526_));
  OAI220     u0504(.A0(men_men_n526_), .A1(men_men_n176_), .B0(men_men_n525_), .B1(men_men_n236_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n44_), .B(i_10_), .Y(men_men_n528_));
  NO2        u0506(.A(men_men_n528_), .B(i_6_), .Y(men_men_n529_));
  NA3        u0507(.A(men_men_n529_), .B(men_men_n527_), .C(men_men_n523_), .Y(men_men_n530_));
  AOI220     u0508(.A0(men_men_n420_), .A1(men_men_n317_), .B0(men_men_n241_), .B1(men_men_n238_), .Y(men_men_n531_));
  OAI220     u0509(.A0(men_men_n531_), .A1(i_12_), .B0(men_men_n459_), .B1(men_men_n129_), .Y(men_men_n532_));
  NA2        u0510(.A(men_men_n532_), .B(men_men_n260_), .Y(men_men_n533_));
  NOi31      u0511(.An(men_men_n285_), .B(men_men_n296_), .C(men_men_n174_), .Y(men_men_n534_));
  NA3        u0512(.A(men_men_n300_), .B(men_men_n167_), .C(men_men_n94_), .Y(men_men_n535_));
  NO2        u0513(.A(men_men_n153_), .B(i_5_), .Y(men_men_n536_));
  NA3        u0514(.A(men_men_n536_), .B(men_men_n396_), .C(men_men_n312_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n537_), .B(men_men_n535_), .Y(men_men_n538_));
  OAI210     u0516(.A0(men_men_n538_), .A1(men_men_n534_), .B0(men_men_n453_), .Y(men_men_n539_));
  NA4        u0517(.A(men_men_n539_), .B(men_men_n533_), .C(men_men_n530_), .D(men_men_n522_), .Y(men_men_n540_));
  NA3        u0518(.A(men_men_n212_), .B(men_men_n69_), .C(men_men_n44_), .Y(men_men_n541_));
  NA2        u0519(.A(men_men_n278_), .B(men_men_n81_), .Y(men_men_n542_));
  AOI210     u0520(.A0(men_men_n541_), .A1(men_men_n339_), .B0(men_men_n542_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n291_), .B(men_men_n281_), .Y(men_men_n544_));
  NO2        u0522(.A(men_men_n544_), .B(men_men_n166_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n440_), .B(men_men_n216_), .Y(men_men_n547_));
  NO2        u0525(.A(men_men_n546_), .B(men_men_n547_), .Y(men_men_n548_));
  AOI210     u0526(.A0(men_men_n358_), .A1(men_men_n46_), .B0(men_men_n362_), .Y(men_men_n549_));
  NA2        u0527(.A(i_0_), .B(men_men_n48_), .Y(men_men_n550_));
  NA3        u0528(.A(men_men_n518_), .B(men_men_n269_), .C(men_men_n550_), .Y(men_men_n551_));
  NO2        u0529(.A(men_men_n549_), .B(men_men_n551_), .Y(men_men_n552_));
  NO4        u0530(.A(men_men_n552_), .B(men_men_n548_), .C(men_men_n545_), .D(men_men_n543_), .Y(men_men_n553_));
  NO4        u0531(.A(men_men_n246_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n554_));
  NO3        u0532(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n555_));
  NO2        u0533(.A(men_men_n228_), .B(men_men_n36_), .Y(men_men_n556_));
  AN2        u0534(.A(men_men_n556_), .B(men_men_n555_), .Y(men_men_n557_));
  OA210      u0535(.A0(men_men_n557_), .A1(men_men_n554_), .B0(men_men_n348_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n407_), .B(i_1_), .Y(men_men_n559_));
  NOi31      u0537(.An(men_men_n559_), .B(men_men_n449_), .C(men_men_n71_), .Y(men_men_n560_));
  AN3        u0538(.A(men_men_n560_), .B(men_men_n404_), .C(i_2_), .Y(men_men_n561_));
  NO2        u0539(.A(men_men_n418_), .B(men_men_n170_), .Y(men_men_n562_));
  NO3        u0540(.A(men_men_n562_), .B(men_men_n561_), .C(men_men_n558_), .Y(men_men_n563_));
  NOi21      u0541(.An(i_10_), .B(i_6_), .Y(men_men_n564_));
  NO2        u0542(.A(men_men_n83_), .B(men_men_n25_), .Y(men_men_n565_));
  NA2        u0543(.A(men_men_n278_), .B(men_men_n565_), .Y(men_men_n566_));
  NO2        u0544(.A(men_men_n566_), .B(men_men_n447_), .Y(men_men_n567_));
  NO2        u0545(.A(men_men_n111_), .B(men_men_n23_), .Y(men_men_n568_));
  NA2        u0546(.A(men_men_n310_), .B(men_men_n160_), .Y(men_men_n569_));
  AOI220     u0547(.A0(men_men_n569_), .A1(men_men_n428_), .B0(men_men_n166_), .B1(men_men_n175_), .Y(men_men_n570_));
  NO2        u0548(.A(men_men_n191_), .B(men_men_n37_), .Y(men_men_n571_));
  NOi31      u0549(.An(men_men_n141_), .B(men_men_n571_), .C(men_men_n325_), .Y(men_men_n572_));
  NO3        u0550(.A(men_men_n572_), .B(men_men_n570_), .C(men_men_n567_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n505_), .B(men_men_n371_), .Y(men_men_n574_));
  INV        u0552(.A(men_men_n312_), .Y(men_men_n575_));
  NO2        u0553(.A(i_12_), .B(men_men_n83_), .Y(men_men_n576_));
  NA3        u0554(.A(men_men_n576_), .B(men_men_n269_), .C(men_men_n550_), .Y(men_men_n577_));
  NA3        u0555(.A(men_men_n379_), .B(men_men_n278_), .C(men_men_n212_), .Y(men_men_n578_));
  AOI210     u0556(.A0(men_men_n578_), .A1(men_men_n577_), .B0(men_men_n575_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n167_), .B(i_0_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n580_), .B(men_men_n296_), .Y(men_men_n581_));
  OR2        u0559(.A(i_2_), .B(i_5_), .Y(men_men_n582_));
  OR2        u0560(.A(men_men_n582_), .B(men_men_n399_), .Y(men_men_n583_));
  NA2        u0561(.A(men_men_n367_), .B(men_men_n238_), .Y(men_men_n584_));
  AOI210     u0562(.A0(men_men_n584_), .A1(men_men_n583_), .B0(men_men_n483_), .Y(men_men_n585_));
  NO4        u0563(.A(men_men_n585_), .B(men_men_n581_), .C(men_men_n579_), .D(men_men_n574_), .Y(men_men_n586_));
  NA4        u0564(.A(men_men_n586_), .B(men_men_n573_), .C(men_men_n563_), .D(men_men_n553_), .Y(men_men_n587_));
  NO4        u0565(.A(men_men_n587_), .B(men_men_n540_), .C(men_men_n517_), .D(men_men_n492_), .Y(men_men_n588_));
  NA4        u0566(.A(men_men_n588_), .B(men_men_n436_), .C(men_men_n347_), .D(men_men_n306_), .Y(men7));
  NO2        u0567(.A(men_men_n104_), .B(men_men_n87_), .Y(men_men_n590_));
  NA2        u0568(.A(men_men_n377_), .B(men_men_n590_), .Y(men_men_n591_));
  NA2        u0569(.A(men_men_n472_), .B(men_men_n81_), .Y(men_men_n592_));
  NA2        u0570(.A(i_11_), .B(men_men_n186_), .Y(men_men_n593_));
  INV        u0571(.A(men_men_n591_), .Y(men_men_n594_));
  NA3        u0572(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n595_));
  NO2        u0573(.A(men_men_n232_), .B(i_4_), .Y(men_men_n596_));
  NA2        u0574(.A(men_men_n596_), .B(i_8_), .Y(men_men_n597_));
  AOI210     u0575(.A0(men_men_n597_), .A1(men_men_n102_), .B0(men_men_n595_), .Y(men_men_n598_));
  NA2        u0576(.A(i_2_), .B(men_men_n83_), .Y(men_men_n599_));
  OAI210     u0577(.A0(men_men_n85_), .A1(men_men_n196_), .B0(men_men_n197_), .Y(men_men_n600_));
  NO2        u0578(.A(i_7_), .B(men_men_n37_), .Y(men_men_n601_));
  NA2        u0579(.A(i_4_), .B(i_8_), .Y(men_men_n602_));
  AOI210     u0580(.A0(men_men_n602_), .A1(men_men_n300_), .B0(men_men_n601_), .Y(men_men_n603_));
  OAI220     u0581(.A0(men_men_n603_), .A1(men_men_n599_), .B0(men_men_n600_), .B1(i_13_), .Y(men_men_n604_));
  NO3        u0582(.A(men_men_n604_), .B(men_men_n598_), .C(men_men_n594_), .Y(men_men_n605_));
  AOI210     u0583(.A0(men_men_n124_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n606_));
  AOI210     u0584(.A0(men_men_n606_), .A1(men_men_n232_), .B0(men_men_n157_), .Y(men_men_n607_));
  OR2        u0585(.A(i_6_), .B(i_10_), .Y(men_men_n608_));
  NO2        u0586(.A(men_men_n608_), .B(men_men_n23_), .Y(men_men_n609_));
  OR3        u0587(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n610_));
  NO3        u0588(.A(men_men_n610_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n611_));
  INV        u0589(.A(men_men_n193_), .Y(men_men_n612_));
  OA220      u0590(.A0(men_men_n610_), .A1(men_men_n575_), .B0(men_men_n607_), .B1(men_men_n262_), .Y(men_men_n613_));
  AOI210     u0591(.A0(men_men_n613_), .A1(men_men_n605_), .B0(men_men_n63_), .Y(men_men_n614_));
  NOi21      u0592(.An(i_11_), .B(i_7_), .Y(men_men_n615_));
  AO210      u0593(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n616_));
  NO2        u0594(.A(men_men_n616_), .B(men_men_n615_), .Y(men_men_n617_));
  NA2        u0595(.A(men_men_n617_), .B(men_men_n200_), .Y(men_men_n618_));
  NA3        u0596(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n619_));
  AOI210     u0597(.A0(men_men_n619_), .A1(men_men_n618_), .B0(men_men_n63_), .Y(men_men_n620_));
  AO210      u0598(.A0(men_men_n84_), .A1(men_men_n371_), .B0(men_men_n40_), .Y(men_men_n621_));
  NO3        u0599(.A(men_men_n254_), .B(men_men_n202_), .C(men_men_n593_), .Y(men_men_n622_));
  OAI210     u0600(.A0(men_men_n622_), .A1(men_men_n221_), .B0(men_men_n63_), .Y(men_men_n623_));
  NA2        u0601(.A(men_men_n400_), .B(men_men_n31_), .Y(men_men_n624_));
  OR2        u0602(.A(men_men_n202_), .B(men_men_n104_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n625_), .B(men_men_n624_), .Y(men_men_n626_));
  NO2        u0604(.A(men_men_n63_), .B(i_9_), .Y(men_men_n627_));
  NO2        u0605(.A(men_men_n627_), .B(i_4_), .Y(men_men_n628_));
  NA2        u0606(.A(men_men_n628_), .B(men_men_n626_), .Y(men_men_n629_));
  NO2        u0607(.A(i_1_), .B(i_12_), .Y(men_men_n630_));
  NA3        u0608(.A(men_men_n630_), .B(men_men_n106_), .C(men_men_n24_), .Y(men_men_n631_));
  NA4        u0609(.A(men_men_n631_), .B(men_men_n629_), .C(men_men_n623_), .D(men_men_n621_), .Y(men_men_n632_));
  OAI210     u0610(.A0(men_men_n632_), .A1(men_men_n620_), .B0(i_6_), .Y(men_men_n633_));
  INV        u0611(.A(men_men_n619_), .Y(men_men_n634_));
  NA2        u0612(.A(men_men_n634_), .B(men_men_n576_), .Y(men_men_n635_));
  NO2        u0613(.A(men_men_n232_), .B(men_men_n83_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n636_), .B(i_11_), .Y(men_men_n637_));
  INV        u0615(.A(men_men_n635_), .Y(men_men_n638_));
  NO4        u0616(.A(men_men_n209_), .B(men_men_n124_), .C(i_13_), .D(men_men_n83_), .Y(men_men_n639_));
  NA2        u0617(.A(men_men_n639_), .B(men_men_n627_), .Y(men_men_n640_));
  NO3        u0618(.A(men_men_n608_), .B(men_men_n228_), .C(men_men_n23_), .Y(men_men_n641_));
  AOI210     u0619(.A0(i_1_), .A1(men_men_n255_), .B0(men_men_n641_), .Y(men_men_n642_));
  OAI210     u0620(.A0(men_men_n642_), .A1(men_men_n44_), .B0(men_men_n640_), .Y(men_men_n643_));
  NA3        u0621(.A(men_men_n523_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n644_));
  NA3        u0622(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n645_));
  NO2        u0623(.A(men_men_n46_), .B(i_1_), .Y(men_men_n646_));
  NA3        u0624(.A(men_men_n646_), .B(men_men_n261_), .C(men_men_n44_), .Y(men_men_n647_));
  NO2        u0625(.A(men_men_n647_), .B(men_men_n645_), .Y(men_men_n648_));
  NA3        u0626(.A(men_men_n627_), .B(men_men_n312_), .C(i_6_), .Y(men_men_n649_));
  NAi21      u0627(.An(men_men_n644_), .B(men_men_n89_), .Y(men_men_n650_));
  NO2        u0628(.A(i_11_), .B(men_men_n37_), .Y(men_men_n651_));
  NA2        u0629(.A(men_men_n651_), .B(men_men_n24_), .Y(men_men_n652_));
  OAI210     u0630(.A0(men_men_n652_), .A1(i_6_), .B0(men_men_n650_), .Y(men_men_n653_));
  OR2        u0631(.A(men_men_n653_), .B(men_men_n648_), .Y(men_men_n654_));
  NO3        u0632(.A(men_men_n654_), .B(men_men_n643_), .C(men_men_n638_), .Y(men_men_n655_));
  NO2        u0633(.A(men_men_n406_), .B(men_men_n83_), .Y(men_men_n656_));
  NA2        u0634(.A(i_3_), .B(men_men_n186_), .Y(men_men_n657_));
  NO2        u0635(.A(men_men_n228_), .B(men_men_n44_), .Y(men_men_n658_));
  NO3        u0636(.A(men_men_n658_), .B(men_men_n303_), .C(i_12_), .Y(men_men_n659_));
  NO2        u0637(.A(men_men_n113_), .B(men_men_n37_), .Y(men_men_n660_));
  NO2        u0638(.A(men_men_n660_), .B(i_6_), .Y(men_men_n661_));
  NO2        u0639(.A(men_men_n83_), .B(i_9_), .Y(men_men_n662_));
  NO2        u0640(.A(men_men_n662_), .B(men_men_n63_), .Y(men_men_n663_));
  NO2        u0641(.A(men_men_n663_), .B(men_men_n630_), .Y(men_men_n664_));
  NO4        u0642(.A(men_men_n664_), .B(men_men_n661_), .C(men_men_n659_), .D(i_4_), .Y(men_men_n665_));
  NA2        u0643(.A(i_1_), .B(i_3_), .Y(men_men_n666_));
  NA2        u0644(.A(men_men_n658_), .B(men_men_n564_), .Y(men_men_n667_));
  NO2        u0645(.A(men_men_n667_), .B(men_men_n666_), .Y(men_men_n668_));
  NO2        u0646(.A(men_men_n668_), .B(men_men_n665_), .Y(men_men_n669_));
  NA3        u0647(.A(men_men_n669_), .B(men_men_n655_), .C(men_men_n633_), .Y(men_men_n670_));
  NO3        u0648(.A(i_11_), .B(i_3_), .C(i_7_), .Y(men_men_n671_));
  OA210      u0649(.A0(men_men_n671_), .A1(men_men_n239_), .B0(men_men_n83_), .Y(men_men_n672_));
  NA2        u0650(.A(men_men_n365_), .B(men_men_n364_), .Y(men_men_n673_));
  NA3        u0651(.A(men_men_n472_), .B(men_men_n508_), .C(men_men_n46_), .Y(men_men_n674_));
  NO3        u0652(.A(men_men_n466_), .B(men_men_n602_), .C(men_men_n83_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n675_), .B(men_men_n25_), .Y(men_men_n676_));
  NA3        u0654(.A(men_men_n676_), .B(men_men_n674_), .C(men_men_n673_), .Y(men_men_n677_));
  OAI210     u0655(.A0(men_men_n677_), .A1(men_men_n672_), .B0(i_1_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n363_), .B(i_2_), .Y(men_men_n679_));
  AOI210     u0657(.A0(men_men_n649_), .A1(men_men_n678_), .B0(i_13_), .Y(men_men_n680_));
  OR2        u0658(.A(i_11_), .B(i_7_), .Y(men_men_n681_));
  NA2        u0659(.A(men_men_n103_), .B(men_men_n133_), .Y(men_men_n682_));
  AOI220     u0660(.A0(men_men_n461_), .A1(men_men_n157_), .B0(men_men_n444_), .B1(men_men_n133_), .Y(men_men_n683_));
  OAI210     u0661(.A0(men_men_n683_), .A1(men_men_n44_), .B0(men_men_n682_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n466_), .B(men_men_n24_), .Y(men_men_n685_));
  AOI210     u0663(.A0(men_men_n685_), .A1(men_men_n656_), .B0(men_men_n239_), .Y(men_men_n686_));
  OAI220     u0664(.A0(men_men_n686_), .A1(men_men_n40_), .B0(men_men_n54_), .B1(men_men_n90_), .Y(men_men_n687_));
  AOI210     u0665(.A0(men_men_n684_), .A1(men_men_n327_), .B0(men_men_n687_), .Y(men_men_n688_));
  AOI220     u0666(.A0(i_12_), .A1(men_men_n70_), .B0(men_men_n379_), .B1(men_men_n646_), .Y(men_men_n689_));
  NO2        u0667(.A(men_men_n689_), .B(men_men_n236_), .Y(men_men_n690_));
  AOI210     u0668(.A0(men_men_n441_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n691_));
  NOi31      u0669(.An(men_men_n691_), .B(men_men_n592_), .C(men_men_n44_), .Y(men_men_n692_));
  NA2        u0670(.A(men_men_n123_), .B(i_13_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n645_), .B(men_men_n111_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n693_), .B(men_men_n1028_), .Y(men_men_n695_));
  NO3        u0673(.A(men_men_n69_), .B(men_men_n32_), .C(men_men_n99_), .Y(men_men_n696_));
  NA2        u0674(.A(i_3_), .B(i_7_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n232_), .B(men_men_n83_), .Y(men_men_n698_));
  AOI210     u0676(.A0(men_men_n698_), .A1(men_men_n697_), .B0(men_men_n696_), .Y(men_men_n699_));
  AOI210     u0677(.A0(men_men_n379_), .A1(men_men_n646_), .B0(men_men_n89_), .Y(men_men_n700_));
  OAI220     u0678(.A0(men_men_n700_), .A1(men_men_n597_), .B0(men_men_n699_), .B1(men_men_n612_), .Y(men_men_n701_));
  NO4        u0679(.A(men_men_n701_), .B(men_men_n695_), .C(men_men_n692_), .D(men_men_n690_), .Y(men_men_n702_));
  NA3        u0680(.A(men_men_n400_), .B(men_men_n601_), .C(men_men_n95_), .Y(men_men_n703_));
  NA2        u0681(.A(men_men_n637_), .B(i_13_), .Y(men_men_n704_));
  NAi21      u0682(.An(i_11_), .B(i_12_), .Y(men_men_n705_));
  NOi41      u0683(.An(men_men_n107_), .B(men_men_n705_), .C(i_13_), .D(men_men_n83_), .Y(men_men_n706_));
  NO2        u0684(.A(men_men_n576_), .B(men_men_n602_), .Y(men_men_n707_));
  AOI210     u0685(.A0(men_men_n707_), .A1(men_men_n307_), .B0(men_men_n706_), .Y(men_men_n708_));
  NA3        u0686(.A(men_men_n708_), .B(men_men_n704_), .C(men_men_n703_), .Y(men_men_n709_));
  OAI210     u0687(.A0(men_men_n709_), .A1(men_men_n694_), .B0(men_men_n63_), .Y(men_men_n710_));
  NA2        u0688(.A(i_8_), .B(men_men_n25_), .Y(men_men_n711_));
  NO3        u0689(.A(men_men_n711_), .B(men_men_n377_), .C(men_men_n596_), .Y(men_men_n712_));
  OAI210     u0690(.A0(men_men_n712_), .A1(men_men_n364_), .B0(men_men_n362_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n124_), .B(i_2_), .Y(men_men_n714_));
  INV        u0692(.A(men_men_n714_), .Y(men_men_n715_));
  NA2        u0693(.A(men_men_n715_), .B(men_men_n713_), .Y(men_men_n716_));
  NA3        u0694(.A(men_men_n716_), .B(men_men_n45_), .C(men_men_n220_), .Y(men_men_n717_));
  NA4        u0695(.A(men_men_n717_), .B(men_men_n710_), .C(men_men_n702_), .D(men_men_n688_), .Y(men_men_n718_));
  OR4        u0696(.A(men_men_n718_), .B(men_men_n680_), .C(men_men_n670_), .D(men_men_n614_), .Y(men5));
  NO2        u0697(.A(men_men_n597_), .B(i_11_), .Y(men_men_n720_));
  NA2        u0698(.A(men_men_n85_), .B(men_men_n720_), .Y(men_men_n721_));
  INV        u0699(.A(men_men_n721_), .Y(men_men_n722_));
  NO3        u0700(.A(i_11_), .B(men_men_n232_), .C(i_13_), .Y(men_men_n723_));
  NO2        u0701(.A(men_men_n120_), .B(men_men_n23_), .Y(men_men_n724_));
  NA2        u0702(.A(i_12_), .B(i_8_), .Y(men_men_n725_));
  OAI210     u0703(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n725_), .Y(men_men_n726_));
  INV        u0704(.A(men_men_n440_), .Y(men_men_n727_));
  AOI220     u0705(.A0(men_men_n312_), .A1(men_men_n568_), .B0(men_men_n726_), .B1(men_men_n724_), .Y(men_men_n728_));
  INV        u0706(.A(men_men_n728_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n729_), .B(men_men_n722_), .Y(men_men_n730_));
  INV        u0708(.A(men_men_n165_), .Y(men_men_n731_));
  INV        u0709(.A(men_men_n239_), .Y(men_men_n732_));
  OAI210     u0710(.A0(men_men_n679_), .A1(men_men_n442_), .B0(men_men_n107_), .Y(men_men_n733_));
  AOI210     u0711(.A0(men_men_n733_), .A1(men_men_n732_), .B0(men_men_n731_), .Y(men_men_n734_));
  NO2        u0712(.A(men_men_n450_), .B(men_men_n26_), .Y(men_men_n735_));
  NO2        u0713(.A(men_men_n735_), .B(men_men_n411_), .Y(men_men_n736_));
  NA2        u0714(.A(men_men_n736_), .B(i_2_), .Y(men_men_n737_));
  INV        u0715(.A(men_men_n737_), .Y(men_men_n738_));
  AOI210     u0716(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n407_), .Y(men_men_n739_));
  AOI210     u0717(.A0(men_men_n739_), .A1(men_men_n738_), .B0(men_men_n734_), .Y(men_men_n740_));
  NO2        u0718(.A(men_men_n183_), .B(men_men_n121_), .Y(men_men_n741_));
  OAI210     u0719(.A0(men_men_n741_), .A1(men_men_n724_), .B0(i_2_), .Y(men_men_n742_));
  NO2        u0720(.A(men_men_n742_), .B(men_men_n186_), .Y(men_men_n743_));
  OA210      u0721(.A0(men_men_n617_), .A1(men_men_n122_), .B0(i_13_), .Y(men_men_n744_));
  NA2        u0722(.A(men_men_n193_), .B(men_men_n196_), .Y(men_men_n745_));
  NO2        u0723(.A(men_men_n745_), .B(men_men_n367_), .Y(men_men_n746_));
  AOI210     u0724(.A0(men_men_n202_), .A1(men_men_n143_), .B0(men_men_n508_), .Y(men_men_n747_));
  NA2        u0725(.A(men_men_n747_), .B(men_men_n411_), .Y(men_men_n748_));
  NO2        u0726(.A(i_2_), .B(men_men_n44_), .Y(men_men_n749_));
  NA3        u0727(.A(men_men_n300_), .B(men_men_n120_), .C(men_men_n42_), .Y(men_men_n750_));
  OAI210     u0728(.A0(men_men_n750_), .A1(men_men_n749_), .B0(men_men_n748_), .Y(men_men_n751_));
  NO4        u0729(.A(men_men_n751_), .B(men_men_n746_), .C(men_men_n744_), .D(men_men_n743_), .Y(men_men_n752_));
  NA2        u0730(.A(men_men_n568_), .B(men_men_n28_), .Y(men_men_n753_));
  NA2        u0731(.A(men_men_n723_), .B(men_men_n270_), .Y(men_men_n754_));
  NA2        u0732(.A(men_men_n754_), .B(men_men_n753_), .Y(men_men_n755_));
  NO2        u0733(.A(men_men_n62_), .B(i_12_), .Y(men_men_n756_));
  NO2        u0734(.A(men_men_n756_), .B(men_men_n122_), .Y(men_men_n757_));
  NO2        u0735(.A(men_men_n757_), .B(men_men_n593_), .Y(men_men_n758_));
  AOI220     u0736(.A0(men_men_n758_), .A1(men_men_n36_), .B0(men_men_n755_), .B1(men_men_n46_), .Y(men_men_n759_));
  NA4        u0737(.A(men_men_n759_), .B(men_men_n752_), .C(men_men_n740_), .D(men_men_n730_), .Y(men6));
  NA2        u0738(.A(men_men_n25_), .B(men_men_n714_), .Y(men_men_n761_));
  NA4        u0739(.A(men_men_n383_), .B(men_men_n471_), .C(men_men_n69_), .D(men_men_n99_), .Y(men_men_n762_));
  INV        u0740(.A(men_men_n762_), .Y(men_men_n763_));
  NO2        u0741(.A(men_men_n215_), .B(men_men_n474_), .Y(men_men_n764_));
  NO2        u0742(.A(i_11_), .B(i_9_), .Y(men_men_n765_));
  NO2        u0743(.A(men_men_n763_), .B(men_men_n322_), .Y(men_men_n766_));
  AO210      u0744(.A0(men_men_n766_), .A1(men_men_n761_), .B0(i_12_), .Y(men_men_n767_));
  NA2        u0745(.A(men_men_n368_), .B(men_men_n329_), .Y(men_men_n768_));
  NA2        u0746(.A(men_men_n576_), .B(men_men_n63_), .Y(men_men_n769_));
  NA2        u0747(.A(men_men_n671_), .B(men_men_n69_), .Y(men_men_n770_));
  NA4        u0748(.A(men_men_n84_), .B(men_men_n770_), .C(men_men_n769_), .D(men_men_n768_), .Y(men_men_n771_));
  AOI220     u0749(.A0(men_men_n189_), .A1(men_men_n765_), .B0(men_men_n771_), .B1(men_men_n71_), .Y(men_men_n772_));
  NA2        u0750(.A(men_men_n1025_), .B(men_men_n756_), .Y(men_men_n773_));
  AOI210     u0751(.A0(men_men_n773_), .A1(men_men_n506_), .B0(men_men_n178_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n32_), .B(i_11_), .Y(men_men_n775_));
  NA3        u0753(.A(men_men_n775_), .B(men_men_n465_), .C(men_men_n383_), .Y(men_men_n776_));
  NAi32      u0754(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n777_));
  AOI210     u0755(.A0(i_6_), .A1(men_men_n84_), .B0(men_men_n777_), .Y(men_men_n778_));
  OAI210     u0756(.A0(men_men_n671_), .A1(men_men_n556_), .B0(men_men_n555_), .Y(men_men_n779_));
  NAi31      u0757(.An(men_men_n778_), .B(men_men_n779_), .C(men_men_n776_), .Y(men_men_n780_));
  OR2        u0758(.A(men_men_n780_), .B(men_men_n774_), .Y(men_men_n781_));
  NA3        u0759(.A(men_men_n343_), .B(men_men_n251_), .C(i_7_), .Y(men_men_n782_));
  NA3        u0760(.A(men_men_n442_), .B(men_men_n142_), .C(men_men_n67_), .Y(men_men_n783_));
  AO210      u0761(.A0(men_men_n481_), .A1(men_men_n727_), .B0(men_men_n36_), .Y(men_men_n784_));
  NA3        u0762(.A(men_men_n784_), .B(men_men_n783_), .C(men_men_n782_), .Y(men_men_n785_));
  AOI210     u0763(.A0(men_men_n1027_), .A1(men_men_n555_), .B0(men_men_n764_), .Y(men_men_n786_));
  NA3        u0764(.A(men_men_n367_), .B(men_men_n233_), .C(men_men_n142_), .Y(men_men_n787_));
  NA2        u0765(.A(men_men_n391_), .B(men_men_n68_), .Y(men_men_n788_));
  NA3        u0766(.A(men_men_n788_), .B(men_men_n787_), .C(men_men_n786_), .Y(men_men_n789_));
  NA3        u0767(.A(men_men_n46_), .B(men_men_n472_), .C(men_men_n212_), .Y(men_men_n790_));
  AOI210     u0768(.A0(men_men_n442_), .A1(men_men_n440_), .B0(men_men_n554_), .Y(men_men_n791_));
  NA2        u0769(.A(men_men_n108_), .B(men_men_n398_), .Y(men_men_n792_));
  NA3        u0770(.A(men_men_n792_), .B(men_men_n791_), .C(men_men_n790_), .Y(men_men_n793_));
  NO4        u0771(.A(men_men_n793_), .B(men_men_n789_), .C(men_men_n785_), .D(men_men_n781_), .Y(men_men_n794_));
  NA4        u0772(.A(men_men_n794_), .B(men_men_n772_), .C(men_men_n767_), .D(men_men_n373_), .Y(men3));
  NA2        u0773(.A(i_12_), .B(i_10_), .Y(men_men_n796_));
  NA2        u0774(.A(i_6_), .B(i_7_), .Y(men_men_n797_));
  NO2        u0775(.A(men_men_n797_), .B(i_0_), .Y(men_men_n798_));
  NO2        u0776(.A(i_11_), .B(men_men_n232_), .Y(men_men_n799_));
  OAI210     u0777(.A0(men_men_n798_), .A1(men_men_n285_), .B0(men_men_n799_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n800_), .B(men_men_n186_), .Y(men_men_n801_));
  NO3        u0779(.A(men_men_n447_), .B(men_men_n87_), .C(men_men_n44_), .Y(men_men_n802_));
  OA210      u0780(.A0(men_men_n802_), .A1(men_men_n801_), .B0(men_men_n167_), .Y(men_men_n803_));
  NA3        u0781(.A(men_men_n787_), .B(men_men_n600_), .C(men_men_n366_), .Y(men_men_n804_));
  NA2        u0782(.A(men_men_n804_), .B(men_men_n39_), .Y(men_men_n805_));
  NOi21      u0783(.An(men_men_n94_), .B(men_men_n736_), .Y(men_men_n806_));
  NO3        u0784(.A(men_men_n625_), .B(men_men_n450_), .C(men_men_n127_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n400_), .B(men_men_n45_), .Y(men_men_n808_));
  AN2        u0786(.A(men_men_n449_), .B(men_men_n55_), .Y(men_men_n809_));
  NO3        u0787(.A(men_men_n809_), .B(men_men_n807_), .C(men_men_n806_), .Y(men_men_n810_));
  AOI210     u0788(.A0(men_men_n810_), .A1(men_men_n805_), .B0(men_men_n48_), .Y(men_men_n811_));
  NA2        u0789(.A(men_men_n178_), .B(men_men_n564_), .Y(men_men_n812_));
  NA2        u0790(.A(men_men_n691_), .B(men_men_n662_), .Y(men_men_n813_));
  NA2        u0791(.A(i_0_), .B(men_men_n430_), .Y(men_men_n814_));
  OAI220     u0792(.A0(men_men_n814_), .A1(men_men_n813_), .B0(men_men_n812_), .B1(men_men_n63_), .Y(men_men_n815_));
  NOi21      u0793(.An(i_5_), .B(i_9_), .Y(men_men_n816_));
  NA2        u0794(.A(men_men_n816_), .B(men_men_n438_), .Y(men_men_n817_));
  NO3        u0795(.A(men_men_n403_), .B(men_men_n261_), .C(men_men_n71_), .Y(men_men_n818_));
  NO2        u0796(.A(men_men_n168_), .B(men_men_n143_), .Y(men_men_n819_));
  AOI210     u0797(.A0(men_men_n819_), .A1(men_men_n238_), .B0(men_men_n818_), .Y(men_men_n820_));
  OAI220     u0798(.A0(men_men_n820_), .A1(men_men_n174_), .B0(men_men_n602_), .B1(men_men_n817_), .Y(men_men_n821_));
  NO4        u0799(.A(men_men_n821_), .B(men_men_n815_), .C(men_men_n811_), .D(men_men_n803_), .Y(men_men_n822_));
  NA2        u0800(.A(men_men_n178_), .B(men_men_n24_), .Y(men_men_n823_));
  NO2        u0801(.A(men_men_n660_), .B(men_men_n590_), .Y(men_men_n824_));
  NO2        u0802(.A(men_men_n824_), .B(men_men_n823_), .Y(men_men_n825_));
  NA2        u0803(.A(men_men_n307_), .B(men_men_n125_), .Y(men_men_n826_));
  NAi21      u0804(.An(men_men_n158_), .B(men_men_n430_), .Y(men_men_n827_));
  OAI220     u0805(.A0(men_men_n827_), .A1(i_2_), .B0(men_men_n826_), .B1(i_10_), .Y(men_men_n828_));
  NO2        u0806(.A(men_men_n828_), .B(men_men_n825_), .Y(men_men_n829_));
  NO2        u0807(.A(men_men_n383_), .B(men_men_n289_), .Y(men_men_n830_));
  NA2        u0808(.A(men_men_n830_), .B(men_men_n694_), .Y(men_men_n831_));
  NA2        u0809(.A(men_men_n565_), .B(i_0_), .Y(men_men_n832_));
  NO3        u0810(.A(men_men_n832_), .B(men_men_n378_), .C(men_men_n85_), .Y(men_men_n833_));
  NO4        u0811(.A(men_men_n582_), .B(men_men_n209_), .C(men_men_n407_), .D(men_men_n399_), .Y(men_men_n834_));
  AOI210     u0812(.A0(men_men_n834_), .A1(i_11_), .B0(men_men_n833_), .Y(men_men_n835_));
  AN2        u0813(.A(men_men_n94_), .B(men_men_n237_), .Y(men_men_n836_));
  NA2        u0814(.A(men_men_n723_), .B(men_men_n322_), .Y(men_men_n837_));
  AOI210     u0815(.A0(men_men_n472_), .A1(men_men_n85_), .B0(men_men_n58_), .Y(men_men_n838_));
  OAI220     u0816(.A0(men_men_n838_), .A1(men_men_n837_), .B0(men_men_n652_), .B1(men_men_n525_), .Y(men_men_n839_));
  NO2        u0817(.A(men_men_n248_), .B(men_men_n149_), .Y(men_men_n840_));
  NA2        u0818(.A(i_0_), .B(i_10_), .Y(men_men_n841_));
  OAI210     u0819(.A0(men_men_n841_), .A1(men_men_n83_), .B0(men_men_n528_), .Y(men_men_n842_));
  NO4        u0820(.A(men_men_n111_), .B(men_men_n58_), .C(men_men_n657_), .D(i_5_), .Y(men_men_n843_));
  AO220      u0821(.A0(men_men_n843_), .A1(men_men_n842_), .B0(men_men_n840_), .B1(i_6_), .Y(men_men_n844_));
  AOI220     u0822(.A0(i_0_), .A1(men_men_n96_), .B0(men_men_n178_), .B1(men_men_n81_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n559_), .B(i_4_), .Y(men_men_n846_));
  OAI220     u0824(.A0(i_1_), .A1(men_men_n837_), .B0(men_men_n846_), .B1(men_men_n845_), .Y(men_men_n847_));
  NO4        u0825(.A(men_men_n847_), .B(men_men_n844_), .C(men_men_n839_), .D(men_men_n836_), .Y(men_men_n848_));
  NA4        u0826(.A(men_men_n848_), .B(men_men_n835_), .C(men_men_n831_), .D(men_men_n829_), .Y(men_men_n849_));
  NO2        u0827(.A(men_men_n100_), .B(men_men_n37_), .Y(men_men_n850_));
  NA2        u0828(.A(i_11_), .B(i_9_), .Y(men_men_n851_));
  NO3        u0829(.A(i_12_), .B(men_men_n851_), .C(men_men_n599_), .Y(men_men_n852_));
  AN2        u0830(.A(men_men_n852_), .B(men_men_n850_), .Y(men_men_n853_));
  NO2        u0831(.A(men_men_n48_), .B(i_7_), .Y(men_men_n854_));
  INV        u0832(.A(men_men_n156_), .Y(men_men_n855_));
  NO2        u0833(.A(men_men_n851_), .B(men_men_n71_), .Y(men_men_n856_));
  NO2        u0834(.A(men_men_n168_), .B(i_0_), .Y(men_men_n857_));
  INV        u0835(.A(men_men_n857_), .Y(men_men_n858_));
  NA2        u0836(.A(men_men_n465_), .B(men_men_n226_), .Y(men_men_n859_));
  INV        u0837(.A(men_men_n397_), .Y(men_men_n860_));
  OAI220     u0838(.A0(men_men_n860_), .A1(men_men_n817_), .B0(men_men_n859_), .B1(men_men_n858_), .Y(men_men_n861_));
  NO3        u0839(.A(men_men_n861_), .B(men_men_n855_), .C(men_men_n853_), .Y(men_men_n862_));
  NA2        u0840(.A(men_men_n651_), .B(men_men_n117_), .Y(men_men_n863_));
  NO2        u0841(.A(i_6_), .B(men_men_n863_), .Y(men_men_n864_));
  AOI210     u0842(.A0(men_men_n441_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n165_), .B(men_men_n100_), .Y(men_men_n866_));
  NOi32      u0844(.An(men_men_n865_), .Bn(men_men_n181_), .C(men_men_n866_), .Y(men_men_n867_));
  AOI210     u0845(.A0(men_men_n601_), .A1(men_men_n322_), .B0(men_men_n237_), .Y(men_men_n868_));
  NO2        u0846(.A(men_men_n868_), .B(men_men_n808_), .Y(men_men_n869_));
  NO3        u0847(.A(men_men_n869_), .B(men_men_n867_), .C(men_men_n864_), .Y(men_men_n870_));
  NOi21      u0848(.An(i_7_), .B(i_5_), .Y(men_men_n871_));
  NOi31      u0849(.An(men_men_n871_), .B(i_0_), .C(men_men_n705_), .Y(men_men_n872_));
  NA3        u0850(.A(men_men_n872_), .B(men_men_n377_), .C(i_6_), .Y(men_men_n873_));
  OA210      u0851(.A0(men_men_n866_), .A1(men_men_n506_), .B0(men_men_n873_), .Y(men_men_n874_));
  NO2        u0852(.A(men_men_n258_), .B(men_men_n313_), .Y(men_men_n875_));
  NO2        u0853(.A(men_men_n705_), .B(men_men_n253_), .Y(men_men_n876_));
  NA2        u0854(.A(men_men_n876_), .B(men_men_n875_), .Y(men_men_n877_));
  NA4        u0855(.A(men_men_n877_), .B(men_men_n874_), .C(men_men_n870_), .D(men_men_n862_), .Y(men_men_n878_));
  NO2        u0856(.A(men_men_n823_), .B(men_men_n234_), .Y(men_men_n879_));
  AN2        u0857(.A(men_men_n327_), .B(men_men_n322_), .Y(men_men_n880_));
  NA2        u0858(.A(men_men_n879_), .B(i_10_), .Y(men_men_n881_));
  NO2        u0859(.A(men_men_n796_), .B(men_men_n312_), .Y(men_men_n882_));
  OA210      u0860(.A0(men_men_n465_), .A1(men_men_n218_), .B0(men_men_n464_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n882_), .B(men_men_n856_), .Y(men_men_n884_));
  NA3        u0862(.A(men_men_n464_), .B(men_men_n400_), .C(men_men_n45_), .Y(men_men_n885_));
  OAI210     u0863(.A0(men_men_n827_), .A1(i_7_), .B0(men_men_n885_), .Y(men_men_n886_));
  NO2        u0864(.A(men_men_n251_), .B(men_men_n46_), .Y(men_men_n887_));
  NA2        u0865(.A(men_men_n856_), .B(men_men_n300_), .Y(men_men_n888_));
  OAI210     u0866(.A0(men_men_n887_), .A1(men_men_n180_), .B0(men_men_n888_), .Y(men_men_n889_));
  AOI220     u0867(.A0(men_men_n889_), .A1(men_men_n465_), .B0(men_men_n886_), .B1(men_men_n71_), .Y(men_men_n890_));
  NA3        u0868(.A(i_5_), .B(men_men_n375_), .C(men_men_n636_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n90_), .B(men_men_n44_), .Y(men_men_n892_));
  NO2        u0870(.A(men_men_n73_), .B(men_men_n725_), .Y(men_men_n893_));
  AOI220     u0871(.A0(men_men_n893_), .A1(men_men_n892_), .B0(men_men_n167_), .B1(men_men_n590_), .Y(men_men_n894_));
  AOI210     u0872(.A0(men_men_n894_), .A1(men_men_n891_), .B0(men_men_n47_), .Y(men_men_n895_));
  NO3        u0873(.A(men_men_n582_), .B(men_men_n350_), .C(men_men_n24_), .Y(men_men_n896_));
  AOI210     u0874(.A0(men_men_n685_), .A1(men_men_n536_), .B0(men_men_n896_), .Y(men_men_n897_));
  NAi21      u0875(.An(i_9_), .B(i_5_), .Y(men_men_n898_));
  NO2        u0876(.A(men_men_n898_), .B(men_men_n394_), .Y(men_men_n899_));
  NO2        u0877(.A(men_men_n595_), .B(men_men_n102_), .Y(men_men_n900_));
  AOI220     u0878(.A0(men_men_n900_), .A1(i_0_), .B0(men_men_n899_), .B1(men_men_n617_), .Y(men_men_n901_));
  OAI220     u0879(.A0(men_men_n901_), .A1(men_men_n83_), .B0(men_men_n897_), .B1(men_men_n166_), .Y(men_men_n902_));
  NO3        u0880(.A(men_men_n902_), .B(men_men_n895_), .C(men_men_n510_), .Y(men_men_n903_));
  NA4        u0881(.A(men_men_n903_), .B(men_men_n890_), .C(men_men_n884_), .D(men_men_n881_), .Y(men_men_n904_));
  NO3        u0882(.A(men_men_n904_), .B(men_men_n878_), .C(men_men_n849_), .Y(men_men_n905_));
  NO2        u0883(.A(i_0_), .B(men_men_n705_), .Y(men_men_n906_));
  NA2        u0884(.A(men_men_n71_), .B(men_men_n44_), .Y(men_men_n907_));
  NO3        u0885(.A(men_men_n102_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n908_));
  AO220      u0886(.A0(men_men_n908_), .A1(men_men_n44_), .B0(men_men_n906_), .B1(men_men_n167_), .Y(men_men_n909_));
  AOI210     u0887(.A0(men_men_n769_), .A1(men_men_n673_), .B0(men_men_n866_), .Y(men_men_n910_));
  AOI210     u0888(.A0(men_men_n909_), .A1(men_men_n340_), .B0(men_men_n910_), .Y(men_men_n911_));
  NA2        u0889(.A(men_men_n714_), .B(men_men_n141_), .Y(men_men_n912_));
  INV        u0890(.A(men_men_n912_), .Y(men_men_n913_));
  NA2        u0891(.A(men_men_n913_), .B(men_men_n662_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n779_), .B(men_men_n394_), .Y(men_men_n915_));
  NA3        u0893(.A(men_men_n798_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n916_));
  NA2        u0894(.A(men_men_n799_), .B(i_9_), .Y(men_men_n917_));
  AOI210     u0895(.A0(men_men_n916_), .A1(men_men_n486_), .B0(men_men_n917_), .Y(men_men_n918_));
  OAI210     u0896(.A0(men_men_n238_), .A1(i_9_), .B0(men_men_n225_), .Y(men_men_n919_));
  AOI210     u0897(.A0(men_men_n919_), .A1(men_men_n832_), .B0(men_men_n149_), .Y(men_men_n920_));
  NO3        u0898(.A(men_men_n920_), .B(men_men_n918_), .C(men_men_n915_), .Y(men_men_n921_));
  NA3        u0899(.A(men_men_n921_), .B(men_men_n914_), .C(men_men_n911_), .Y(men_men_n922_));
  NA2        u0900(.A(men_men_n880_), .B(men_men_n367_), .Y(men_men_n923_));
  AOI210     u0901(.A0(men_men_n296_), .A1(men_men_n158_), .B0(men_men_n923_), .Y(men_men_n924_));
  INV        u0902(.A(men_men_n924_), .Y(men_men_n925_));
  NO3        u0903(.A(men_men_n841_), .B(men_men_n816_), .C(men_men_n183_), .Y(men_men_n926_));
  NA2        u0904(.A(men_men_n926_), .B(i_11_), .Y(men_men_n927_));
  NO3        u0905(.A(men_men_n204_), .B(men_men_n376_), .C(i_0_), .Y(men_men_n928_));
  OAI210     u0906(.A0(men_men_n928_), .A1(men_men_n74_), .B0(i_13_), .Y(men_men_n929_));
  INV        u0907(.A(men_men_n212_), .Y(men_men_n930_));
  NO2        u0908(.A(i_12_), .B(men_men_n612_), .Y(men_men_n931_));
  NA3        u0909(.A(men_men_n931_), .B(men_men_n392_), .C(men_men_n930_), .Y(men_men_n932_));
  NA4        u0910(.A(men_men_n932_), .B(men_men_n929_), .C(men_men_n927_), .D(men_men_n925_), .Y(men_men_n933_));
  NO2        u0911(.A(men_men_n236_), .B(men_men_n90_), .Y(men_men_n934_));
  AOI210     u0912(.A0(men_men_n934_), .A1(men_men_n906_), .B0(men_men_n105_), .Y(men_men_n935_));
  AOI220     u0913(.A0(men_men_n871_), .A1(men_men_n475_), .B0(men_men_n798_), .B1(men_men_n159_), .Y(men_men_n936_));
  NA2        u0914(.A(men_men_n343_), .B(men_men_n169_), .Y(men_men_n937_));
  OA220      u0915(.A0(men_men_n937_), .A1(men_men_n936_), .B0(men_men_n935_), .B1(i_5_), .Y(men_men_n938_));
  AOI210     u0916(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n168_), .Y(men_men_n939_));
  NA2        u0917(.A(men_men_n939_), .B(men_men_n883_), .Y(men_men_n940_));
  NA3        u0918(.A(men_men_n609_), .B(men_men_n178_), .C(men_men_n81_), .Y(men_men_n941_));
  NA2        u0919(.A(men_men_n941_), .B(men_men_n535_), .Y(men_men_n942_));
  NO3        u0920(.A(men_men_n808_), .B(men_men_n54_), .C(men_men_n48_), .Y(men_men_n943_));
  NA3        u0921(.A(men_men_n480_), .B(men_men_n473_), .C(men_men_n462_), .Y(men_men_n944_));
  NO3        u0922(.A(men_men_n944_), .B(men_men_n943_), .C(men_men_n942_), .Y(men_men_n945_));
  NA3        u0923(.A(men_men_n383_), .B(men_men_n165_), .C(men_men_n164_), .Y(men_men_n946_));
  NA3        u0924(.A(men_men_n383_), .B(men_men_n328_), .C(men_men_n216_), .Y(men_men_n947_));
  INV        u0925(.A(men_men_n947_), .Y(men_men_n948_));
  NOi31      u0926(.An(men_men_n382_), .B(men_men_n907_), .C(men_men_n234_), .Y(men_men_n949_));
  NO3        u0927(.A(men_men_n949_), .B(men_men_n948_), .C(men_men_n1024_), .Y(men_men_n950_));
  NA4        u0928(.A(men_men_n950_), .B(men_men_n945_), .C(men_men_n940_), .D(men_men_n938_), .Y(men_men_n951_));
  INV        u0929(.A(men_men_n611_), .Y(men_men_n952_));
  NO3        u0930(.A(men_men_n952_), .B(men_men_n550_), .C(i_3_), .Y(men_men_n953_));
  NO2        u0931(.A(men_men_n83_), .B(i_5_), .Y(men_men_n954_));
  NA3        u0932(.A(men_men_n799_), .B(men_men_n106_), .C(men_men_n120_), .Y(men_men_n955_));
  INV        u0933(.A(men_men_n955_), .Y(men_men_n956_));
  AOI210     u0934(.A0(men_men_n956_), .A1(men_men_n954_), .B0(men_men_n953_), .Y(men_men_n957_));
  NA3        u0935(.A(men_men_n300_), .B(i_5_), .C(men_men_n186_), .Y(men_men_n958_));
  NO4        u0936(.A(men_men_n234_), .B(men_men_n204_), .C(i_0_), .D(i_12_), .Y(men_men_n959_));
  AOI220     u0937(.A0(men_men_n959_), .A1(i_10_), .B0(men_men_n763_), .B1(men_men_n169_), .Y(men_men_n960_));
  AN2        u0938(.A(men_men_n841_), .B(men_men_n149_), .Y(men_men_n961_));
  NO4        u0939(.A(men_men_n961_), .B(i_12_), .C(men_men_n644_), .D(men_men_n127_), .Y(men_men_n962_));
  NA2        u0940(.A(men_men_n962_), .B(men_men_n212_), .Y(men_men_n963_));
  NA3        u0941(.A(men_men_n96_), .B(men_men_n564_), .C(i_11_), .Y(men_men_n964_));
  NO2        u0942(.A(men_men_n964_), .B(men_men_n151_), .Y(men_men_n965_));
  NA2        u0943(.A(men_men_n871_), .B(men_men_n461_), .Y(men_men_n966_));
  INV        u0944(.A(men_men_n64_), .Y(men_men_n967_));
  OAI220     u0945(.A0(men_men_n967_), .A1(men_men_n958_), .B0(men_men_n966_), .B1(men_men_n663_), .Y(men_men_n968_));
  AOI210     u0946(.A0(men_men_n968_), .A1(men_men_n857_), .B0(men_men_n965_), .Y(men_men_n969_));
  NA4        u0947(.A(men_men_n969_), .B(men_men_n963_), .C(men_men_n960_), .D(men_men_n957_), .Y(men_men_n970_));
  NO4        u0948(.A(men_men_n970_), .B(men_men_n951_), .C(men_men_n933_), .D(men_men_n922_), .Y(men_men_n971_));
  NA2        u0949(.A(men_men_n775_), .B(men_men_n37_), .Y(men_men_n972_));
  NA3        u0950(.A(men_men_n865_), .B(men_men_n362_), .C(i_5_), .Y(men_men_n973_));
  NA3        u0951(.A(men_men_n973_), .B(men_men_n972_), .C(men_men_n607_), .Y(men_men_n974_));
  NA2        u0952(.A(men_men_n974_), .B(men_men_n200_), .Y(men_men_n975_));
  AN2        u0953(.A(men_men_n681_), .B(men_men_n363_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n179_), .B(men_men_n181_), .Y(men_men_n977_));
  AO210      u0955(.A0(men_men_n976_), .A1(men_men_n33_), .B0(men_men_n977_), .Y(men_men_n978_));
  OAI210     u0956(.A0(men_men_n611_), .A1(men_men_n609_), .B0(men_men_n312_), .Y(men_men_n979_));
  NAi31      u0957(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n980_));
  NO2        u0958(.A(men_men_n68_), .B(men_men_n980_), .Y(men_men_n981_));
  NO2        u0959(.A(men_men_n981_), .B(men_men_n641_), .Y(men_men_n982_));
  NA3        u0960(.A(men_men_n982_), .B(men_men_n979_), .C(men_men_n978_), .Y(men_men_n983_));
  NO2        u0961(.A(men_men_n454_), .B(men_men_n261_), .Y(men_men_n984_));
  NO4        u0962(.A(men_men_n228_), .B(men_men_n140_), .C(men_men_n666_), .D(men_men_n37_), .Y(men_men_n985_));
  NO3        u0963(.A(men_men_n985_), .B(men_men_n984_), .C(men_men_n834_), .Y(men_men_n986_));
  OAI210     u0964(.A0(men_men_n964_), .A1(men_men_n143_), .B0(men_men_n986_), .Y(men_men_n987_));
  AOI210     u0965(.A0(men_men_n983_), .A1(men_men_n48_), .B0(men_men_n987_), .Y(men_men_n988_));
  AOI210     u0966(.A0(men_men_n988_), .A1(men_men_n975_), .B0(men_men_n71_), .Y(men_men_n989_));
  NO2        u0967(.A(men_men_n557_), .B(men_men_n372_), .Y(men_men_n990_));
  NO2        u0968(.A(men_men_n990_), .B(men_men_n731_), .Y(men_men_n991_));
  OAI210     u0969(.A0(men_men_n78_), .A1(men_men_n54_), .B0(men_men_n104_), .Y(men_men_n992_));
  NA2        u0970(.A(men_men_n992_), .B(men_men_n74_), .Y(men_men_n993_));
  AOI210     u0971(.A0(men_men_n939_), .A1(men_men_n854_), .B0(men_men_n872_), .Y(men_men_n994_));
  AOI210     u0972(.A0(men_men_n994_), .A1(men_men_n993_), .B0(men_men_n666_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n258_), .B(men_men_n57_), .Y(men_men_n996_));
  AOI220     u0974(.A0(men_men_n996_), .A1(men_men_n74_), .B0(men_men_n338_), .B1(men_men_n250_), .Y(men_men_n997_));
  NO2        u0975(.A(men_men_n997_), .B(men_men_n232_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n94_), .B(men_men_n302_), .C(men_men_n31_), .Y(men_men_n999_));
  INV        u0977(.A(men_men_n999_), .Y(men_men_n1000_));
  NO3        u0978(.A(men_men_n1000_), .B(men_men_n998_), .C(men_men_n995_), .Y(men_men_n1001_));
  OAI210     u0979(.A0(men_men_n263_), .A1(men_men_n154_), .B0(men_men_n85_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n735_), .B(men_men_n285_), .C(men_men_n78_), .Y(men_men_n1003_));
  AOI210     u0981(.A0(men_men_n1003_), .A1(men_men_n1002_), .B0(i_11_), .Y(men_men_n1004_));
  NA2        u0982(.A(men_men_n602_), .B(men_men_n209_), .Y(men_men_n1005_));
  OAI210     u0983(.A0(men_men_n1005_), .A1(men_men_n865_), .B0(men_men_n200_), .Y(men_men_n1006_));
  NA2        u0984(.A(men_men_n160_), .B(i_5_), .Y(men_men_n1007_));
  NO2        u0985(.A(men_men_n1006_), .B(men_men_n1007_), .Y(men_men_n1008_));
  NO3        u0986(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1009_));
  OAI210     u0987(.A0(men_men_n875_), .A1(men_men_n302_), .B0(men_men_n1009_), .Y(men_men_n1010_));
  NO2        u0988(.A(men_men_n1010_), .B(men_men_n705_), .Y(men_men_n1011_));
  NO4        u0989(.A(men_men_n898_), .B(i_11_), .C(men_men_n247_), .D(men_men_n246_), .Y(men_men_n1012_));
  NO2        u0990(.A(men_men_n1012_), .B(men_men_n554_), .Y(men_men_n1013_));
  NO2        u0991(.A(men_men_n778_), .B(men_men_n355_), .Y(men_men_n1014_));
  AOI210     u0992(.A0(men_men_n1014_), .A1(men_men_n1013_), .B0(men_men_n40_), .Y(men_men_n1015_));
  NO4        u0993(.A(men_men_n1015_), .B(men_men_n1011_), .C(men_men_n1008_), .D(men_men_n1004_), .Y(men_men_n1016_));
  OAI210     u0994(.A0(men_men_n1001_), .A1(i_4_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  NO3        u0995(.A(men_men_n1017_), .B(men_men_n991_), .C(men_men_n989_), .Y(men_men_n1018_));
  NA4        u0996(.A(men_men_n1018_), .B(men_men_n971_), .C(men_men_n905_), .D(men_men_n822_), .Y(men4));
  INV        u0997(.A(i_5_), .Y(men_men_n1022_));
  INV        u0998(.A(i_3_), .Y(men_men_n1023_));
  INV        u0999(.A(men_men_n946_), .Y(men_men_n1024_));
  INV        u1000(.A(i_9_), .Y(men_men_n1025_));
  INV        u1001(.A(i_1_), .Y(men_men_n1026_));
  INV        u1002(.A(i_11_), .Y(men_men_n1027_));
  INV        u1003(.A(i_1_), .Y(men_men_n1028_));
  INV        u1004(.A(i_10_), .Y(men_men_n1029_));
  INV        u1005(.A(men_men_n191_), .Y(men_men_n1030_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule