//Benchmark atmr_max1024_476_0.0313

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n62_), .B(ori_ori_n36_), .Y(ori_ori_n63_));
  NO2        o047(.A(x7), .B(x6), .Y(ori_ori_n64_));
  NO2        o048(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n65_));
  NO2        o049(.A(x8), .B(x2), .Y(ori_ori_n66_));
  INV        o050(.A(ori_ori_n66_), .Y(ori_ori_n67_));
  AN2        o051(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  NA2        o055(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n74_));
  NA2        o058(.A(x5), .B(x3), .Y(ori_ori_n75_));
  NO2        o059(.A(x8), .B(x6), .Y(ori_ori_n76_));
  NO4        o060(.A(ori_ori_n76_), .B(ori_ori_n75_), .C(ori_ori_n64_), .D(ori_ori_n54_), .Y(ori_ori_n77_));
  NAi21      o061(.An(x4), .B(x3), .Y(ori_ori_n78_));
  INV        o062(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n22_), .Y(ori_ori_n80_));
  NO2        o064(.A(x4), .B(x2), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n82_));
  NO3        o066(.A(ori_ori_n82_), .B(ori_ori_n80_), .C(ori_ori_n18_), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n84_));
  NA2        o068(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n86_));
  INV        o070(.A(x8), .Y(ori_ori_n87_));
  NA2        o071(.A(x2), .B(x1), .Y(ori_ori_n88_));
  INV        o072(.A(ori_ori_n86_), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n89_), .B(ori_ori_n26_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n91_));
  OAI210     o075(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n92_));
  NO3        o076(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(ori_ori_n90_), .Y(ori_ori_n93_));
  NA2        o077(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n95_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n96_));
  AOI210     o080(.A0(ori_ori_n94_), .A1(ori_ori_n52_), .B0(ori_ori_n96_), .Y(ori_ori_n97_));
  NO2        o081(.A(x3), .B(x2), .Y(ori_ori_n98_));
  NA3        o082(.A(ori_ori_n98_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n99_));
  AOI210     o083(.A0(x8), .A1(x6), .B0(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n101_));
  OAI210     o085(.A0(ori_ori_n101_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n102_));
  NO4        o086(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n97_), .D(ori_ori_n93_), .Y(ori_ori_n103_));
  AO210      o087(.A0(ori_ori_n84_), .A1(ori_ori_n72_), .B0(ori_ori_n103_), .Y(ori02));
  NO2        o088(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n105_));
  NO2        o089(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n108_));
  INV        o092(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  AOI220     o093(.A0(ori_ori_n109_), .A1(ori_ori_n106_), .B0(ori_ori_n105_), .B1(x4), .Y(ori_ori_n110_));
  NO3        o094(.A(ori_ori_n110_), .B(x7), .C(x5), .Y(ori_ori_n111_));
  OR2        o095(.A(x8), .B(x0), .Y(ori_ori_n112_));
  INV        o096(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NAi21      o097(.An(x2), .B(x8), .Y(ori_ori_n114_));
  INV        o098(.A(ori_ori_n114_), .Y(ori_ori_n115_));
  NO2        o099(.A(x4), .B(x1), .Y(ori_ori_n116_));
  NA3        o100(.A(ori_ori_n116_), .B(x2), .C(ori_ori_n60_), .Y(ori_ori_n117_));
  NOi21      o101(.An(x0), .B(x1), .Y(ori_ori_n118_));
  NO3        o102(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n119_));
  NOi21      o103(.An(x0), .B(x4), .Y(ori_ori_n120_));
  NAi21      o104(.An(x8), .B(x7), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n121_), .B(ori_ori_n62_), .Y(ori_ori_n122_));
  AOI220     o106(.A0(ori_ori_n122_), .A1(ori_ori_n120_), .B0(ori_ori_n119_), .B1(ori_ori_n118_), .Y(ori_ori_n123_));
  AOI210     o107(.A0(ori_ori_n123_), .A1(ori_ori_n117_), .B0(ori_ori_n75_), .Y(ori_ori_n124_));
  NO2        o108(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n125_));
  NA2        o109(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n126_));
  AOI210     o110(.A0(ori_ori_n126_), .A1(ori_ori_n101_), .B0(ori_ori_n108_), .Y(ori_ori_n127_));
  OAI210     o111(.A0(ori_ori_n127_), .A1(ori_ori_n35_), .B0(ori_ori_n125_), .Y(ori_ori_n128_));
  NAi21      o112(.An(x0), .B(x4), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n129_), .B(x1), .Y(ori_ori_n130_));
  NO2        o114(.A(x7), .B(x0), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n81_), .B(ori_ori_n95_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n132_), .B(x3), .Y(ori_ori_n133_));
  OAI210     o117(.A0(ori_ori_n131_), .A1(ori_ori_n130_), .B0(ori_ori_n133_), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n135_));
  NA2        o119(.A(x5), .B(x0), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n137_));
  NA3        o121(.A(ori_ori_n137_), .B(ori_ori_n136_), .C(ori_ori_n135_), .Y(ori_ori_n138_));
  NA4        o122(.A(ori_ori_n138_), .B(ori_ori_n134_), .C(ori_ori_n128_), .D(ori_ori_n36_), .Y(ori_ori_n139_));
  NO3        o123(.A(ori_ori_n139_), .B(ori_ori_n124_), .C(ori_ori_n111_), .Y(ori_ori_n140_));
  NO3        o124(.A(ori_ori_n75_), .B(ori_ori_n73_), .C(ori_ori_n24_), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n142_));
  NA2        o126(.A(x7), .B(x3), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n94_), .B(x5), .Y(ori_ori_n144_));
  NO2        o128(.A(x9), .B(x7), .Y(ori_ori_n145_));
  NOi21      o129(.An(x8), .B(x0), .Y(ori_ori_n146_));
  OA210      o130(.A0(ori_ori_n145_), .A1(x1), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n148_));
  INV        o132(.A(x7), .Y(ori_ori_n149_));
  NA2        o133(.A(ori_ori_n149_), .B(ori_ori_n18_), .Y(ori_ori_n150_));
  AOI220     o134(.A0(ori_ori_n150_), .A1(ori_ori_n148_), .B0(ori_ori_n105_), .B1(ori_ori_n38_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n152_), .B(ori_ori_n120_), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n153_), .B(ori_ori_n151_), .Y(ori_ori_n154_));
  AOI210     o138(.A0(ori_ori_n147_), .A1(ori_ori_n144_), .B0(ori_ori_n154_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n143_), .A1(ori_ori_n50_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o140(.A(x5), .B(x1), .Y(ori_ori_n157_));
  INV        o141(.A(ori_ori_n157_), .Y(ori_ori_n158_));
  AOI210     o142(.A0(ori_ori_n158_), .A1(ori_ori_n120_), .B0(ori_ori_n36_), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n62_), .B(ori_ori_n87_), .Y(ori_ori_n160_));
  NAi21      o144(.An(x2), .B(x7), .Y(ori_ori_n161_));
  NO2        o145(.A(ori_ori_n161_), .B(ori_ori_n48_), .Y(ori_ori_n162_));
  NA2        o146(.A(ori_ori_n162_), .B(ori_ori_n65_), .Y(ori_ori_n163_));
  NAi31      o147(.An(ori_ori_n75_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n164_));
  NA3        o148(.A(ori_ori_n164_), .B(ori_ori_n163_), .C(ori_ori_n159_), .Y(ori_ori_n165_));
  NO3        o149(.A(ori_ori_n165_), .B(ori_ori_n156_), .C(ori_ori_n141_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n166_), .B(ori_ori_n140_), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n136_), .B(ori_ori_n132_), .Y(ori_ori_n168_));
  NA2        o152(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n169_));
  NA2        o153(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n170_));
  NA3        o154(.A(ori_ori_n170_), .B(ori_ori_n169_), .C(ori_ori_n24_), .Y(ori_ori_n171_));
  AN2        o155(.A(ori_ori_n171_), .B(ori_ori_n137_), .Y(ori_ori_n172_));
  NA2        o156(.A(x8), .B(x0), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n149_), .B(ori_ori_n25_), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n118_), .B(x4), .Y(ori_ori_n175_));
  NA2        o159(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  AOI210     o160(.A0(ori_ori_n173_), .A1(ori_ori_n126_), .B0(ori_ori_n176_), .Y(ori_ori_n177_));
  NA2        o161(.A(x2), .B(x0), .Y(ori_ori_n178_));
  NA2        o162(.A(x4), .B(x1), .Y(ori_ori_n179_));
  NAi21      o163(.An(ori_ori_n116_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NOi31      o164(.An(ori_ori_n180_), .B(ori_ori_n152_), .C(ori_ori_n178_), .Y(ori_ori_n181_));
  NO4        o165(.A(ori_ori_n181_), .B(ori_ori_n177_), .C(ori_ori_n172_), .D(ori_ori_n168_), .Y(ori_ori_n182_));
  NO2        o166(.A(ori_ori_n182_), .B(ori_ori_n43_), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n171_), .B(ori_ori_n73_), .Y(ori_ori_n184_));
  INV        o168(.A(ori_ori_n125_), .Y(ori_ori_n185_));
  NO2        o169(.A(ori_ori_n101_), .B(ori_ori_n17_), .Y(ori_ori_n186_));
  AOI210     o170(.A0(ori_ori_n35_), .A1(ori_ori_n87_), .B0(ori_ori_n186_), .Y(ori_ori_n187_));
  NO3        o171(.A(ori_ori_n187_), .B(ori_ori_n185_), .C(x7), .Y(ori_ori_n188_));
  NA3        o172(.A(ori_ori_n180_), .B(ori_ori_n185_), .C(ori_ori_n42_), .Y(ori_ori_n189_));
  OAI210     o173(.A0(ori_ori_n170_), .A1(ori_ori_n132_), .B0(ori_ori_n189_), .Y(ori_ori_n190_));
  NO3        o174(.A(ori_ori_n190_), .B(ori_ori_n188_), .C(ori_ori_n184_), .Y(ori_ori_n191_));
  NO2        o175(.A(ori_ori_n191_), .B(x3), .Y(ori_ori_n192_));
  NO3        o176(.A(ori_ori_n192_), .B(ori_ori_n183_), .C(ori_ori_n167_), .Y(ori03));
  NO2        o177(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n194_));
  NO2        o178(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n196_));
  NO2        o180(.A(ori_ori_n75_), .B(x6), .Y(ori_ori_n197_));
  NA2        o181(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n198_));
  NO2        o182(.A(ori_ori_n198_), .B(x4), .Y(ori_ori_n199_));
  NO2        o183(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n200_));
  AO220      o184(.A0(ori_ori_n200_), .A1(ori_ori_n199_), .B0(ori_ori_n197_), .B1(ori_ori_n55_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n201_), .B(ori_ori_n62_), .Y(ori_ori_n202_));
  NA2        o186(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n203_), .B(ori_ori_n198_), .Y(ori_ori_n204_));
  NA2        o188(.A(x9), .B(ori_ori_n54_), .Y(ori_ori_n205_));
  NA2        o189(.A(ori_ori_n205_), .B(x4), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n198_), .B(ori_ori_n78_), .Y(ori_ori_n207_));
  AOI210     o191(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n178_), .Y(ori_ori_n208_));
  AOI220     o192(.A0(ori_ori_n208_), .A1(ori_ori_n207_), .B0(ori_ori_n206_), .B1(ori_ori_n204_), .Y(ori_ori_n209_));
  NO3        o193(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n210_));
  NO2        o194(.A(x5), .B(x1), .Y(ori_ori_n211_));
  NO2        o195(.A(ori_ori_n203_), .B(ori_ori_n169_), .Y(ori_ori_n212_));
  NO3        o196(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n213_));
  NO2        o197(.A(ori_ori_n213_), .B(ori_ori_n212_), .Y(ori_ori_n214_));
  INV        o198(.A(ori_ori_n214_), .Y(ori_ori_n215_));
  AOI220     o199(.A0(ori_ori_n215_), .A1(ori_ori_n48_), .B0(ori_ori_n210_), .B1(ori_ori_n125_), .Y(ori_ori_n216_));
  NA3        o200(.A(ori_ori_n216_), .B(ori_ori_n209_), .C(ori_ori_n202_), .Y(ori_ori_n217_));
  NO2        o201(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n218_));
  NA2        o202(.A(ori_ori_n218_), .B(ori_ori_n19_), .Y(ori_ori_n219_));
  NO2        o203(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n220_));
  NO2        o204(.A(ori_ori_n220_), .B(x6), .Y(ori_ori_n221_));
  NOi21      o205(.An(ori_ori_n81_), .B(ori_ori_n221_), .Y(ori_ori_n222_));
  NA2        o206(.A(ori_ori_n62_), .B(ori_ori_n87_), .Y(ori_ori_n223_));
  NA3        o207(.A(ori_ori_n223_), .B(ori_ori_n220_), .C(x6), .Y(ori_ori_n224_));
  AOI210     o208(.A0(ori_ori_n224_), .A1(ori_ori_n222_), .B0(ori_ori_n149_), .Y(ori_ori_n225_));
  AO210      o209(.A0(ori_ori_n225_), .A1(ori_ori_n219_), .B0(ori_ori_n174_), .Y(ori_ori_n226_));
  NA2        o210(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n227_));
  NA2        o211(.A(ori_ori_n137_), .B(ori_ori_n86_), .Y(ori_ori_n228_));
  NA2        o212(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n229_));
  OAI210     o213(.A0(ori_ori_n113_), .A1(ori_ori_n76_), .B0(x4), .Y(ori_ori_n230_));
  AOI210     o214(.A0(ori_ori_n230_), .A1(ori_ori_n229_), .B0(ori_ori_n75_), .Y(ori_ori_n231_));
  NO2        o215(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n232_));
  NO2        o216(.A(ori_ori_n157_), .B(ori_ori_n43_), .Y(ori_ori_n233_));
  OAI210     o217(.A0(ori_ori_n233_), .A1(ori_ori_n212_), .B0(ori_ori_n232_), .Y(ori_ori_n234_));
  NA2        o218(.A(ori_ori_n195_), .B(ori_ori_n130_), .Y(ori_ori_n235_));
  NA3        o219(.A(ori_ori_n203_), .B(ori_ori_n125_), .C(x6), .Y(ori_ori_n236_));
  OAI210     o220(.A0(ori_ori_n87_), .A1(ori_ori_n36_), .B0(ori_ori_n65_), .Y(ori_ori_n237_));
  NA4        o221(.A(ori_ori_n237_), .B(ori_ori_n236_), .C(ori_ori_n235_), .D(ori_ori_n234_), .Y(ori_ori_n238_));
  OAI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n231_), .B0(x2), .Y(ori_ori_n239_));
  NA3        o223(.A(ori_ori_n239_), .B(ori_ori_n228_), .C(ori_ori_n226_), .Y(ori_ori_n240_));
  AOI210     o224(.A0(ori_ori_n217_), .A1(x8), .B0(ori_ori_n240_), .Y(ori_ori_n241_));
  NO2        o225(.A(ori_ori_n87_), .B(x3), .Y(ori_ori_n242_));
  NA2        o226(.A(ori_ori_n242_), .B(ori_ori_n199_), .Y(ori_ori_n243_));
  NO3        o227(.A(ori_ori_n85_), .B(ori_ori_n76_), .C(ori_ori_n25_), .Y(ori_ori_n244_));
  AOI210     o228(.A0(ori_ori_n221_), .A1(ori_ori_n152_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  AOI210     o229(.A0(ori_ori_n245_), .A1(ori_ori_n243_), .B0(x2), .Y(ori_ori_n246_));
  NO2        o230(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n247_));
  AOI220     o231(.A0(ori_ori_n199_), .A1(ori_ori_n186_), .B0(ori_ori_n247_), .B1(ori_ori_n65_), .Y(ori_ori_n248_));
  NA2        o232(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n249_));
  NA3        o233(.A(ori_ori_n25_), .B(x3), .C(x2), .Y(ori_ori_n250_));
  NO2        o234(.A(ori_ori_n250_), .B(ori_ori_n249_), .Y(ori_ori_n251_));
  NA2        o235(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n252_));
  NO2        o236(.A(ori_ori_n252_), .B(ori_ori_n25_), .Y(ori_ori_n253_));
  OAI210     o237(.A0(ori_ori_n253_), .A1(ori_ori_n251_), .B0(ori_ori_n116_), .Y(ori_ori_n254_));
  NA2        o238(.A(ori_ori_n203_), .B(x6), .Y(ori_ori_n255_));
  NO2        o239(.A(ori_ori_n203_), .B(x6), .Y(ori_ori_n256_));
  NAi21      o240(.An(ori_ori_n160_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  NA3        o241(.A(ori_ori_n257_), .B(ori_ori_n255_), .C(ori_ori_n142_), .Y(ori_ori_n258_));
  NA4        o242(.A(ori_ori_n258_), .B(ori_ori_n254_), .C(ori_ori_n248_), .D(ori_ori_n149_), .Y(ori_ori_n259_));
  NA2        o243(.A(ori_ori_n195_), .B(ori_ori_n220_), .Y(ori_ori_n260_));
  NAi21      o244(.An(x1), .B(x4), .Y(ori_ori_n261_));
  AOI210     o245(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n262_));
  OAI210     o246(.A0(ori_ori_n136_), .A1(x3), .B0(ori_ori_n262_), .Y(ori_ori_n263_));
  NA2        o247(.A(ori_ori_n263_), .B(ori_ori_n261_), .Y(ori_ori_n264_));
  NA2        o248(.A(ori_ori_n264_), .B(ori_ori_n260_), .Y(ori_ori_n265_));
  NA2        o249(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n266_));
  NA2        o250(.A(x6), .B(x2), .Y(ori_ori_n267_));
  NO2        o251(.A(ori_ori_n175_), .B(ori_ori_n46_), .Y(ori_ori_n268_));
  NA2        o252(.A(ori_ori_n268_), .B(ori_ori_n265_), .Y(ori_ori_n269_));
  NA2        o253(.A(x9), .B(ori_ori_n43_), .Y(ori_ori_n270_));
  NO2        o254(.A(ori_ori_n270_), .B(ori_ori_n198_), .Y(ori_ori_n271_));
  OR3        o255(.A(ori_ori_n271_), .B(ori_ori_n197_), .C(ori_ori_n144_), .Y(ori_ori_n272_));
  NA2        o256(.A(x4), .B(x0), .Y(ori_ori_n273_));
  NA2        o257(.A(ori_ori_n272_), .B(ori_ori_n42_), .Y(ori_ori_n274_));
  AOI210     o258(.A0(ori_ori_n274_), .A1(ori_ori_n269_), .B0(x8), .Y(ori_ori_n275_));
  INV        o259(.A(ori_ori_n249_), .Y(ori_ori_n276_));
  NA2        o260(.A(ori_ori_n211_), .B(ori_ori_n276_), .Y(ori_ori_n277_));
  INV        o261(.A(ori_ori_n173_), .Y(ori_ori_n278_));
  OAI210     o262(.A0(ori_ori_n278_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n279_));
  AOI210     o263(.A0(ori_ori_n279_), .A1(ori_ori_n277_), .B0(ori_ori_n227_), .Y(ori_ori_n280_));
  NO4        o264(.A(ori_ori_n280_), .B(ori_ori_n275_), .C(ori_ori_n259_), .D(ori_ori_n246_), .Y(ori_ori_n281_));
  NO2        o265(.A(ori_ori_n160_), .B(x1), .Y(ori_ori_n282_));
  NO3        o266(.A(ori_ori_n282_), .B(x3), .C(ori_ori_n36_), .Y(ori_ori_n283_));
  OAI210     o267(.A0(ori_ori_n283_), .A1(ori_ori_n256_), .B0(x2), .Y(ori_ori_n284_));
  OAI210     o268(.A0(ori_ori_n278_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n285_));
  AOI210     o269(.A0(ori_ori_n285_), .A1(ori_ori_n284_), .B0(ori_ori_n185_), .Y(ori_ori_n286_));
  NOi21      o270(.An(ori_ori_n267_), .B(ori_ori_n17_), .Y(ori_ori_n287_));
  NA3        o271(.A(ori_ori_n287_), .B(ori_ori_n211_), .C(ori_ori_n40_), .Y(ori_ori_n288_));
  AOI210     o272(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n289_));
  NA3        o273(.A(ori_ori_n289_), .B(ori_ori_n158_), .C(ori_ori_n32_), .Y(ori_ori_n290_));
  NA2        o274(.A(x3), .B(x2), .Y(ori_ori_n291_));
  AOI220     o275(.A0(ori_ori_n291_), .A1(ori_ori_n227_), .B0(ori_ori_n290_), .B1(ori_ori_n288_), .Y(ori_ori_n292_));
  NAi21      o276(.An(x4), .B(x0), .Y(ori_ori_n293_));
  NO3        o277(.A(ori_ori_n293_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n294_));
  OAI210     o278(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  OAI220     o279(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n296_));
  NO2        o280(.A(x9), .B(x8), .Y(ori_ori_n297_));
  NO2        o281(.A(ori_ori_n289_), .B(ori_ori_n287_), .Y(ori_ori_n298_));
  AOI220     o282(.A0(ori_ori_n298_), .A1(ori_ori_n79_), .B0(ori_ori_n296_), .B1(ori_ori_n31_), .Y(ori_ori_n299_));
  AOI210     o283(.A0(ori_ori_n299_), .A1(ori_ori_n295_), .B0(ori_ori_n25_), .Y(ori_ori_n300_));
  NA3        o284(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n301_));
  OAI210     o285(.A0(ori_ori_n289_), .A1(ori_ori_n287_), .B0(ori_ori_n301_), .Y(ori_ori_n302_));
  INV        o286(.A(ori_ori_n212_), .Y(ori_ori_n303_));
  NA2        o287(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n304_));
  OR2        o288(.A(ori_ori_n304_), .B(ori_ori_n273_), .Y(ori_ori_n305_));
  OAI220     o289(.A0(ori_ori_n305_), .A1(ori_ori_n157_), .B0(ori_ori_n229_), .B1(ori_ori_n303_), .Y(ori_ori_n306_));
  AO210      o290(.A0(ori_ori_n302_), .A1(ori_ori_n144_), .B0(ori_ori_n306_), .Y(ori_ori_n307_));
  NO4        o291(.A(ori_ori_n307_), .B(ori_ori_n300_), .C(ori_ori_n292_), .D(ori_ori_n286_), .Y(ori_ori_n308_));
  OAI210     o292(.A0(ori_ori_n281_), .A1(ori_ori_n241_), .B0(ori_ori_n308_), .Y(ori04));
  NO2        o293(.A(x2), .B(x1), .Y(ori_ori_n310_));
  OAI210     o294(.A0(ori_ori_n252_), .A1(ori_ori_n310_), .B0(ori_ori_n36_), .Y(ori_ori_n311_));
  NO2        o295(.A(ori_ori_n310_), .B(ori_ori_n293_), .Y(ori_ori_n312_));
  AOI210     o296(.A0(ori_ori_n62_), .A1(x4), .B0(ori_ori_n107_), .Y(ori_ori_n313_));
  OAI210     o297(.A0(ori_ori_n313_), .A1(ori_ori_n312_), .B0(ori_ori_n242_), .Y(ori_ori_n314_));
  NO2        o298(.A(ori_ori_n266_), .B(ori_ori_n85_), .Y(ori_ori_n315_));
  NO2        o299(.A(ori_ori_n315_), .B(ori_ori_n36_), .Y(ori_ori_n316_));
  NO2        o300(.A(ori_ori_n291_), .B(ori_ori_n200_), .Y(ori_ori_n317_));
  NA2        o301(.A(x9), .B(x0), .Y(ori_ori_n318_));
  AOI210     o302(.A0(ori_ori_n85_), .A1(ori_ori_n73_), .B0(ori_ori_n318_), .Y(ori_ori_n319_));
  OAI210     o303(.A0(ori_ori_n319_), .A1(ori_ori_n317_), .B0(ori_ori_n87_), .Y(ori_ori_n320_));
  NA3        o304(.A(ori_ori_n320_), .B(ori_ori_n316_), .C(ori_ori_n314_), .Y(ori_ori_n321_));
  NA2        o305(.A(ori_ori_n321_), .B(ori_ori_n311_), .Y(ori_ori_n322_));
  NO2        o306(.A(ori_ori_n205_), .B(ori_ori_n108_), .Y(ori_ori_n323_));
  NO3        o307(.A(ori_ori_n249_), .B(ori_ori_n114_), .C(ori_ori_n18_), .Y(ori_ori_n324_));
  NO2        o308(.A(ori_ori_n324_), .B(ori_ori_n323_), .Y(ori_ori_n325_));
  OAI210     o309(.A0(ori_ori_n112_), .A1(ori_ori_n101_), .B0(ori_ori_n173_), .Y(ori_ori_n326_));
  NA3        o310(.A(ori_ori_n326_), .B(x6), .C(x3), .Y(ori_ori_n327_));
  NOi21      o311(.An(ori_ori_n146_), .B(ori_ori_n126_), .Y(ori_ori_n328_));
  AOI210     o312(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n329_));
  OAI220     o313(.A0(ori_ori_n329_), .A1(ori_ori_n304_), .B0(ori_ori_n266_), .B1(ori_ori_n301_), .Y(ori_ori_n330_));
  AOI210     o314(.A0(ori_ori_n328_), .A1(ori_ori_n63_), .B0(ori_ori_n330_), .Y(ori_ori_n331_));
  NA2        o315(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n332_));
  OAI210     o316(.A0(ori_ori_n101_), .A1(ori_ori_n17_), .B0(ori_ori_n332_), .Y(ori_ori_n333_));
  NA2        o317(.A(ori_ori_n333_), .B(ori_ori_n76_), .Y(ori_ori_n334_));
  NA4        o318(.A(ori_ori_n334_), .B(ori_ori_n331_), .C(ori_ori_n327_), .D(ori_ori_n325_), .Y(ori_ori_n335_));
  OAI210     o319(.A0(ori_ori_n106_), .A1(x3), .B0(ori_ori_n294_), .Y(ori_ori_n336_));
  NA2        o320(.A(ori_ori_n210_), .B(ori_ori_n81_), .Y(ori_ori_n337_));
  NA3        o321(.A(ori_ori_n337_), .B(ori_ori_n336_), .C(ori_ori_n149_), .Y(ori_ori_n338_));
  AOI210     o322(.A0(ori_ori_n335_), .A1(x4), .B0(ori_ori_n338_), .Y(ori_ori_n339_));
  NA3        o323(.A(ori_ori_n312_), .B(ori_ori_n205_), .C(ori_ori_n87_), .Y(ori_ori_n340_));
  NOi21      o324(.An(x4), .B(x0), .Y(ori_ori_n341_));
  XO2        o325(.A(x4), .B(x0), .Y(ori_ori_n342_));
  INV        o326(.A(ori_ori_n261_), .Y(ori_ori_n343_));
  AOI220     o327(.A0(ori_ori_n343_), .A1(x8), .B0(ori_ori_n341_), .B1(ori_ori_n88_), .Y(ori_ori_n344_));
  AOI210     o328(.A0(ori_ori_n344_), .A1(ori_ori_n340_), .B0(x3), .Y(ori_ori_n345_));
  INV        o329(.A(ori_ori_n88_), .Y(ori_ori_n346_));
  NO2        o330(.A(ori_ori_n87_), .B(x4), .Y(ori_ori_n347_));
  AOI220     o331(.A0(ori_ori_n347_), .A1(ori_ori_n44_), .B0(ori_ori_n120_), .B1(ori_ori_n346_), .Y(ori_ori_n348_));
  NO3        o332(.A(ori_ori_n342_), .B(ori_ori_n160_), .C(x2), .Y(ori_ori_n349_));
  INV        o333(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NA4        o334(.A(ori_ori_n350_), .B(ori_ori_n348_), .C(ori_ori_n219_), .D(x6), .Y(ori_ori_n351_));
  OAI220     o335(.A0(ori_ori_n293_), .A1(ori_ori_n85_), .B0(ori_ori_n178_), .B1(ori_ori_n87_), .Y(ori_ori_n352_));
  NO2        o336(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n353_));
  NA2        o337(.A(ori_ori_n352_), .B(ori_ori_n61_), .Y(ori_ori_n354_));
  NO2        o338(.A(ori_ori_n146_), .B(ori_ori_n78_), .Y(ori_ori_n355_));
  NO2        o339(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n356_));
  NOi21      o340(.An(ori_ori_n116_), .B(ori_ori_n27_), .Y(ori_ori_n357_));
  AOI210     o341(.A0(ori_ori_n356_), .A1(ori_ori_n355_), .B0(ori_ori_n357_), .Y(ori_ori_n358_));
  OAI210     o342(.A0(ori_ori_n354_), .A1(ori_ori_n62_), .B0(ori_ori_n358_), .Y(ori_ori_n359_));
  OAI220     o343(.A0(ori_ori_n359_), .A1(x6), .B0(ori_ori_n351_), .B1(ori_ori_n345_), .Y(ori_ori_n360_));
  OAI210     o344(.A0(ori_ori_n63_), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n361_));
  OAI210     o345(.A0(ori_ori_n361_), .A1(ori_ori_n87_), .B0(ori_ori_n305_), .Y(ori_ori_n362_));
  AOI210     o346(.A0(ori_ori_n362_), .A1(ori_ori_n18_), .B0(ori_ori_n149_), .Y(ori_ori_n363_));
  AO220      o347(.A0(ori_ori_n363_), .A1(ori_ori_n360_), .B0(ori_ori_n339_), .B1(ori_ori_n322_), .Y(ori_ori_n364_));
  NA2        o348(.A(ori_ori_n356_), .B(x6), .Y(ori_ori_n365_));
  AOI210     o349(.A0(x6), .A1(x1), .B0(ori_ori_n148_), .Y(ori_ori_n366_));
  NA2        o350(.A(ori_ori_n347_), .B(x0), .Y(ori_ori_n367_));
  NA2        o351(.A(ori_ori_n81_), .B(x6), .Y(ori_ori_n368_));
  OAI210     o352(.A0(ori_ori_n367_), .A1(ori_ori_n366_), .B0(ori_ori_n368_), .Y(ori_ori_n369_));
  AOI220     o353(.A0(ori_ori_n369_), .A1(ori_ori_n365_), .B0(ori_ori_n213_), .B1(ori_ori_n49_), .Y(ori_ori_n370_));
  NA2        o354(.A(ori_ori_n370_), .B(ori_ori_n364_), .Y(ori_ori_n371_));
  AOI210     o355(.A0(ori_ori_n196_), .A1(x8), .B0(ori_ori_n106_), .Y(ori_ori_n372_));
  NA2        o356(.A(ori_ori_n372_), .B(ori_ori_n332_), .Y(ori_ori_n373_));
  NA3        o357(.A(ori_ori_n373_), .B(ori_ori_n194_), .C(ori_ori_n149_), .Y(ori_ori_n374_));
  OAI210     o358(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n227_), .Y(ori_ori_n375_));
  AO220      o359(.A0(ori_ori_n375_), .A1(ori_ori_n145_), .B0(ori_ori_n105_), .B1(x4), .Y(ori_ori_n376_));
  NA3        o360(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n377_));
  NA2        o361(.A(ori_ori_n218_), .B(x0), .Y(ori_ori_n378_));
  OAI220     o362(.A0(ori_ori_n378_), .A1(ori_ori_n205_), .B0(ori_ori_n377_), .B1(ori_ori_n346_), .Y(ori_ori_n379_));
  AOI210     o363(.A0(ori_ori_n376_), .A1(ori_ori_n113_), .B0(ori_ori_n379_), .Y(ori_ori_n380_));
  AOI210     o364(.A0(ori_ori_n380_), .A1(ori_ori_n374_), .B0(ori_ori_n25_), .Y(ori_ori_n381_));
  NA3        o365(.A(ori_ori_n115_), .B(ori_ori_n218_), .C(x0), .Y(ori_ori_n382_));
  AOI210     o366(.A0(ori_ori_n114_), .A1(ori_ori_n112_), .B0(ori_ori_n42_), .Y(ori_ori_n383_));
  NAi31      o367(.An(ori_ori_n50_), .B(ori_ori_n282_), .C(ori_ori_n174_), .Y(ori_ori_n384_));
  NA2        o368(.A(ori_ori_n384_), .B(ori_ori_n382_), .Y(ori_ori_n385_));
  OAI210     o369(.A0(ori_ori_n385_), .A1(ori_ori_n381_), .B0(x6), .Y(ori_ori_n386_));
  OAI210     o370(.A0(ori_ori_n160_), .A1(ori_ori_n48_), .B0(ori_ori_n131_), .Y(ori_ori_n387_));
  NA3        o371(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n388_));
  AOI220     o372(.A0(ori_ori_n388_), .A1(ori_ori_n387_), .B0(ori_ori_n40_), .B1(ori_ori_n32_), .Y(ori_ori_n389_));
  NO2        o373(.A(ori_ori_n149_), .B(x0), .Y(ori_ori_n390_));
  AOI220     o374(.A0(ori_ori_n390_), .A1(ori_ori_n218_), .B0(ori_ori_n194_), .B1(ori_ori_n149_), .Y(ori_ori_n391_));
  AOI210     o375(.A0(ori_ori_n122_), .A1(ori_ori_n247_), .B0(x1), .Y(ori_ori_n392_));
  OAI210     o376(.A0(ori_ori_n391_), .A1(x8), .B0(ori_ori_n392_), .Y(ori_ori_n393_));
  NAi31      o377(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n394_));
  OAI210     o378(.A0(ori_ori_n394_), .A1(x4), .B0(ori_ori_n161_), .Y(ori_ori_n395_));
  NA3        o379(.A(ori_ori_n395_), .B(ori_ori_n143_), .C(x9), .Y(ori_ori_n396_));
  NO3        o380(.A(x9), .B(ori_ori_n149_), .C(x0), .Y(ori_ori_n397_));
  AOI220     o381(.A0(ori_ori_n397_), .A1(ori_ori_n242_), .B0(ori_ori_n355_), .B1(ori_ori_n149_), .Y(ori_ori_n398_));
  NA4        o382(.A(ori_ori_n398_), .B(x1), .C(ori_ori_n396_), .D(ori_ori_n50_), .Y(ori_ori_n399_));
  OAI210     o383(.A0(ori_ori_n393_), .A1(ori_ori_n389_), .B0(ori_ori_n399_), .Y(ori_ori_n400_));
  NOi31      o384(.An(ori_ori_n390_), .B(ori_ori_n32_), .C(x8), .Y(ori_ori_n401_));
  AOI210     o385(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n129_), .Y(ori_ori_n402_));
  NO3        o386(.A(ori_ori_n402_), .B(ori_ori_n119_), .C(ori_ori_n43_), .Y(ori_ori_n403_));
  NOi31      o387(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n404_));
  AOI220     o388(.A0(ori_ori_n404_), .A1(ori_ori_n341_), .B0(ori_ori_n120_), .B1(x3), .Y(ori_ori_n405_));
  AOI210     o389(.A0(ori_ori_n261_), .A1(ori_ori_n60_), .B0(ori_ori_n118_), .Y(ori_ori_n406_));
  OAI210     o390(.A0(ori_ori_n406_), .A1(x3), .B0(ori_ori_n405_), .Y(ori_ori_n407_));
  NO3        o391(.A(ori_ori_n407_), .B(ori_ori_n403_), .C(x2), .Y(ori_ori_n408_));
  OAI220     o392(.A0(ori_ori_n342_), .A1(ori_ori_n297_), .B0(ori_ori_n293_), .B1(ori_ori_n43_), .Y(ori_ori_n409_));
  AOI210     o393(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n377_), .Y(ori_ori_n410_));
  AOI220     o394(.A0(ori_ori_n410_), .A1(ori_ori_n87_), .B0(ori_ori_n409_), .B1(ori_ori_n149_), .Y(ori_ori_n411_));
  NO2        o395(.A(ori_ori_n411_), .B(ori_ori_n54_), .Y(ori_ori_n412_));
  NO3        o396(.A(ori_ori_n412_), .B(ori_ori_n408_), .C(ori_ori_n401_), .Y(ori_ori_n413_));
  AOI210     o397(.A0(ori_ori_n413_), .A1(ori_ori_n400_), .B0(ori_ori_n25_), .Y(ori_ori_n414_));
  NA4        o398(.A(ori_ori_n31_), .B(ori_ori_n87_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n415_));
  NO3        o399(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n416_));
  NO3        o400(.A(ori_ori_n66_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n417_));
  AOI220     o401(.A0(ori_ori_n417_), .A1(ori_ori_n262_), .B0(ori_ori_n416_), .B1(ori_ori_n383_), .Y(ori_ori_n418_));
  NO2        o402(.A(ori_ori_n418_), .B(ori_ori_n98_), .Y(ori_ori_n419_));
  NO3        o403(.A(ori_ori_n266_), .B(ori_ori_n173_), .C(ori_ori_n40_), .Y(ori_ori_n420_));
  OAI210     o404(.A0(ori_ori_n420_), .A1(ori_ori_n419_), .B0(x7), .Y(ori_ori_n421_));
  NA2        o405(.A(ori_ori_n223_), .B(x7), .Y(ori_ori_n422_));
  NA3        o406(.A(ori_ori_n422_), .B(ori_ori_n148_), .C(ori_ori_n130_), .Y(ori_ori_n423_));
  NA3        o407(.A(ori_ori_n423_), .B(ori_ori_n421_), .C(ori_ori_n415_), .Y(ori_ori_n424_));
  OAI210     o408(.A0(ori_ori_n424_), .A1(ori_ori_n414_), .B0(ori_ori_n36_), .Y(ori_ori_n425_));
  NO2        o409(.A(ori_ori_n397_), .B(ori_ori_n200_), .Y(ori_ori_n426_));
  NO4        o410(.A(ori_ori_n426_), .B(ori_ori_n75_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n427_));
  NA2        o411(.A(ori_ori_n252_), .B(ori_ori_n21_), .Y(ori_ori_n428_));
  NO2        o412(.A(ori_ori_n157_), .B(ori_ori_n131_), .Y(ori_ori_n429_));
  NA2        o413(.A(ori_ori_n429_), .B(ori_ori_n428_), .Y(ori_ori_n430_));
  AOI210     o414(.A0(ori_ori_n430_), .A1(ori_ori_n164_), .B0(ori_ori_n28_), .Y(ori_ori_n431_));
  AOI220     o415(.A0(ori_ori_n353_), .A1(ori_ori_n87_), .B0(ori_ori_n146_), .B1(ori_ori_n196_), .Y(ori_ori_n432_));
  NA3        o416(.A(ori_ori_n432_), .B(ori_ori_n394_), .C(ori_ori_n85_), .Y(ori_ori_n433_));
  NA2        o417(.A(ori_ori_n433_), .B(ori_ori_n174_), .Y(ori_ori_n434_));
  OAI220     o418(.A0(ori_ori_n270_), .A1(ori_ori_n67_), .B0(ori_ori_n157_), .B1(ori_ori_n43_), .Y(ori_ori_n435_));
  NA2        o419(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n436_));
  OAI210     o420(.A0(ori_ori_n145_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n437_));
  NO3        o421(.A(ori_ori_n404_), .B(x3), .C(ori_ori_n54_), .Y(ori_ori_n438_));
  NA2        o422(.A(ori_ori_n438_), .B(ori_ori_n437_), .Y(ori_ori_n439_));
  OAI210     o423(.A0(ori_ori_n150_), .A1(ori_ori_n436_), .B0(ori_ori_n439_), .Y(ori_ori_n440_));
  AOI220     o424(.A0(ori_ori_n440_), .A1(x0), .B0(ori_ori_n435_), .B1(ori_ori_n131_), .Y(ori_ori_n441_));
  AOI210     o425(.A0(ori_ori_n441_), .A1(ori_ori_n434_), .B0(ori_ori_n229_), .Y(ori_ori_n442_));
  NO3        o426(.A(ori_ori_n442_), .B(ori_ori_n431_), .C(ori_ori_n427_), .Y(ori_ori_n443_));
  NA3        o427(.A(ori_ori_n443_), .B(ori_ori_n425_), .C(ori_ori_n386_), .Y(ori_ori_n444_));
  AOI210     o428(.A0(ori_ori_n371_), .A1(ori_ori_n25_), .B0(ori_ori_n444_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n24_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  OA210      m015(.A0(mai_mai_n31_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n23_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n25_), .Y(mai_mai_n36_));
  AN2        m020(.A(x8), .B(x7), .Y(mai_mai_n37_));
  NA2        m021(.A(x4), .B(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n23_), .B(mai_mai_n38_), .Y(mai_mai_n39_));
  NO2        m023(.A(x2), .B(x0), .Y(mai_mai_n40_));
  INV        m024(.A(x3), .Y(mai_mai_n41_));
  NO2        m025(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n42_));
  INV        m026(.A(mai_mai_n42_), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n44_));
  OAI210     m028(.A0(mai_mai_n44_), .A1(mai_mai_n43_), .B0(mai_mai_n40_), .Y(mai_mai_n45_));
  INV        m029(.A(x4), .Y(mai_mai_n46_));
  NO2        m030(.A(mai_mai_n46_), .B(mai_mai_n17_), .Y(mai_mai_n47_));
  NA2        m031(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n48_));
  OAI210     m032(.A0(mai_mai_n48_), .A1(mai_mai_n20_), .B0(mai_mai_n45_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n50_));
  AOI220     m034(.A0(mai_mai_n50_), .A1(mai_mai_n34_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n51_));
  INV        m035(.A(x2), .Y(mai_mai_n52_));
  NO2        m036(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n55_));
  OAI210     m039(.A0(mai_mai_n51_), .A1(mai_mai_n31_), .B0(mai_mai_n55_), .Y(mai_mai_n56_));
  NO3        m040(.A(mai_mai_n56_), .B(mai_mai_n49_), .C(mai_mai_n39_), .Y(mai01));
  NA2        m041(.A(x8), .B(x7), .Y(mai_mai_n58_));
  NA2        m042(.A(mai_mai_n41_), .B(x1), .Y(mai_mai_n59_));
  INV        m043(.A(x9), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n60_), .B(mai_mai_n35_), .Y(mai_mai_n61_));
  INV        m045(.A(mai_mai_n61_), .Y(mai_mai_n62_));
  NO3        m046(.A(mai_mai_n62_), .B(mai_mai_n59_), .C(mai_mai_n58_), .Y(mai_mai_n63_));
  NO2        m047(.A(x7), .B(x6), .Y(mai_mai_n64_));
  NO2        m048(.A(mai_mai_n59_), .B(x5), .Y(mai_mai_n65_));
  NO2        m049(.A(x8), .B(x2), .Y(mai_mai_n66_));
  INV        m050(.A(mai_mai_n66_), .Y(mai_mai_n67_));
  NO2        m051(.A(mai_mai_n67_), .B(x1), .Y(mai_mai_n68_));
  OA210      m052(.A0(mai_mai_n68_), .A1(mai_mai_n65_), .B0(mai_mai_n64_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n42_), .A1(mai_mai_n25_), .B0(mai_mai_n52_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n54_), .A1(mai_mai_n20_), .B0(mai_mai_n70_), .Y(mai_mai_n71_));
  NAi31      m055(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n72_));
  NO2        m056(.A(mai_mai_n71_), .B(mai_mai_n69_), .Y(mai_mai_n73_));
  OAI210     m057(.A0(mai_mai_n73_), .A1(mai_mai_n63_), .B0(x4), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n75_));
  OAI210     m059(.A0(mai_mai_n75_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n76_));
  NA2        m060(.A(x5), .B(x3), .Y(mai_mai_n77_));
  NO2        m061(.A(x8), .B(x6), .Y(mai_mai_n78_));
  NO4        m062(.A(mai_mai_n78_), .B(mai_mai_n77_), .C(mai_mai_n64_), .D(mai_mai_n52_), .Y(mai_mai_n79_));
  NAi21      m063(.An(x4), .B(x3), .Y(mai_mai_n80_));
  INV        m064(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m065(.A(mai_mai_n81_), .B(mai_mai_n22_), .Y(mai_mai_n82_));
  NO2        m066(.A(x4), .B(x2), .Y(mai_mai_n83_));
  NO2        m067(.A(mai_mai_n83_), .B(x3), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n82_), .C(mai_mai_n18_), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n79_), .C(mai_mai_n76_), .Y(mai_mai_n86_));
  NO4        m070(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n41_), .D(x1), .Y(mai_mai_n87_));
  NA2        m071(.A(mai_mai_n60_), .B(mai_mai_n46_), .Y(mai_mai_n88_));
  INV        m072(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OAI210     m073(.A0(mai_mai_n87_), .A1(mai_mai_n65_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NA2        m074(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n91_));
  NO2        m075(.A(mai_mai_n91_), .B(mai_mai_n25_), .Y(mai_mai_n92_));
  INV        m076(.A(x8), .Y(mai_mai_n93_));
  NA2        m077(.A(x2), .B(x1), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n92_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n96_), .B(mai_mai_n26_), .Y(mai_mai_n97_));
  AOI210     m081(.A0(mai_mai_n54_), .A1(mai_mai_n25_), .B0(mai_mai_n52_), .Y(mai_mai_n98_));
  OAI210     m082(.A0(mai_mai_n43_), .A1(mai_mai_n36_), .B0(mai_mai_n46_), .Y(mai_mai_n99_));
  NO3        m083(.A(mai_mai_n99_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n100_));
  NA2        m084(.A(x4), .B(mai_mai_n41_), .Y(mai_mai_n101_));
  NO2        m085(.A(mai_mai_n46_), .B(mai_mai_n52_), .Y(mai_mai_n102_));
  OAI210     m086(.A0(mai_mai_n102_), .A1(mai_mai_n41_), .B0(mai_mai_n18_), .Y(mai_mai_n103_));
  AOI210     m087(.A0(mai_mai_n101_), .A1(mai_mai_n50_), .B0(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m088(.A(x3), .B(x2), .Y(mai_mai_n105_));
  NA3        m089(.A(mai_mai_n105_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n106_));
  AOI210     m090(.A0(x8), .A1(x6), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  NA2        m091(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n108_));
  OAI210     m092(.A0(mai_mai_n108_), .A1(mai_mai_n38_), .B0(mai_mai_n17_), .Y(mai_mai_n109_));
  NO4        m093(.A(mai_mai_n109_), .B(mai_mai_n107_), .C(mai_mai_n104_), .D(mai_mai_n100_), .Y(mai_mai_n110_));
  AO220      m094(.A0(mai_mai_n110_), .A1(mai_mai_n90_), .B0(mai_mai_n86_), .B1(mai_mai_n74_), .Y(mai02));
  NO2        m095(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n112_));
  NO2        m096(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n113_));
  NA2        m097(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n114_));
  NA2        m098(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n115_));
  OAI210     m099(.A0(mai_mai_n88_), .A1(mai_mai_n114_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  AOI220     m100(.A0(mai_mai_n116_), .A1(mai_mai_n113_), .B0(mai_mai_n112_), .B1(x4), .Y(mai_mai_n117_));
  NO3        m101(.A(mai_mai_n117_), .B(x7), .C(x5), .Y(mai_mai_n118_));
  NA2        m102(.A(x9), .B(x2), .Y(mai_mai_n119_));
  OR2        m103(.A(x8), .B(x0), .Y(mai_mai_n120_));
  INV        m104(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NAi21      m105(.An(x2), .B(x8), .Y(mai_mai_n122_));
  INV        m106(.A(mai_mai_n122_), .Y(mai_mai_n123_));
  OAI220     m107(.A0(mai_mai_n123_), .A1(mai_mai_n121_), .B0(mai_mai_n119_), .B1(x7), .Y(mai_mai_n124_));
  NO2        m108(.A(x4), .B(x1), .Y(mai_mai_n125_));
  NA3        m109(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(mai_mai_n58_), .Y(mai_mai_n126_));
  NOi21      m110(.An(x0), .B(x1), .Y(mai_mai_n127_));
  NO3        m111(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n128_));
  NOi21      m112(.An(x0), .B(x4), .Y(mai_mai_n129_));
  NAi21      m113(.An(x8), .B(x7), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n130_), .B(mai_mai_n60_), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n126_), .B(mai_mai_n77_), .Y(mai_mai_n132_));
  NO2        m116(.A(x5), .B(mai_mai_n46_), .Y(mai_mai_n133_));
  NA2        m117(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n134_));
  AOI210     m118(.A0(mai_mai_n134_), .A1(mai_mai_n108_), .B0(mai_mai_n115_), .Y(mai_mai_n135_));
  OAI210     m119(.A0(mai_mai_n135_), .A1(mai_mai_n34_), .B0(mai_mai_n133_), .Y(mai_mai_n136_));
  NAi21      m120(.An(x0), .B(x4), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n137_), .B(x1), .Y(mai_mai_n138_));
  NO2        m122(.A(x7), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n83_), .B(mai_mai_n102_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n140_), .B(x3), .Y(mai_mai_n141_));
  OAI210     m125(.A0(mai_mai_n139_), .A1(mai_mai_n138_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n21_), .B(mai_mai_n41_), .Y(mai_mai_n143_));
  NA2        m127(.A(x5), .B(x0), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n145_));
  NA3        m129(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(mai_mai_n143_), .Y(mai_mai_n146_));
  NA4        m130(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n136_), .D(mai_mai_n35_), .Y(mai_mai_n147_));
  NO3        m131(.A(mai_mai_n147_), .B(mai_mai_n132_), .C(mai_mai_n118_), .Y(mai_mai_n148_));
  NO3        m132(.A(mai_mai_n77_), .B(mai_mai_n75_), .C(mai_mai_n24_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n150_));
  AOI220     m134(.A0(mai_mai_n127_), .A1(mai_mai_n150_), .B0(mai_mai_n65_), .B1(mai_mai_n17_), .Y(mai_mai_n151_));
  NO3        m135(.A(mai_mai_n151_), .B(mai_mai_n58_), .C(mai_mai_n60_), .Y(mai_mai_n152_));
  NA2        m136(.A(x7), .B(x3), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n101_), .B(x5), .Y(mai_mai_n154_));
  NO2        m138(.A(x9), .B(x7), .Y(mai_mai_n155_));
  NOi21      m139(.An(x8), .B(x0), .Y(mai_mai_n156_));
  OA210      m140(.A0(mai_mai_n155_), .A1(x1), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NO2        m141(.A(mai_mai_n41_), .B(x2), .Y(mai_mai_n158_));
  INV        m142(.A(x7), .Y(mai_mai_n159_));
  NA2        m143(.A(mai_mai_n159_), .B(mai_mai_n18_), .Y(mai_mai_n160_));
  AOI220     m144(.A0(mai_mai_n160_), .A1(mai_mai_n158_), .B0(mai_mai_n112_), .B1(mai_mai_n37_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n162_));
  NO2        m146(.A(mai_mai_n162_), .B(mai_mai_n129_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n163_), .B(mai_mai_n161_), .Y(mai_mai_n164_));
  AOI210     m148(.A0(mai_mai_n157_), .A1(mai_mai_n154_), .B0(mai_mai_n164_), .Y(mai_mai_n165_));
  OAI210     m149(.A0(mai_mai_n153_), .A1(mai_mai_n48_), .B0(mai_mai_n165_), .Y(mai_mai_n166_));
  NA2        m150(.A(x5), .B(x1), .Y(mai_mai_n167_));
  INV        m151(.A(mai_mai_n167_), .Y(mai_mai_n168_));
  AOI210     m152(.A0(mai_mai_n168_), .A1(mai_mai_n129_), .B0(mai_mai_n35_), .Y(mai_mai_n169_));
  NO2        m153(.A(mai_mai_n60_), .B(mai_mai_n93_), .Y(mai_mai_n170_));
  NAi21      m154(.An(x2), .B(x7), .Y(mai_mai_n171_));
  NO3        m155(.A(mai_mai_n171_), .B(mai_mai_n170_), .C(mai_mai_n46_), .Y(mai_mai_n172_));
  NA2        m156(.A(mai_mai_n172_), .B(mai_mai_n65_), .Y(mai_mai_n173_));
  NA2        m157(.A(mai_mai_n173_), .B(mai_mai_n169_), .Y(mai_mai_n174_));
  NO4        m158(.A(mai_mai_n174_), .B(mai_mai_n166_), .C(mai_mai_n152_), .D(mai_mai_n149_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n175_), .B(mai_mai_n148_), .Y(mai_mai_n176_));
  NO2        m160(.A(mai_mai_n144_), .B(mai_mai_n140_), .Y(mai_mai_n177_));
  NA2        m161(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n178_));
  NA2        m162(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n179_));
  NA3        m163(.A(mai_mai_n179_), .B(mai_mai_n178_), .C(mai_mai_n24_), .Y(mai_mai_n180_));
  AN2        m164(.A(mai_mai_n180_), .B(mai_mai_n145_), .Y(mai_mai_n181_));
  NA2        m165(.A(x8), .B(x0), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n159_), .B(mai_mai_n25_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n127_), .B(x4), .Y(mai_mai_n184_));
  NA2        m168(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  AOI210     m169(.A0(mai_mai_n182_), .A1(mai_mai_n134_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NA2        m170(.A(x2), .B(x0), .Y(mai_mai_n187_));
  NA2        m171(.A(x4), .B(x1), .Y(mai_mai_n188_));
  NAi21      m172(.An(mai_mai_n125_), .B(mai_mai_n188_), .Y(mai_mai_n189_));
  NOi31      m173(.An(mai_mai_n189_), .B(mai_mai_n162_), .C(mai_mai_n187_), .Y(mai_mai_n190_));
  NO4        m174(.A(mai_mai_n190_), .B(mai_mai_n186_), .C(mai_mai_n181_), .D(mai_mai_n177_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n191_), .B(mai_mai_n41_), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n180_), .B(mai_mai_n75_), .Y(mai_mai_n193_));
  INV        m177(.A(mai_mai_n133_), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n108_), .B(mai_mai_n17_), .Y(mai_mai_n195_));
  AOI210     m179(.A0(mai_mai_n34_), .A1(mai_mai_n93_), .B0(mai_mai_n195_), .Y(mai_mai_n196_));
  NO3        m180(.A(mai_mai_n196_), .B(mai_mai_n194_), .C(x7), .Y(mai_mai_n197_));
  NA3        m181(.A(mai_mai_n189_), .B(mai_mai_n194_), .C(mai_mai_n40_), .Y(mai_mai_n198_));
  OAI210     m182(.A0(mai_mai_n179_), .A1(mai_mai_n140_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  NO3        m183(.A(mai_mai_n199_), .B(mai_mai_n197_), .C(mai_mai_n193_), .Y(mai_mai_n200_));
  NO2        m184(.A(mai_mai_n200_), .B(x3), .Y(mai_mai_n201_));
  NO3        m185(.A(mai_mai_n201_), .B(mai_mai_n192_), .C(mai_mai_n176_), .Y(mai03));
  NO2        m186(.A(mai_mai_n46_), .B(x3), .Y(mai_mai_n203_));
  NO2        m187(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n204_));
  INV        m188(.A(mai_mai_n204_), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n206_));
  OAI210     m190(.A0(mai_mai_n206_), .A1(mai_mai_n25_), .B0(mai_mai_n61_), .Y(mai_mai_n207_));
  OAI220     m191(.A0(mai_mai_n207_), .A1(mai_mai_n17_), .B0(mai_mai_n205_), .B1(mai_mai_n108_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n203_), .Y(mai_mai_n209_));
  NO2        m193(.A(mai_mai_n77_), .B(x6), .Y(mai_mai_n210_));
  NA2        m194(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n211_));
  NO2        m195(.A(mai_mai_n211_), .B(x4), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n213_));
  AO220      m197(.A0(mai_mai_n213_), .A1(mai_mai_n212_), .B0(mai_mai_n210_), .B1(mai_mai_n53_), .Y(mai_mai_n214_));
  NA2        m198(.A(mai_mai_n214_), .B(mai_mai_n60_), .Y(mai_mai_n215_));
  NA2        m199(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n216_));
  NA2        m200(.A(mai_mai_n211_), .B(mai_mai_n80_), .Y(mai_mai_n217_));
  AOI210     m201(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n187_), .Y(mai_mai_n218_));
  NA2        m202(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n219_));
  NO2        m203(.A(x5), .B(x1), .Y(mai_mai_n220_));
  AOI220     m204(.A0(mai_mai_n220_), .A1(mai_mai_n17_), .B0(mai_mai_n105_), .B1(x5), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n216_), .B(mai_mai_n178_), .Y(mai_mai_n222_));
  NO3        m206(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n223_));
  NO2        m207(.A(mai_mai_n223_), .B(mai_mai_n222_), .Y(mai_mai_n224_));
  OAI210     m208(.A0(mai_mai_n221_), .A1(mai_mai_n62_), .B0(mai_mai_n224_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n225_), .B(mai_mai_n46_), .Y(mai_mai_n226_));
  NA4        m210(.A(mai_mai_n226_), .B(mai_mai_n219_), .C(mai_mai_n215_), .D(mai_mai_n209_), .Y(mai_mai_n227_));
  NO2        m211(.A(mai_mai_n46_), .B(mai_mai_n41_), .Y(mai_mai_n228_));
  NA2        m212(.A(mai_mai_n228_), .B(mai_mai_n19_), .Y(mai_mai_n229_));
  NO2        m213(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n230_));
  NO2        m214(.A(mai_mai_n230_), .B(x6), .Y(mai_mai_n231_));
  NOi21      m215(.An(mai_mai_n83_), .B(mai_mai_n231_), .Y(mai_mai_n232_));
  NA2        m216(.A(mai_mai_n60_), .B(mai_mai_n93_), .Y(mai_mai_n233_));
  NA3        m217(.A(mai_mai_n233_), .B(mai_mai_n230_), .C(x6), .Y(mai_mai_n234_));
  AOI210     m218(.A0(mai_mai_n234_), .A1(mai_mai_n232_), .B0(mai_mai_n159_), .Y(mai_mai_n235_));
  AO210      m219(.A0(mai_mai_n235_), .A1(mai_mai_n229_), .B0(mai_mai_n183_), .Y(mai_mai_n236_));
  NA2        m220(.A(mai_mai_n41_), .B(mai_mai_n52_), .Y(mai_mai_n237_));
  OAI210     m221(.A0(mai_mai_n237_), .A1(mai_mai_n25_), .B0(mai_mai_n179_), .Y(mai_mai_n238_));
  NO3        m222(.A(mai_mai_n188_), .B(mai_mai_n60_), .C(x6), .Y(mai_mai_n239_));
  AOI220     m223(.A0(mai_mai_n239_), .A1(mai_mai_n238_), .B0(mai_mai_n145_), .B1(mai_mai_n92_), .Y(mai_mai_n240_));
  NA2        m224(.A(x6), .B(mai_mai_n46_), .Y(mai_mai_n241_));
  OAI210     m225(.A0(mai_mai_n121_), .A1(mai_mai_n78_), .B0(x4), .Y(mai_mai_n242_));
  AOI210     m226(.A0(mai_mai_n242_), .A1(mai_mai_n241_), .B0(mai_mai_n77_), .Y(mai_mai_n243_));
  NA2        m227(.A(mai_mai_n204_), .B(mai_mai_n138_), .Y(mai_mai_n244_));
  NA3        m228(.A(mai_mai_n216_), .B(mai_mai_n133_), .C(x6), .Y(mai_mai_n245_));
  OAI210     m229(.A0(mai_mai_n93_), .A1(mai_mai_n35_), .B0(mai_mai_n65_), .Y(mai_mai_n246_));
  NA3        m230(.A(mai_mai_n246_), .B(mai_mai_n245_), .C(mai_mai_n244_), .Y(mai_mai_n247_));
  OAI210     m231(.A0(mai_mai_n247_), .A1(mai_mai_n243_), .B0(x2), .Y(mai_mai_n248_));
  NA3        m232(.A(mai_mai_n248_), .B(mai_mai_n240_), .C(mai_mai_n236_), .Y(mai_mai_n249_));
  AOI210     m233(.A0(mai_mai_n227_), .A1(x8), .B0(mai_mai_n249_), .Y(mai_mai_n250_));
  NO2        m234(.A(mai_mai_n93_), .B(x3), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n251_), .B(mai_mai_n212_), .Y(mai_mai_n252_));
  NO2        m236(.A(mai_mai_n91_), .B(mai_mai_n25_), .Y(mai_mai_n253_));
  AOI210     m237(.A0(mai_mai_n231_), .A1(mai_mai_n162_), .B0(mai_mai_n253_), .Y(mai_mai_n254_));
  AOI210     m238(.A0(mai_mai_n254_), .A1(mai_mai_n252_), .B0(x2), .Y(mai_mai_n255_));
  NO2        m239(.A(x4), .B(mai_mai_n52_), .Y(mai_mai_n256_));
  AOI220     m240(.A0(mai_mai_n212_), .A1(mai_mai_n195_), .B0(mai_mai_n256_), .B1(mai_mai_n65_), .Y(mai_mai_n257_));
  NA2        m241(.A(mai_mai_n60_), .B(x6), .Y(mai_mai_n258_));
  NA3        m242(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n259_));
  AOI210     m243(.A0(mai_mai_n259_), .A1(mai_mai_n144_), .B0(mai_mai_n258_), .Y(mai_mai_n260_));
  NA2        m244(.A(mai_mai_n41_), .B(mai_mai_n17_), .Y(mai_mai_n261_));
  NO2        m245(.A(mai_mai_n261_), .B(mai_mai_n25_), .Y(mai_mai_n262_));
  OAI210     m246(.A0(mai_mai_n262_), .A1(mai_mai_n260_), .B0(mai_mai_n125_), .Y(mai_mai_n263_));
  NA2        m247(.A(mai_mai_n216_), .B(x6), .Y(mai_mai_n264_));
  NO2        m248(.A(mai_mai_n216_), .B(x6), .Y(mai_mai_n265_));
  NAi21      m249(.An(mai_mai_n170_), .B(mai_mai_n265_), .Y(mai_mai_n266_));
  NA3        m250(.A(mai_mai_n266_), .B(mai_mai_n264_), .C(mai_mai_n150_), .Y(mai_mai_n267_));
  NA4        m251(.A(mai_mai_n267_), .B(mai_mai_n263_), .C(mai_mai_n257_), .D(mai_mai_n159_), .Y(mai_mai_n268_));
  NA2        m252(.A(mai_mai_n204_), .B(mai_mai_n230_), .Y(mai_mai_n269_));
  NO2        m253(.A(x9), .B(x6), .Y(mai_mai_n270_));
  NO2        m254(.A(mai_mai_n144_), .B(mai_mai_n18_), .Y(mai_mai_n271_));
  NAi21      m255(.An(mai_mai_n271_), .B(mai_mai_n259_), .Y(mai_mai_n272_));
  NAi21      m256(.An(x1), .B(x4), .Y(mai_mai_n273_));
  AOI210     m257(.A0(x3), .A1(x2), .B0(mai_mai_n46_), .Y(mai_mai_n274_));
  OAI210     m258(.A0(mai_mai_n144_), .A1(x3), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  AOI220     m259(.A0(mai_mai_n275_), .A1(mai_mai_n273_), .B0(mai_mai_n272_), .B1(mai_mai_n270_), .Y(mai_mai_n276_));
  NA2        m260(.A(mai_mai_n276_), .B(mai_mai_n269_), .Y(mai_mai_n277_));
  NA2        m261(.A(mai_mai_n60_), .B(x2), .Y(mai_mai_n278_));
  NO2        m262(.A(mai_mai_n278_), .B(mai_mai_n269_), .Y(mai_mai_n279_));
  NO3        m263(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n280_));
  NA2        m264(.A(mai_mai_n108_), .B(mai_mai_n25_), .Y(mai_mai_n281_));
  NA2        m265(.A(x6), .B(x2), .Y(mai_mai_n282_));
  NO2        m266(.A(mai_mai_n282_), .B(mai_mai_n178_), .Y(mai_mai_n283_));
  AOI210     m267(.A0(mai_mai_n281_), .A1(mai_mai_n280_), .B0(mai_mai_n283_), .Y(mai_mai_n284_));
  OAI220     m268(.A0(mai_mai_n284_), .A1(mai_mai_n41_), .B0(mai_mai_n184_), .B1(mai_mai_n44_), .Y(mai_mai_n285_));
  OAI210     m269(.A0(mai_mai_n285_), .A1(mai_mai_n279_), .B0(mai_mai_n277_), .Y(mai_mai_n286_));
  NA2        m270(.A(x9), .B(mai_mai_n41_), .Y(mai_mai_n287_));
  NO2        m271(.A(mai_mai_n287_), .B(mai_mai_n211_), .Y(mai_mai_n288_));
  OR3        m272(.A(mai_mai_n288_), .B(mai_mai_n210_), .C(mai_mai_n154_), .Y(mai_mai_n289_));
  NA2        m273(.A(x4), .B(x0), .Y(mai_mai_n290_));
  NO3        m274(.A(mai_mai_n72_), .B(mai_mai_n290_), .C(x6), .Y(mai_mai_n291_));
  AOI210     m275(.A0(mai_mai_n289_), .A1(mai_mai_n40_), .B0(mai_mai_n291_), .Y(mai_mai_n292_));
  AOI210     m276(.A0(mai_mai_n292_), .A1(mai_mai_n286_), .B0(x8), .Y(mai_mai_n293_));
  INV        m277(.A(mai_mai_n258_), .Y(mai_mai_n294_));
  OAI210     m278(.A0(mai_mai_n271_), .A1(mai_mai_n220_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  INV        m279(.A(mai_mai_n182_), .Y(mai_mai_n296_));
  OAI210     m280(.A0(mai_mai_n296_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n297_), .A1(mai_mai_n295_), .B0(mai_mai_n237_), .Y(mai_mai_n298_));
  NO4        m282(.A(mai_mai_n298_), .B(mai_mai_n293_), .C(mai_mai_n268_), .D(mai_mai_n255_), .Y(mai_mai_n299_));
  NO2        m283(.A(mai_mai_n170_), .B(x1), .Y(mai_mai_n300_));
  NO3        m284(.A(mai_mai_n300_), .B(x3), .C(mai_mai_n35_), .Y(mai_mai_n301_));
  OAI210     m285(.A0(mai_mai_n301_), .A1(mai_mai_n265_), .B0(x2), .Y(mai_mai_n302_));
  OAI210     m286(.A0(mai_mai_n296_), .A1(x6), .B0(mai_mai_n42_), .Y(mai_mai_n303_));
  AOI210     m287(.A0(mai_mai_n303_), .A1(mai_mai_n302_), .B0(mai_mai_n194_), .Y(mai_mai_n304_));
  NOi21      m288(.An(mai_mai_n282_), .B(mai_mai_n17_), .Y(mai_mai_n305_));
  NA3        m289(.A(mai_mai_n305_), .B(mai_mai_n220_), .C(mai_mai_n38_), .Y(mai_mai_n306_));
  AOI210     m290(.A0(mai_mai_n35_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n307_));
  NA3        m291(.A(mai_mai_n307_), .B(mai_mai_n168_), .C(mai_mai_n31_), .Y(mai_mai_n308_));
  NA2        m292(.A(x3), .B(x2), .Y(mai_mai_n309_));
  AOI220     m293(.A0(mai_mai_n309_), .A1(mai_mai_n237_), .B0(mai_mai_n308_), .B1(mai_mai_n306_), .Y(mai_mai_n310_));
  NAi21      m294(.An(x4), .B(x0), .Y(mai_mai_n311_));
  NO3        m295(.A(mai_mai_n311_), .B(mai_mai_n42_), .C(x2), .Y(mai_mai_n312_));
  OAI210     m296(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n312_), .Y(mai_mai_n313_));
  OAI220     m297(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n314_));
  NO2        m298(.A(x9), .B(x8), .Y(mai_mai_n315_));
  NA3        m299(.A(mai_mai_n315_), .B(mai_mai_n35_), .C(mai_mai_n52_), .Y(mai_mai_n316_));
  OAI210     m300(.A0(mai_mai_n307_), .A1(mai_mai_n305_), .B0(mai_mai_n316_), .Y(mai_mai_n317_));
  AOI220     m301(.A0(mai_mai_n317_), .A1(mai_mai_n81_), .B0(mai_mai_n314_), .B1(mai_mai_n30_), .Y(mai_mai_n318_));
  AOI210     m302(.A0(mai_mai_n318_), .A1(mai_mai_n313_), .B0(mai_mai_n25_), .Y(mai_mai_n319_));
  NA3        m303(.A(mai_mai_n35_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n320_));
  OAI210     m304(.A0(mai_mai_n307_), .A1(mai_mai_n305_), .B0(mai_mai_n320_), .Y(mai_mai_n321_));
  INV        m305(.A(mai_mai_n222_), .Y(mai_mai_n322_));
  NA2        m306(.A(mai_mai_n35_), .B(mai_mai_n41_), .Y(mai_mai_n323_));
  OR2        m307(.A(mai_mai_n323_), .B(mai_mai_n290_), .Y(mai_mai_n324_));
  OAI220     m308(.A0(mai_mai_n324_), .A1(mai_mai_n167_), .B0(mai_mai_n241_), .B1(mai_mai_n322_), .Y(mai_mai_n325_));
  AO210      m309(.A0(mai_mai_n321_), .A1(mai_mai_n154_), .B0(mai_mai_n325_), .Y(mai_mai_n326_));
  NO4        m310(.A(mai_mai_n326_), .B(mai_mai_n319_), .C(mai_mai_n310_), .D(mai_mai_n304_), .Y(mai_mai_n327_));
  OAI210     m311(.A0(mai_mai_n299_), .A1(mai_mai_n250_), .B0(mai_mai_n327_), .Y(mai04));
  OAI210     m312(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n329_));
  NA3        m313(.A(mai_mai_n329_), .B(mai_mai_n280_), .C(mai_mai_n84_), .Y(mai_mai_n330_));
  NO2        m314(.A(x2), .B(x1), .Y(mai_mai_n331_));
  OAI210     m315(.A0(mai_mai_n261_), .A1(mai_mai_n331_), .B0(mai_mai_n35_), .Y(mai_mai_n332_));
  NO2        m316(.A(mai_mai_n331_), .B(mai_mai_n311_), .Y(mai_mai_n333_));
  AOI210     m317(.A0(mai_mai_n60_), .A1(x4), .B0(mai_mai_n114_), .Y(mai_mai_n334_));
  OAI210     m318(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n251_), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n278_), .B(mai_mai_n91_), .Y(mai_mai_n336_));
  NO2        m320(.A(mai_mai_n336_), .B(mai_mai_n35_), .Y(mai_mai_n337_));
  NO2        m321(.A(mai_mai_n309_), .B(mai_mai_n213_), .Y(mai_mai_n338_));
  NA2        m322(.A(mai_mai_n338_), .B(mai_mai_n93_), .Y(mai_mai_n339_));
  NA3        m323(.A(mai_mai_n339_), .B(mai_mai_n337_), .C(mai_mai_n335_), .Y(mai_mai_n340_));
  NA2        m324(.A(mai_mai_n340_), .B(mai_mai_n332_), .Y(mai_mai_n341_));
  NO3        m325(.A(mai_mai_n258_), .B(mai_mai_n122_), .C(mai_mai_n18_), .Y(mai_mai_n342_));
  INV        m326(.A(mai_mai_n342_), .Y(mai_mai_n343_));
  OAI210     m327(.A0(mai_mai_n120_), .A1(mai_mai_n108_), .B0(mai_mai_n182_), .Y(mai_mai_n344_));
  NA3        m328(.A(mai_mai_n344_), .B(x6), .C(x3), .Y(mai_mai_n345_));
  AOI210     m329(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n346_));
  OAI220     m330(.A0(mai_mai_n346_), .A1(mai_mai_n323_), .B0(mai_mai_n278_), .B1(mai_mai_n320_), .Y(mai_mai_n347_));
  INV        m331(.A(mai_mai_n347_), .Y(mai_mai_n348_));
  NA2        m332(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n349_));
  OAI210     m333(.A0(mai_mai_n108_), .A1(mai_mai_n17_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  AOI220     m334(.A0(mai_mai_n350_), .A1(mai_mai_n78_), .B0(mai_mai_n336_), .B1(mai_mai_n93_), .Y(mai_mai_n351_));
  NA4        m335(.A(mai_mai_n351_), .B(mai_mai_n348_), .C(mai_mai_n345_), .D(mai_mai_n343_), .Y(mai_mai_n352_));
  OAI210     m336(.A0(mai_mai_n113_), .A1(x3), .B0(mai_mai_n312_), .Y(mai_mai_n353_));
  NA2        m337(.A(mai_mai_n353_), .B(mai_mai_n159_), .Y(mai_mai_n354_));
  AOI210     m338(.A0(mai_mai_n352_), .A1(x4), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NA2        m339(.A(mai_mai_n333_), .B(mai_mai_n93_), .Y(mai_mai_n356_));
  NOi21      m340(.An(x4), .B(x0), .Y(mai_mai_n357_));
  XO2        m341(.A(x4), .B(x0), .Y(mai_mai_n358_));
  OAI210     m342(.A0(mai_mai_n358_), .A1(mai_mai_n119_), .B0(mai_mai_n273_), .Y(mai_mai_n359_));
  AOI220     m343(.A0(mai_mai_n359_), .A1(x8), .B0(mai_mai_n357_), .B1(mai_mai_n94_), .Y(mai_mai_n360_));
  AOI210     m344(.A0(mai_mai_n360_), .A1(mai_mai_n356_), .B0(x3), .Y(mai_mai_n361_));
  INV        m345(.A(mai_mai_n94_), .Y(mai_mai_n362_));
  NO2        m346(.A(mai_mai_n93_), .B(x4), .Y(mai_mai_n363_));
  AOI220     m347(.A0(mai_mai_n363_), .A1(mai_mai_n42_), .B0(mai_mai_n129_), .B1(mai_mai_n362_), .Y(mai_mai_n364_));
  NO3        m348(.A(mai_mai_n358_), .B(mai_mai_n170_), .C(x2), .Y(mai_mai_n365_));
  NO3        m349(.A(mai_mai_n233_), .B(mai_mai_n28_), .C(mai_mai_n24_), .Y(mai_mai_n366_));
  NO2        m350(.A(mai_mai_n366_), .B(mai_mai_n365_), .Y(mai_mai_n367_));
  NA4        m351(.A(mai_mai_n367_), .B(mai_mai_n364_), .C(mai_mai_n229_), .D(x6), .Y(mai_mai_n368_));
  OAI220     m352(.A0(mai_mai_n311_), .A1(mai_mai_n91_), .B0(mai_mai_n187_), .B1(mai_mai_n93_), .Y(mai_mai_n369_));
  NO2        m353(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n370_));
  OR2        m354(.A(mai_mai_n363_), .B(mai_mai_n370_), .Y(mai_mai_n371_));
  NO2        m355(.A(mai_mai_n156_), .B(mai_mai_n108_), .Y(mai_mai_n372_));
  AOI220     m356(.A0(mai_mai_n372_), .A1(mai_mai_n371_), .B0(mai_mai_n369_), .B1(mai_mai_n59_), .Y(mai_mai_n373_));
  NO2        m357(.A(mai_mai_n156_), .B(mai_mai_n80_), .Y(mai_mai_n374_));
  NO2        m358(.A(mai_mai_n34_), .B(x2), .Y(mai_mai_n375_));
  NOi21      m359(.An(mai_mai_n125_), .B(mai_mai_n27_), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n375_), .A1(mai_mai_n374_), .B0(mai_mai_n376_), .Y(mai_mai_n377_));
  OAI210     m361(.A0(mai_mai_n373_), .A1(mai_mai_n60_), .B0(mai_mai_n377_), .Y(mai_mai_n378_));
  OAI220     m362(.A0(mai_mai_n378_), .A1(x6), .B0(mai_mai_n368_), .B1(mai_mai_n361_), .Y(mai_mai_n379_));
  NA2        m363(.A(mai_mai_n46_), .B(mai_mai_n40_), .Y(mai_mai_n380_));
  OAI210     m364(.A0(mai_mai_n380_), .A1(mai_mai_n93_), .B0(mai_mai_n324_), .Y(mai_mai_n381_));
  AOI210     m365(.A0(mai_mai_n381_), .A1(mai_mai_n18_), .B0(mai_mai_n159_), .Y(mai_mai_n382_));
  AO220      m366(.A0(mai_mai_n382_), .A1(mai_mai_n379_), .B0(mai_mai_n355_), .B1(mai_mai_n341_), .Y(mai_mai_n383_));
  NA2        m367(.A(mai_mai_n375_), .B(x6), .Y(mai_mai_n384_));
  AOI210     m368(.A0(x6), .A1(x1), .B0(mai_mai_n158_), .Y(mai_mai_n385_));
  NA2        m369(.A(mai_mai_n363_), .B(x0), .Y(mai_mai_n386_));
  NA2        m370(.A(mai_mai_n83_), .B(x6), .Y(mai_mai_n387_));
  OAI210     m371(.A0(mai_mai_n386_), .A1(mai_mai_n385_), .B0(mai_mai_n387_), .Y(mai_mai_n388_));
  AOI220     m372(.A0(mai_mai_n388_), .A1(mai_mai_n384_), .B0(mai_mai_n223_), .B1(mai_mai_n47_), .Y(mai_mai_n389_));
  NA3        m373(.A(mai_mai_n389_), .B(mai_mai_n383_), .C(mai_mai_n330_), .Y(mai_mai_n390_));
  AOI210     m374(.A0(mai_mai_n206_), .A1(x8), .B0(mai_mai_n113_), .Y(mai_mai_n391_));
  NA2        m375(.A(mai_mai_n391_), .B(mai_mai_n349_), .Y(mai_mai_n392_));
  NA3        m376(.A(mai_mai_n392_), .B(mai_mai_n203_), .C(mai_mai_n159_), .Y(mai_mai_n393_));
  OAI210     m377(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n237_), .Y(mai_mai_n394_));
  AO220      m378(.A0(mai_mai_n394_), .A1(mai_mai_n155_), .B0(mai_mai_n112_), .B1(x4), .Y(mai_mai_n395_));
  NA3        m379(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n396_));
  NO2        m380(.A(mai_mai_n396_), .B(mai_mai_n362_), .Y(mai_mai_n397_));
  AOI210     m381(.A0(mai_mai_n395_), .A1(mai_mai_n121_), .B0(mai_mai_n397_), .Y(mai_mai_n398_));
  AOI210     m382(.A0(mai_mai_n398_), .A1(mai_mai_n393_), .B0(mai_mai_n25_), .Y(mai_mai_n399_));
  NA3        m383(.A(mai_mai_n123_), .B(mai_mai_n228_), .C(x0), .Y(mai_mai_n400_));
  OAI210     m384(.A0(mai_mai_n203_), .A1(mai_mai_n66_), .B0(mai_mai_n213_), .Y(mai_mai_n401_));
  NA3        m385(.A(mai_mai_n206_), .B(mai_mai_n230_), .C(x8), .Y(mai_mai_n402_));
  AOI210     m386(.A0(mai_mai_n402_), .A1(mai_mai_n401_), .B0(mai_mai_n25_), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n122_), .A1(mai_mai_n120_), .B0(mai_mai_n40_), .Y(mai_mai_n404_));
  NOi31      m388(.An(mai_mai_n404_), .B(mai_mai_n370_), .C(mai_mai_n188_), .Y(mai_mai_n405_));
  OAI210     m389(.A0(mai_mai_n405_), .A1(mai_mai_n403_), .B0(mai_mai_n155_), .Y(mai_mai_n406_));
  NAi31      m390(.An(mai_mai_n48_), .B(mai_mai_n300_), .C(mai_mai_n183_), .Y(mai_mai_n407_));
  NA3        m391(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(mai_mai_n400_), .Y(mai_mai_n408_));
  OAI210     m392(.A0(mai_mai_n408_), .A1(mai_mai_n399_), .B0(x6), .Y(mai_mai_n409_));
  OAI210     m393(.A0(mai_mai_n170_), .A1(mai_mai_n46_), .B0(mai_mai_n139_), .Y(mai_mai_n410_));
  NA3        m394(.A(mai_mai_n53_), .B(mai_mai_n37_), .C(mai_mai_n30_), .Y(mai_mai_n411_));
  AOI220     m395(.A0(mai_mai_n411_), .A1(mai_mai_n410_), .B0(mai_mai_n38_), .B1(mai_mai_n31_), .Y(mai_mai_n412_));
  NO2        m396(.A(mai_mai_n159_), .B(x0), .Y(mai_mai_n413_));
  AOI220     m397(.A0(mai_mai_n413_), .A1(mai_mai_n228_), .B0(mai_mai_n203_), .B1(mai_mai_n159_), .Y(mai_mai_n414_));
  AOI210     m398(.A0(mai_mai_n131_), .A1(mai_mai_n256_), .B0(x1), .Y(mai_mai_n415_));
  OAI210     m399(.A0(mai_mai_n414_), .A1(x8), .B0(mai_mai_n415_), .Y(mai_mai_n416_));
  INV        m400(.A(mai_mai_n171_), .Y(mai_mai_n417_));
  NA3        m401(.A(mai_mai_n417_), .B(mai_mai_n153_), .C(x9), .Y(mai_mai_n418_));
  NO4        m402(.A(mai_mai_n130_), .B(mai_mai_n311_), .C(x9), .D(x2), .Y(mai_mai_n419_));
  NOi21      m403(.An(mai_mai_n128_), .B(mai_mai_n187_), .Y(mai_mai_n420_));
  NO3        m404(.A(mai_mai_n420_), .B(mai_mai_n419_), .C(mai_mai_n18_), .Y(mai_mai_n421_));
  NO3        m405(.A(x9), .B(mai_mai_n159_), .C(x0), .Y(mai_mai_n422_));
  AOI220     m406(.A0(mai_mai_n422_), .A1(mai_mai_n251_), .B0(mai_mai_n374_), .B1(mai_mai_n159_), .Y(mai_mai_n423_));
  NA4        m407(.A(mai_mai_n423_), .B(mai_mai_n421_), .C(mai_mai_n418_), .D(mai_mai_n48_), .Y(mai_mai_n424_));
  OAI210     m408(.A0(mai_mai_n416_), .A1(mai_mai_n412_), .B0(mai_mai_n424_), .Y(mai_mai_n425_));
  NOi31      m409(.An(mai_mai_n413_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n426_));
  AOI210     m410(.A0(mai_mai_n37_), .A1(x9), .B0(mai_mai_n137_), .Y(mai_mai_n427_));
  NO3        m411(.A(mai_mai_n427_), .B(mai_mai_n128_), .C(mai_mai_n41_), .Y(mai_mai_n428_));
  NOi31      m412(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n429_));
  AOI220     m413(.A0(mai_mai_n429_), .A1(mai_mai_n357_), .B0(mai_mai_n129_), .B1(x3), .Y(mai_mai_n430_));
  AOI210     m414(.A0(mai_mai_n273_), .A1(mai_mai_n58_), .B0(mai_mai_n127_), .Y(mai_mai_n431_));
  OAI210     m415(.A0(mai_mai_n431_), .A1(x3), .B0(mai_mai_n430_), .Y(mai_mai_n432_));
  NO3        m416(.A(mai_mai_n432_), .B(mai_mai_n428_), .C(x2), .Y(mai_mai_n433_));
  OAI220     m417(.A0(mai_mai_n358_), .A1(mai_mai_n315_), .B0(mai_mai_n311_), .B1(mai_mai_n41_), .Y(mai_mai_n434_));
  INV        m418(.A(mai_mai_n396_), .Y(mai_mai_n435_));
  AOI220     m419(.A0(mai_mai_n435_), .A1(mai_mai_n93_), .B0(mai_mai_n434_), .B1(mai_mai_n159_), .Y(mai_mai_n436_));
  NO2        m420(.A(mai_mai_n436_), .B(mai_mai_n52_), .Y(mai_mai_n437_));
  NO3        m421(.A(mai_mai_n437_), .B(mai_mai_n433_), .C(mai_mai_n426_), .Y(mai_mai_n438_));
  AOI210     m422(.A0(mai_mai_n438_), .A1(mai_mai_n425_), .B0(mai_mai_n25_), .Y(mai_mai_n439_));
  NA4        m423(.A(mai_mai_n30_), .B(mai_mai_n93_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n440_));
  NO3        m424(.A(mai_mai_n66_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n441_));
  NA2        m425(.A(mai_mai_n441_), .B(mai_mai_n274_), .Y(mai_mai_n442_));
  NO2        m426(.A(mai_mai_n442_), .B(mai_mai_n105_), .Y(mai_mai_n443_));
  NO3        m427(.A(mai_mai_n278_), .B(mai_mai_n182_), .C(mai_mai_n38_), .Y(mai_mai_n444_));
  OAI210     m428(.A0(mai_mai_n444_), .A1(mai_mai_n443_), .B0(x7), .Y(mai_mai_n445_));
  NA2        m429(.A(mai_mai_n233_), .B(x7), .Y(mai_mai_n446_));
  NA3        m430(.A(mai_mai_n446_), .B(mai_mai_n158_), .C(mai_mai_n138_), .Y(mai_mai_n447_));
  NA3        m431(.A(mai_mai_n447_), .B(mai_mai_n445_), .C(mai_mai_n440_), .Y(mai_mai_n448_));
  OAI210     m432(.A0(mai_mai_n448_), .A1(mai_mai_n439_), .B0(mai_mai_n35_), .Y(mai_mai_n449_));
  NO2        m433(.A(mai_mai_n422_), .B(mai_mai_n213_), .Y(mai_mai_n450_));
  NO4        m434(.A(mai_mai_n450_), .B(mai_mai_n77_), .C(x4), .D(mai_mai_n52_), .Y(mai_mai_n451_));
  AOI220     m435(.A0(mai_mai_n370_), .A1(mai_mai_n93_), .B0(mai_mai_n156_), .B1(mai_mai_n206_), .Y(mai_mai_n452_));
  NA2        m436(.A(mai_mai_n452_), .B(mai_mai_n91_), .Y(mai_mai_n453_));
  NA2        m437(.A(mai_mai_n453_), .B(mai_mai_n183_), .Y(mai_mai_n454_));
  OAI220     m438(.A0(mai_mai_n287_), .A1(mai_mai_n67_), .B0(mai_mai_n167_), .B1(mai_mai_n41_), .Y(mai_mai_n455_));
  NA2        m439(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n456_));
  AOI210     m440(.A0(mai_mai_n171_), .A1(mai_mai_n27_), .B0(mai_mai_n72_), .Y(mai_mai_n457_));
  OAI210     m441(.A0(mai_mai_n155_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n458_));
  NO3        m442(.A(mai_mai_n429_), .B(x3), .C(mai_mai_n52_), .Y(mai_mai_n459_));
  AOI210     m443(.A0(mai_mai_n459_), .A1(mai_mai_n458_), .B0(mai_mai_n457_), .Y(mai_mai_n460_));
  OAI210     m444(.A0(mai_mai_n160_), .A1(mai_mai_n456_), .B0(mai_mai_n460_), .Y(mai_mai_n461_));
  AOI220     m445(.A0(mai_mai_n461_), .A1(x0), .B0(mai_mai_n455_), .B1(mai_mai_n139_), .Y(mai_mai_n462_));
  AOI210     m446(.A0(mai_mai_n462_), .A1(mai_mai_n454_), .B0(mai_mai_n241_), .Y(mai_mai_n463_));
  NA2        m447(.A(x9), .B(x5), .Y(mai_mai_n464_));
  NO4        m448(.A(mai_mai_n108_), .B(mai_mai_n464_), .C(mai_mai_n58_), .D(mai_mai_n31_), .Y(mai_mai_n465_));
  NO3        m449(.A(mai_mai_n465_), .B(mai_mai_n463_), .C(mai_mai_n451_), .Y(mai_mai_n466_));
  NA3        m450(.A(mai_mai_n466_), .B(mai_mai_n449_), .C(mai_mai_n409_), .Y(mai_mai_n467_));
  AOI210     m451(.A0(mai_mai_n390_), .A1(mai_mai_n25_), .B0(mai_mai_n467_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  INV        u005(.A(men_men_n19_), .Y(men_men_n22_));
  NA2        u006(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n23_));
  INV        u007(.A(x5), .Y(men_men_n24_));
  NA2        u008(.A(x7), .B(x6), .Y(men_men_n25_));
  NA2        u009(.A(x8), .B(x3), .Y(men_men_n26_));
  NA2        u010(.A(x4), .B(x2), .Y(men_men_n27_));
  NO4        u011(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .D(men_men_n24_), .Y(men_men_n28_));
  NO2        u012(.A(men_men_n28_), .B(men_men_n23_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n22_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n24_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA3        u020(.A(men_men_n36_), .B(men_men_n35_), .C(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n22_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n35_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n50_), .B(men_men_n33_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n34_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO3        u046(.A(men_men_n62_), .B(men_men_n59_), .C(men_men_n58_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NO2        u051(.A(men_men_n67_), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n42_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n41_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n46_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO4        u062(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(x4), .B(x2), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(x3), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n80_), .B(men_men_n18_), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n85_));
  NO4        u069(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n86_));
  NA2        u070(.A(men_men_n60_), .B(men_men_n46_), .Y(men_men_n87_));
  INV        u071(.A(men_men_n87_), .Y(men_men_n88_));
  OAI210     u072(.A0(men_men_n86_), .A1(men_men_n65_), .B0(men_men_n88_), .Y(men_men_n89_));
  NA2        u073(.A(x3), .B(men_men_n18_), .Y(men_men_n90_));
  NO2        u074(.A(men_men_n90_), .B(men_men_n24_), .Y(men_men_n91_));
  INV        u075(.A(x8), .Y(men_men_n92_));
  NA2        u076(.A(x2), .B(x1), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n91_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n25_), .Y(men_men_n96_));
  AOI210     u080(.A0(men_men_n54_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n43_), .A1(men_men_n35_), .B0(men_men_n46_), .Y(men_men_n98_));
  NO3        u082(.A(men_men_n98_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n99_));
  NA2        u083(.A(x4), .B(men_men_n41_), .Y(men_men_n100_));
  NO2        u084(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n101_));
  OAI210     u085(.A0(men_men_n101_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n102_));
  AOI210     u086(.A0(men_men_n100_), .A1(men_men_n50_), .B0(men_men_n102_), .Y(men_men_n103_));
  NO2        u087(.A(x3), .B(x2), .Y(men_men_n104_));
  NA3        u088(.A(men_men_n104_), .B(men_men_n25_), .C(men_men_n24_), .Y(men_men_n105_));
  AOI210     u089(.A0(x8), .A1(x6), .B0(men_men_n105_), .Y(men_men_n106_));
  NA2        u090(.A(men_men_n52_), .B(x1), .Y(men_men_n107_));
  OAI210     u091(.A0(men_men_n107_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n108_));
  NO4        u092(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n103_), .D(men_men_n99_), .Y(men_men_n109_));
  AO220      u093(.A0(men_men_n109_), .A1(men_men_n89_), .B0(men_men_n85_), .B1(men_men_n74_), .Y(men02));
  NO2        u094(.A(x3), .B(men_men_n52_), .Y(men_men_n111_));
  NO2        u095(.A(x8), .B(men_men_n18_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n41_), .B(x0), .Y(men_men_n114_));
  OAI210     u098(.A0(men_men_n87_), .A1(men_men_n113_), .B0(men_men_n114_), .Y(men_men_n115_));
  AOI220     u099(.A0(men_men_n115_), .A1(men_men_n112_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n116_));
  NO3        u100(.A(men_men_n116_), .B(x7), .C(x5), .Y(men_men_n117_));
  NA2        u101(.A(x9), .B(x2), .Y(men_men_n118_));
  OR2        u102(.A(x8), .B(x0), .Y(men_men_n119_));
  INV        u103(.A(men_men_n119_), .Y(men_men_n120_));
  NAi21      u104(.An(x2), .B(x8), .Y(men_men_n121_));
  INV        u105(.A(men_men_n121_), .Y(men_men_n122_));
  OAI220     u106(.A0(men_men_n122_), .A1(men_men_n120_), .B0(men_men_n118_), .B1(x7), .Y(men_men_n123_));
  NO2        u107(.A(x4), .B(x1), .Y(men_men_n124_));
  NA3        u108(.A(men_men_n124_), .B(men_men_n123_), .C(men_men_n58_), .Y(men_men_n125_));
  NOi21      u109(.An(x0), .B(x1), .Y(men_men_n126_));
  NO3        u110(.A(x9), .B(x8), .C(x7), .Y(men_men_n127_));
  NOi21      u111(.An(x0), .B(x4), .Y(men_men_n128_));
  NAi21      u112(.An(x8), .B(x7), .Y(men_men_n129_));
  NO2        u113(.A(men_men_n129_), .B(men_men_n60_), .Y(men_men_n130_));
  AOI220     u114(.A0(men_men_n130_), .A1(men_men_n128_), .B0(men_men_n127_), .B1(men_men_n126_), .Y(men_men_n131_));
  AOI210     u115(.A0(men_men_n131_), .A1(men_men_n125_), .B0(men_men_n77_), .Y(men_men_n132_));
  NO2        u116(.A(x5), .B(men_men_n46_), .Y(men_men_n133_));
  NA2        u117(.A(x2), .B(men_men_n18_), .Y(men_men_n134_));
  AOI210     u118(.A0(men_men_n134_), .A1(men_men_n107_), .B0(men_men_n114_), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n135_), .A1(men_men_n33_), .B0(men_men_n133_), .Y(men_men_n136_));
  NAi21      u120(.An(x0), .B(x4), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x1), .Y(men_men_n138_));
  NO2        u122(.A(x7), .B(x0), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n82_), .B(men_men_n101_), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n140_), .B(x3), .Y(men_men_n141_));
  OAI210     u125(.A0(men_men_n139_), .A1(men_men_n138_), .B0(men_men_n141_), .Y(men_men_n142_));
  NA2        u126(.A(x5), .B(x0), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n46_), .B(x2), .Y(men_men_n144_));
  NA3        u128(.A(men_men_n142_), .B(men_men_n136_), .C(men_men_n34_), .Y(men_men_n145_));
  NO3        u129(.A(men_men_n145_), .B(men_men_n132_), .C(men_men_n117_), .Y(men_men_n146_));
  NO3        u130(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n23_), .Y(men_men_n147_));
  NO2        u131(.A(men_men_n27_), .B(men_men_n24_), .Y(men_men_n148_));
  AOI220     u132(.A0(men_men_n126_), .A1(men_men_n148_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n149_));
  NO3        u133(.A(men_men_n149_), .B(men_men_n58_), .C(men_men_n60_), .Y(men_men_n150_));
  NA2        u134(.A(x7), .B(x3), .Y(men_men_n151_));
  NO2        u135(.A(men_men_n100_), .B(x5), .Y(men_men_n152_));
  NO2        u136(.A(x9), .B(x7), .Y(men_men_n153_));
  NOi21      u137(.An(x8), .B(x0), .Y(men_men_n154_));
  NO2        u138(.A(men_men_n41_), .B(x2), .Y(men_men_n155_));
  INV        u139(.A(x7), .Y(men_men_n156_));
  NA2        u140(.A(men_men_n156_), .B(men_men_n18_), .Y(men_men_n157_));
  AOI220     u141(.A0(men_men_n157_), .A1(men_men_n155_), .B0(men_men_n111_), .B1(men_men_n36_), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n24_), .B(x4), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n159_), .B(men_men_n128_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n160_), .B(men_men_n158_), .Y(men_men_n161_));
  INV        u145(.A(men_men_n161_), .Y(men_men_n162_));
  OAI210     u146(.A0(men_men_n151_), .A1(men_men_n48_), .B0(men_men_n162_), .Y(men_men_n163_));
  NA2        u147(.A(x5), .B(x1), .Y(men_men_n164_));
  INV        u148(.A(men_men_n164_), .Y(men_men_n165_));
  AOI210     u149(.A0(men_men_n165_), .A1(men_men_n128_), .B0(men_men_n34_), .Y(men_men_n166_));
  NO2        u150(.A(men_men_n60_), .B(men_men_n92_), .Y(men_men_n167_));
  NAi21      u151(.An(x2), .B(x7), .Y(men_men_n168_));
  NO3        u152(.A(men_men_n168_), .B(men_men_n167_), .C(men_men_n46_), .Y(men_men_n169_));
  NA2        u153(.A(men_men_n169_), .B(men_men_n65_), .Y(men_men_n170_));
  NAi31      u154(.An(men_men_n77_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n171_));
  NA3        u155(.A(men_men_n171_), .B(men_men_n170_), .C(men_men_n166_), .Y(men_men_n172_));
  NO4        u156(.A(men_men_n172_), .B(men_men_n163_), .C(men_men_n150_), .D(men_men_n147_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n173_), .B(men_men_n146_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n143_), .B(men_men_n140_), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n176_));
  NA2        u160(.A(men_men_n24_), .B(men_men_n17_), .Y(men_men_n177_));
  NA3        u161(.A(men_men_n177_), .B(men_men_n176_), .C(men_men_n23_), .Y(men_men_n178_));
  AN2        u162(.A(men_men_n178_), .B(men_men_n144_), .Y(men_men_n179_));
  NA2        u163(.A(x8), .B(x0), .Y(men_men_n180_));
  NO2        u164(.A(men_men_n156_), .B(men_men_n24_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n126_), .B(x4), .Y(men_men_n182_));
  NA2        u166(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  AOI210     u167(.A0(men_men_n180_), .A1(men_men_n134_), .B0(men_men_n183_), .Y(men_men_n184_));
  NA2        u168(.A(x2), .B(x0), .Y(men_men_n185_));
  NA2        u169(.A(x4), .B(x1), .Y(men_men_n186_));
  NAi21      u170(.An(men_men_n124_), .B(men_men_n186_), .Y(men_men_n187_));
  NOi31      u171(.An(men_men_n187_), .B(men_men_n159_), .C(men_men_n185_), .Y(men_men_n188_));
  NO4        u172(.A(men_men_n188_), .B(men_men_n184_), .C(men_men_n179_), .D(men_men_n175_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n189_), .B(men_men_n41_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n178_), .B(men_men_n75_), .Y(men_men_n191_));
  INV        u175(.A(men_men_n133_), .Y(men_men_n192_));
  NO2        u176(.A(men_men_n107_), .B(men_men_n17_), .Y(men_men_n193_));
  AOI210     u177(.A0(men_men_n33_), .A1(men_men_n92_), .B0(men_men_n193_), .Y(men_men_n194_));
  NO3        u178(.A(men_men_n194_), .B(men_men_n192_), .C(x7), .Y(men_men_n195_));
  NA3        u179(.A(men_men_n187_), .B(men_men_n192_), .C(men_men_n40_), .Y(men_men_n196_));
  OAI210     u180(.A0(men_men_n177_), .A1(men_men_n140_), .B0(men_men_n196_), .Y(men_men_n197_));
  NO3        u181(.A(men_men_n197_), .B(men_men_n195_), .C(men_men_n191_), .Y(men_men_n198_));
  NO2        u182(.A(men_men_n198_), .B(x3), .Y(men_men_n199_));
  NO3        u183(.A(men_men_n199_), .B(men_men_n190_), .C(men_men_n174_), .Y(men03));
  NO2        u184(.A(men_men_n46_), .B(x3), .Y(men_men_n201_));
  NO2        u185(.A(x6), .B(men_men_n24_), .Y(men_men_n202_));
  INV        u186(.A(men_men_n202_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n52_), .B(x1), .Y(men_men_n204_));
  OAI210     u188(.A0(men_men_n204_), .A1(men_men_n24_), .B0(men_men_n61_), .Y(men_men_n205_));
  OAI220     u189(.A0(men_men_n205_), .A1(men_men_n17_), .B0(men_men_n203_), .B1(men_men_n107_), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n206_), .B(men_men_n201_), .Y(men_men_n207_));
  NA2        u191(.A(x6), .B(men_men_n24_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n208_), .B(x4), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n18_), .B(x0), .Y(men_men_n210_));
  NA2        u194(.A(x3), .B(men_men_n17_), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n211_), .B(men_men_n208_), .Y(men_men_n212_));
  NA2        u196(.A(x9), .B(men_men_n52_), .Y(men_men_n213_));
  NA2        u197(.A(men_men_n213_), .B(x4), .Y(men_men_n214_));
  NA2        u198(.A(men_men_n208_), .B(men_men_n80_), .Y(men_men_n215_));
  AOI210     u199(.A0(men_men_n24_), .A1(x3), .B0(men_men_n185_), .Y(men_men_n216_));
  AOI220     u200(.A0(men_men_n216_), .A1(men_men_n215_), .B0(men_men_n214_), .B1(men_men_n212_), .Y(men_men_n217_));
  NO3        u201(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n218_));
  NO2        u202(.A(x5), .B(x1), .Y(men_men_n219_));
  AOI220     u203(.A0(men_men_n219_), .A1(men_men_n17_), .B0(men_men_n104_), .B1(x5), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n211_), .B(men_men_n176_), .Y(men_men_n221_));
  NO3        u205(.A(x3), .B(x2), .C(x1), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n222_), .B(men_men_n221_), .Y(men_men_n223_));
  OAI210     u207(.A0(men_men_n220_), .A1(men_men_n62_), .B0(men_men_n223_), .Y(men_men_n224_));
  AOI220     u208(.A0(men_men_n224_), .A1(men_men_n46_), .B0(men_men_n218_), .B1(men_men_n133_), .Y(men_men_n225_));
  NA3        u209(.A(men_men_n225_), .B(men_men_n217_), .C(men_men_n207_), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n227_));
  NA2        u211(.A(men_men_n227_), .B(men_men_n19_), .Y(men_men_n228_));
  NO2        u212(.A(x3), .B(men_men_n17_), .Y(men_men_n229_));
  NO2        u213(.A(men_men_n229_), .B(x6), .Y(men_men_n230_));
  NOi21      u214(.An(men_men_n82_), .B(men_men_n230_), .Y(men_men_n231_));
  NA2        u215(.A(men_men_n60_), .B(men_men_n92_), .Y(men_men_n232_));
  NA3        u216(.A(men_men_n232_), .B(men_men_n229_), .C(x6), .Y(men_men_n233_));
  AOI210     u217(.A0(men_men_n233_), .A1(men_men_n231_), .B0(men_men_n156_), .Y(men_men_n234_));
  AO210      u218(.A0(men_men_n234_), .A1(men_men_n228_), .B0(men_men_n181_), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n236_));
  OAI210     u220(.A0(men_men_n236_), .A1(men_men_n24_), .B0(men_men_n177_), .Y(men_men_n237_));
  NO3        u221(.A(men_men_n186_), .B(men_men_n60_), .C(x6), .Y(men_men_n238_));
  AOI220     u222(.A0(men_men_n238_), .A1(men_men_n237_), .B0(men_men_n144_), .B1(men_men_n91_), .Y(men_men_n239_));
  NA2        u223(.A(x6), .B(men_men_n46_), .Y(men_men_n240_));
  OAI210     u224(.A0(men_men_n120_), .A1(men_men_n78_), .B0(x4), .Y(men_men_n241_));
  AOI210     u225(.A0(men_men_n241_), .A1(men_men_n240_), .B0(men_men_n77_), .Y(men_men_n242_));
  NO2        u226(.A(men_men_n60_), .B(x6), .Y(men_men_n243_));
  NO2        u227(.A(men_men_n164_), .B(men_men_n41_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n221_), .B0(men_men_n243_), .Y(men_men_n245_));
  NA2        u229(.A(men_men_n202_), .B(men_men_n138_), .Y(men_men_n246_));
  NA3        u230(.A(men_men_n211_), .B(men_men_n133_), .C(x6), .Y(men_men_n247_));
  OAI210     u231(.A0(men_men_n92_), .A1(men_men_n34_), .B0(men_men_n65_), .Y(men_men_n248_));
  NA4        u232(.A(men_men_n248_), .B(men_men_n247_), .C(men_men_n246_), .D(men_men_n245_), .Y(men_men_n249_));
  OAI210     u233(.A0(men_men_n249_), .A1(men_men_n242_), .B0(x2), .Y(men_men_n250_));
  NA3        u234(.A(men_men_n250_), .B(men_men_n239_), .C(men_men_n235_), .Y(men_men_n251_));
  AOI210     u235(.A0(men_men_n226_), .A1(x8), .B0(men_men_n251_), .Y(men_men_n252_));
  NO2        u236(.A(men_men_n92_), .B(x3), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n253_), .B(men_men_n209_), .Y(men_men_n254_));
  NO3        u238(.A(men_men_n90_), .B(men_men_n78_), .C(men_men_n24_), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n230_), .A1(men_men_n159_), .B0(men_men_n255_), .Y(men_men_n256_));
  AOI210     u240(.A0(men_men_n256_), .A1(men_men_n254_), .B0(x2), .Y(men_men_n257_));
  NO2        u241(.A(x4), .B(men_men_n52_), .Y(men_men_n258_));
  AOI220     u242(.A0(men_men_n209_), .A1(men_men_n193_), .B0(men_men_n258_), .B1(men_men_n65_), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n60_), .B(x6), .Y(men_men_n260_));
  NA3        u244(.A(men_men_n24_), .B(x3), .C(x2), .Y(men_men_n261_));
  AOI210     u245(.A0(men_men_n261_), .A1(men_men_n143_), .B0(men_men_n260_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n263_), .B(men_men_n24_), .Y(men_men_n264_));
  OAI210     u248(.A0(men_men_n264_), .A1(men_men_n262_), .B0(men_men_n124_), .Y(men_men_n265_));
  NA2        u249(.A(men_men_n211_), .B(x6), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n211_), .B(x6), .Y(men_men_n267_));
  NAi21      u251(.An(men_men_n167_), .B(men_men_n267_), .Y(men_men_n268_));
  NA3        u252(.A(men_men_n268_), .B(men_men_n266_), .C(men_men_n148_), .Y(men_men_n269_));
  NA4        u253(.A(men_men_n269_), .B(men_men_n265_), .C(men_men_n259_), .D(men_men_n156_), .Y(men_men_n270_));
  NA2        u254(.A(men_men_n202_), .B(men_men_n229_), .Y(men_men_n271_));
  NO2        u255(.A(x9), .B(x6), .Y(men_men_n272_));
  NO2        u256(.A(men_men_n143_), .B(men_men_n18_), .Y(men_men_n273_));
  NAi21      u257(.An(men_men_n273_), .B(men_men_n261_), .Y(men_men_n274_));
  NAi21      u258(.An(x1), .B(x4), .Y(men_men_n275_));
  AOI210     u259(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n276_));
  OAI210     u260(.A0(men_men_n143_), .A1(x3), .B0(men_men_n276_), .Y(men_men_n277_));
  AOI220     u261(.A0(men_men_n277_), .A1(men_men_n275_), .B0(men_men_n274_), .B1(men_men_n272_), .Y(men_men_n278_));
  NA2        u262(.A(men_men_n278_), .B(men_men_n271_), .Y(men_men_n279_));
  NA2        u263(.A(men_men_n60_), .B(x2), .Y(men_men_n280_));
  NO2        u264(.A(men_men_n280_), .B(men_men_n271_), .Y(men_men_n281_));
  NO3        u265(.A(x9), .B(x6), .C(x0), .Y(men_men_n282_));
  NA2        u266(.A(men_men_n107_), .B(men_men_n24_), .Y(men_men_n283_));
  NA2        u267(.A(x6), .B(x2), .Y(men_men_n284_));
  NO2        u268(.A(men_men_n284_), .B(men_men_n176_), .Y(men_men_n285_));
  AOI210     u269(.A0(men_men_n283_), .A1(men_men_n282_), .B0(men_men_n285_), .Y(men_men_n286_));
  OAI220     u270(.A0(men_men_n286_), .A1(men_men_n41_), .B0(men_men_n182_), .B1(men_men_n44_), .Y(men_men_n287_));
  OAI210     u271(.A0(men_men_n287_), .A1(men_men_n281_), .B0(men_men_n279_), .Y(men_men_n288_));
  NO2        u272(.A(x3), .B(men_men_n208_), .Y(men_men_n289_));
  NA2        u273(.A(x4), .B(x0), .Y(men_men_n290_));
  NO3        u274(.A(men_men_n72_), .B(men_men_n290_), .C(x6), .Y(men_men_n291_));
  AOI210     u275(.A0(men_men_n289_), .A1(men_men_n40_), .B0(men_men_n291_), .Y(men_men_n292_));
  AOI210     u276(.A0(men_men_n292_), .A1(men_men_n288_), .B0(x8), .Y(men_men_n293_));
  INV        u277(.A(men_men_n260_), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n273_), .A1(men_men_n219_), .B0(men_men_n294_), .Y(men_men_n295_));
  OAI210     u279(.A0(x0), .A1(x4), .B0(men_men_n20_), .Y(men_men_n296_));
  AOI210     u280(.A0(men_men_n296_), .A1(men_men_n295_), .B0(men_men_n236_), .Y(men_men_n297_));
  NO4        u281(.A(men_men_n297_), .B(men_men_n293_), .C(men_men_n270_), .D(men_men_n257_), .Y(men_men_n298_));
  NO2        u282(.A(men_men_n167_), .B(x1), .Y(men_men_n299_));
  NO3        u283(.A(men_men_n299_), .B(x3), .C(men_men_n34_), .Y(men_men_n300_));
  OAI210     u284(.A0(men_men_n300_), .A1(men_men_n267_), .B0(x2), .Y(men_men_n301_));
  OAI210     u285(.A0(x0), .A1(x6), .B0(men_men_n42_), .Y(men_men_n302_));
  AOI210     u286(.A0(men_men_n302_), .A1(men_men_n301_), .B0(men_men_n192_), .Y(men_men_n303_));
  NOi21      u287(.An(men_men_n284_), .B(men_men_n17_), .Y(men_men_n304_));
  NA3        u288(.A(men_men_n304_), .B(men_men_n219_), .C(men_men_n38_), .Y(men_men_n305_));
  AOI210     u289(.A0(men_men_n34_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n306_));
  NA3        u290(.A(men_men_n306_), .B(men_men_n165_), .C(men_men_n31_), .Y(men_men_n307_));
  NA2        u291(.A(x3), .B(x2), .Y(men_men_n308_));
  AOI220     u292(.A0(men_men_n308_), .A1(men_men_n236_), .B0(men_men_n307_), .B1(men_men_n305_), .Y(men_men_n309_));
  NAi21      u293(.An(x4), .B(x0), .Y(men_men_n310_));
  NO3        u294(.A(men_men_n310_), .B(men_men_n42_), .C(x2), .Y(men_men_n311_));
  OAI210     u295(.A0(x6), .A1(men_men_n18_), .B0(men_men_n311_), .Y(men_men_n312_));
  OAI220     u296(.A0(men_men_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n313_));
  NO2        u297(.A(x9), .B(x8), .Y(men_men_n314_));
  NA3        u298(.A(men_men_n314_), .B(men_men_n34_), .C(men_men_n52_), .Y(men_men_n315_));
  OAI210     u299(.A0(men_men_n306_), .A1(men_men_n304_), .B0(men_men_n315_), .Y(men_men_n316_));
  AOI220     u300(.A0(men_men_n316_), .A1(men_men_n81_), .B0(men_men_n313_), .B1(men_men_n30_), .Y(men_men_n317_));
  AOI210     u301(.A0(men_men_n317_), .A1(men_men_n312_), .B0(men_men_n24_), .Y(men_men_n318_));
  NA3        u302(.A(men_men_n34_), .B(x1), .C(men_men_n17_), .Y(men_men_n319_));
  OAI210     u303(.A0(men_men_n306_), .A1(men_men_n304_), .B0(men_men_n319_), .Y(men_men_n320_));
  INV        u304(.A(men_men_n221_), .Y(men_men_n321_));
  NA2        u305(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n322_));
  OR2        u306(.A(men_men_n322_), .B(men_men_n290_), .Y(men_men_n323_));
  OAI220     u307(.A0(men_men_n323_), .A1(men_men_n164_), .B0(men_men_n240_), .B1(men_men_n321_), .Y(men_men_n324_));
  AO210      u308(.A0(men_men_n320_), .A1(men_men_n152_), .B0(men_men_n324_), .Y(men_men_n325_));
  NO4        u309(.A(men_men_n325_), .B(men_men_n318_), .C(men_men_n309_), .D(men_men_n303_), .Y(men_men_n326_));
  OAI210     u310(.A0(men_men_n298_), .A1(men_men_n252_), .B0(men_men_n326_), .Y(men04));
  OAI210     u311(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n328_));
  NA3        u312(.A(men_men_n328_), .B(men_men_n282_), .C(men_men_n83_), .Y(men_men_n329_));
  NO2        u313(.A(x2), .B(x1), .Y(men_men_n330_));
  OAI210     u314(.A0(men_men_n263_), .A1(men_men_n330_), .B0(men_men_n34_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n330_), .B(men_men_n310_), .Y(men_men_n332_));
  AOI210     u316(.A0(men_men_n60_), .A1(x4), .B0(men_men_n113_), .Y(men_men_n333_));
  OAI210     u317(.A0(men_men_n333_), .A1(men_men_n332_), .B0(men_men_n253_), .Y(men_men_n334_));
  NO2        u318(.A(men_men_n280_), .B(men_men_n90_), .Y(men_men_n335_));
  NO2        u319(.A(men_men_n335_), .B(men_men_n34_), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n308_), .B(men_men_n210_), .Y(men_men_n337_));
  NA2        u321(.A(x9), .B(x0), .Y(men_men_n338_));
  AOI210     u322(.A0(men_men_n90_), .A1(men_men_n75_), .B0(men_men_n338_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n339_), .A1(men_men_n337_), .B0(men_men_n92_), .Y(men_men_n340_));
  NA3        u324(.A(men_men_n340_), .B(men_men_n336_), .C(men_men_n334_), .Y(men_men_n341_));
  NA2        u325(.A(men_men_n341_), .B(men_men_n331_), .Y(men_men_n342_));
  NO2        u326(.A(men_men_n213_), .B(men_men_n114_), .Y(men_men_n343_));
  INV        u327(.A(men_men_n343_), .Y(men_men_n344_));
  OAI210     u328(.A0(men_men_n119_), .A1(men_men_n107_), .B0(men_men_n180_), .Y(men_men_n345_));
  NA3        u329(.A(men_men_n345_), .B(x6), .C(x3), .Y(men_men_n346_));
  NOi21      u330(.An(men_men_n154_), .B(men_men_n134_), .Y(men_men_n347_));
  AOI210     u331(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n348_));
  OAI220     u332(.A0(men_men_n348_), .A1(men_men_n322_), .B0(men_men_n280_), .B1(men_men_n319_), .Y(men_men_n349_));
  AOI210     u333(.A0(men_men_n347_), .A1(men_men_n61_), .B0(men_men_n349_), .Y(men_men_n350_));
  NA2        u334(.A(x2), .B(men_men_n17_), .Y(men_men_n351_));
  NA2        u335(.A(men_men_n335_), .B(men_men_n92_), .Y(men_men_n352_));
  NA4        u336(.A(men_men_n352_), .B(men_men_n350_), .C(men_men_n346_), .D(men_men_n344_), .Y(men_men_n353_));
  OAI210     u337(.A0(men_men_n112_), .A1(x3), .B0(men_men_n311_), .Y(men_men_n354_));
  NA3        u338(.A(men_men_n232_), .B(men_men_n218_), .C(men_men_n82_), .Y(men_men_n355_));
  NA3        u339(.A(men_men_n355_), .B(men_men_n354_), .C(men_men_n156_), .Y(men_men_n356_));
  AOI210     u340(.A0(men_men_n353_), .A1(x4), .B0(men_men_n356_), .Y(men_men_n357_));
  NA3        u341(.A(men_men_n332_), .B(men_men_n213_), .C(men_men_n92_), .Y(men_men_n358_));
  NOi21      u342(.An(x4), .B(x0), .Y(men_men_n359_));
  XO2        u343(.A(x4), .B(x0), .Y(men_men_n360_));
  OAI210     u344(.A0(men_men_n360_), .A1(men_men_n118_), .B0(men_men_n275_), .Y(men_men_n361_));
  AOI220     u345(.A0(men_men_n361_), .A1(x8), .B0(men_men_n359_), .B1(men_men_n93_), .Y(men_men_n362_));
  AOI210     u346(.A0(men_men_n362_), .A1(men_men_n358_), .B0(x3), .Y(men_men_n363_));
  INV        u347(.A(men_men_n93_), .Y(men_men_n364_));
  NO2        u348(.A(men_men_n92_), .B(x4), .Y(men_men_n365_));
  AOI220     u349(.A0(men_men_n365_), .A1(men_men_n42_), .B0(men_men_n128_), .B1(men_men_n364_), .Y(men_men_n366_));
  NO3        u350(.A(men_men_n360_), .B(men_men_n167_), .C(x2), .Y(men_men_n367_));
  NO3        u351(.A(men_men_n232_), .B(men_men_n27_), .C(men_men_n23_), .Y(men_men_n368_));
  NO2        u352(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n369_));
  NA4        u353(.A(men_men_n369_), .B(men_men_n366_), .C(men_men_n228_), .D(x6), .Y(men_men_n370_));
  OAI220     u354(.A0(men_men_n310_), .A1(men_men_n90_), .B0(men_men_n185_), .B1(men_men_n92_), .Y(men_men_n371_));
  NO2        u355(.A(men_men_n41_), .B(x0), .Y(men_men_n372_));
  OR2        u356(.A(men_men_n365_), .B(men_men_n372_), .Y(men_men_n373_));
  NO2        u357(.A(men_men_n154_), .B(men_men_n107_), .Y(men_men_n374_));
  AOI220     u358(.A0(men_men_n374_), .A1(men_men_n373_), .B0(men_men_n371_), .B1(men_men_n59_), .Y(men_men_n375_));
  NO2        u359(.A(men_men_n154_), .B(men_men_n80_), .Y(men_men_n376_));
  NO2        u360(.A(men_men_n33_), .B(x2), .Y(men_men_n377_));
  NOi21      u361(.An(men_men_n124_), .B(men_men_n26_), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n377_), .A1(men_men_n376_), .B0(men_men_n378_), .Y(men_men_n379_));
  OAI210     u363(.A0(men_men_n375_), .A1(men_men_n60_), .B0(men_men_n379_), .Y(men_men_n380_));
  OAI220     u364(.A0(men_men_n380_), .A1(x6), .B0(men_men_n370_), .B1(men_men_n363_), .Y(men_men_n381_));
  OAI210     u365(.A0(men_men_n61_), .A1(men_men_n46_), .B0(men_men_n40_), .Y(men_men_n382_));
  OAI210     u366(.A0(men_men_n382_), .A1(men_men_n92_), .B0(men_men_n323_), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n383_), .A1(men_men_n18_), .B0(men_men_n156_), .Y(men_men_n384_));
  AO220      u368(.A0(men_men_n384_), .A1(men_men_n381_), .B0(men_men_n357_), .B1(men_men_n342_), .Y(men_men_n385_));
  NA2        u369(.A(men_men_n377_), .B(x6), .Y(men_men_n386_));
  AOI210     u370(.A0(x6), .A1(x1), .B0(men_men_n155_), .Y(men_men_n387_));
  NA2        u371(.A(men_men_n365_), .B(x0), .Y(men_men_n388_));
  NA2        u372(.A(men_men_n82_), .B(x6), .Y(men_men_n389_));
  OAI210     u373(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n389_), .Y(men_men_n390_));
  AOI220     u374(.A0(men_men_n390_), .A1(men_men_n386_), .B0(men_men_n222_), .B1(men_men_n47_), .Y(men_men_n391_));
  NA3        u375(.A(men_men_n391_), .B(men_men_n385_), .C(men_men_n329_), .Y(men_men_n392_));
  AOI210     u376(.A0(men_men_n204_), .A1(x8), .B0(men_men_n112_), .Y(men_men_n393_));
  NA2        u377(.A(men_men_n393_), .B(men_men_n351_), .Y(men_men_n394_));
  NA3        u378(.A(men_men_n394_), .B(men_men_n201_), .C(men_men_n156_), .Y(men_men_n395_));
  NA3        u379(.A(x7), .B(x3), .C(x0), .Y(men_men_n396_));
  NA2        u380(.A(men_men_n227_), .B(x0), .Y(men_men_n397_));
  OAI220     u381(.A0(men_men_n397_), .A1(men_men_n213_), .B0(men_men_n396_), .B1(men_men_n364_), .Y(men_men_n398_));
  INV        u382(.A(men_men_n398_), .Y(men_men_n399_));
  AOI210     u383(.A0(men_men_n399_), .A1(men_men_n395_), .B0(men_men_n24_), .Y(men_men_n400_));
  OAI210     u384(.A0(men_men_n201_), .A1(men_men_n66_), .B0(men_men_n210_), .Y(men_men_n401_));
  NA3        u385(.A(men_men_n204_), .B(men_men_n229_), .C(x8), .Y(men_men_n402_));
  AOI210     u386(.A0(men_men_n402_), .A1(men_men_n401_), .B0(men_men_n24_), .Y(men_men_n403_));
  AOI210     u387(.A0(men_men_n121_), .A1(men_men_n119_), .B0(men_men_n40_), .Y(men_men_n404_));
  NOi31      u388(.An(men_men_n404_), .B(men_men_n372_), .C(men_men_n186_), .Y(men_men_n405_));
  OAI210     u389(.A0(men_men_n405_), .A1(men_men_n403_), .B0(men_men_n153_), .Y(men_men_n406_));
  NAi31      u390(.An(men_men_n48_), .B(men_men_n299_), .C(men_men_n181_), .Y(men_men_n407_));
  NA2        u391(.A(men_men_n407_), .B(men_men_n406_), .Y(men_men_n408_));
  OAI210     u392(.A0(men_men_n408_), .A1(men_men_n400_), .B0(x6), .Y(men_men_n409_));
  OAI210     u393(.A0(men_men_n167_), .A1(men_men_n46_), .B0(men_men_n139_), .Y(men_men_n410_));
  NA3        u394(.A(men_men_n53_), .B(men_men_n36_), .C(men_men_n30_), .Y(men_men_n411_));
  AOI220     u395(.A0(men_men_n411_), .A1(men_men_n410_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n412_));
  NO2        u396(.A(men_men_n156_), .B(x0), .Y(men_men_n413_));
  AOI220     u397(.A0(men_men_n413_), .A1(men_men_n227_), .B0(men_men_n201_), .B1(men_men_n156_), .Y(men_men_n414_));
  AOI210     u398(.A0(men_men_n130_), .A1(men_men_n258_), .B0(x1), .Y(men_men_n415_));
  OAI210     u399(.A0(men_men_n414_), .A1(x8), .B0(men_men_n415_), .Y(men_men_n416_));
  NAi31      u400(.An(x2), .B(x8), .C(x0), .Y(men_men_n417_));
  OAI210     u401(.A0(men_men_n417_), .A1(x4), .B0(men_men_n168_), .Y(men_men_n418_));
  NA3        u402(.A(men_men_n418_), .B(men_men_n151_), .C(x9), .Y(men_men_n419_));
  NO4        u403(.A(men_men_n129_), .B(men_men_n310_), .C(x9), .D(x2), .Y(men_men_n420_));
  NOi21      u404(.An(men_men_n127_), .B(men_men_n185_), .Y(men_men_n421_));
  NO3        u405(.A(men_men_n421_), .B(men_men_n420_), .C(men_men_n18_), .Y(men_men_n422_));
  NA2        u406(.A(men_men_n376_), .B(men_men_n156_), .Y(men_men_n423_));
  NA4        u407(.A(men_men_n423_), .B(men_men_n422_), .C(men_men_n419_), .D(men_men_n48_), .Y(men_men_n424_));
  OAI210     u408(.A0(men_men_n416_), .A1(men_men_n412_), .B0(men_men_n424_), .Y(men_men_n425_));
  NOi31      u409(.An(men_men_n413_), .B(men_men_n31_), .C(x8), .Y(men_men_n426_));
  AOI210     u410(.A0(men_men_n36_), .A1(x9), .B0(men_men_n137_), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n427_), .B(men_men_n127_), .C(men_men_n41_), .Y(men_men_n428_));
  NOi31      u412(.An(x1), .B(x8), .C(x7), .Y(men_men_n429_));
  AOI210     u413(.A0(men_men_n275_), .A1(men_men_n58_), .B0(men_men_n126_), .Y(men_men_n430_));
  NO2        u414(.A(men_men_n430_), .B(x3), .Y(men_men_n431_));
  NO3        u415(.A(men_men_n431_), .B(men_men_n428_), .C(x2), .Y(men_men_n432_));
  OAI220     u416(.A0(men_men_n360_), .A1(men_men_n314_), .B0(men_men_n310_), .B1(men_men_n41_), .Y(men_men_n433_));
  AOI210     u417(.A0(x9), .A1(men_men_n46_), .B0(men_men_n396_), .Y(men_men_n434_));
  AOI220     u418(.A0(men_men_n434_), .A1(men_men_n92_), .B0(men_men_n433_), .B1(men_men_n156_), .Y(men_men_n435_));
  NO2        u419(.A(men_men_n435_), .B(men_men_n52_), .Y(men_men_n436_));
  NO3        u420(.A(men_men_n436_), .B(men_men_n432_), .C(men_men_n426_), .Y(men_men_n437_));
  AOI210     u421(.A0(men_men_n437_), .A1(men_men_n425_), .B0(men_men_n24_), .Y(men_men_n438_));
  NO3        u422(.A(men_men_n60_), .B(x4), .C(x1), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n440_));
  AOI220     u424(.A0(men_men_n440_), .A1(men_men_n276_), .B0(men_men_n439_), .B1(men_men_n404_), .Y(men_men_n441_));
  NO2        u425(.A(men_men_n441_), .B(men_men_n104_), .Y(men_men_n442_));
  NA2        u426(.A(men_men_n442_), .B(x7), .Y(men_men_n443_));
  NA2        u427(.A(men_men_n232_), .B(x7), .Y(men_men_n444_));
  NA3        u428(.A(men_men_n444_), .B(men_men_n155_), .C(men_men_n138_), .Y(men_men_n445_));
  NA2        u429(.A(men_men_n445_), .B(men_men_n443_), .Y(men_men_n446_));
  OAI210     u430(.A0(men_men_n446_), .A1(men_men_n438_), .B0(men_men_n34_), .Y(men_men_n447_));
  INV        u431(.A(men_men_n210_), .Y(men_men_n448_));
  NO4        u432(.A(men_men_n448_), .B(men_men_n77_), .C(x4), .D(men_men_n52_), .Y(men_men_n449_));
  NA2        u433(.A(men_men_n263_), .B(men_men_n21_), .Y(men_men_n450_));
  NO2        u434(.A(men_men_n164_), .B(men_men_n139_), .Y(men_men_n451_));
  NA2        u435(.A(men_men_n451_), .B(men_men_n450_), .Y(men_men_n452_));
  AOI210     u436(.A0(men_men_n452_), .A1(men_men_n171_), .B0(men_men_n27_), .Y(men_men_n453_));
  AOI220     u437(.A0(men_men_n372_), .A1(men_men_n92_), .B0(men_men_n154_), .B1(men_men_n204_), .Y(men_men_n454_));
  NA3        u438(.A(men_men_n454_), .B(men_men_n417_), .C(men_men_n90_), .Y(men_men_n455_));
  NA2        u439(.A(men_men_n455_), .B(men_men_n181_), .Y(men_men_n456_));
  OAI220     u440(.A0(x3), .A1(men_men_n67_), .B0(men_men_n164_), .B1(men_men_n41_), .Y(men_men_n457_));
  NA2        u441(.A(x3), .B(men_men_n52_), .Y(men_men_n458_));
  AOI210     u442(.A0(men_men_n168_), .A1(men_men_n26_), .B0(men_men_n72_), .Y(men_men_n459_));
  OAI210     u443(.A0(men_men_n153_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n460_));
  NO3        u444(.A(men_men_n429_), .B(x3), .C(men_men_n52_), .Y(men_men_n461_));
  AOI210     u445(.A0(men_men_n461_), .A1(men_men_n460_), .B0(men_men_n459_), .Y(men_men_n462_));
  OAI210     u446(.A0(men_men_n157_), .A1(men_men_n458_), .B0(men_men_n462_), .Y(men_men_n463_));
  AOI220     u447(.A0(men_men_n463_), .A1(x0), .B0(men_men_n457_), .B1(men_men_n139_), .Y(men_men_n464_));
  AOI210     u448(.A0(men_men_n464_), .A1(men_men_n456_), .B0(men_men_n240_), .Y(men_men_n465_));
  NA2        u449(.A(x9), .B(x5), .Y(men_men_n466_));
  NO4        u450(.A(men_men_n107_), .B(men_men_n466_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n467_));
  NO4        u451(.A(men_men_n467_), .B(men_men_n465_), .C(men_men_n453_), .D(men_men_n449_), .Y(men_men_n468_));
  NA3        u452(.A(men_men_n468_), .B(men_men_n447_), .C(men_men_n409_), .Y(men_men_n469_));
  AOI210     u453(.A0(men_men_n392_), .A1(men_men_n24_), .B0(men_men_n469_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule