// Benchmark "top" written by ABC on Fri Jun 21 17:49:26 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1058_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO2        g0062(.A(new_new_n83_), .B(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  NO2        g0064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  OAI210     g0066(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n88_), .Y(new_new_n89_));
  NAi21      g0067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g0068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g0069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n63_), .Y(new_new_n92_));
  NA2        g0070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  INV        g0071(.A(new_new_n92_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n89_), .B0(new_new_n80_), .Y(new_new_n95_));
  AN3        g0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g0074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g0075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g0076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g0077(.A0(new_new_n99_), .A1(new_new_n62_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g0078(.A(i_7_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n47_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g0080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(new_new_n86_), .Y(new_new_n104_));
  NA2        g0082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g0083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g0084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g0085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  NO3        g0086(.A(new_new_n108_), .B(new_new_n90_), .C(new_new_n54_), .Y(new_new_n109_));
  AN2        g0087(.A(i_2_), .B(i_10_), .Y(new_new_n110_));
  NO2        g0088(.A(new_new_n110_), .B(i_7_), .Y(new_new_n111_));
  OR2        g0089(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n112_));
  NO2        g0090(.A(i_8_), .B(new_new_n101_), .Y(new_new_n113_));
  NO3        g0091(.A(new_new_n113_), .B(new_new_n112_), .C(new_new_n111_), .Y(new_new_n114_));
  NA2        g0092(.A(i_12_), .B(i_7_), .Y(new_new_n115_));
  NO2        g0093(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  INV        g0095(.A(new_new_n117_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n118_), .B(new_new_n114_), .Y(new_new_n119_));
  NAi41      g0097(.An(new_new_n109_), .B(new_new_n119_), .C(new_new_n107_), .D(new_new_n100_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n47_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NOi31      g0107(.An(new_new_n129_), .B(new_new_n127_), .C(new_new_n126_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n86_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n48_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n108_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n95_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g0127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(new_new_n27_), .Y(new_new_n152_));
  NA2        g0130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n36_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  NO2        g0144(.A(new_new_n166_), .B(new_new_n156_), .Y(new_new_n167_));
  AOI210     g0145(.A0(new_new_n167_), .A1(new_new_n150_), .B0(new_new_n143_), .Y(new_new_n168_));
  NA3        g0146(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n169_));
  NA2        g0147(.A(i_3_), .B(new_new_n49_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_4_), .B(i_9_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_11_), .B(i_13_), .Y(new_new_n172_));
  NA2        g0150(.A(new_new_n172_), .B(new_new_n171_), .Y(new_new_n173_));
  OR2        g0151(.A(new_new_n173_), .B(new_new_n170_), .Y(new_new_n174_));
  NO2        g0152(.A(i_4_), .B(i_5_), .Y(new_new_n175_));
  NAi21      g0153(.An(i_12_), .B(i_11_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n176_), .B(i_13_), .Y(new_new_n177_));
  NA3        g0155(.A(new_new_n177_), .B(new_new_n175_), .C(new_new_n83_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(new_new_n169_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n180_));
  NA2        g0158(.A(new_new_n180_), .B(new_new_n47_), .Y(new_new_n181_));
  NAi31      g0159(.An(i_4_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n182_));
  NA2        g0160(.A(i_3_), .B(i_5_), .Y(new_new_n183_));
  OR2        g0161(.A(new_new_n183_), .B(new_new_n173_), .Y(new_new_n184_));
  AOI210     g0162(.A0(new_new_n184_), .A1(new_new_n182_), .B0(new_new_n181_), .Y(new_new_n185_));
  NO2        g0163(.A(new_new_n73_), .B(i_5_), .Y(new_new_n186_));
  NO2        g0164(.A(i_13_), .B(i_10_), .Y(new_new_n187_));
  NA3        g0165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n45_), .Y(new_new_n188_));
  NO2        g0166(.A(i_2_), .B(i_1_), .Y(new_new_n189_));
  NA2        g0167(.A(new_new_n189_), .B(i_3_), .Y(new_new_n190_));
  NAi21      g0168(.An(i_4_), .B(i_12_), .Y(new_new_n191_));
  NO4        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n188_), .D(new_new_n25_), .Y(new_new_n192_));
  NO3        g0170(.A(new_new_n192_), .B(new_new_n185_), .C(new_new_n179_), .Y(new_new_n193_));
  INV        g0171(.A(i_8_), .Y(new_new_n194_));
  NO2        g0172(.A(new_new_n194_), .B(i_7_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(i_6_), .Y(new_new_n196_));
  NO3        g0174(.A(i_3_), .B(new_new_n86_), .C(new_new_n49_), .Y(new_new_n197_));
  NA2        g0175(.A(new_new_n197_), .B(new_new_n113_), .Y(new_new_n198_));
  NO3        g0176(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n199_));
  NA3        g0177(.A(new_new_n199_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n200_));
  NO3        g0178(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n201_));
  OAI210     g0179(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n201_), .Y(new_new_n202_));
  AOI210     g0180(.A0(new_new_n202_), .A1(new_new_n200_), .B0(new_new_n198_), .Y(new_new_n203_));
  NO2        g0181(.A(i_3_), .B(i_8_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n205_));
  NA3        g0183(.A(new_new_n205_), .B(new_new_n204_), .C(new_new_n40_), .Y(new_new_n206_));
  NO2        g0184(.A(new_new_n103_), .B(new_new_n58_), .Y(new_new_n207_));
  INV        g0185(.A(new_new_n207_), .Y(new_new_n208_));
  NO2        g0186(.A(i_13_), .B(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(i_6_), .C(new_new_n194_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_3_), .Y(new_new_n211_));
  NO2        g0189(.A(new_new_n45_), .B(i_5_), .Y(new_new_n212_));
  NO3        g0190(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n213_));
  NA3        g0191(.A(new_new_n213_), .B(new_new_n212_), .C(i_10_), .Y(new_new_n214_));
  OAI220     g0192(.A0(new_new_n214_), .A1(new_new_n210_), .B0(new_new_n208_), .B1(new_new_n206_), .Y(new_new_n215_));
  AOI210     g0193(.A0(new_new_n215_), .A1(i_7_), .B0(new_new_n203_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(i_4_), .B0(new_new_n196_), .B1(new_new_n193_), .Y(new_new_n217_));
  NAi21      g0195(.An(i_12_), .B(i_7_), .Y(new_new_n218_));
  NA3        g0196(.A(i_13_), .B(new_new_n194_), .C(i_10_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n220_));
  NA2        g0198(.A(i_0_), .B(i_5_), .Y(new_new_n221_));
  NA2        g0199(.A(new_new_n221_), .B(new_new_n104_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(new_new_n190_), .B0(new_new_n181_), .B1(new_new_n133_), .Y(new_new_n223_));
  NAi31      g0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n36_), .B(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n226_), .C(new_new_n225_), .Y(new_new_n228_));
  INV        g0206(.A(i_13_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n229_), .Y(new_new_n230_));
  NA3        g0208(.A(new_new_n230_), .B(new_new_n199_), .C(new_new_n197_), .Y(new_new_n231_));
  OAI210     g0209(.A0(new_new_n228_), .A1(new_new_n224_), .B0(new_new_n231_), .Y(new_new_n232_));
  AOI220     g0210(.A0(new_new_n232_), .A1(new_new_n142_), .B0(new_new_n223_), .B1(new_new_n220_), .Y(new_new_n233_));
  NO2        g0211(.A(i_12_), .B(new_new_n37_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n183_), .B(i_4_), .Y(new_new_n235_));
  NA2        g0213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  OR2        g0214(.A(i_8_), .B(i_7_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n237_), .B(new_new_n86_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n54_), .B(i_1_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  INV        g0218(.A(i_12_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n45_), .B(new_new_n241_), .Y(new_new_n242_));
  NO3        g0220(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(i_2_), .B(i_1_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n240_), .B(new_new_n236_), .Y(new_new_n245_));
  NO3        g0223(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_4_), .B(i_3_), .Y(new_new_n247_));
  NO2        g0225(.A(i_0_), .B(i_6_), .Y(new_new_n248_));
  NOi41      g0226(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n249_));
  NA2        g0227(.A(new_new_n249_), .B(new_new_n248_), .Y(new_new_n250_));
  NO2        g0228(.A(new_new_n244_), .B(new_new_n183_), .Y(new_new_n251_));
  NAi21      g0229(.An(new_new_n250_), .B(new_new_n251_), .Y(new_new_n252_));
  INV        g0230(.A(new_new_n252_), .Y(new_new_n253_));
  AOI210     g0231(.A0(new_new_n253_), .A1(new_new_n40_), .B0(new_new_n245_), .Y(new_new_n254_));
  NO2        g0232(.A(i_11_), .B(new_new_n229_), .Y(new_new_n255_));
  NOi21      g0233(.An(i_1_), .B(i_6_), .Y(new_new_n256_));
  NAi21      g0234(.An(i_3_), .B(i_7_), .Y(new_new_n257_));
  NA2        g0235(.A(new_new_n241_), .B(i_9_), .Y(new_new_n258_));
  OR4        g0236(.A(new_new_n258_), .B(new_new_n257_), .C(new_new_n256_), .D(new_new_n186_), .Y(new_new_n259_));
  NO2        g0237(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n260_));
  NO2        g0238(.A(i_12_), .B(i_3_), .Y(new_new_n261_));
  NA2        g0239(.A(new_new_n73_), .B(i_5_), .Y(new_new_n262_));
  NA2        g0240(.A(i_3_), .B(i_9_), .Y(new_new_n263_));
  NAi21      g0241(.An(i_7_), .B(i_10_), .Y(new_new_n264_));
  NO2        g0242(.A(new_new_n264_), .B(new_new_n263_), .Y(new_new_n265_));
  NA3        g0243(.A(new_new_n265_), .B(new_new_n262_), .C(new_new_n64_), .Y(new_new_n266_));
  NA2        g0244(.A(new_new_n266_), .B(new_new_n259_), .Y(new_new_n267_));
  NA3        g0245(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n268_));
  INV        g0246(.A(new_new_n143_), .Y(new_new_n269_));
  NA2        g0247(.A(new_new_n241_), .B(i_13_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n270_), .B(new_new_n75_), .Y(new_new_n271_));
  AOI220     g0249(.A0(new_new_n271_), .A1(new_new_n269_), .B0(new_new_n267_), .B1(new_new_n255_), .Y(new_new_n272_));
  NO2        g0250(.A(new_new_n237_), .B(new_new_n37_), .Y(new_new_n273_));
  NA2        g0251(.A(i_12_), .B(i_6_), .Y(new_new_n274_));
  OR2        g0252(.A(i_13_), .B(i_9_), .Y(new_new_n275_));
  NO2        g0253(.A(new_new_n247_), .B(i_2_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n255_), .B(i_9_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n154_), .B(new_new_n63_), .Y(new_new_n278_));
  NO3        g0256(.A(i_11_), .B(new_new_n229_), .C(new_new_n25_), .Y(new_new_n279_));
  NO2        g0257(.A(new_new_n257_), .B(i_8_), .Y(new_new_n280_));
  NO2        g0258(.A(i_6_), .B(new_new_n49_), .Y(new_new_n281_));
  NA3        g0259(.A(new_new_n281_), .B(new_new_n280_), .C(new_new_n279_), .Y(new_new_n282_));
  NO3        g0260(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n283_));
  NA3        g0261(.A(new_new_n283_), .B(new_new_n273_), .C(new_new_n230_), .Y(new_new_n284_));
  AOI210     g0262(.A0(new_new_n284_), .A1(new_new_n282_), .B0(new_new_n278_), .Y(new_new_n285_));
  INV        g0263(.A(new_new_n285_), .Y(new_new_n286_));
  NA4        g0264(.A(new_new_n286_), .B(new_new_n272_), .C(new_new_n254_), .D(new_new_n233_), .Y(new_new_n287_));
  NO3        g0265(.A(i_12_), .B(new_new_n229_), .C(new_new_n37_), .Y(new_new_n288_));
  INV        g0266(.A(new_new_n288_), .Y(new_new_n289_));
  NA2        g0267(.A(i_8_), .B(new_new_n101_), .Y(new_new_n290_));
  NOi21      g0268(.An(new_new_n163_), .B(new_new_n86_), .Y(new_new_n291_));
  NO3        g0269(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n292_));
  AOI220     g0270(.A0(new_new_n292_), .A1(new_new_n197_), .B0(new_new_n291_), .B1(new_new_n239_), .Y(new_new_n293_));
  NO2        g0271(.A(new_new_n293_), .B(new_new_n290_), .Y(new_new_n294_));
  NO3        g0272(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n244_), .B(i_0_), .Y(new_new_n296_));
  AOI220     g0274(.A0(new_new_n296_), .A1(new_new_n195_), .B0(new_new_n295_), .B1(new_new_n142_), .Y(new_new_n297_));
  NA2        g0275(.A(new_new_n281_), .B(new_new_n26_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n298_), .B(new_new_n297_), .Y(new_new_n299_));
  NA2        g0277(.A(i_0_), .B(i_1_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n300_), .B(i_2_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n59_), .B(i_6_), .Y(new_new_n302_));
  NA3        g0280(.A(new_new_n302_), .B(new_new_n301_), .C(new_new_n163_), .Y(new_new_n303_));
  OAI210     g0281(.A0(new_new_n165_), .A1(new_new_n143_), .B0(new_new_n303_), .Y(new_new_n304_));
  NO3        g0282(.A(new_new_n304_), .B(new_new_n299_), .C(new_new_n294_), .Y(new_new_n305_));
  NO2        g0283(.A(i_3_), .B(i_10_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n307_));
  NO2        g0285(.A(i_2_), .B(new_new_n101_), .Y(new_new_n308_));
  NA2        g0286(.A(i_1_), .B(new_new_n36_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n309_), .B(i_8_), .Y(new_new_n310_));
  NOi21      g0288(.An(new_new_n221_), .B(new_new_n103_), .Y(new_new_n311_));
  NA3        g0289(.A(new_new_n311_), .B(new_new_n310_), .C(new_new_n308_), .Y(new_new_n312_));
  AN2        g0290(.A(i_3_), .B(i_10_), .Y(new_new_n313_));
  NA4        g0291(.A(new_new_n313_), .B(new_new_n199_), .C(new_new_n177_), .D(new_new_n175_), .Y(new_new_n314_));
  NO2        g0292(.A(i_5_), .B(new_new_n37_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n316_));
  OR2        g0294(.A(new_new_n312_), .B(new_new_n307_), .Y(new_new_n317_));
  OAI220     g0295(.A0(new_new_n317_), .A1(i_6_), .B0(new_new_n305_), .B1(new_new_n289_), .Y(new_new_n318_));
  NO4        g0296(.A(new_new_n318_), .B(new_new_n287_), .C(new_new_n217_), .D(new_new_n168_), .Y(new_new_n319_));
  NO3        g0297(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n320_));
  NO2        g0298(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n296_), .B(new_new_n321_), .Y(new_new_n322_));
  NO3        g0300(.A(i_6_), .B(new_new_n194_), .C(i_7_), .Y(new_new_n323_));
  NA2        g0301(.A(new_new_n323_), .B(new_new_n199_), .Y(new_new_n324_));
  AOI210     g0302(.A0(new_new_n324_), .A1(new_new_n322_), .B0(new_new_n170_), .Y(new_new_n325_));
  NO2        g0303(.A(i_2_), .B(i_3_), .Y(new_new_n326_));
  OR2        g0304(.A(i_0_), .B(i_5_), .Y(new_new_n327_));
  NA2        g0305(.A(new_new_n221_), .B(new_new_n327_), .Y(new_new_n328_));
  NA4        g0306(.A(new_new_n328_), .B(new_new_n238_), .C(new_new_n326_), .D(i_1_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n296_), .B(new_new_n291_), .C(new_new_n113_), .Y(new_new_n330_));
  NAi21      g0308(.An(i_8_), .B(i_7_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n331_), .B(i_6_), .Y(new_new_n332_));
  NO2        g0310(.A(new_new_n157_), .B(new_new_n47_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n333_), .B(new_new_n332_), .C(new_new_n163_), .Y(new_new_n334_));
  NA3        g0312(.A(new_new_n334_), .B(new_new_n330_), .C(new_new_n329_), .Y(new_new_n335_));
  OAI210     g0313(.A0(new_new_n335_), .A1(new_new_n325_), .B0(i_4_), .Y(new_new_n336_));
  NO2        g0314(.A(i_12_), .B(i_10_), .Y(new_new_n337_));
  NOi21      g0315(.An(i_5_), .B(i_0_), .Y(new_new_n338_));
  NO3        g0316(.A(new_new_n309_), .B(new_new_n338_), .C(new_new_n128_), .Y(new_new_n339_));
  NA2        g0317(.A(new_new_n339_), .B(new_new_n337_), .Y(new_new_n340_));
  NO2        g0318(.A(i_6_), .B(i_8_), .Y(new_new_n341_));
  NOi21      g0319(.An(i_0_), .B(i_2_), .Y(new_new_n342_));
  AN2        g0320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NO2        g0321(.A(i_1_), .B(i_7_), .Y(new_new_n344_));
  AO220      g0322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(new_new_n332_), .B1(new_new_n239_), .Y(new_new_n345_));
  NA2        g0323(.A(new_new_n345_), .B(new_new_n42_), .Y(new_new_n346_));
  NA3        g0324(.A(new_new_n346_), .B(new_new_n340_), .C(new_new_n336_), .Y(new_new_n347_));
  NO3        g0325(.A(new_new_n237_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n348_));
  NO3        g0326(.A(new_new_n331_), .B(i_2_), .C(i_1_), .Y(new_new_n349_));
  OAI210     g0327(.A0(new_new_n349_), .A1(new_new_n348_), .B0(i_6_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n256_), .B(new_new_n308_), .C(new_new_n194_), .Y(new_new_n351_));
  AOI210     g0329(.A0(new_new_n351_), .A1(new_new_n350_), .B0(new_new_n328_), .Y(new_new_n352_));
  NOi21      g0330(.An(new_new_n153_), .B(new_new_n104_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n353_), .B(new_new_n124_), .Y(new_new_n354_));
  OAI210     g0332(.A0(new_new_n354_), .A1(new_new_n352_), .B0(i_3_), .Y(new_new_n355_));
  INV        g0333(.A(new_new_n84_), .Y(new_new_n356_));
  NO2        g0334(.A(new_new_n300_), .B(new_new_n81_), .Y(new_new_n357_));
  NA2        g0335(.A(new_new_n357_), .B(new_new_n132_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n93_), .B(new_new_n194_), .Y(new_new_n359_));
  NA3        g0337(.A(new_new_n311_), .B(new_new_n359_), .C(new_new_n63_), .Y(new_new_n360_));
  AOI210     g0338(.A0(new_new_n360_), .A1(new_new_n358_), .B0(new_new_n356_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n194_), .B(i_9_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n207_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n363_), .B(new_new_n47_), .Y(new_new_n364_));
  NO3        g0342(.A(new_new_n364_), .B(new_new_n361_), .C(new_new_n299_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n365_), .A1(new_new_n355_), .B0(new_new_n162_), .Y(new_new_n366_));
  AOI210     g0344(.A0(new_new_n347_), .A1(new_new_n320_), .B0(new_new_n366_), .Y(new_new_n367_));
  NOi32      g0345(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n368_));
  INV        g0346(.A(new_new_n368_), .Y(new_new_n369_));
  NAi21      g0347(.An(i_0_), .B(i_6_), .Y(new_new_n370_));
  NAi21      g0348(.An(i_1_), .B(i_5_), .Y(new_new_n371_));
  NA2        g0349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  NA2        g0350(.A(new_new_n372_), .B(new_new_n25_), .Y(new_new_n373_));
  OAI210     g0351(.A0(new_new_n373_), .A1(new_new_n159_), .B0(new_new_n250_), .Y(new_new_n374_));
  NAi41      g0352(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n375_));
  OAI220     g0353(.A0(new_new_n375_), .A1(new_new_n371_), .B0(new_new_n224_), .B1(new_new_n159_), .Y(new_new_n376_));
  AOI210     g0354(.A0(new_new_n375_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n377_));
  NOi32      g0355(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n378_));
  NAi21      g0356(.An(i_6_), .B(i_1_), .Y(new_new_n379_));
  NA3        g0357(.A(new_new_n379_), .B(new_new_n378_), .C(new_new_n47_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n380_), .B(i_0_), .Y(new_new_n381_));
  OR3        g0359(.A(new_new_n381_), .B(new_new_n377_), .C(new_new_n376_), .Y(new_new_n382_));
  NO2        g0360(.A(i_1_), .B(new_new_n101_), .Y(new_new_n383_));
  NAi21      g0361(.An(i_3_), .B(i_4_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n384_), .B(i_9_), .Y(new_new_n385_));
  AN2        g0363(.A(i_6_), .B(i_7_), .Y(new_new_n386_));
  OAI210     g0364(.A0(new_new_n386_), .A1(new_new_n383_), .B0(new_new_n385_), .Y(new_new_n387_));
  NA2        g0365(.A(i_2_), .B(i_7_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n384_), .B(i_10_), .Y(new_new_n389_));
  NA3        g0367(.A(new_new_n389_), .B(new_new_n388_), .C(new_new_n248_), .Y(new_new_n390_));
  AOI210     g0368(.A0(new_new_n390_), .A1(new_new_n387_), .B0(new_new_n186_), .Y(new_new_n391_));
  AOI210     g0369(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n392_));
  OAI210     g0370(.A0(new_new_n392_), .A1(new_new_n189_), .B0(new_new_n389_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n393_), .B(i_5_), .Y(new_new_n394_));
  NO4        g0372(.A(new_new_n394_), .B(new_new_n391_), .C(new_new_n382_), .D(new_new_n374_), .Y(new_new_n395_));
  NO2        g0373(.A(new_new_n395_), .B(new_new_n369_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n397_));
  AN2        g0375(.A(i_12_), .B(i_5_), .Y(new_new_n398_));
  NA2        g0376(.A(i_3_), .B(new_new_n398_), .Y(new_new_n399_));
  NO2        g0377(.A(i_11_), .B(i_6_), .Y(new_new_n400_));
  NA3        g0378(.A(new_new_n400_), .B(new_new_n333_), .C(new_new_n229_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n401_), .B(new_new_n399_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n247_), .B(i_5_), .Y(new_new_n403_));
  NO2        g0381(.A(i_5_), .B(i_10_), .Y(new_new_n404_));
  AOI220     g0382(.A0(new_new_n404_), .A1(new_new_n276_), .B0(new_new_n403_), .B1(new_new_n199_), .Y(new_new_n405_));
  NA2        g0383(.A(new_new_n144_), .B(new_new_n46_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n406_), .B(new_new_n405_), .Y(new_new_n407_));
  OAI210     g0385(.A0(new_new_n407_), .A1(new_new_n402_), .B0(new_new_n397_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n150_), .B(new_new_n86_), .Y(new_new_n410_));
  OAI210     g0388(.A0(new_new_n410_), .A1(new_new_n402_), .B0(new_new_n409_), .Y(new_new_n411_));
  NO3        g0389(.A(new_new_n86_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n412_));
  NO2        g0390(.A(i_3_), .B(new_new_n101_), .Y(new_new_n413_));
  NA2        g0391(.A(new_new_n306_), .B(new_new_n91_), .Y(new_new_n414_));
  NO2        g0392(.A(i_11_), .B(i_12_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n415_), .B(new_new_n36_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n414_), .B(new_new_n416_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n404_), .B(new_new_n241_), .Y(new_new_n418_));
  NA3        g0396(.A(new_new_n113_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n224_), .Y(new_new_n420_));
  NAi21      g0398(.An(i_13_), .B(i_0_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n421_), .B(new_new_n244_), .Y(new_new_n422_));
  OAI210     g0400(.A0(new_new_n420_), .A1(new_new_n417_), .B0(new_new_n422_), .Y(new_new_n423_));
  NA3        g0401(.A(new_new_n423_), .B(new_new_n411_), .C(new_new_n408_), .Y(new_new_n424_));
  NO3        g0402(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n425_));
  NO2        g0403(.A(i_0_), .B(i_11_), .Y(new_new_n426_));
  INV        g0404(.A(i_5_), .Y(new_new_n427_));
  AN2        g0405(.A(i_1_), .B(i_6_), .Y(new_new_n428_));
  NOi21      g0406(.An(i_2_), .B(i_12_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n430_), .B(new_new_n427_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n142_), .B(i_9_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n432_), .B(i_4_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n431_), .B(new_new_n433_), .Y(new_new_n434_));
  NAi21      g0412(.An(i_9_), .B(i_4_), .Y(new_new_n435_));
  OR2        g0413(.A(i_13_), .B(i_10_), .Y(new_new_n436_));
  NO3        g0414(.A(new_new_n436_), .B(new_new_n117_), .C(new_new_n435_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n173_), .B(new_new_n123_), .Y(new_new_n438_));
  OR2        g0416(.A(new_new_n219_), .B(new_new_n218_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n288_), .B(new_new_n440_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n281_), .B(new_new_n213_), .Y(new_new_n442_));
  OAI220     g0420(.A0(new_new_n442_), .A1(new_new_n439_), .B0(new_new_n441_), .B1(new_new_n353_), .Y(new_new_n443_));
  INV        g0421(.A(new_new_n443_), .Y(new_new_n444_));
  AOI210     g0422(.A0(new_new_n444_), .A1(new_new_n434_), .B0(new_new_n26_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n330_), .B(new_new_n329_), .Y(new_new_n446_));
  AOI220     g0424(.A0(new_new_n302_), .A1(new_new_n292_), .B0(new_new_n296_), .B1(new_new_n321_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(new_new_n170_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n183_), .B(new_new_n86_), .Y(new_new_n449_));
  AOI220     g0427(.A0(new_new_n449_), .A1(new_new_n301_), .B0(new_new_n283_), .B1(new_new_n213_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n450_), .B(new_new_n290_), .Y(new_new_n451_));
  NO3        g0429(.A(new_new_n451_), .B(new_new_n448_), .C(new_new_n446_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n197_), .B(new_new_n96_), .Y(new_new_n453_));
  NA3        g0431(.A(new_new_n333_), .B(new_new_n163_), .C(new_new_n86_), .Y(new_new_n454_));
  AOI210     g0432(.A0(new_new_n454_), .A1(new_new_n453_), .B0(new_new_n331_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n194_), .B(i_10_), .Y(new_new_n456_));
  NA3        g0434(.A(new_new_n262_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n302_), .B(new_new_n239_), .Y(new_new_n458_));
  OAI220     g0436(.A0(new_new_n458_), .A1(new_new_n183_), .B0(new_new_n457_), .B1(new_new_n456_), .Y(new_new_n459_));
  NO2        g0437(.A(i_3_), .B(new_new_n49_), .Y(new_new_n460_));
  NA3        g0438(.A(new_new_n344_), .B(new_new_n343_), .C(new_new_n460_), .Y(new_new_n461_));
  NA2        g0439(.A(new_new_n323_), .B(new_new_n328_), .Y(new_new_n462_));
  OAI210     g0440(.A0(new_new_n462_), .A1(new_new_n190_), .B0(new_new_n461_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n463_), .B(new_new_n459_), .C(new_new_n455_), .Y(new_new_n464_));
  AOI210     g0442(.A0(new_new_n464_), .A1(new_new_n452_), .B0(new_new_n277_), .Y(new_new_n465_));
  NO4        g0443(.A(new_new_n465_), .B(new_new_n445_), .C(new_new_n424_), .D(new_new_n396_), .Y(new_new_n466_));
  NO2        g0444(.A(new_new_n63_), .B(i_4_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n73_), .B(i_13_), .Y(new_new_n468_));
  NO2        g0446(.A(i_10_), .B(i_9_), .Y(new_new_n469_));
  NAi21      g0447(.An(i_12_), .B(i_8_), .Y(new_new_n470_));
  NO2        g0448(.A(new_new_n470_), .B(i_3_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n47_), .B(i_4_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n472_), .B(new_new_n104_), .Y(new_new_n473_));
  NO2        g0451(.A(new_new_n473_), .B(new_new_n206_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n316_), .B(i_0_), .Y(new_new_n475_));
  NO3        g0453(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n274_), .B(new_new_n97_), .Y(new_new_n477_));
  NA2        g0455(.A(new_new_n477_), .B(new_new_n476_), .Y(new_new_n478_));
  NA2        g0456(.A(i_8_), .B(i_9_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n255_), .B(new_new_n315_), .Y(new_new_n480_));
  NO3        g0458(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n481_));
  INV        g0459(.A(new_new_n481_), .Y(new_new_n482_));
  NA3        g0460(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n483_));
  NA4        g0461(.A(new_new_n145_), .B(new_new_n116_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n484_));
  OAI220     g0462(.A0(new_new_n484_), .A1(new_new_n483_), .B0(new_new_n482_), .B1(new_new_n480_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n485_), .B(new_new_n474_), .Y(new_new_n486_));
  INV        g0464(.A(new_new_n301_), .Y(new_new_n487_));
  OR2        g0465(.A(new_new_n487_), .B(new_new_n210_), .Y(new_new_n488_));
  OA210      g0466(.A0(new_new_n363_), .A1(new_new_n101_), .B0(new_new_n303_), .Y(new_new_n489_));
  OA220      g0467(.A0(new_new_n489_), .A1(new_new_n162_), .B0(new_new_n488_), .B1(new_new_n236_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n96_), .B(i_13_), .Y(new_new_n491_));
  NA2        g0469(.A(new_new_n449_), .B(new_new_n397_), .Y(new_new_n492_));
  NO2        g0470(.A(i_2_), .B(i_13_), .Y(new_new_n493_));
  NA3        g0471(.A(new_new_n493_), .B(new_new_n161_), .C(new_new_n99_), .Y(new_new_n494_));
  OAI220     g0472(.A0(new_new_n494_), .A1(new_new_n241_), .B0(new_new_n492_), .B1(new_new_n491_), .Y(new_new_n495_));
  NO3        g0473(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n496_));
  NO2        g0474(.A(i_6_), .B(i_7_), .Y(new_new_n497_));
  NA2        g0475(.A(new_new_n497_), .B(new_new_n496_), .Y(new_new_n498_));
  NO2        g0476(.A(i_11_), .B(i_1_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n73_), .B(i_3_), .Y(new_new_n500_));
  OR2        g0478(.A(i_11_), .B(i_8_), .Y(new_new_n501_));
  NOi21      g0479(.An(i_2_), .B(i_7_), .Y(new_new_n502_));
  NAi31      g0480(.An(new_new_n501_), .B(new_new_n502_), .C(new_new_n500_), .Y(new_new_n503_));
  NO2        g0481(.A(new_new_n436_), .B(i_6_), .Y(new_new_n504_));
  NA2        g0482(.A(new_new_n504_), .B(new_new_n467_), .Y(new_new_n505_));
  NO2        g0483(.A(new_new_n505_), .B(new_new_n503_), .Y(new_new_n506_));
  NO2        g0484(.A(i_3_), .B(new_new_n194_), .Y(new_new_n507_));
  NO2        g0485(.A(i_6_), .B(i_10_), .Y(new_new_n508_));
  NA4        g0486(.A(new_new_n508_), .B(new_new_n320_), .C(new_new_n507_), .D(new_new_n241_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n509_), .B(new_new_n155_), .Y(new_new_n510_));
  NA3        g0488(.A(new_new_n249_), .B(new_new_n172_), .C(new_new_n132_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n512_));
  NO2        g0490(.A(new_new_n157_), .B(i_3_), .Y(new_new_n513_));
  NAi31      g0491(.An(new_new_n512_), .B(new_new_n513_), .C(new_new_n230_), .Y(new_new_n514_));
  NA3        g0492(.A(new_new_n409_), .B(new_new_n180_), .C(new_new_n149_), .Y(new_new_n515_));
  NA3        g0493(.A(new_new_n515_), .B(new_new_n514_), .C(new_new_n511_), .Y(new_new_n516_));
  NO4        g0494(.A(new_new_n516_), .B(new_new_n510_), .C(new_new_n506_), .D(new_new_n495_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n476_), .B(new_new_n398_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n481_), .B(new_new_n404_), .Y(new_new_n519_));
  NO2        g0497(.A(new_new_n519_), .B(new_new_n228_), .Y(new_new_n520_));
  NAi21      g0498(.An(new_new_n219_), .B(new_new_n415_), .Y(new_new_n521_));
  NO2        g0499(.A(new_new_n26_), .B(i_5_), .Y(new_new_n522_));
  NO2        g0500(.A(i_0_), .B(new_new_n86_), .Y(new_new_n523_));
  NA3        g0501(.A(new_new_n523_), .B(new_new_n522_), .C(new_new_n142_), .Y(new_new_n524_));
  OR3        g0502(.A(new_new_n309_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n524_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n27_), .B(i_10_), .Y(new_new_n527_));
  NO2        g0505(.A(new_new_n527_), .B(new_new_n491_), .Y(new_new_n528_));
  NA4        g0506(.A(new_new_n313_), .B(new_new_n227_), .C(new_new_n73_), .D(new_new_n241_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n529_), .B(new_new_n498_), .Y(new_new_n530_));
  NO4        g0508(.A(new_new_n530_), .B(new_new_n528_), .C(new_new_n526_), .D(new_new_n520_), .Y(new_new_n531_));
  NA4        g0509(.A(new_new_n531_), .B(new_new_n517_), .C(new_new_n490_), .D(new_new_n486_), .Y(new_new_n532_));
  NA3        g0510(.A(new_new_n313_), .B(new_new_n177_), .C(new_new_n175_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n307_), .A1(i_4_), .B0(new_new_n533_), .Y(new_new_n534_));
  AN2        g0512(.A(new_new_n292_), .B(new_new_n238_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n535_), .B(new_new_n534_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n320_), .B(new_new_n164_), .Y(new_new_n537_));
  OAI210     g0515(.A0(new_new_n537_), .A1(new_new_n236_), .B0(new_new_n314_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n538_), .B(new_new_n332_), .Y(new_new_n539_));
  NA2        g0517(.A(new_new_n398_), .B(new_new_n229_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n386_), .B(new_new_n378_), .Y(new_new_n541_));
  OR2        g0519(.A(new_new_n540_), .B(new_new_n541_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n36_), .B(i_8_), .Y(new_new_n543_));
  AOI210     g0521(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n437_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n544_), .B(new_new_n542_), .Y(new_new_n545_));
  INV        g0523(.A(new_new_n545_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n262_), .B(new_new_n64_), .Y(new_new_n547_));
  OAI210     g0525(.A0(i_8_), .A1(new_new_n547_), .B0(new_new_n134_), .Y(new_new_n548_));
  AOI210     g0526(.A0(new_new_n195_), .A1(i_9_), .B0(new_new_n273_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n549_), .B(new_new_n200_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n183_), .B(new_new_n86_), .Y(new_new_n551_));
  AOI220     g0529(.A0(new_new_n551_), .A1(new_new_n550_), .B0(new_new_n548_), .B1(new_new_n438_), .Y(new_new_n552_));
  NA4        g0530(.A(new_new_n552_), .B(new_new_n546_), .C(new_new_n539_), .D(new_new_n536_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n403_), .B(new_new_n301_), .Y(new_new_n554_));
  OAI210     g0532(.A0(new_new_n399_), .A1(new_new_n169_), .B0(new_new_n554_), .Y(new_new_n555_));
  NO2        g0533(.A(i_12_), .B(new_new_n194_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n556_), .B(new_new_n229_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n508_), .B(new_new_n27_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n558_), .B(new_new_n557_), .Y(new_new_n559_));
  NOi31      g0537(.An(new_new_n323_), .B(new_new_n436_), .C(new_new_n38_), .Y(new_new_n560_));
  OAI210     g0538(.A0(new_new_n560_), .A1(new_new_n559_), .B0(new_new_n555_), .Y(new_new_n561_));
  NO2        g0539(.A(i_8_), .B(i_7_), .Y(new_new_n562_));
  OAI210     g0540(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n563_), .B(new_new_n227_), .Y(new_new_n564_));
  AOI220     g0542(.A0(new_new_n333_), .A1(new_new_n40_), .B0(new_new_n239_), .B1(new_new_n209_), .Y(new_new_n565_));
  OAI220     g0543(.A0(new_new_n565_), .A1(new_new_n183_), .B0(new_new_n564_), .B1(new_new_n247_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n45_), .B(i_10_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n567_), .B(i_6_), .Y(new_new_n568_));
  NA3        g0546(.A(new_new_n568_), .B(new_new_n566_), .C(new_new_n562_), .Y(new_new_n569_));
  NA2        g0547(.A(new_new_n449_), .B(new_new_n333_), .Y(new_new_n570_));
  OAI220     g0548(.A0(new_new_n570_), .A1(new_new_n270_), .B0(new_new_n491_), .B1(new_new_n133_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n571_), .B(new_new_n273_), .Y(new_new_n572_));
  NOi31      g0550(.An(new_new_n296_), .B(new_new_n307_), .C(i_4_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n157_), .B(i_5_), .Y(new_new_n574_));
  NA2        g0552(.A(new_new_n573_), .B(new_new_n481_), .Y(new_new_n575_));
  NA4        g0553(.A(new_new_n575_), .B(new_new_n572_), .C(new_new_n569_), .D(new_new_n561_), .Y(new_new_n576_));
  NA3        g0554(.A(new_new_n221_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n577_));
  NA2        g0555(.A(new_new_n288_), .B(new_new_n84_), .Y(new_new_n578_));
  AOI210     g0556(.A0(new_new_n577_), .A1(new_new_n358_), .B0(new_new_n578_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n302_), .B(new_new_n292_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n580_), .B(new_new_n174_), .Y(new_new_n581_));
  NA2        g0559(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n582_));
  NA2        g0560(.A(new_new_n469_), .B(new_new_n225_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n582_), .B(new_new_n583_), .Y(new_new_n584_));
  AOI210     g0562(.A0(new_new_n379_), .A1(new_new_n47_), .B0(new_new_n383_), .Y(new_new_n585_));
  NA2        g0563(.A(i_0_), .B(new_new_n49_), .Y(new_new_n586_));
  NA3        g0564(.A(new_new_n556_), .B(new_new_n279_), .C(new_new_n586_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n585_), .B(new_new_n587_), .Y(new_new_n588_));
  NO4        g0566(.A(new_new_n588_), .B(new_new_n584_), .C(new_new_n581_), .D(new_new_n579_), .Y(new_new_n589_));
  NO4        g0567(.A(new_new_n256_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n590_));
  NO3        g0568(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n237_), .B(new_new_n36_), .Y(new_new_n592_));
  AN2        g0570(.A(new_new_n592_), .B(new_new_n591_), .Y(new_new_n593_));
  OA210      g0571(.A0(new_new_n593_), .A1(new_new_n590_), .B0(new_new_n368_), .Y(new_new_n594_));
  NO2        g0572(.A(new_new_n436_), .B(i_1_), .Y(new_new_n595_));
  NOi31      g0573(.An(new_new_n595_), .B(new_new_n477_), .C(new_new_n73_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n447_), .B(new_new_n178_), .Y(new_new_n597_));
  NO2        g0575(.A(new_new_n597_), .B(new_new_n594_), .Y(new_new_n598_));
  NOi21      g0576(.An(i_10_), .B(i_6_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n600_));
  NO2        g0578(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n601_));
  NA2        g0579(.A(new_new_n323_), .B(new_new_n164_), .Y(new_new_n602_));
  AOI220     g0580(.A0(new_new_n602_), .A1(new_new_n458_), .B0(new_new_n184_), .B1(new_new_n182_), .Y(new_new_n603_));
  INV        g0581(.A(new_new_n603_), .Y(new_new_n604_));
  INV        g0582(.A(new_new_n326_), .Y(new_new_n605_));
  NO2        g0583(.A(i_12_), .B(new_new_n86_), .Y(new_new_n606_));
  NA3        g0584(.A(new_new_n606_), .B(new_new_n279_), .C(new_new_n586_), .Y(new_new_n607_));
  NA3        g0585(.A(new_new_n400_), .B(new_new_n288_), .C(new_new_n221_), .Y(new_new_n608_));
  AOI210     g0586(.A0(new_new_n608_), .A1(new_new_n607_), .B0(new_new_n605_), .Y(new_new_n609_));
  NO3        g0587(.A(i_4_), .B(new_new_n350_), .C(new_new_n307_), .Y(new_new_n610_));
  OR2        g0588(.A(i_2_), .B(i_5_), .Y(new_new_n611_));
  OR2        g0589(.A(new_new_n611_), .B(new_new_n428_), .Y(new_new_n612_));
  AOI210     g0590(.A0(new_new_n388_), .A1(new_new_n248_), .B0(new_new_n199_), .Y(new_new_n613_));
  AOI210     g0591(.A0(new_new_n613_), .A1(new_new_n612_), .B0(new_new_n521_), .Y(new_new_n614_));
  NO3        g0592(.A(new_new_n614_), .B(new_new_n610_), .C(new_new_n609_), .Y(new_new_n615_));
  NA4        g0593(.A(new_new_n615_), .B(new_new_n604_), .C(new_new_n598_), .D(new_new_n589_), .Y(new_new_n616_));
  NO4        g0594(.A(new_new_n616_), .B(new_new_n576_), .C(new_new_n553_), .D(new_new_n532_), .Y(new_new_n617_));
  NA4        g0595(.A(new_new_n617_), .B(new_new_n466_), .C(new_new_n367_), .D(new_new_n319_), .Y(men7));
  NO2        g0596(.A(new_new_n93_), .B(new_new_n55_), .Y(new_new_n619_));
  NA2        g0597(.A(new_new_n508_), .B(new_new_n84_), .Y(new_new_n620_));
  NA2        g0598(.A(i_11_), .B(new_new_n194_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n144_), .B(new_new_n621_), .Y(new_new_n622_));
  NO2        g0600(.A(new_new_n622_), .B(new_new_n620_), .Y(new_new_n623_));
  NA3        g0601(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n241_), .B(i_4_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n625_), .B(i_8_), .Y(new_new_n626_));
  NO2        g0604(.A(new_new_n105_), .B(new_new_n624_), .Y(new_new_n627_));
  NA2        g0605(.A(i_2_), .B(new_new_n86_), .Y(new_new_n628_));
  OAI210     g0606(.A0(new_new_n87_), .A1(new_new_n204_), .B0(new_new_n205_), .Y(new_new_n629_));
  NO2        g0607(.A(i_7_), .B(new_new_n37_), .Y(new_new_n630_));
  NA2        g0608(.A(i_4_), .B(i_8_), .Y(new_new_n631_));
  AOI210     g0609(.A0(new_new_n631_), .A1(new_new_n313_), .B0(new_new_n630_), .Y(new_new_n632_));
  OAI220     g0610(.A0(new_new_n632_), .A1(new_new_n628_), .B0(new_new_n629_), .B1(i_13_), .Y(new_new_n633_));
  NO4        g0611(.A(new_new_n633_), .B(new_new_n627_), .C(new_new_n623_), .D(new_new_n619_), .Y(new_new_n634_));
  AOI210     g0612(.A0(new_new_n128_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n635_));
  AOI210     g0613(.A0(new_new_n635_), .A1(new_new_n241_), .B0(new_new_n161_), .Y(new_new_n636_));
  OR2        g0614(.A(i_6_), .B(i_10_), .Y(new_new_n637_));
  NO2        g0615(.A(new_new_n637_), .B(new_new_n23_), .Y(new_new_n638_));
  OR3        g0616(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n639_));
  NO3        g0617(.A(new_new_n639_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n640_));
  INV        g0618(.A(new_new_n201_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n640_), .B(new_new_n638_), .Y(new_new_n642_));
  OA220      g0620(.A0(new_new_n642_), .A1(new_new_n605_), .B0(new_new_n636_), .B1(new_new_n275_), .Y(new_new_n643_));
  AOI210     g0621(.A0(new_new_n643_), .A1(new_new_n634_), .B0(new_new_n63_), .Y(new_new_n644_));
  NOi21      g0622(.An(i_11_), .B(i_7_), .Y(new_new_n645_));
  AO210      g0623(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n647_), .B(new_new_n209_), .Y(new_new_n648_));
  NA3        g0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n649_));
  NAi31      g0627(.An(new_new_n649_), .B(new_new_n218_), .C(i_11_), .Y(new_new_n650_));
  AOI210     g0628(.A0(new_new_n650_), .A1(new_new_n648_), .B0(new_new_n63_), .Y(new_new_n651_));
  NA2        g0629(.A(new_new_n230_), .B(new_new_n63_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n63_), .B(i_9_), .Y(new_new_n653_));
  NO2        g0631(.A(i_1_), .B(i_12_), .Y(new_new_n654_));
  INV        g0632(.A(new_new_n652_), .Y(new_new_n655_));
  OAI210     g0633(.A0(new_new_n655_), .A1(new_new_n651_), .B0(i_6_), .Y(new_new_n656_));
  NO2        g0634(.A(new_new_n649_), .B(new_new_n108_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(new_new_n606_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n241_), .B(new_new_n86_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n659_), .B(i_11_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n658_), .B(new_new_n478_), .Y(new_new_n661_));
  NO4        g0639(.A(new_new_n218_), .B(new_new_n128_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(new_new_n653_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n241_), .B(i_6_), .Y(new_new_n664_));
  NO3        g0642(.A(new_new_n637_), .B(new_new_n237_), .C(new_new_n23_), .Y(new_new_n665_));
  AOI210     g0643(.A0(i_1_), .A1(new_new_n265_), .B0(new_new_n665_), .Y(new_new_n666_));
  OAI210     g0644(.A0(new_new_n666_), .A1(new_new_n45_), .B0(new_new_n663_), .Y(new_new_n667_));
  NA3        g0645(.A(new_new_n562_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n138_), .B(i_9_), .Y(new_new_n669_));
  NA3        g0647(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n47_), .B(i_1_), .Y(new_new_n671_));
  NA3        g0649(.A(new_new_n671_), .B(new_new_n274_), .C(new_new_n45_), .Y(new_new_n672_));
  OAI220     g0650(.A0(new_new_n672_), .A1(new_new_n670_), .B0(new_new_n669_), .B1(new_new_n1058_), .Y(new_new_n673_));
  NA3        g0651(.A(new_new_n653_), .B(new_new_n326_), .C(i_6_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n23_), .Y(new_new_n675_));
  AOI210     g0653(.A0(new_new_n499_), .A1(new_new_n440_), .B0(new_new_n246_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n676_), .B(new_new_n628_), .Y(new_new_n677_));
  NAi21      g0655(.An(new_new_n668_), .B(new_new_n92_), .Y(new_new_n678_));
  NA2        g0656(.A(new_new_n671_), .B(new_new_n274_), .Y(new_new_n679_));
  NO2        g0657(.A(i_11_), .B(new_new_n37_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n680_), .B(new_new_n24_), .Y(new_new_n681_));
  OAI210     g0659(.A0(new_new_n681_), .A1(new_new_n679_), .B0(new_new_n678_), .Y(new_new_n682_));
  OR4        g0660(.A(new_new_n682_), .B(new_new_n677_), .C(new_new_n675_), .D(new_new_n673_), .Y(new_new_n683_));
  NO3        g0661(.A(new_new_n683_), .B(new_new_n667_), .C(new_new_n661_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n241_), .B(new_new_n101_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n685_), .B(new_new_n645_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n686_), .B(i_1_), .Y(new_new_n687_));
  NO2        g0665(.A(new_new_n687_), .B(new_new_n639_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n435_), .B(new_new_n86_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n688_), .B(new_new_n47_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n237_), .B(new_new_n45_), .Y(new_new_n691_));
  NO3        g0669(.A(new_new_n691_), .B(new_new_n316_), .C(new_new_n242_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n693_), .B(i_6_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n86_), .B(i_9_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n63_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n654_), .Y(new_new_n697_));
  NO4        g0675(.A(new_new_n697_), .B(new_new_n694_), .C(new_new_n692_), .D(i_4_), .Y(new_new_n698_));
  NA2        g0676(.A(i_1_), .B(i_3_), .Y(new_new_n699_));
  INV        g0677(.A(new_new_n698_), .Y(new_new_n700_));
  NA4        g0678(.A(new_new_n700_), .B(new_new_n690_), .C(new_new_n684_), .D(new_new_n656_), .Y(new_new_n701_));
  NA2        g0679(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n702_));
  NA3        g0680(.A(new_new_n508_), .B(new_new_n543_), .C(new_new_n47_), .Y(new_new_n703_));
  NO3        g0681(.A(new_new_n502_), .B(new_new_n631_), .C(new_new_n86_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n704_), .B(new_new_n25_), .Y(new_new_n705_));
  NA3        g0683(.A(new_new_n161_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n706_));
  NA4        g0684(.A(new_new_n706_), .B(new_new_n705_), .C(new_new_n703_), .D(new_new_n702_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n707_), .B(i_1_), .Y(new_new_n708_));
  AOI210     g0686(.A0(new_new_n274_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n709_));
  NO2        g0687(.A(new_new_n384_), .B(i_2_), .Y(new_new_n710_));
  NA2        g0688(.A(new_new_n710_), .B(new_new_n709_), .Y(new_new_n711_));
  OAI210     g0689(.A0(new_new_n674_), .A1(new_new_n470_), .B0(new_new_n711_), .Y(new_new_n712_));
  INV        g0690(.A(new_new_n712_), .Y(new_new_n713_));
  AOI210     g0691(.A0(new_new_n713_), .A1(new_new_n708_), .B0(i_13_), .Y(new_new_n714_));
  OR2        g0692(.A(i_11_), .B(i_7_), .Y(new_new_n715_));
  NA3        g0693(.A(new_new_n715_), .B(new_new_n106_), .C(new_new_n138_), .Y(new_new_n716_));
  AOI220     g0694(.A0(new_new_n493_), .A1(new_new_n161_), .B0(new_new_n472_), .B1(new_new_n138_), .Y(new_new_n717_));
  OAI210     g0695(.A0(new_new_n717_), .A1(new_new_n45_), .B0(new_new_n716_), .Y(new_new_n718_));
  NO2        g0696(.A(new_new_n55_), .B(i_12_), .Y(new_new_n719_));
  INV        g0697(.A(new_new_n719_), .Y(new_new_n720_));
  NO2        g0698(.A(new_new_n502_), .B(new_new_n24_), .Y(new_new_n721_));
  AOI220     g0699(.A0(new_new_n721_), .A1(new_new_n689_), .B0(new_new_n249_), .B1(new_new_n131_), .Y(new_new_n722_));
  OAI220     g0700(.A0(new_new_n722_), .A1(new_new_n41_), .B0(new_new_n720_), .B1(new_new_n93_), .Y(new_new_n723_));
  AOI210     g0701(.A0(new_new_n718_), .A1(new_new_n341_), .B0(new_new_n723_), .Y(new_new_n724_));
  INV        g0702(.A(new_new_n115_), .Y(new_new_n725_));
  AOI220     g0703(.A0(new_new_n725_), .A1(new_new_n72_), .B0(new_new_n400_), .B1(new_new_n671_), .Y(new_new_n726_));
  NO2        g0704(.A(new_new_n726_), .B(new_new_n247_), .Y(new_new_n727_));
  AOI210     g0705(.A0(new_new_n470_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n728_));
  NA2        g0706(.A(new_new_n127_), .B(i_13_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n670_), .B(new_new_n115_), .Y(new_new_n730_));
  INV        g0708(.A(new_new_n730_), .Y(new_new_n731_));
  OAI220     g0709(.A0(new_new_n731_), .A1(new_new_n71_), .B0(new_new_n729_), .B1(new_new_n709_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n26_), .B(new_new_n194_), .Y(new_new_n733_));
  NA2        g0711(.A(new_new_n733_), .B(i_7_), .Y(new_new_n734_));
  NO3        g0712(.A(new_new_n502_), .B(new_new_n241_), .C(new_new_n86_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(new_new_n734_), .Y(new_new_n736_));
  AOI220     g0714(.A0(new_new_n400_), .A1(new_new_n671_), .B0(new_new_n92_), .B1(new_new_n102_), .Y(new_new_n737_));
  OAI220     g0715(.A0(new_new_n737_), .A1(new_new_n626_), .B0(new_new_n736_), .B1(new_new_n641_), .Y(new_new_n738_));
  NO3        g0716(.A(new_new_n738_), .B(new_new_n732_), .C(new_new_n727_), .Y(new_new_n739_));
  OR2        g0717(.A(i_11_), .B(i_6_), .Y(new_new_n740_));
  NA3        g0718(.A(new_new_n625_), .B(new_new_n733_), .C(i_7_), .Y(new_new_n741_));
  AOI210     g0719(.A0(new_new_n741_), .A1(new_new_n731_), .B0(new_new_n740_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n429_), .B(new_new_n630_), .C(new_new_n97_), .Y(new_new_n743_));
  NA2        g0721(.A(new_new_n660_), .B(i_13_), .Y(new_new_n744_));
  NAi21      g0722(.An(i_11_), .B(i_12_), .Y(new_new_n745_));
  NOi41      g0723(.An(new_new_n111_), .B(new_new_n745_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n746_));
  NO3        g0724(.A(new_new_n502_), .B(new_new_n606_), .C(new_new_n631_), .Y(new_new_n747_));
  AOI220     g0725(.A0(new_new_n747_), .A1(new_new_n320_), .B0(new_new_n746_), .B1(new_new_n47_), .Y(new_new_n748_));
  NA3        g0726(.A(new_new_n748_), .B(new_new_n744_), .C(new_new_n743_), .Y(new_new_n749_));
  OAI210     g0727(.A0(new_new_n749_), .A1(new_new_n742_), .B0(new_new_n63_), .Y(new_new_n750_));
  NO2        g0728(.A(i_2_), .B(i_12_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n383_), .B(new_new_n751_), .Y(new_new_n752_));
  NA2        g0730(.A(i_8_), .B(new_new_n25_), .Y(new_new_n753_));
  NO3        g0731(.A(new_new_n753_), .B(i_3_), .C(new_new_n625_), .Y(new_new_n754_));
  OAI210     g0732(.A0(new_new_n754_), .A1(new_new_n385_), .B0(new_new_n383_), .Y(new_new_n755_));
  NO2        g0733(.A(new_new_n128_), .B(i_2_), .Y(new_new_n756_));
  NA2        g0734(.A(new_new_n756_), .B(new_new_n654_), .Y(new_new_n757_));
  NA3        g0735(.A(new_new_n757_), .B(new_new_n755_), .C(new_new_n752_), .Y(new_new_n758_));
  NA3        g0736(.A(new_new_n758_), .B(new_new_n46_), .C(new_new_n229_), .Y(new_new_n759_));
  NA4        g0737(.A(new_new_n759_), .B(new_new_n750_), .C(new_new_n739_), .D(new_new_n724_), .Y(new_new_n760_));
  OR4        g0738(.A(new_new_n760_), .B(new_new_n714_), .C(new_new_n701_), .D(new_new_n644_), .Y(men5));
  NA2        g0739(.A(new_new_n686_), .B(new_new_n276_), .Y(new_new_n762_));
  AN2        g0740(.A(new_new_n24_), .B(i_10_), .Y(new_new_n763_));
  NA3        g0741(.A(new_new_n763_), .B(new_new_n751_), .C(new_new_n108_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n626_), .B(i_11_), .Y(new_new_n765_));
  NA2        g0743(.A(new_new_n87_), .B(new_new_n765_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n764_), .C(new_new_n762_), .Y(new_new_n767_));
  NO3        g0745(.A(i_11_), .B(new_new_n241_), .C(i_13_), .Y(new_new_n768_));
  NO2        g0746(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n769_));
  NA2        g0747(.A(i_12_), .B(i_8_), .Y(new_new_n770_));
  OAI210     g0748(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n770_), .Y(new_new_n771_));
  INV        g0749(.A(new_new_n469_), .Y(new_new_n772_));
  AOI220     g0750(.A0(new_new_n326_), .A1(new_new_n601_), .B0(new_new_n771_), .B1(new_new_n769_), .Y(new_new_n773_));
  INV        g0751(.A(new_new_n773_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n774_), .B(new_new_n767_), .Y(new_new_n775_));
  INV        g0753(.A(new_new_n172_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n249_), .Y(new_new_n777_));
  OAI210     g0755(.A0(new_new_n710_), .A1(new_new_n471_), .B0(new_new_n111_), .Y(new_new_n778_));
  AOI210     g0756(.A0(new_new_n778_), .A1(new_new_n777_), .B0(new_new_n776_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n479_), .B(new_new_n26_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n780_), .B(new_new_n440_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n781_), .B(i_2_), .Y(new_new_n782_));
  INV        g0760(.A(new_new_n782_), .Y(new_new_n783_));
  AOI210     g0761(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n436_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n784_), .A1(new_new_n783_), .B0(new_new_n779_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n191_), .B(new_new_n125_), .Y(new_new_n786_));
  OAI210     g0764(.A0(new_new_n786_), .A1(new_new_n769_), .B0(i_2_), .Y(new_new_n787_));
  INV        g0765(.A(new_new_n173_), .Y(new_new_n788_));
  NO3        g0766(.A(new_new_n646_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n789_));
  AOI210     g0767(.A0(new_new_n788_), .A1(new_new_n87_), .B0(new_new_n789_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n790_), .A1(new_new_n787_), .B0(new_new_n194_), .Y(new_new_n791_));
  OA210      g0769(.A0(new_new_n647_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n201_), .B(new_new_n204_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n151_), .B(new_new_n621_), .Y(new_new_n794_));
  AOI210     g0772(.A0(new_new_n794_), .A1(new_new_n793_), .B0(new_new_n388_), .Y(new_new_n795_));
  AOI210     g0773(.A0(new_new_n211_), .A1(new_new_n148_), .B0(new_new_n543_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n796_), .B(new_new_n440_), .Y(new_new_n797_));
  NO2        g0775(.A(new_new_n102_), .B(new_new_n45_), .Y(new_new_n798_));
  INV        g0776(.A(new_new_n308_), .Y(new_new_n799_));
  NA4        g0777(.A(new_new_n799_), .B(new_new_n313_), .C(new_new_n124_), .D(new_new_n43_), .Y(new_new_n800_));
  OAI210     g0778(.A0(new_new_n800_), .A1(new_new_n798_), .B0(new_new_n797_), .Y(new_new_n801_));
  NO4        g0779(.A(new_new_n801_), .B(new_new_n795_), .C(new_new_n792_), .D(new_new_n791_), .Y(new_new_n802_));
  NA2        g0780(.A(new_new_n601_), .B(new_new_n28_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n768_), .B(new_new_n280_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n804_), .B(new_new_n803_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n62_), .B(i_12_), .Y(new_new_n806_));
  NO2        g0784(.A(new_new_n806_), .B(new_new_n126_), .Y(new_new_n807_));
  NO2        g0785(.A(new_new_n807_), .B(new_new_n621_), .Y(new_new_n808_));
  AOI220     g0786(.A0(new_new_n808_), .A1(new_new_n36_), .B0(new_new_n805_), .B1(new_new_n47_), .Y(new_new_n809_));
  NA4        g0787(.A(new_new_n809_), .B(new_new_n802_), .C(new_new_n785_), .D(new_new_n775_), .Y(men6));
  NO3        g0788(.A(new_new_n260_), .B(new_new_n315_), .C(i_1_), .Y(new_new_n811_));
  NO2        g0789(.A(new_new_n186_), .B(new_new_n139_), .Y(new_new_n812_));
  OAI210     g0790(.A0(new_new_n812_), .A1(new_new_n811_), .B0(new_new_n756_), .Y(new_new_n813_));
  NO2        g0791(.A(new_new_n224_), .B(new_new_n512_), .Y(new_new_n814_));
  NO2        g0792(.A(i_11_), .B(i_9_), .Y(new_new_n815_));
  INV        g0793(.A(new_new_n338_), .Y(new_new_n816_));
  AO210      g0794(.A0(new_new_n816_), .A1(new_new_n813_), .B0(i_12_), .Y(new_new_n817_));
  NA2        g0795(.A(new_new_n389_), .B(new_new_n344_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n606_), .B(new_new_n63_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n819_), .B(new_new_n818_), .Y(new_new_n820_));
  INV        g0798(.A(new_new_n198_), .Y(new_new_n821_));
  AOI220     g0799(.A0(new_new_n821_), .A1(new_new_n815_), .B0(new_new_n820_), .B1(new_new_n73_), .Y(new_new_n822_));
  INV        g0800(.A(new_new_n337_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n75_), .B(new_new_n131_), .Y(new_new_n824_));
  INV        g0802(.A(new_new_n124_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n825_), .B(new_new_n47_), .Y(new_new_n826_));
  AOI210     g0804(.A0(new_new_n826_), .A1(new_new_n824_), .B0(new_new_n823_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n256_), .B(i_9_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n828_), .B(new_new_n806_), .Y(new_new_n829_));
  AOI210     g0807(.A0(new_new_n829_), .A1(new_new_n541_), .B0(new_new_n186_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n32_), .B(i_11_), .Y(new_new_n831_));
  NAi32      g0809(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n740_), .B(new_new_n832_), .Y(new_new_n833_));
  OR3        g0811(.A(new_new_n833_), .B(new_new_n830_), .C(new_new_n827_), .Y(new_new_n834_));
  NO2        g0812(.A(new_new_n715_), .B(i_2_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n836_));
  NO2        g0814(.A(new_new_n836_), .B(new_new_n428_), .Y(new_new_n837_));
  NA2        g0815(.A(new_new_n837_), .B(new_new_n835_), .Y(new_new_n838_));
  AO220      g0816(.A0(new_new_n372_), .A1(new_new_n362_), .B0(new_new_n412_), .B1(new_new_n621_), .Y(new_new_n839_));
  NA3        g0817(.A(new_new_n839_), .B(new_new_n261_), .C(i_7_), .Y(new_new_n840_));
  OR2        g0818(.A(new_new_n647_), .B(new_new_n471_), .Y(new_new_n841_));
  NA3        g0819(.A(new_new_n841_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n842_));
  AO210      g0820(.A0(new_new_n519_), .A1(new_new_n772_), .B0(new_new_n36_), .Y(new_new_n843_));
  NA4        g0821(.A(new_new_n843_), .B(new_new_n842_), .C(new_new_n840_), .D(new_new_n838_), .Y(new_new_n844_));
  NO2        g0822(.A(new_new_n659_), .B(i_11_), .Y(new_new_n845_));
  AOI220     g0823(.A0(new_new_n845_), .A1(new_new_n591_), .B0(new_new_n814_), .B1(new_new_n734_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n388_), .B(new_new_n243_), .C(new_new_n147_), .Y(new_new_n847_));
  NA2        g0825(.A(new_new_n412_), .B(new_new_n70_), .Y(new_new_n848_));
  NA4        g0826(.A(new_new_n848_), .B(new_new_n847_), .C(new_new_n846_), .D(new_new_n629_), .Y(new_new_n849_));
  AOI210     g0827(.A0(new_new_n471_), .A1(new_new_n469_), .B0(new_new_n590_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n112_), .B(new_new_n426_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n248_), .B(new_new_n47_), .Y(new_new_n852_));
  INV        g0830(.A(new_new_n612_), .Y(new_new_n853_));
  NA3        g0831(.A(new_new_n853_), .B(new_new_n337_), .C(i_7_), .Y(new_new_n854_));
  NA3        g0832(.A(new_new_n854_), .B(new_new_n851_), .C(new_new_n850_), .Y(new_new_n855_));
  NO4        g0833(.A(new_new_n855_), .B(new_new_n849_), .C(new_new_n844_), .D(new_new_n834_), .Y(new_new_n856_));
  NA4        g0834(.A(new_new_n856_), .B(new_new_n822_), .C(new_new_n817_), .D(new_new_n395_), .Y(men3));
  NA2        g0835(.A(i_12_), .B(i_10_), .Y(new_new_n858_));
  NA2        g0836(.A(i_6_), .B(i_7_), .Y(new_new_n859_));
  NO2        g0837(.A(new_new_n859_), .B(i_0_), .Y(new_new_n860_));
  NO2        g0838(.A(i_11_), .B(new_new_n241_), .Y(new_new_n861_));
  OAI210     g0839(.A0(new_new_n860_), .A1(new_new_n296_), .B0(new_new_n861_), .Y(new_new_n862_));
  NO2        g0840(.A(new_new_n862_), .B(new_new_n194_), .Y(new_new_n863_));
  NO3        g0841(.A(new_new_n475_), .B(new_new_n90_), .C(new_new_n45_), .Y(new_new_n864_));
  OA210      g0842(.A0(new_new_n864_), .A1(new_new_n863_), .B0(new_new_n175_), .Y(new_new_n865_));
  NA3        g0843(.A(new_new_n847_), .B(new_new_n629_), .C(new_new_n387_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n866_), .B(new_new_n40_), .Y(new_new_n867_));
  NOi21      g0845(.An(new_new_n96_), .B(new_new_n781_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n429_), .B(new_new_n46_), .Y(new_new_n869_));
  INV        g0847(.A(new_new_n868_), .Y(new_new_n870_));
  AOI210     g0848(.A0(new_new_n870_), .A1(new_new_n867_), .B0(new_new_n49_), .Y(new_new_n871_));
  NO4        g0849(.A(new_new_n392_), .B(new_new_n398_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n186_), .B(new_new_n599_), .Y(new_new_n873_));
  NOi21      g0851(.An(new_new_n873_), .B(new_new_n872_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n728_), .B(new_new_n695_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n342_), .B(new_new_n460_), .Y(new_new_n876_));
  OAI220     g0854(.A0(new_new_n876_), .A1(new_new_n875_), .B0(new_new_n874_), .B1(new_new_n63_), .Y(new_new_n877_));
  NOi21      g0855(.An(i_5_), .B(i_9_), .Y(new_new_n878_));
  NA2        g0856(.A(new_new_n878_), .B(new_new_n468_), .Y(new_new_n879_));
  BUFFER     g0857(.A(new_new_n274_), .Y(new_new_n880_));
  AOI210     g0858(.A0(new_new_n880_), .A1(new_new_n499_), .B0(new_new_n704_), .Y(new_new_n881_));
  NO2        g0859(.A(new_new_n176_), .B(new_new_n148_), .Y(new_new_n882_));
  NO2        g0860(.A(new_new_n881_), .B(new_new_n879_), .Y(new_new_n883_));
  NO4        g0861(.A(new_new_n883_), .B(new_new_n877_), .C(new_new_n871_), .D(new_new_n865_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n186_), .B(new_new_n24_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n320_), .B(new_new_n129_), .Y(new_new_n886_));
  NAi21      g0864(.An(new_new_n162_), .B(new_new_n460_), .Y(new_new_n887_));
  OAI220     g0865(.A0(new_new_n887_), .A1(new_new_n852_), .B0(new_new_n886_), .B1(new_new_n418_), .Y(new_new_n888_));
  INV        g0866(.A(new_new_n888_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n404_), .B(new_new_n300_), .Y(new_new_n890_));
  NA2        g0868(.A(new_new_n890_), .B(new_new_n730_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n600_), .B(i_0_), .Y(new_new_n892_));
  NO4        g0870(.A(new_new_n611_), .B(new_new_n218_), .C(new_new_n436_), .D(new_new_n428_), .Y(new_new_n893_));
  INV        g0871(.A(new_new_n497_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n768_), .B(new_new_n338_), .Y(new_new_n895_));
  INV        g0873(.A(new_new_n58_), .Y(new_new_n896_));
  OAI220     g0874(.A0(new_new_n896_), .A1(new_new_n895_), .B0(new_new_n681_), .B1(new_new_n564_), .Y(new_new_n897_));
  NO2        g0875(.A(new_new_n258_), .B(new_new_n153_), .Y(new_new_n898_));
  NA2        g0876(.A(i_0_), .B(i_10_), .Y(new_new_n899_));
  AN2        g0877(.A(new_new_n898_), .B(i_6_), .Y(new_new_n900_));
  AOI220     g0878(.A0(new_new_n342_), .A1(new_new_n98_), .B0(new_new_n186_), .B1(new_new_n84_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n595_), .B(i_4_), .Y(new_new_n902_));
  NO2        g0880(.A(new_new_n902_), .B(new_new_n901_), .Y(new_new_n903_));
  NO3        g0881(.A(new_new_n903_), .B(new_new_n900_), .C(new_new_n897_), .Y(new_new_n904_));
  NA3        g0882(.A(new_new_n904_), .B(new_new_n891_), .C(new_new_n889_), .Y(new_new_n905_));
  NA2        g0883(.A(i_11_), .B(i_9_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n409_), .B(new_new_n180_), .Y(new_new_n907_));
  NA2        g0885(.A(new_new_n907_), .B(new_new_n160_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n906_), .B(new_new_n73_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n176_), .B(i_0_), .Y(new_new_n910_));
  INV        g0888(.A(new_new_n910_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n497_), .B(new_new_n235_), .Y(new_new_n912_));
  AOI210     g0890(.A0(new_new_n386_), .A1(new_new_n42_), .B0(new_new_n425_), .Y(new_new_n913_));
  OAI220     g0891(.A0(new_new_n913_), .A1(new_new_n879_), .B0(new_new_n912_), .B1(new_new_n911_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n914_), .B(new_new_n908_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n680_), .B(new_new_n121_), .Y(new_new_n916_));
  NO2        g0894(.A(i_6_), .B(new_new_n916_), .Y(new_new_n917_));
  AOI210     g0895(.A0(new_new_n470_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n172_), .B(new_new_n103_), .Y(new_new_n919_));
  NOi32      g0897(.An(new_new_n918_), .Bn(new_new_n189_), .C(new_new_n919_), .Y(new_new_n920_));
  NA2        g0898(.A(new_new_n630_), .B(new_new_n338_), .Y(new_new_n921_));
  NO2        g0899(.A(new_new_n921_), .B(new_new_n869_), .Y(new_new_n922_));
  NO3        g0900(.A(new_new_n922_), .B(new_new_n920_), .C(new_new_n917_), .Y(new_new_n923_));
  NOi21      g0901(.An(i_7_), .B(i_5_), .Y(new_new_n924_));
  OR2        g0902(.A(new_new_n919_), .B(new_new_n541_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n421_), .B(new_new_n375_), .C(new_new_n371_), .Y(new_new_n926_));
  NO2        g0904(.A(new_new_n268_), .B(new_new_n327_), .Y(new_new_n927_));
  NO2        g0905(.A(new_new_n745_), .B(new_new_n263_), .Y(new_new_n928_));
  AOI210     g0906(.A0(new_new_n928_), .A1(new_new_n927_), .B0(new_new_n926_), .Y(new_new_n929_));
  NA4        g0907(.A(new_new_n929_), .B(new_new_n925_), .C(new_new_n923_), .D(new_new_n915_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n885_), .B(new_new_n244_), .Y(new_new_n931_));
  AN2        g0909(.A(new_new_n341_), .B(new_new_n338_), .Y(new_new_n932_));
  AN2        g0910(.A(new_new_n932_), .B(new_new_n882_), .Y(new_new_n933_));
  OAI210     g0911(.A0(new_new_n933_), .A1(new_new_n931_), .B0(i_10_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n858_), .B(new_new_n326_), .Y(new_new_n935_));
  NA2        g0913(.A(new_new_n935_), .B(new_new_n909_), .Y(new_new_n936_));
  NA3        g0914(.A(new_new_n496_), .B(new_new_n429_), .C(new_new_n46_), .Y(new_new_n937_));
  OAI210     g0915(.A0(new_new_n887_), .A1(new_new_n894_), .B0(new_new_n937_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n261_), .B(new_new_n47_), .Y(new_new_n939_));
  NA2        g0917(.A(new_new_n909_), .B(new_new_n313_), .Y(new_new_n940_));
  OAI210     g0918(.A0(new_new_n939_), .A1(new_new_n188_), .B0(new_new_n940_), .Y(new_new_n941_));
  AOI220     g0919(.A0(new_new_n941_), .A1(new_new_n497_), .B0(new_new_n938_), .B1(new_new_n73_), .Y(new_new_n942_));
  NA3        g0920(.A(new_new_n836_), .B(new_new_n397_), .C(new_new_n659_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n943_), .B(new_new_n48_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n611_), .B(new_new_n370_), .C(new_new_n24_), .Y(new_new_n945_));
  AOI210     g0923(.A0(new_new_n721_), .A1(new_new_n574_), .B0(new_new_n945_), .Y(new_new_n946_));
  NAi21      g0924(.An(i_9_), .B(i_5_), .Y(new_new_n947_));
  NO2        g0925(.A(new_new_n947_), .B(new_new_n421_), .Y(new_new_n948_));
  NO2        g0926(.A(new_new_n624_), .B(new_new_n105_), .Y(new_new_n949_));
  AOI220     g0927(.A0(new_new_n949_), .A1(i_0_), .B0(new_new_n948_), .B1(new_new_n647_), .Y(new_new_n950_));
  OAI220     g0928(.A0(new_new_n950_), .A1(new_new_n86_), .B0(new_new_n946_), .B1(new_new_n173_), .Y(new_new_n951_));
  NO3        g0929(.A(new_new_n951_), .B(new_new_n944_), .C(new_new_n545_), .Y(new_new_n952_));
  NA4        g0930(.A(new_new_n952_), .B(new_new_n942_), .C(new_new_n936_), .D(new_new_n934_), .Y(new_new_n953_));
  NO3        g0931(.A(new_new_n953_), .B(new_new_n930_), .C(new_new_n905_), .Y(new_new_n954_));
  NA2        g0932(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n899_), .B(new_new_n955_), .Y(new_new_n956_));
  NO3        g0934(.A(new_new_n105_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n957_));
  AN2        g0935(.A(new_new_n957_), .B(new_new_n956_), .Y(new_new_n958_));
  AOI210     g0936(.A0(new_new_n819_), .A1(new_new_n702_), .B0(new_new_n919_), .Y(new_new_n959_));
  AOI210     g0937(.A0(new_new_n958_), .A1(new_new_n359_), .B0(new_new_n959_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n756_), .B(new_new_n146_), .Y(new_new_n961_));
  INV        g0939(.A(new_new_n961_), .Y(new_new_n962_));
  NA3        g0940(.A(new_new_n962_), .B(new_new_n695_), .C(new_new_n73_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n860_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n964_));
  NA2        g0942(.A(new_new_n861_), .B(i_9_), .Y(new_new_n965_));
  AOI210     g0943(.A0(new_new_n964_), .A1(new_new_n524_), .B0(new_new_n965_), .Y(new_new_n966_));
  OAI210     g0944(.A0(new_new_n248_), .A1(i_9_), .B0(new_new_n234_), .Y(new_new_n967_));
  AOI210     g0945(.A0(new_new_n967_), .A1(new_new_n892_), .B0(new_new_n153_), .Y(new_new_n968_));
  NO2        g0946(.A(new_new_n968_), .B(new_new_n966_), .Y(new_new_n969_));
  NA3        g0947(.A(new_new_n969_), .B(new_new_n963_), .C(new_new_n960_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n932_), .B(new_new_n388_), .Y(new_new_n971_));
  AOI210     g0949(.A0(new_new_n307_), .A1(new_new_n162_), .B0(new_new_n971_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n973_));
  NA2        g0951(.A(i_5_), .B(new_new_n513_), .Y(new_new_n974_));
  AOI210     g0952(.A0(new_new_n973_), .A1(new_new_n162_), .B0(new_new_n974_), .Y(new_new_n975_));
  NO2        g0953(.A(new_new_n975_), .B(new_new_n972_), .Y(new_new_n976_));
  NO3        g0954(.A(new_new_n899_), .B(new_new_n878_), .C(new_new_n191_), .Y(new_new_n977_));
  AOI220     g0955(.A0(new_new_n977_), .A1(i_11_), .B0(new_new_n596_), .B1(new_new_n75_), .Y(new_new_n978_));
  NO3        g0956(.A(new_new_n212_), .B(new_new_n398_), .C(i_0_), .Y(new_new_n979_));
  OAI210     g0957(.A0(new_new_n979_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n980_));
  INV        g0958(.A(new_new_n221_), .Y(new_new_n981_));
  OAI220     g0959(.A0(new_new_n557_), .A1(new_new_n139_), .B0(new_new_n664_), .B1(new_new_n641_), .Y(new_new_n982_));
  NA3        g0960(.A(new_new_n982_), .B(new_new_n413_), .C(new_new_n981_), .Y(new_new_n983_));
  NA4        g0961(.A(new_new_n983_), .B(new_new_n980_), .C(new_new_n978_), .D(new_new_n976_), .Y(new_new_n984_));
  INV        g0962(.A(new_new_n109_), .Y(new_new_n985_));
  AOI220     g0963(.A0(new_new_n924_), .A1(new_new_n513_), .B0(new_new_n860_), .B1(new_new_n163_), .Y(new_new_n986_));
  NA2        g0964(.A(new_new_n362_), .B(new_new_n177_), .Y(new_new_n987_));
  OA220      g0965(.A0(new_new_n987_), .A1(new_new_n986_), .B0(new_new_n985_), .B1(i_5_), .Y(new_new_n988_));
  NA3        g0966(.A(new_new_n638_), .B(new_new_n186_), .C(new_new_n84_), .Y(new_new_n989_));
  INV        g0967(.A(new_new_n989_), .Y(new_new_n990_));
  NO3        g0968(.A(new_new_n869_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n991_));
  NA2        g0969(.A(new_new_n518_), .B(new_new_n494_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n992_), .B(new_new_n991_), .C(new_new_n990_), .Y(new_new_n993_));
  NA3        g0971(.A(new_new_n404_), .B(new_new_n343_), .C(new_new_n225_), .Y(new_new_n994_));
  INV        g0972(.A(new_new_n994_), .Y(new_new_n995_));
  NOi31      g0973(.An(new_new_n403_), .B(new_new_n955_), .C(new_new_n244_), .Y(new_new_n996_));
  NO3        g0974(.A(new_new_n906_), .B(new_new_n221_), .C(new_new_n191_), .Y(new_new_n997_));
  NO3        g0975(.A(new_new_n997_), .B(new_new_n996_), .C(new_new_n995_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n998_), .B(new_new_n993_), .C(new_new_n988_), .Y(new_new_n999_));
  INV        g0977(.A(new_new_n640_), .Y(new_new_n1000_));
  NO3        g0978(.A(new_new_n1000_), .B(new_new_n586_), .C(new_new_n356_), .Y(new_new_n1001_));
  NO2        g0979(.A(new_new_n86_), .B(i_5_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n861_), .B(new_new_n110_), .C(new_new_n124_), .Y(new_new_n1003_));
  INV        g0981(.A(new_new_n1003_), .Y(new_new_n1004_));
  AOI210     g0982(.A0(new_new_n1004_), .A1(new_new_n1002_), .B0(new_new_n1001_), .Y(new_new_n1005_));
  AN2        g0983(.A(new_new_n899_), .B(new_new_n153_), .Y(new_new_n1006_));
  NO4        g0984(.A(new_new_n1006_), .B(i_12_), .C(new_new_n668_), .D(new_new_n131_), .Y(new_new_n1007_));
  NA2        g0985(.A(new_new_n1007_), .B(new_new_n221_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n98_), .B(new_new_n599_), .C(i_11_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n1009_), .B(new_new_n155_), .Y(new_new_n1010_));
  INV        g0988(.A(new_new_n1010_), .Y(new_new_n1011_));
  NA3        g0989(.A(new_new_n1011_), .B(new_new_n1008_), .C(new_new_n1005_), .Y(new_new_n1012_));
  NO4        g0990(.A(new_new_n1012_), .B(new_new_n999_), .C(new_new_n984_), .D(new_new_n970_), .Y(new_new_n1013_));
  OAI210     g0991(.A0(new_new_n835_), .A1(new_new_n831_), .B0(new_new_n37_), .Y(new_new_n1014_));
  NA3        g0992(.A(new_new_n918_), .B(new_new_n383_), .C(i_5_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n1015_), .B(new_new_n1014_), .C(new_new_n636_), .Y(new_new_n1016_));
  NA2        g0994(.A(new_new_n1016_), .B(new_new_n209_), .Y(new_new_n1017_));
  NA2        g0995(.A(new_new_n187_), .B(new_new_n189_), .Y(new_new_n1018_));
  AO210      g0996(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1018_), .Y(new_new_n1019_));
  OAI210     g0997(.A0(new_new_n640_), .A1(new_new_n638_), .B0(new_new_n326_), .Y(new_new_n1020_));
  NAi31      g0998(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1021_));
  NO2        g0999(.A(new_new_n70_), .B(new_new_n1021_), .Y(new_new_n1022_));
  NO2        g1000(.A(new_new_n1022_), .B(new_new_n665_), .Y(new_new_n1023_));
  NA3        g1001(.A(new_new_n1023_), .B(new_new_n1020_), .C(new_new_n1019_), .Y(new_new_n1024_));
  NO2        g1002(.A(new_new_n483_), .B(new_new_n274_), .Y(new_new_n1025_));
  NO4        g1003(.A(new_new_n237_), .B(new_new_n145_), .C(new_new_n699_), .D(new_new_n37_), .Y(new_new_n1026_));
  NO3        g1004(.A(new_new_n1026_), .B(new_new_n1025_), .C(new_new_n893_), .Y(new_new_n1027_));
  OAI210     g1005(.A0(new_new_n1009_), .A1(new_new_n148_), .B0(new_new_n1027_), .Y(new_new_n1028_));
  AOI210     g1006(.A0(new_new_n1024_), .A1(new_new_n49_), .B0(new_new_n1028_), .Y(new_new_n1029_));
  AOI210     g1007(.A0(new_new_n1029_), .A1(new_new_n1017_), .B0(new_new_n73_), .Y(new_new_n1030_));
  NO2        g1008(.A(new_new_n593_), .B(new_new_n394_), .Y(new_new_n1031_));
  NO2        g1009(.A(new_new_n1031_), .B(new_new_n776_), .Y(new_new_n1032_));
  INV        g1010(.A(new_new_n76_), .Y(new_new_n1033_));
  NO2        g1011(.A(new_new_n1033_), .B(new_new_n699_), .Y(new_new_n1034_));
  NA2        g1012(.A(new_new_n268_), .B(new_new_n57_), .Y(new_new_n1035_));
  AOI220     g1013(.A0(new_new_n1035_), .A1(new_new_n76_), .B0(new_new_n357_), .B1(new_new_n260_), .Y(new_new_n1036_));
  NO2        g1014(.A(new_new_n1036_), .B(new_new_n241_), .Y(new_new_n1037_));
  NA3        g1015(.A(new_new_n96_), .B(new_new_n315_), .C(new_new_n31_), .Y(new_new_n1038_));
  INV        g1016(.A(new_new_n1038_), .Y(new_new_n1039_));
  NO3        g1017(.A(new_new_n1039_), .B(new_new_n1037_), .C(new_new_n1034_), .Y(new_new_n1040_));
  NA2        g1018(.A(new_new_n158_), .B(new_new_n87_), .Y(new_new_n1041_));
  NA3        g1019(.A(new_new_n780_), .B(new_new_n296_), .C(new_new_n80_), .Y(new_new_n1042_));
  AOI210     g1020(.A0(new_new_n1042_), .A1(new_new_n1041_), .B0(i_11_), .Y(new_new_n1043_));
  NA2        g1021(.A(new_new_n631_), .B(new_new_n218_), .Y(new_new_n1044_));
  OAI210     g1022(.A0(new_new_n1044_), .A1(new_new_n918_), .B0(new_new_n209_), .Y(new_new_n1045_));
  NA2        g1023(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n1045_), .B(new_new_n1046_), .Y(new_new_n1047_));
  NO4        g1025(.A(new_new_n947_), .B(new_new_n501_), .C(new_new_n257_), .D(new_new_n256_), .Y(new_new_n1048_));
  NO2        g1026(.A(new_new_n1048_), .B(new_new_n590_), .Y(new_new_n1049_));
  INV        g1027(.A(new_new_n376_), .Y(new_new_n1050_));
  AOI210     g1028(.A0(new_new_n1050_), .A1(new_new_n1049_), .B0(new_new_n41_), .Y(new_new_n1051_));
  NO3        g1029(.A(new_new_n1051_), .B(new_new_n1047_), .C(new_new_n1043_), .Y(new_new_n1052_));
  OAI210     g1030(.A0(new_new_n1040_), .A1(i_4_), .B0(new_new_n1052_), .Y(new_new_n1053_));
  NO3        g1031(.A(new_new_n1053_), .B(new_new_n1032_), .C(new_new_n1030_), .Y(new_new_n1054_));
  NA4        g1032(.A(new_new_n1054_), .B(new_new_n1013_), .C(new_new_n954_), .D(new_new_n884_), .Y(men4));
  INV        g1033(.A(i_2_), .Y(new_new_n1058_));
endmodule


