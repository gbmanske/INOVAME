//Benchmark atmr_intb_466_0.5

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n88_, ori_ori_n92_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n146_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n156_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n478_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o00(.A(x11), .Y(ori_ori_n23_));
  NA2        o01(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o02(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o03(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o04(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o05(.A(x02), .Y(ori_ori_n28_));
  INV        o06(.A(x10), .Y(ori_ori_n29_));
  NA2        o07(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o08(.A(x03), .Y(ori_ori_n31_));
  NA2        o09(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o10(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o11(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o12(.A(x04), .Y(ori_ori_n35_));
  INV        o13(.A(x08), .Y(ori_ori_n36_));
  NA2        o14(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o15(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o16(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o17(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o18(.A(x05), .Y(ori_ori_n41_));
  NO2        o19(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o20(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o21(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o22(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o23(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o24(.A(x01), .Y(ori_ori_n47_));
  INV        o25(.A(x06), .Y(ori_ori_n48_));
  INV        o26(.A(x09), .Y(ori_ori_n49_));
  NO2        o27(.A(x10), .B(x02), .Y(ori_ori_n50_));
  INV        o28(.A(x00), .Y(ori_ori_n51_));
  INV        o29(.A(x07), .Y(ori_ori_n52_));
  NO2        o30(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n53_));
  NO2        o31(.A(x08), .B(x01), .Y(ori_ori_n54_));
  OAI210     o32(.A0(ori_ori_n54_), .A1(ori_ori_n53_), .B0(ori_ori_n35_), .Y(ori_ori_n55_));
  INV        o33(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NA2        o34(.A(x11), .B(x00), .Y(ori_ori_n57_));
  NO2        o35(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n58_));
  NOi21      o36(.An(ori_ori_n57_), .B(ori_ori_n58_), .Y(ori_ori_n59_));
  INV        o37(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NO2        o38(.A(ori_ori_n60_), .B(x07), .Y(ori_ori_n61_));
  INV        o39(.A(ori_ori_n61_), .Y(ori01));
  INV        o40(.A(x12), .Y(ori_ori_n63_));
  NA2        o41(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n64_));
  NA2        o42(.A(x10), .B(ori_ori_n51_), .Y(ori_ori_n65_));
  NA2        o43(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  NO2        o44(.A(x09), .B(x05), .Y(ori_ori_n67_));
  NA2        o45(.A(ori_ori_n67_), .B(ori_ori_n47_), .Y(ori_ori_n68_));
  NO2        o46(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n69_));
  NA2        o47(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n70_));
  NO2        o48(.A(ori_ori_n49_), .B(x03), .Y(ori_ori_n71_));
  NA2        o49(.A(x13), .B(ori_ori_n63_), .Y(ori_ori_n72_));
  INV        o50(.A(ori_ori_n59_), .Y(ori_ori_n73_));
  NO2        o51(.A(ori_ori_n73_), .B(x07), .Y(ori_ori_n74_));
  INV        o52(.A(ori_ori_n74_), .Y(ori_ori_n75_));
  OAI210     o53(.A0(ori_ori_n92_), .A1(ori_ori_n52_), .B0(ori_ori_n75_), .Y(ori02));
  INV        o54(.A(ori_ori_n66_), .Y(ori_ori_n77_));
  NA2        o55(.A(ori_ori_n77_), .B(ori_ori_n48_), .Y(ori_ori_n78_));
  NO2        o56(.A(ori_ori_n69_), .B(ori_ori_n50_), .Y(ori_ori_n79_));
  INV        o57(.A(ori_ori_n79_), .Y(ori_ori_n80_));
  NA2        o58(.A(ori_ori_n80_), .B(x06), .Y(ori_ori_n81_));
  NA2        o59(.A(ori_ori_n81_), .B(ori_ori_n78_), .Y(ori_ori_n82_));
  INV        o60(.A(ori_ori_n82_), .Y(ori03));
  OR2        o61(.A(ori_ori_n42_), .B(ori_ori_n71_), .Y(ori_ori_n84_));
  AOI210     o62(.A0(ori_ori_n35_), .A1(ori_ori_n63_), .B0(ori_ori_n84_), .Y(ori_ori_n85_));
  NA2        o63(.A(ori_ori_n85_), .B(x05), .Y(ori_ori_n86_));
  NA2        o64(.A(ori_ori_n68_), .B(ori_ori_n86_), .Y(ori04));
  NO2        o65(.A(ori_ori_n56_), .B(ori_ori_n39_), .Y(ori_ori_n88_));
  XO2        o66(.A(ori_ori_n88_), .B(ori_ori_n72_), .Y(ori05));
  INV        o67(.A(ori_ori_n70_), .Y(ori_ori_n92_));
  ZERO       o68(.Y(ori06));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  INV        m017(.A(x05), .Y(mai_mai_n40_));
  NO2        m018(.A(x09), .B(x02), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n41_), .B(mai_mai_n40_), .Y(mai_mai_n42_));
  NA2        m020(.A(mai_mai_n42_), .B(x03), .Y(mai_mai_n43_));
  INV        m021(.A(mai_mai_n43_), .Y(mai_mai_n44_));
  NO3        m022(.A(mai_mai_n44_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m023(.A(x01), .Y(mai_mai_n46_));
  INV        m024(.A(x06), .Y(mai_mai_n47_));
  NO2        m025(.A(x02), .B(x11), .Y(mai_mai_n48_));
  INV        m026(.A(x09), .Y(mai_mai_n49_));
  NO2        m027(.A(x10), .B(x02), .Y(mai_mai_n50_));
  NA2        m028(.A(mai_mai_n48_), .B(mai_mai_n46_), .Y(mai_mai_n51_));
  NOi21      m029(.An(x01), .B(x09), .Y(mai_mai_n52_));
  INV        m030(.A(x00), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n49_), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  NO2        m032(.A(mai_mai_n54_), .B(mai_mai_n52_), .Y(mai_mai_n55_));
  NA2        m033(.A(x09), .B(mai_mai_n53_), .Y(mai_mai_n56_));
  INV        m034(.A(x07), .Y(mai_mai_n57_));
  OAI210     m035(.A0(mai_mai_n30_), .A1(x11), .B0(x07), .Y(mai_mai_n58_));
  AOI220     m036(.A0(mai_mai_n58_), .A1(mai_mai_n55_), .B0(mai_mai_n55_), .B1(mai_mai_n31_), .Y(mai_mai_n59_));
  AOI210     m037(.A0(mai_mai_n59_), .A1(mai_mai_n51_), .B0(x05), .Y(mai_mai_n60_));
  NA2        m038(.A(x11), .B(x03), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n24_), .Y(mai_mai_n62_));
  NO2        m040(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n63_));
  NO2        m041(.A(x08), .B(x01), .Y(mai_mai_n64_));
  OAI210     m042(.A0(mai_mai_n64_), .A1(mai_mai_n63_), .B0(mai_mai_n35_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n49_), .B(mai_mai_n36_), .Y(mai_mai_n66_));
  NO2        m044(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n67_));
  AN2        m045(.A(mai_mai_n67_), .B(mai_mai_n61_), .Y(mai_mai_n68_));
  INV        m046(.A(mai_mai_n65_), .Y(mai_mai_n69_));
  NA2        m047(.A(x11), .B(x00), .Y(mai_mai_n70_));
  NO2        m048(.A(x11), .B(mai_mai_n46_), .Y(mai_mai_n71_));
  NOi21      m049(.An(mai_mai_n70_), .B(mai_mai_n71_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n69_), .B(mai_mai_n72_), .Y(mai_mai_n73_));
  NOi21      m051(.An(x01), .B(x10), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n29_), .B(mai_mai_n53_), .Y(mai_mai_n75_));
  NO3        m053(.A(mai_mai_n75_), .B(mai_mai_n74_), .C(x06), .Y(mai_mai_n76_));
  NA2        m054(.A(mai_mai_n76_), .B(mai_mai_n27_), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n73_), .A1(x07), .B0(mai_mai_n77_), .Y(mai_mai_n78_));
  NO3        m056(.A(mai_mai_n78_), .B(mai_mai_n68_), .C(mai_mai_n60_), .Y(mai01));
  INV        m057(.A(x12), .Y(mai_mai_n80_));
  NA2        m058(.A(mai_mai_n29_), .B(mai_mai_n46_), .Y(mai_mai_n81_));
  NA2        m059(.A(x10), .B(mai_mai_n53_), .Y(mai_mai_n82_));
  NA2        m060(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n49_), .B(x05), .Y(mai_mai_n84_));
  NO2        m062(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n85_));
  NO2        m063(.A(mai_mai_n49_), .B(mai_mai_n40_), .Y(mai_mai_n86_));
  NA2        m064(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n87_));
  NO2        m065(.A(x09), .B(x05), .Y(mai_mai_n88_));
  NA2        m066(.A(mai_mai_n88_), .B(mai_mai_n46_), .Y(mai_mai_n89_));
  NO2        m067(.A(x03), .B(x02), .Y(mai_mai_n90_));
  OR2        m068(.A(x02), .B(x11), .Y(mai_mai_n91_));
  OAI210     m069(.A0(x03), .A1(mai_mai_n23_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NO2        m070(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n94_), .B(x12), .Y(mai_mai_n95_));
  INV        m073(.A(mai_mai_n95_), .Y(mai_mai_n96_));
  AOI210     m074(.A0(mai_mai_n92_), .A1(mai_mai_n80_), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  AOI210     m075(.A0(x06), .A1(x02), .B0(x12), .Y(mai_mai_n98_));
  NO2        m076(.A(mai_mai_n53_), .B(mai_mai_n23_), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n98_), .B(mai_mai_n99_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n49_), .B(x03), .Y(mai_mai_n101_));
  INV        m079(.A(mai_mai_n71_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(x12), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n49_), .B(mai_mai_n36_), .Y(mai_mai_n104_));
  NA2        m082(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n105_));
  NA2        m083(.A(x13), .B(mai_mai_n80_), .Y(mai_mai_n106_));
  NA2        m084(.A(x12), .B(mai_mai_n72_), .Y(mai_mai_n107_));
  INV        m085(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n103_), .B(mai_mai_n108_), .Y(mai_mai_n109_));
  AOI210     m087(.A0(mai_mai_n109_), .A1(mai_mai_n100_), .B0(x07), .Y(mai_mai_n110_));
  NA2        m088(.A(mai_mai_n49_), .B(mai_mai_n40_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n111_), .B(x01), .Y(mai_mai_n112_));
  NO3        m090(.A(mai_mai_n70_), .B(x12), .C(x03), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n113_), .B(mai_mai_n110_), .Y(mai_mai_n114_));
  OAI210     m092(.A0(mai_mai_n97_), .A1(mai_mai_n57_), .B0(mai_mai_n114_), .Y(mai02));
  NO2        m093(.A(mai_mai_n32_), .B(mai_mai_n47_), .Y(mai_mai_n116_));
  NO2        m094(.A(x02), .B(mai_mai_n87_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n105_), .B(mai_mai_n46_), .Y(mai_mai_n118_));
  INV        m096(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  INV        m097(.A(x06), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n120_), .B(mai_mai_n75_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(mai_mai_n119_), .Y(mai_mai_n122_));
  NO3        m100(.A(mai_mai_n122_), .B(mai_mai_n117_), .C(mai_mai_n116_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n86_), .B(x03), .Y(mai_mai_n124_));
  NA2        m102(.A(x12), .B(mai_mai_n83_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(mai_mai_n47_), .Y(mai_mai_n126_));
  INV        m104(.A(mai_mai_n104_), .Y(mai_mai_n127_));
  NO2        m105(.A(mai_mai_n93_), .B(mai_mai_n50_), .Y(mai_mai_n128_));
  NA2        m106(.A(x12), .B(mai_mai_n128_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n129_), .B(x06), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n126_), .Y(mai_mai_n131_));
  OAI210     m109(.A0(mai_mai_n123_), .A1(x12), .B0(mai_mai_n131_), .Y(mai03));
  OR2        m110(.A(mai_mai_n41_), .B(mai_mai_n101_), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n80_), .B(mai_mai_n133_), .Y(mai_mai_n134_));
  AO210      m112(.A0(mai_mai_n127_), .A1(mai_mai_n66_), .B0(x12), .Y(mai_mai_n135_));
  NA2        m113(.A(mai_mai_n156_), .B(mai_mai_n90_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n136_), .B(mai_mai_n135_), .Y(mai_mai_n137_));
  OAI210     m115(.A0(mai_mai_n137_), .A1(mai_mai_n134_), .B0(x05), .Y(mai_mai_n138_));
  INV        m116(.A(x05), .Y(mai_mai_n139_));
  NO2        m117(.A(x04), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m118(.A(x05), .B(mai_mai_n55_), .Y(mai_mai_n141_));
  OAI210     m119(.A0(mai_mai_n141_), .A1(mai_mai_n140_), .B0(mai_mai_n80_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n80_), .B(mai_mai_n89_), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n85_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  NA3        m122(.A(mai_mai_n144_), .B(mai_mai_n142_), .C(mai_mai_n138_), .Y(mai04));
  NO2        m123(.A(mai_mai_n69_), .B(mai_mai_n39_), .Y(mai_mai_n146_));
  XO2        m124(.A(mai_mai_n146_), .B(mai_mai_n106_), .Y(mai05));
  NOi21      m125(.An(mai_mai_n124_), .B(mai_mai_n85_), .Y(mai_mai_n148_));
  NO2        m126(.A(mai_mai_n84_), .B(mai_mai_n28_), .Y(mai_mai_n149_));
  NO2        m127(.A(mai_mai_n149_), .B(mai_mai_n112_), .Y(mai_mai_n150_));
  NA3        m128(.A(mai_mai_n150_), .B(mai_mai_n148_), .C(x12), .Y(mai_mai_n151_));
  NA2        m129(.A(x14), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  INV        m130(.A(mai_mai_n152_), .Y(mai06));
  INV        m131(.A(x12), .Y(mai_mai_n156_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men05));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men05), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  INV        u030(.A(men_men_n52_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n54_), .B(men_men_n50_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI220     u039(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n61_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  OAI220     u042(.A0(men_men_n64_), .A1(men_men_n58_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  NO2        u044(.A(men_men_n30_), .B(x11), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  NA3        u050(.A(men_men_n72_), .B(men_men_n71_), .C(men_men_n28_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n74_));
  NA2        u052(.A(men_men_n73_), .B(x03), .Y(men_men_n75_));
  NOi31      u053(.An(x08), .B(x04), .C(x00), .Y(men_men_n76_));
  NO2        u054(.A(x10), .B(x09), .Y(men_men_n77_));
  NO2        u055(.A(men_men_n478_), .B(men_men_n24_), .Y(men_men_n78_));
  NO2        u056(.A(x09), .B(men_men_n41_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n79_), .B(men_men_n36_), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n79_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n81_));
  AOI210     u059(.A0(men_men_n80_), .A1(men_men_n48_), .B0(men_men_n81_), .Y(men_men_n82_));
  NO2        u060(.A(men_men_n36_), .B(x00), .Y(men_men_n83_));
  NO2        u061(.A(x08), .B(x01), .Y(men_men_n84_));
  OAI210     u062(.A0(men_men_n84_), .A1(men_men_n83_), .B0(men_men_n35_), .Y(men_men_n85_));
  NA2        u063(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n86_));
  NO3        u064(.A(men_men_n85_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n87_));
  AN2        u065(.A(men_men_n87_), .B(men_men_n75_), .Y(men_men_n88_));
  NO2        u066(.A(x06), .B(x05), .Y(men_men_n89_));
  NA2        u067(.A(x11), .B(x00), .Y(men_men_n90_));
  NO2        u068(.A(x11), .B(men_men_n47_), .Y(men_men_n91_));
  NOi21      u069(.An(men_men_n90_), .B(men_men_n91_), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n89_), .B(men_men_n92_), .Y(men_men_n93_));
  NOi21      u071(.An(x01), .B(x10), .Y(men_men_n94_));
  NO2        u072(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n94_), .C(x06), .Y(men_men_n96_));
  NA2        u074(.A(men_men_n96_), .B(men_men_n27_), .Y(men_men_n97_));
  OAI210     u075(.A0(men_men_n93_), .A1(x07), .B0(men_men_n97_), .Y(men_men_n98_));
  NO3        u076(.A(men_men_n98_), .B(men_men_n88_), .C(men_men_n69_), .Y(men01));
  INV        u077(.A(x12), .Y(men_men_n100_));
  INV        u078(.A(x13), .Y(men_men_n101_));
  NA2        u079(.A(men_men_n89_), .B(x01), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n102_), .B(men_men_n70_), .Y(men_men_n103_));
  NA2        u081(.A(x08), .B(x04), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n57_), .Y(men_men_n105_));
  NA2        u083(.A(men_men_n105_), .B(men_men_n103_), .Y(men_men_n106_));
  NA2        u084(.A(men_men_n94_), .B(men_men_n28_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n71_), .Y(men_men_n108_));
  NO2        u086(.A(x10), .B(x01), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n29_), .B(x00), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n110_), .B(men_men_n109_), .Y(men_men_n111_));
  NA2        u089(.A(x04), .B(men_men_n28_), .Y(men_men_n112_));
  NO3        u090(.A(men_men_n112_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n113_));
  AOI210     u091(.A0(men_men_n113_), .A1(men_men_n111_), .B0(men_men_n108_), .Y(men_men_n114_));
  AOI210     u092(.A0(men_men_n114_), .A1(men_men_n106_), .B0(men_men_n101_), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n56_), .B(x05), .Y(men_men_n116_));
  NOi21      u094(.An(men_men_n116_), .B(men_men_n58_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n35_), .B(x02), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n101_), .B(men_men_n36_), .Y(men_men_n119_));
  NA3        u097(.A(men_men_n119_), .B(men_men_n118_), .C(x06), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(men_men_n117_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n84_), .B(x13), .Y(men_men_n122_));
  NA2        u100(.A(x09), .B(men_men_n35_), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n123_), .B(men_men_n122_), .Y(men_men_n124_));
  NA2        u102(.A(x13), .B(men_men_n35_), .Y(men_men_n125_));
  NO2        u103(.A(men_men_n125_), .B(x05), .Y(men_men_n126_));
  NO2        u104(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n128_), .B(men_men_n101_), .Y(men_men_n129_));
  AOI210     u107(.A0(men_men_n129_), .A1(men_men_n80_), .B0(men_men_n117_), .Y(men_men_n130_));
  AOI210     u108(.A0(men_men_n130_), .A1(men_men_n127_), .B0(men_men_n72_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n132_));
  NA2        u110(.A(x10), .B(men_men_n57_), .Y(men_men_n133_));
  NA2        u111(.A(men_men_n133_), .B(men_men_n132_), .Y(men_men_n134_));
  NA2        u112(.A(men_men_n51_), .B(x05), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n36_), .B(x04), .Y(men_men_n136_));
  NA3        u114(.A(men_men_n136_), .B(men_men_n135_), .C(x13), .Y(men_men_n137_));
  NO3        u115(.A(men_men_n128_), .B(men_men_n79_), .C(men_men_n36_), .Y(men_men_n138_));
  NO2        u116(.A(men_men_n60_), .B(x05), .Y(men_men_n139_));
  NOi41      u117(.An(men_men_n137_), .B(men_men_n139_), .C(men_men_n138_), .D(men_men_n134_), .Y(men_men_n140_));
  NO3        u118(.A(men_men_n140_), .B(x06), .C(x03), .Y(men_men_n141_));
  NO4        u119(.A(men_men_n141_), .B(men_men_n131_), .C(men_men_n121_), .D(men_men_n115_), .Y(men_men_n142_));
  NA2        u120(.A(x13), .B(men_men_n36_), .Y(men_men_n143_));
  OAI210     u121(.A0(men_men_n84_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n145_));
  NOi21      u123(.An(men_men_n89_), .B(men_men_n57_), .Y(men_men_n146_));
  NO2        u124(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n147_));
  OA210      u125(.A0(men_men_n146_), .A1(men_men_n77_), .B0(men_men_n147_), .Y(men_men_n148_));
  NO2        u126(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n149_));
  NA2        u127(.A(men_men_n29_), .B(x06), .Y(men_men_n150_));
  AOI210     u128(.A0(men_men_n150_), .A1(men_men_n49_), .B0(men_men_n149_), .Y(men_men_n151_));
  OA210      u129(.A0(men_men_n151_), .A1(men_men_n148_), .B0(men_men_n145_), .Y(men_men_n152_));
  NO2        u130(.A(x09), .B(x05), .Y(men_men_n153_));
  NA2        u131(.A(men_men_n153_), .B(men_men_n47_), .Y(men_men_n154_));
  AOI210     u132(.A0(men_men_n154_), .A1(men_men_n111_), .B0(men_men_n49_), .Y(men_men_n155_));
  NA2        u133(.A(x09), .B(x00), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n116_), .B(men_men_n156_), .Y(men_men_n157_));
  NA2        u135(.A(men_men_n76_), .B(men_men_n51_), .Y(men_men_n158_));
  AOI210     u136(.A0(men_men_n158_), .A1(men_men_n157_), .B0(men_men_n150_), .Y(men_men_n159_));
  NO3        u137(.A(men_men_n159_), .B(men_men_n155_), .C(men_men_n152_), .Y(men_men_n160_));
  NO2        u138(.A(x03), .B(x02), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n85_), .B(men_men_n101_), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n162_), .A1(men_men_n117_), .B0(men_men_n161_), .Y(men_men_n163_));
  OA210      u141(.A0(men_men_n160_), .A1(x11), .B0(men_men_n163_), .Y(men_men_n164_));
  OAI210     u142(.A0(men_men_n142_), .A1(men_men_n23_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u143(.A(men_men_n111_), .B(men_men_n40_), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n167_));
  NAi21      u145(.An(x06), .B(x10), .Y(men_men_n168_));
  NOi21      u146(.An(x01), .B(x13), .Y(men_men_n169_));
  NA2        u147(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  OR2        u148(.A(men_men_n170_), .B(men_men_n167_), .Y(men_men_n171_));
  AOI210     u149(.A0(men_men_n171_), .A1(men_men_n166_), .B0(men_men_n41_), .Y(men_men_n172_));
  NO2        u150(.A(men_men_n29_), .B(x03), .Y(men_men_n173_));
  NA2        u151(.A(men_men_n101_), .B(x01), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n174_), .B(x08), .Y(men_men_n175_));
  OAI210     u153(.A0(x05), .A1(men_men_n175_), .B0(men_men_n51_), .Y(men_men_n176_));
  AOI210     u154(.A0(men_men_n176_), .A1(men_men_n173_), .B0(men_men_n48_), .Y(men_men_n177_));
  AOI210     u155(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n177_), .A1(men_men_n172_), .B0(men_men_n178_), .Y(men_men_n179_));
  NA2        u157(.A(x04), .B(x02), .Y(men_men_n180_));
  NA2        u158(.A(x10), .B(x05), .Y(men_men_n181_));
  NA2        u159(.A(x09), .B(x06), .Y(men_men_n182_));
  AOI210     u160(.A0(men_men_n182_), .A1(men_men_n181_), .B0(men_men_n167_), .Y(men_men_n183_));
  NO2        u161(.A(x09), .B(x01), .Y(men_men_n184_));
  NO3        u162(.A(men_men_n184_), .B(men_men_n109_), .C(men_men_n31_), .Y(men_men_n185_));
  OAI210     u163(.A0(men_men_n185_), .A1(men_men_n183_), .B0(x00), .Y(men_men_n186_));
  NO2        u164(.A(men_men_n116_), .B(x08), .Y(men_men_n187_));
  NA3        u165(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n51_), .Y(men_men_n188_));
  NA2        u166(.A(men_men_n94_), .B(x05), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n119_), .B0(men_men_n188_), .Y(men_men_n190_));
  AOI210     u168(.A0(men_men_n187_), .A1(x06), .B0(men_men_n190_), .Y(men_men_n191_));
  OAI210     u169(.A0(men_men_n191_), .A1(x11), .B0(men_men_n186_), .Y(men_men_n192_));
  NAi21      u170(.An(men_men_n180_), .B(men_men_n192_), .Y(men_men_n193_));
  INV        u171(.A(men_men_n25_), .Y(men_men_n194_));
  NAi21      u172(.An(x13), .B(x00), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n195_), .Y(men_men_n196_));
  AOI220     u174(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n197_));
  OAI210     u175(.A0(men_men_n181_), .A1(men_men_n35_), .B0(men_men_n197_), .Y(men_men_n198_));
  AN2        u176(.A(men_men_n198_), .B(men_men_n196_), .Y(men_men_n199_));
  AN2        u177(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n200_));
  NO2        u178(.A(men_men_n95_), .B(x06), .Y(men_men_n201_));
  NO2        u179(.A(men_men_n195_), .B(men_men_n36_), .Y(men_men_n202_));
  INV        u180(.A(men_men_n202_), .Y(men_men_n203_));
  OAI220     u181(.A0(men_men_n203_), .A1(men_men_n182_), .B0(men_men_n201_), .B1(men_men_n200_), .Y(men_men_n204_));
  OAI210     u182(.A0(men_men_n204_), .A1(men_men_n199_), .B0(men_men_n194_), .Y(men_men_n205_));
  NOi21      u183(.An(x09), .B(x00), .Y(men_men_n206_));
  NO3        u184(.A(men_men_n83_), .B(men_men_n206_), .C(men_men_n47_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(men_men_n133_), .Y(men_men_n208_));
  NA2        u186(.A(x10), .B(x08), .Y(men_men_n209_));
  INV        u187(.A(men_men_n209_), .Y(men_men_n210_));
  NA2        u188(.A(x06), .B(x05), .Y(men_men_n211_));
  OAI210     u189(.A0(men_men_n211_), .A1(men_men_n35_), .B0(men_men_n100_), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n210_), .A1(men_men_n58_), .B0(men_men_n212_), .Y(men_men_n213_));
  NA2        u191(.A(men_men_n213_), .B(men_men_n208_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n101_), .B(x12), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n215_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n94_), .B(men_men_n51_), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n218_), .B(x02), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n219_), .B(men_men_n217_), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n216_), .A1(men_men_n214_), .B0(men_men_n220_), .Y(men_men_n221_));
  NA4        u199(.A(men_men_n221_), .B(men_men_n205_), .C(men_men_n193_), .D(men_men_n179_), .Y(men_men_n222_));
  AOI210     u200(.A0(men_men_n165_), .A1(men_men_n100_), .B0(men_men_n222_), .Y(men_men_n223_));
  AOI210     u201(.A0(men_men_n143_), .A1(x09), .B0(men_men_n73_), .Y(men_men_n224_));
  NA2        u202(.A(men_men_n224_), .B(men_men_n145_), .Y(men_men_n225_));
  NA2        u203(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n226_), .B(men_men_n144_), .Y(men_men_n227_));
  AOI210     u205(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n132_), .B(x06), .Y(men_men_n229_));
  AOI210     u207(.A0(men_men_n228_), .A1(men_men_n227_), .B0(men_men_n229_), .Y(men_men_n230_));
  AOI210     u208(.A0(men_men_n230_), .A1(men_men_n225_), .B0(x12), .Y(men_men_n231_));
  INV        u209(.A(men_men_n76_), .Y(men_men_n232_));
  AOI210     u210(.A0(men_men_n209_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n233_));
  OAI210     u211(.A0(men_men_n233_), .A1(men_men_n170_), .B0(men_men_n57_), .Y(men_men_n234_));
  NA2        u212(.A(men_men_n234_), .B(men_men_n232_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n94_), .B(x06), .Y(men_men_n236_));
  AOI210     u214(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n237_));
  NO3        u215(.A(men_men_n237_), .B(men_men_n236_), .C(men_men_n41_), .Y(men_men_n238_));
  NA4        u216(.A(men_men_n168_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n239_), .B(men_men_n150_), .Y(men_men_n240_));
  OAI210     u218(.A0(men_men_n240_), .A1(men_men_n238_), .B0(x02), .Y(men_men_n241_));
  AOI210     u219(.A0(men_men_n241_), .A1(men_men_n235_), .B0(men_men_n23_), .Y(men_men_n242_));
  OAI210     u220(.A0(men_men_n231_), .A1(men_men_n57_), .B0(men_men_n242_), .Y(men_men_n243_));
  INV        u221(.A(men_men_n150_), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n51_), .B(x03), .Y(men_men_n245_));
  OAI210     u223(.A0(men_men_n79_), .A1(men_men_n36_), .B0(men_men_n123_), .Y(men_men_n246_));
  NO2        u224(.A(men_men_n101_), .B(x03), .Y(men_men_n247_));
  AOI220     u225(.A0(men_men_n247_), .A1(men_men_n246_), .B0(men_men_n76_), .B1(men_men_n245_), .Y(men_men_n248_));
  NA2        u226(.A(men_men_n32_), .B(x06), .Y(men_men_n249_));
  INV        u227(.A(men_men_n168_), .Y(men_men_n250_));
  NOi21      u228(.An(x13), .B(x04), .Y(men_men_n251_));
  NO3        u229(.A(men_men_n251_), .B(men_men_n76_), .C(men_men_n206_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(x05), .Y(men_men_n253_));
  AOI220     u231(.A0(men_men_n253_), .A1(men_men_n249_), .B0(men_men_n250_), .B1(men_men_n57_), .Y(men_men_n254_));
  OAI210     u232(.A0(men_men_n248_), .A1(men_men_n244_), .B0(men_men_n254_), .Y(men_men_n255_));
  INV        u233(.A(men_men_n91_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n257_));
  NO2        u235(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n258_));
  OAI210     u236(.A0(men_men_n258_), .A1(men_men_n198_), .B0(men_men_n196_), .Y(men_men_n259_));
  AOI210     u237(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n260_));
  NO2        u238(.A(x06), .B(x00), .Y(men_men_n261_));
  NO3        u239(.A(men_men_n261_), .B(men_men_n260_), .C(men_men_n41_), .Y(men_men_n262_));
  OAI210     u240(.A0(men_men_n104_), .A1(men_men_n156_), .B0(men_men_n72_), .Y(men_men_n263_));
  NO2        u241(.A(men_men_n263_), .B(men_men_n262_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n265_));
  NA2        u243(.A(men_men_n265_), .B(x03), .Y(men_men_n266_));
  OA210      u244(.A0(men_men_n266_), .A1(men_men_n264_), .B0(men_men_n259_), .Y(men_men_n267_));
  NA2        u245(.A(x13), .B(men_men_n100_), .Y(men_men_n268_));
  NA3        u246(.A(men_men_n268_), .B(men_men_n212_), .C(men_men_n92_), .Y(men_men_n269_));
  OAI210     u247(.A0(men_men_n267_), .A1(men_men_n257_), .B0(men_men_n269_), .Y(men_men_n270_));
  AOI210     u248(.A0(men_men_n91_), .A1(men_men_n255_), .B0(men_men_n270_), .Y(men_men_n271_));
  AOI210     u249(.A0(men_men_n271_), .A1(men_men_n243_), .B0(x07), .Y(men_men_n272_));
  NA2        u250(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n273_));
  NOi31      u251(.An(men_men_n143_), .B(men_men_n251_), .C(men_men_n206_), .Y(men_men_n274_));
  AOI210     u252(.A0(men_men_n274_), .A1(men_men_n158_), .B0(men_men_n273_), .Y(men_men_n275_));
  NO2        u253(.A(men_men_n101_), .B(x06), .Y(men_men_n276_));
  INV        u254(.A(men_men_n276_), .Y(men_men_n277_));
  NO2        u255(.A(x08), .B(x05), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n278_), .B(men_men_n260_), .Y(men_men_n279_));
  OAI210     u257(.A0(men_men_n76_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n280_));
  OAI210     u258(.A0(men_men_n279_), .A1(men_men_n277_), .B0(men_men_n280_), .Y(men_men_n281_));
  NO2        u259(.A(x12), .B(x02), .Y(men_men_n282_));
  INV        u260(.A(men_men_n282_), .Y(men_men_n283_));
  NO2        u261(.A(men_men_n283_), .B(men_men_n256_), .Y(men_men_n284_));
  OA210      u262(.A0(men_men_n281_), .A1(men_men_n275_), .B0(men_men_n284_), .Y(men_men_n285_));
  NA2        u263(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n286_));
  NO2        u264(.A(men_men_n286_), .B(x01), .Y(men_men_n287_));
  NOi21      u265(.An(men_men_n84_), .B(men_men_n123_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n288_), .B(men_men_n287_), .Y(men_men_n289_));
  AOI210     u267(.A0(men_men_n289_), .A1(men_men_n137_), .B0(men_men_n29_), .Y(men_men_n290_));
  NA2        u268(.A(men_men_n276_), .B(men_men_n246_), .Y(men_men_n291_));
  NA2        u269(.A(men_men_n101_), .B(x04), .Y(men_men_n292_));
  NA2        u270(.A(men_men_n292_), .B(men_men_n28_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n293_), .A1(men_men_n122_), .B0(men_men_n291_), .Y(men_men_n294_));
  NO3        u272(.A(men_men_n90_), .B(x12), .C(x03), .Y(men_men_n295_));
  OAI210     u273(.A0(men_men_n294_), .A1(men_men_n290_), .B0(men_men_n295_), .Y(men_men_n296_));
  AOI210     u274(.A0(men_men_n217_), .A1(men_men_n211_), .B0(men_men_n104_), .Y(men_men_n297_));
  NOi21      u275(.An(men_men_n273_), .B(men_men_n236_), .Y(men_men_n298_));
  NO2        u276(.A(men_men_n25_), .B(x00), .Y(men_men_n299_));
  OAI210     u277(.A0(men_men_n298_), .A1(men_men_n297_), .B0(men_men_n299_), .Y(men_men_n300_));
  NO2        u278(.A(men_men_n58_), .B(x05), .Y(men_men_n301_));
  NO3        u279(.A(men_men_n301_), .B(men_men_n237_), .C(men_men_n201_), .Y(men_men_n302_));
  NO2        u280(.A(men_men_n257_), .B(men_men_n28_), .Y(men_men_n303_));
  OAI210     u281(.A0(men_men_n302_), .A1(men_men_n244_), .B0(men_men_n303_), .Y(men_men_n304_));
  NA3        u282(.A(men_men_n304_), .B(men_men_n300_), .C(men_men_n296_), .Y(men_men_n305_));
  NO3        u283(.A(men_men_n305_), .B(men_men_n285_), .C(men_men_n272_), .Y(men_men_n306_));
  OAI210     u284(.A0(men_men_n223_), .A1(men_men_n61_), .B0(men_men_n306_), .Y(men02));
  AOI210     u285(.A0(men_men_n143_), .A1(men_men_n85_), .B0(men_men_n135_), .Y(men_men_n308_));
  NOi21      u286(.An(men_men_n252_), .B(men_men_n184_), .Y(men_men_n309_));
  NO2        u287(.A(men_men_n101_), .B(men_men_n35_), .Y(men_men_n310_));
  NA3        u288(.A(men_men_n310_), .B(men_men_n210_), .C(men_men_n56_), .Y(men_men_n311_));
  OAI210     u289(.A0(men_men_n309_), .A1(men_men_n32_), .B0(men_men_n311_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n312_), .A1(men_men_n308_), .B0(men_men_n181_), .Y(men_men_n313_));
  INV        u291(.A(men_men_n181_), .Y(men_men_n314_));
  AOI210     u292(.A0(men_men_n118_), .A1(men_men_n86_), .B0(men_men_n237_), .Y(men_men_n315_));
  OAI220     u293(.A0(men_men_n315_), .A1(men_men_n101_), .B0(men_men_n85_), .B1(men_men_n51_), .Y(men_men_n316_));
  AOI220     u294(.A0(men_men_n316_), .A1(men_men_n314_), .B0(men_men_n162_), .B1(men_men_n161_), .Y(men_men_n317_));
  AOI210     u295(.A0(men_men_n317_), .A1(men_men_n313_), .B0(men_men_n48_), .Y(men_men_n318_));
  NO2        u296(.A(x05), .B(x02), .Y(men_men_n319_));
  OAI210     u297(.A0(men_men_n227_), .A1(men_men_n206_), .B0(men_men_n319_), .Y(men_men_n320_));
  AOI220     u298(.A0(men_men_n278_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n321_));
  NOi21      u299(.An(men_men_n310_), .B(men_men_n321_), .Y(men_men_n322_));
  AOI210     u300(.A0(men_men_n251_), .A1(men_men_n79_), .B0(men_men_n322_), .Y(men_men_n323_));
  AOI210     u301(.A0(men_men_n323_), .A1(men_men_n320_), .B0(men_men_n150_), .Y(men_men_n324_));
  NAi21      u302(.An(men_men_n253_), .B(men_men_n248_), .Y(men_men_n325_));
  NO2        u303(.A(men_men_n265_), .B(men_men_n47_), .Y(men_men_n326_));
  NA2        u304(.A(men_men_n326_), .B(men_men_n325_), .Y(men_men_n327_));
  AN2        u305(.A(men_men_n247_), .B(men_men_n246_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n329_));
  NA2        u307(.A(x13), .B(men_men_n28_), .Y(men_men_n330_));
  OA210      u308(.A0(men_men_n330_), .A1(x08), .B0(men_men_n154_), .Y(men_men_n331_));
  AOI210     u309(.A0(men_men_n331_), .A1(men_men_n144_), .B0(men_men_n329_), .Y(men_men_n332_));
  OAI210     u310(.A0(men_men_n332_), .A1(men_men_n328_), .B0(men_men_n95_), .Y(men_men_n333_));
  NA3        u311(.A(men_men_n95_), .B(men_men_n84_), .C(men_men_n245_), .Y(men_men_n334_));
  NA3        u312(.A(men_men_n94_), .B(men_men_n83_), .C(men_men_n42_), .Y(men_men_n335_));
  AOI210     u313(.A0(men_men_n335_), .A1(men_men_n334_), .B0(x04), .Y(men_men_n336_));
  INV        u314(.A(men_men_n161_), .Y(men_men_n337_));
  OAI220     u315(.A0(men_men_n279_), .A1(men_men_n107_), .B0(men_men_n337_), .B1(men_men_n134_), .Y(men_men_n338_));
  AOI210     u316(.A0(men_men_n338_), .A1(x13), .B0(men_men_n336_), .Y(men_men_n339_));
  NA3        u317(.A(men_men_n339_), .B(men_men_n333_), .C(men_men_n327_), .Y(men_men_n340_));
  NO3        u318(.A(men_men_n340_), .B(men_men_n324_), .C(men_men_n318_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n149_), .B(x03), .Y(men_men_n342_));
  INV        u320(.A(men_men_n195_), .Y(men_men_n343_));
  OAI210     u321(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n344_));
  AOI220     u322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n218_), .B1(x08), .Y(men_men_n345_));
  OAI210     u323(.A0(men_men_n345_), .A1(men_men_n301_), .B0(men_men_n342_), .Y(men_men_n346_));
  NA2        u324(.A(men_men_n346_), .B(men_men_n109_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n180_), .B(men_men_n174_), .Y(men_men_n348_));
  AN2        u326(.A(men_men_n348_), .B(men_men_n187_), .Y(men_men_n349_));
  INV        u327(.A(men_men_n56_), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n292_), .A1(men_men_n350_), .B0(men_men_n135_), .B1(men_men_n28_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n351_), .A1(men_men_n349_), .B0(men_men_n110_), .Y(men_men_n352_));
  NA2        u330(.A(men_men_n292_), .B(men_men_n100_), .Y(men_men_n353_));
  NA2        u331(.A(men_men_n100_), .B(men_men_n41_), .Y(men_men_n354_));
  NA3        u332(.A(men_men_n354_), .B(men_men_n353_), .C(men_men_n134_), .Y(men_men_n355_));
  NA4        u333(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n347_), .D(men_men_n48_), .Y(men_men_n356_));
  INV        u334(.A(men_men_n218_), .Y(men_men_n357_));
  NO2        u335(.A(men_men_n175_), .B(men_men_n40_), .Y(men_men_n358_));
  NA2        u336(.A(men_men_n32_), .B(x05), .Y(men_men_n359_));
  OAI220     u337(.A0(men_men_n359_), .A1(men_men_n358_), .B0(men_men_n357_), .B1(men_men_n59_), .Y(men_men_n360_));
  NA2        u338(.A(men_men_n360_), .B(x02), .Y(men_men_n361_));
  INV        u339(.A(men_men_n258_), .Y(men_men_n362_));
  NA2        u340(.A(men_men_n215_), .B(x04), .Y(men_men_n363_));
  NO2        u341(.A(men_men_n363_), .B(men_men_n362_), .Y(men_men_n364_));
  NO3        u342(.A(men_men_n197_), .B(x13), .C(men_men_n31_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n364_), .B0(men_men_n95_), .Y(men_men_n366_));
  NO3        u344(.A(men_men_n215_), .B(men_men_n173_), .C(men_men_n52_), .Y(men_men_n367_));
  OAI210     u345(.A0(men_men_n156_), .A1(men_men_n36_), .B0(men_men_n100_), .Y(men_men_n368_));
  OAI210     u346(.A0(men_men_n368_), .A1(men_men_n207_), .B0(men_men_n367_), .Y(men_men_n369_));
  NA4        u347(.A(men_men_n369_), .B(men_men_n366_), .C(men_men_n361_), .D(x06), .Y(men_men_n370_));
  NA2        u348(.A(x09), .B(x03), .Y(men_men_n371_));
  OAI220     u349(.A0(men_men_n371_), .A1(men_men_n133_), .B0(men_men_n226_), .B1(men_men_n63_), .Y(men_men_n372_));
  OAI220     u350(.A0(men_men_n174_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n373_));
  NO3        u351(.A(men_men_n301_), .B(men_men_n132_), .C(x08), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n373_), .A1(men_men_n244_), .B0(men_men_n374_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n376_));
  NO3        u354(.A(men_men_n116_), .B(men_men_n133_), .C(men_men_n38_), .Y(men_men_n377_));
  AOI210     u355(.A0(men_men_n367_), .A1(men_men_n376_), .B0(men_men_n377_), .Y(men_men_n378_));
  OAI210     u356(.A0(men_men_n375_), .A1(men_men_n28_), .B0(men_men_n378_), .Y(men_men_n379_));
  AO220      u357(.A0(men_men_n379_), .A1(x04), .B0(men_men_n372_), .B1(x05), .Y(men_men_n380_));
  AOI210     u358(.A0(men_men_n370_), .A1(men_men_n356_), .B0(men_men_n380_), .Y(men_men_n381_));
  OAI210     u359(.A0(men_men_n341_), .A1(x12), .B0(men_men_n381_), .Y(men03));
  OR2        u360(.A(men_men_n42_), .B(men_men_n245_), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n162_), .A1(men_men_n100_), .B0(men_men_n383_), .Y(men_men_n384_));
  AO210      u362(.A0(men_men_n362_), .A1(men_men_n86_), .B0(men_men_n363_), .Y(men_men_n385_));
  NA2        u363(.A(men_men_n215_), .B(men_men_n161_), .Y(men_men_n386_));
  NA3        u364(.A(men_men_n386_), .B(men_men_n385_), .C(men_men_n219_), .Y(men_men_n387_));
  OAI210     u365(.A0(men_men_n387_), .A1(men_men_n384_), .B0(x05), .Y(men_men_n388_));
  NA2        u366(.A(men_men_n383_), .B(x05), .Y(men_men_n389_));
  AOI210     u367(.A0(men_men_n144_), .A1(men_men_n232_), .B0(men_men_n389_), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n247_), .A1(men_men_n80_), .B0(men_men_n126_), .Y(men_men_n391_));
  OAI220     u369(.A0(men_men_n391_), .A1(men_men_n59_), .B0(men_men_n330_), .B1(men_men_n321_), .Y(men_men_n392_));
  OAI210     u370(.A0(men_men_n392_), .A1(men_men_n390_), .B0(men_men_n100_), .Y(men_men_n393_));
  AOI210     u371(.A0(men_men_n154_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n394_));
  NO2        u372(.A(men_men_n184_), .B(men_men_n139_), .Y(men_men_n395_));
  OAI220     u373(.A0(men_men_n395_), .A1(men_men_n37_), .B0(men_men_n157_), .B1(x13), .Y(men_men_n396_));
  OAI210     u374(.A0(men_men_n396_), .A1(men_men_n394_), .B0(x04), .Y(men_men_n397_));
  NO3        u375(.A(men_men_n354_), .B(men_men_n85_), .C(men_men_n59_), .Y(men_men_n398_));
  NO2        u376(.A(men_men_n203_), .B(men_men_n154_), .Y(men_men_n399_));
  OA210      u377(.A0(men_men_n175_), .A1(x12), .B0(men_men_n139_), .Y(men_men_n400_));
  NO3        u378(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n398_), .Y(men_men_n401_));
  NA4        u379(.A(men_men_n401_), .B(men_men_n397_), .C(men_men_n393_), .D(men_men_n388_), .Y(men04));
  AOI210     u380(.A0(men_men_n71_), .A1(men_men_n52_), .B0(men_men_n229_), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n403_), .A1(men_men_n329_), .B0(men_men_n25_), .Y(men_men_n404_));
  NA3        u382(.A(men_men_n150_), .B(men_men_n135_), .C(men_men_n31_), .Y(men_men_n405_));
  AOI210     u383(.A0(men_men_n250_), .A1(men_men_n57_), .B0(men_men_n89_), .Y(men_men_n406_));
  AOI210     u384(.A0(men_men_n406_), .A1(men_men_n405_), .B0(men_men_n24_), .Y(men_men_n407_));
  OAI210     u385(.A0(men_men_n407_), .A1(men_men_n404_), .B0(men_men_n100_), .Y(men_men_n408_));
  NA2        u386(.A(x11), .B(men_men_n31_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n410_));
  NA2        u388(.A(men_men_n273_), .B(x03), .Y(men_men_n411_));
  OAI220     u389(.A0(men_men_n411_), .A1(men_men_n410_), .B0(men_men_n409_), .B1(men_men_n81_), .Y(men_men_n412_));
  OAI210     u390(.A0(men_men_n26_), .A1(men_men_n100_), .B0(x07), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n412_), .A1(x06), .B0(men_men_n413_), .Y(men_men_n414_));
  AOI220     u392(.A0(men_men_n81_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n415_));
  NO3        u393(.A(men_men_n415_), .B(men_men_n23_), .C(x00), .Y(men_men_n416_));
  NA2        u394(.A(men_men_n70_), .B(x02), .Y(men_men_n417_));
  AOI210     u395(.A0(men_men_n417_), .A1(men_men_n411_), .B0(men_men_n276_), .Y(men_men_n418_));
  OR2        u396(.A(men_men_n418_), .B(men_men_n257_), .Y(men_men_n419_));
  NA2        u397(.A(men_men_n169_), .B(x05), .Y(men_men_n420_));
  NA3        u398(.A(men_men_n420_), .B(men_men_n261_), .C(men_men_n256_), .Y(men_men_n421_));
  NO2        u399(.A(men_men_n23_), .B(x10), .Y(men_men_n422_));
  OAI210     u400(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n423_));
  OR3        u401(.A(men_men_n423_), .B(men_men_n422_), .C(men_men_n44_), .Y(men_men_n424_));
  NA3        u402(.A(men_men_n424_), .B(men_men_n421_), .C(men_men_n419_), .Y(men_men_n425_));
  OAI210     u403(.A0(men_men_n425_), .A1(men_men_n416_), .B0(men_men_n100_), .Y(men_men_n426_));
  NA2        u404(.A(men_men_n33_), .B(men_men_n100_), .Y(men_men_n427_));
  AOI210     u405(.A0(men_men_n427_), .A1(men_men_n91_), .B0(x07), .Y(men_men_n428_));
  AOI220     u406(.A0(men_men_n428_), .A1(men_men_n426_), .B0(men_men_n414_), .B1(men_men_n408_), .Y(men_men_n429_));
  NA3        u407(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n430_));
  AO210      u408(.A0(men_men_n430_), .A1(men_men_n286_), .B0(men_men_n283_), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n422_), .A1(men_men_n74_), .B0(men_men_n149_), .Y(men_men_n432_));
  OR2        u410(.A(men_men_n432_), .B(x03), .Y(men_men_n433_));
  NA2        u411(.A(men_men_n376_), .B(men_men_n61_), .Y(men_men_n434_));
  NO2        u412(.A(men_men_n434_), .B(x11), .Y(men_men_n435_));
  NO3        u413(.A(men_men_n435_), .B(men_men_n153_), .C(men_men_n28_), .Y(men_men_n436_));
  AOI220     u414(.A0(men_men_n436_), .A1(men_men_n433_), .B0(men_men_n431_), .B1(men_men_n47_), .Y(men_men_n437_));
  NO4        u415(.A(men_men_n354_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n438_));
  OAI210     u416(.A0(men_men_n438_), .A1(men_men_n437_), .B0(men_men_n101_), .Y(men_men_n439_));
  AOI210     u417(.A0(men_men_n363_), .A1(men_men_n112_), .B0(men_men_n282_), .Y(men_men_n440_));
  NOi21      u418(.An(men_men_n342_), .B(men_men_n139_), .Y(men_men_n441_));
  NO2        u419(.A(men_men_n441_), .B(men_men_n283_), .Y(men_men_n442_));
  OAI210     u420(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n443_));
  AOI210     u421(.A0(men_men_n268_), .A1(men_men_n47_), .B0(men_men_n443_), .Y(men_men_n444_));
  NO4        u422(.A(men_men_n444_), .B(men_men_n442_), .C(men_men_n440_), .D(x08), .Y(men_men_n445_));
  AOI210     u423(.A0(men_men_n422_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n446_));
  NA2        u424(.A(x09), .B(men_men_n41_), .Y(men_men_n447_));
  OAI220     u425(.A0(men_men_n447_), .A1(men_men_n446_), .B0(men_men_n409_), .B1(men_men_n66_), .Y(men_men_n448_));
  NO2        u426(.A(x13), .B(x12), .Y(men_men_n449_));
  NO2        u427(.A(men_men_n135_), .B(men_men_n28_), .Y(men_men_n450_));
  NO2        u428(.A(men_men_n450_), .B(men_men_n287_), .Y(men_men_n451_));
  OR3        u429(.A(men_men_n451_), .B(x12), .C(x03), .Y(men_men_n452_));
  NA3        u430(.A(men_men_n357_), .B(men_men_n128_), .C(x12), .Y(men_men_n453_));
  AO210      u431(.A0(men_men_n357_), .A1(men_men_n128_), .B0(men_men_n268_), .Y(men_men_n454_));
  NA4        u432(.A(men_men_n454_), .B(men_men_n453_), .C(men_men_n452_), .D(x08), .Y(men_men_n455_));
  AOI210     u433(.A0(men_men_n449_), .A1(men_men_n448_), .B0(men_men_n455_), .Y(men_men_n456_));
  AOI210     u434(.A0(men_men_n445_), .A1(men_men_n439_), .B0(men_men_n456_), .Y(men_men_n457_));
  OAI210     u435(.A0(men_men_n434_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n458_));
  NA2        u436(.A(men_men_n314_), .B(x07), .Y(men_men_n459_));
  OAI220     u437(.A0(men_men_n459_), .A1(men_men_n410_), .B0(men_men_n153_), .B1(men_men_n43_), .Y(men_men_n460_));
  OAI210     u438(.A0(men_men_n460_), .A1(men_men_n458_), .B0(men_men_n202_), .Y(men_men_n461_));
  NA3        u439(.A(men_men_n451_), .B(men_men_n441_), .C(men_men_n353_), .Y(men_men_n462_));
  NO3        u440(.A(men_men_n342_), .B(men_men_n107_), .C(x11), .Y(men_men_n463_));
  NO3        u441(.A(men_men_n174_), .B(men_men_n74_), .C(men_men_n57_), .Y(men_men_n464_));
  NO3        u442(.A(men_men_n430_), .B(men_men_n354_), .C(men_men_n195_), .Y(men_men_n465_));
  NO3        u443(.A(men_men_n465_), .B(men_men_n464_), .C(men_men_n463_), .Y(men_men_n466_));
  NA3        u444(.A(men_men_n466_), .B(men_men_n462_), .C(men_men_n461_), .Y(men_men_n467_));
  AOI220     u445(.A0(men_men_n427_), .A1(men_men_n61_), .B0(men_men_n450_), .B1(men_men_n173_), .Y(men_men_n468_));
  NOi21      u446(.An(men_men_n292_), .B(men_men_n157_), .Y(men_men_n469_));
  NO3        u447(.A(men_men_n132_), .B(men_men_n24_), .C(x06), .Y(men_men_n470_));
  AOI210     u448(.A0(men_men_n299_), .A1(men_men_n250_), .B0(men_men_n470_), .Y(men_men_n471_));
  OAI210     u449(.A0(men_men_n44_), .A1(x04), .B0(men_men_n471_), .Y(men_men_n472_));
  OAI210     u450(.A0(men_men_n472_), .A1(men_men_n469_), .B0(men_men_n100_), .Y(men_men_n473_));
  OAI210     u451(.A0(men_men_n468_), .A1(men_men_n90_), .B0(men_men_n473_), .Y(men_men_n474_));
  NO4        u452(.A(men_men_n474_), .B(men_men_n467_), .C(men_men_n457_), .D(men_men_n429_), .Y(men06));
  INV        u453(.A(x07), .Y(men_men_n478_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule