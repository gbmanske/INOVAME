library verilog;
use verilog.vl_types.all;
entity interp_vlg_vec_tst is
end interp_vlg_vec_tst;
