//Benchmark atmr_9sym_175_0.5

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m00(.A(i_3_), .Y(mai_mai_n11_));
  INV        m01(.A(i_6_), .Y(mai_mai_n12_));
  INV        m02(.A(i_5_), .Y(mai_mai_n13_));
  INV        m03(.A(i_0_), .Y(mai_mai_n14_));
  INV        m04(.A(i_4_), .Y(mai_mai_n15_));
  NA2        m05(.A(i_0_), .B(mai_mai_n15_), .Y(mai_mai_n16_));
  INV        m06(.A(i_7_), .Y(mai_mai_n17_));
  NA3        m07(.A(i_6_), .B(i_5_), .C(mai_mai_n17_), .Y(mai_mai_n18_));
  NO2        m08(.A(mai_mai_n18_), .B(mai_mai_n16_), .Y(mai_mai_n19_));
  NA2        m09(.A(mai_mai_n19_), .B(mai_mai_n11_), .Y(mai_mai_n20_));
  NA2        m10(.A(mai_mai_n14_), .B(i_5_), .Y(mai_mai_n21_));
  INV        m11(.A(i_2_), .Y(mai_mai_n22_));
  NOi21      m12(.An(i_5_), .B(i_0_), .Y(mai_mai_n23_));
  NOi21      m13(.An(i_6_), .B(i_8_), .Y(mai_mai_n24_));
  NOi21      m14(.An(i_7_), .B(i_1_), .Y(mai_mai_n25_));
  NOi21      m15(.An(i_5_), .B(i_6_), .Y(mai_mai_n26_));
  AOI220     m16(.A0(mai_mai_n26_), .A1(mai_mai_n25_), .B0(mai_mai_n24_), .B1(mai_mai_n23_), .Y(mai_mai_n27_));
  NO3        m17(.A(mai_mai_n27_), .B(mai_mai_n22_), .C(i_4_), .Y(mai_mai_n28_));
  NOi21      m18(.An(i_0_), .B(i_4_), .Y(mai_mai_n29_));
  XO2        m19(.A(i_1_), .B(i_3_), .Y(mai_mai_n30_));
  NOi21      m20(.An(i_7_), .B(i_5_), .Y(mai_mai_n31_));
  AN3        m21(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  INV        m22(.A(i_1_), .Y(mai_mai_n33_));
  NOi21      m23(.An(i_3_), .B(i_0_), .Y(mai_mai_n34_));
  NA2        m24(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  NA3        m25(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n36_));
  AOI210     m26(.A0(mai_mai_n36_), .A1(mai_mai_n18_), .B0(mai_mai_n35_), .Y(mai_mai_n37_));
  NO3        m27(.A(mai_mai_n37_), .B(mai_mai_n32_), .C(mai_mai_n28_), .Y(mai_mai_n38_));
  NOi21      m28(.An(i_2_), .B(i_8_), .Y(mai_mai_n39_));
  NOi21      m29(.An(i_4_), .B(i_3_), .Y(mai_mai_n40_));
  NOi21      m30(.An(i_1_), .B(i_4_), .Y(mai_mai_n41_));
  OAI210     m31(.A0(mai_mai_n41_), .A1(mai_mai_n40_), .B0(mai_mai_n39_), .Y(mai_mai_n42_));
  INV        m32(.A(mai_mai_n42_), .Y(mai_mai_n43_));
  NOi21      m33(.An(i_8_), .B(i_7_), .Y(mai_mai_n44_));
  NA3        m34(.A(mai_mai_n44_), .B(mai_mai_n40_), .C(i_6_), .Y(mai_mai_n45_));
  INV        m35(.A(mai_mai_n45_), .Y(mai_mai_n46_));
  AOI220     m36(.A0(mai_mai_n46_), .A1(mai_mai_n22_), .B0(mai_mai_n43_), .B1(mai_mai_n26_), .Y(mai_mai_n47_));
  NA3        m37(.A(mai_mai_n47_), .B(mai_mai_n38_), .C(mai_mai_n20_), .Y(mai_mai_n48_));
  NA2        m38(.A(i_8_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  AOI220     m39(.A0(mai_mai_n34_), .A1(i_1_), .B0(mai_mai_n30_), .B1(i_2_), .Y(mai_mai_n50_));
  NOi21      m40(.An(i_1_), .B(i_2_), .Y(mai_mai_n51_));
  NO2        m41(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n52_));
  NA2        m42(.A(mai_mai_n52_), .B(mai_mai_n13_), .Y(mai_mai_n53_));
  NA3        m43(.A(mai_mai_n44_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n54_));
  INV        m44(.A(mai_mai_n53_), .Y(mai_mai_n55_));
  NA2        m45(.A(mai_mai_n24_), .B(mai_mai_n23_), .Y(mai_mai_n56_));
  INV        m46(.A(mai_mai_n56_), .Y(mai_mai_n57_));
  NA2        m47(.A(mai_mai_n57_), .B(mai_mai_n51_), .Y(mai_mai_n58_));
  NA3        m48(.A(mai_mai_n44_), .B(mai_mai_n22_), .C(i_3_), .Y(mai_mai_n59_));
  NO2        m49(.A(mai_mai_n16_), .B(mai_mai_n59_), .Y(mai_mai_n60_));
  NOi21      m50(.An(i_4_), .B(i_6_), .Y(mai_mai_n61_));
  INV        m51(.A(mai_mai_n60_), .Y(mai_mai_n62_));
  NA2        m52(.A(mai_mai_n62_), .B(mai_mai_n58_), .Y(mai_mai_n63_));
  NA2        m53(.A(mai_mai_n40_), .B(mai_mai_n25_), .Y(mai_mai_n64_));
  AOI210     m54(.A0(mai_mai_n64_), .A1(mai_mai_n54_), .B0(mai_mai_n21_), .Y(mai_mai_n65_));
  NOi21      m55(.An(i_0_), .B(i_2_), .Y(mai_mai_n66_));
  NA3        m56(.A(mai_mai_n66_), .B(mai_mai_n25_), .C(mai_mai_n61_), .Y(mai_mai_n67_));
  NA3        m57(.A(mai_mai_n66_), .B(mai_mai_n40_), .C(mai_mai_n24_), .Y(mai_mai_n68_));
  NA2        m58(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NO2        m59(.A(mai_mai_n69_), .B(mai_mai_n65_), .Y(mai_mai_n70_));
  NA3        m60(.A(mai_mai_n66_), .B(mai_mai_n44_), .C(mai_mai_n61_), .Y(mai_mai_n71_));
  OAI210     m61(.A0(mai_mai_n59_), .A1(mai_mai_n21_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  INV        m62(.A(mai_mai_n72_), .Y(mai_mai_n73_));
  NA2        m63(.A(mai_mai_n73_), .B(mai_mai_n70_), .Y(mai_mai_n74_));
  OR4        m64(.A(mai_mai_n74_), .B(mai_mai_n63_), .C(mai_mai_n55_), .D(mai_mai_n48_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  NO2        u016(.A(men_men_n26_), .B(men_men_n22_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n28_));
  NA2        u018(.A(i_0_), .B(men_men_n14_), .Y(men_men_n29_));
  NA2        u019(.A(men_men_n17_), .B(i_5_), .Y(men_men_n30_));
  NO2        u020(.A(i_2_), .B(i_4_), .Y(men_men_n31_));
  NA3        u021(.A(men_men_n31_), .B(i_6_), .C(i_8_), .Y(men_men_n32_));
  AOI210     u022(.A0(men_men_n30_), .A1(men_men_n29_), .B0(men_men_n32_), .Y(men_men_n33_));
  INV        u023(.A(i_2_), .Y(men_men_n34_));
  NOi21      u024(.An(i_5_), .B(i_0_), .Y(men_men_n35_));
  NOi21      u025(.An(i_6_), .B(i_8_), .Y(men_men_n36_));
  NOi21      u026(.An(i_5_), .B(i_6_), .Y(men_men_n37_));
  NOi21      u027(.An(i_0_), .B(i_4_), .Y(men_men_n38_));
  NOi21      u028(.An(i_7_), .B(i_5_), .Y(men_men_n39_));
  INV        u029(.A(i_1_), .Y(men_men_n40_));
  NOi21      u030(.An(i_3_), .B(i_0_), .Y(men_men_n41_));
  INV        u031(.A(men_men_n33_), .Y(men_men_n42_));
  INV        u032(.A(i_8_), .Y(men_men_n43_));
  NA2        u033(.A(i_1_), .B(men_men_n11_), .Y(men_men_n44_));
  NO4        u034(.A(men_men_n44_), .B(men_men_n29_), .C(i_2_), .D(men_men_n43_), .Y(men_men_n45_));
  NOi21      u035(.An(i_4_), .B(i_0_), .Y(men_men_n46_));
  AOI210     u036(.A0(men_men_n46_), .A1(men_men_n24_), .B0(men_men_n15_), .Y(men_men_n47_));
  NA2        u037(.A(i_1_), .B(men_men_n14_), .Y(men_men_n48_));
  NOi21      u038(.An(i_2_), .B(i_8_), .Y(men_men_n49_));
  NO3        u039(.A(men_men_n49_), .B(men_men_n46_), .C(men_men_n38_), .Y(men_men_n50_));
  NO3        u040(.A(men_men_n50_), .B(men_men_n48_), .C(men_men_n47_), .Y(men_men_n51_));
  NO2        u041(.A(men_men_n51_), .B(men_men_n45_), .Y(men_men_n52_));
  NOi31      u042(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n53_));
  NA2        u043(.A(men_men_n53_), .B(i_0_), .Y(men_men_n54_));
  NOi21      u044(.An(i_4_), .B(i_3_), .Y(men_men_n55_));
  NOi21      u045(.An(i_1_), .B(i_4_), .Y(men_men_n56_));
  INV        u046(.A(men_men_n54_), .Y(men_men_n57_));
  AN2        u047(.A(i_8_), .B(i_7_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(men_men_n12_), .Y(men_men_n59_));
  NOi21      u049(.An(i_8_), .B(i_7_), .Y(men_men_n60_));
  NO2        u050(.A(men_men_n59_), .B(men_men_n48_), .Y(men_men_n61_));
  AOI220     u051(.A0(men_men_n61_), .A1(men_men_n34_), .B0(men_men_n57_), .B1(men_men_n37_), .Y(men_men_n62_));
  NA4        u052(.A(men_men_n62_), .B(men_men_n52_), .C(men_men_n42_), .D(men_men_n28_), .Y(men_men_n63_));
  NA2        u053(.A(i_8_), .B(i_7_), .Y(men_men_n64_));
  NO3        u054(.A(men_men_n64_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n65_));
  NOi21      u055(.An(i_1_), .B(i_2_), .Y(men_men_n66_));
  NA3        u056(.A(men_men_n66_), .B(men_men_n46_), .C(i_6_), .Y(men_men_n67_));
  INV        u057(.A(men_men_n67_), .Y(men_men_n68_));
  OAI210     u058(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n14_), .Y(men_men_n69_));
  NA3        u059(.A(men_men_n60_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n70_));
  NA3        u060(.A(men_men_n25_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n71_));
  NA2        u061(.A(men_men_n71_), .B(men_men_n70_), .Y(men_men_n72_));
  NOi32      u062(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n73_));
  NA2        u063(.A(men_men_n73_), .B(i_3_), .Y(men_men_n74_));
  NA3        u064(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n75_));
  NA2        u065(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NO2        u066(.A(i_0_), .B(i_4_), .Y(men_men_n77_));
  AOI220     u067(.A0(men_men_n77_), .A1(men_men_n76_), .B0(men_men_n72_), .B1(men_men_n55_), .Y(men_men_n78_));
  NA2        u068(.A(men_men_n78_), .B(men_men_n69_), .Y(men_men_n79_));
  NAi21      u069(.An(i_3_), .B(i_6_), .Y(men_men_n80_));
  NO3        u070(.A(men_men_n80_), .B(i_0_), .C(men_men_n43_), .Y(men_men_n81_));
  NOi21      u071(.An(i_7_), .B(i_8_), .Y(men_men_n82_));
  NOi31      u072(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n83_));
  AOI210     u073(.A0(men_men_n82_), .A1(men_men_n12_), .B0(men_men_n83_), .Y(men_men_n84_));
  NO2        u074(.A(men_men_n84_), .B(men_men_n11_), .Y(men_men_n85_));
  OAI210     u075(.A0(men_men_n85_), .A1(men_men_n81_), .B0(men_men_n66_), .Y(men_men_n86_));
  NA3        u076(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n87_));
  AOI210     u077(.A0(men_men_n22_), .A1(men_men_n44_), .B0(men_men_n87_), .Y(men_men_n88_));
  AOI220     u078(.A0(men_men_n41_), .A1(men_men_n40_), .B0(men_men_n18_), .B1(men_men_n34_), .Y(men_men_n89_));
  NA3        u079(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n90_));
  OAI210     u080(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n91_));
  NA3        u081(.A(men_men_n64_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n92_));
  OAI220     u082(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n90_), .B1(men_men_n89_), .Y(men_men_n93_));
  NO2        u083(.A(men_men_n93_), .B(men_men_n88_), .Y(men_men_n94_));
  NA3        u084(.A(men_men_n60_), .B(men_men_n34_), .C(i_3_), .Y(men_men_n95_));
  NA2        u085(.A(men_men_n40_), .B(i_6_), .Y(men_men_n96_));
  NO2        u086(.A(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  NOi21      u087(.An(i_2_), .B(i_1_), .Y(men_men_n98_));
  AN3        u088(.A(men_men_n82_), .B(men_men_n98_), .C(men_men_n46_), .Y(men_men_n99_));
  NAi21      u089(.An(i_6_), .B(i_0_), .Y(men_men_n100_));
  NA3        u090(.A(men_men_n56_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n101_));
  NOi21      u091(.An(i_4_), .B(i_6_), .Y(men_men_n102_));
  NOi21      u092(.An(i_5_), .B(i_3_), .Y(men_men_n103_));
  NA3        u093(.A(men_men_n103_), .B(men_men_n66_), .C(men_men_n102_), .Y(men_men_n104_));
  OAI210     u094(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n104_), .Y(men_men_n105_));
  NA2        u095(.A(men_men_n66_), .B(men_men_n36_), .Y(men_men_n106_));
  NOi21      u096(.An(men_men_n39_), .B(men_men_n106_), .Y(men_men_n107_));
  NO4        u097(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n99_), .D(men_men_n97_), .Y(men_men_n108_));
  NOi21      u098(.An(i_6_), .B(i_1_), .Y(men_men_n109_));
  AOI220     u099(.A0(men_men_n109_), .A1(i_7_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n110_));
  NOi31      u100(.An(men_men_n46_), .B(men_men_n110_), .C(i_2_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n60_), .B(men_men_n12_), .Y(men_men_n112_));
  NA2        u102(.A(men_men_n36_), .B(men_men_n14_), .Y(men_men_n113_));
  NOi21      u103(.An(i_3_), .B(i_1_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n114_), .B(i_4_), .Y(men_men_n115_));
  AOI210     u105(.A0(men_men_n113_), .A1(men_men_n112_), .B0(men_men_n115_), .Y(men_men_n116_));
  AOI220     u106(.A0(men_men_n82_), .A1(men_men_n14_), .B0(men_men_n102_), .B1(men_men_n23_), .Y(men_men_n117_));
  NOi31      u107(.An(men_men_n41_), .B(men_men_n117_), .C(men_men_n34_), .Y(men_men_n118_));
  NO3        u108(.A(men_men_n118_), .B(men_men_n116_), .C(men_men_n111_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n119_), .B(men_men_n108_), .C(men_men_n94_), .D(men_men_n86_), .Y(men_men_n120_));
  NA2        u110(.A(men_men_n49_), .B(men_men_n15_), .Y(men_men_n121_));
  NOi31      u111(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n122_));
  NOi31      u112(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n123_));
  OAI210     u113(.A0(men_men_n123_), .A1(men_men_n122_), .B0(i_7_), .Y(men_men_n124_));
  NA3        u114(.A(men_men_n36_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n125_));
  NA4        u115(.A(men_men_n125_), .B(men_men_n124_), .C(men_men_n121_), .D(men_men_n106_), .Y(men_men_n126_));
  NA2        u116(.A(men_men_n126_), .B(men_men_n38_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n58_), .B(men_men_n98_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n128_));
  NAi31      u118(.An(men_men_n100_), .B(men_men_n82_), .C(men_men_n98_), .Y(men_men_n129_));
  NA3        u119(.A(men_men_n60_), .B(men_men_n53_), .C(i_6_), .Y(men_men_n130_));
  NA3        u120(.A(men_men_n130_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n131_));
  NA3        u121(.A(men_men_n46_), .B(men_men_n39_), .C(men_men_n18_), .Y(men_men_n132_));
  NOi32      u122(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n133_));
  NA2        u123(.A(men_men_n133_), .B(men_men_n122_), .Y(men_men_n134_));
  NA2        u124(.A(men_men_n134_), .B(men_men_n132_), .Y(men_men_n135_));
  NA4        u125(.A(men_men_n53_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n136_));
  NA4        u126(.A(men_men_n56_), .B(men_men_n37_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n137_));
  NA4        u127(.A(men_men_n56_), .B(men_men_n41_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n138_));
  NA3        u128(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NO3        u129(.A(men_men_n139_), .B(men_men_n135_), .C(men_men_n131_), .Y(men_men_n140_));
  NOi21      u130(.An(i_5_), .B(i_2_), .Y(men_men_n141_));
  AOI220     u131(.A0(men_men_n141_), .A1(men_men_n82_), .B0(men_men_n58_), .B1(men_men_n31_), .Y(men_men_n142_));
  AOI210     u132(.A0(men_men_n142_), .A1(men_men_n121_), .B0(men_men_n96_), .Y(men_men_n143_));
  NO4        u133(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n144_));
  NA2        u134(.A(i_2_), .B(i_4_), .Y(men_men_n145_));
  AOI210     u135(.A0(men_men_n100_), .A1(men_men_n80_), .B0(men_men_n145_), .Y(men_men_n146_));
  NO2        u136(.A(i_8_), .B(i_7_), .Y(men_men_n147_));
  OA210      u137(.A0(men_men_n146_), .A1(men_men_n144_), .B0(men_men_n147_), .Y(men_men_n148_));
  NA4        u138(.A(men_men_n114_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n149_));
  NO2        u139(.A(men_men_n149_), .B(i_4_), .Y(men_men_n150_));
  NO3        u140(.A(men_men_n150_), .B(men_men_n148_), .C(men_men_n143_), .Y(men_men_n151_));
  NA2        u141(.A(men_men_n82_), .B(men_men_n12_), .Y(men_men_n152_));
  NA3        u142(.A(i_2_), .B(i_1_), .C(men_men_n14_), .Y(men_men_n153_));
  NA2        u143(.A(men_men_n46_), .B(i_3_), .Y(men_men_n154_));
  AOI210     u144(.A0(men_men_n154_), .A1(men_men_n153_), .B0(men_men_n152_), .Y(men_men_n155_));
  NA4        u145(.A(men_men_n103_), .B(men_men_n58_), .C(men_men_n40_), .D(men_men_n21_), .Y(men_men_n156_));
  NA3        u146(.A(men_men_n83_), .B(men_men_n114_), .C(i_0_), .Y(men_men_n157_));
  NA3        u147(.A(men_men_n49_), .B(men_men_n35_), .C(men_men_n15_), .Y(men_men_n158_));
  NOi31      u148(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n159_));
  OAI210     u149(.A0(men_men_n133_), .A1(men_men_n73_), .B0(men_men_n159_), .Y(men_men_n160_));
  NA4        u150(.A(men_men_n160_), .B(men_men_n158_), .C(men_men_n157_), .D(men_men_n156_), .Y(men_men_n161_));
  NO2        u151(.A(men_men_n161_), .B(men_men_n155_), .Y(men_men_n162_));
  NA4        u152(.A(men_men_n162_), .B(men_men_n151_), .C(men_men_n140_), .D(men_men_n127_), .Y(men_men_n163_));
  OR4        u153(.A(men_men_n163_), .B(men_men_n120_), .C(men_men_n79_), .D(men_men_n63_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule