module test;
reg [7:0] a = 10;
initial
begin
$display("%b", a);
end
endmodule