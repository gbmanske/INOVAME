`ifndef empty_if__sv
`define empty_if__sv

interface empty_if (input clk);
  logic [7:0]   var0;
endinterface : empty_if

`endif



