//Benchmark atmr_alu4_1266_0.0313

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1033_, mai_mai_n1034_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1080_, men_men_n1081_, men_men_n1082_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NA2        o032(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n55_));
  NO2        o033(.A(i_1_), .B(i_6_), .Y(ori_ori_n56_));
  NA2        o034(.A(i_8_), .B(i_7_), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(i_12_), .Y(ori_ori_n59_));
  NAi21      o037(.An(i_2_), .B(i_7_), .Y(ori_ori_n60_));
  INV        o038(.A(i_1_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n61_), .B(i_6_), .Y(ori_ori_n62_));
  NA3        o040(.A(ori_ori_n62_), .B(ori_ori_n60_), .C(ori_ori_n31_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_1_), .B(i_10_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(i_6_), .Y(ori_ori_n65_));
  NAi31      o043(.An(ori_ori_n65_), .B(ori_ori_n63_), .C(ori_ori_n59_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n67_));
  AOI210     o045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n68_));
  NA2        o046(.A(i_1_), .B(i_6_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n25_), .Y(ori_ori_n70_));
  INV        o048(.A(i_0_), .Y(ori_ori_n71_));
  NAi21      o049(.An(i_5_), .B(i_10_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_5_), .B(i_9_), .Y(ori_ori_n73_));
  AOI210     o051(.A0(ori_ori_n73_), .A1(ori_ori_n72_), .B0(ori_ori_n71_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n74_), .B(ori_ori_n70_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n68_), .A1(ori_ori_n67_), .B0(ori_ori_n75_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n76_), .A1(ori_ori_n66_), .B0(i_0_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_12_), .B(i_5_), .Y(ori_ori_n78_));
  NA2        o056(.A(i_2_), .B(i_8_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n56_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_3_), .B(i_9_), .Y(ori_ori_n81_));
  NO2        o059(.A(i_3_), .B(i_7_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n81_), .B(ori_ori_n61_), .Y(ori_ori_n83_));
  INV        o061(.A(i_6_), .Y(ori_ori_n84_));
  OR4        o062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n85_));
  INV        o063(.A(ori_ori_n85_), .Y(ori_ori_n86_));
  NO2        o064(.A(i_2_), .B(i_7_), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n86_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  OAI210     o066(.A0(ori_ori_n83_), .A1(ori_ori_n80_), .B0(ori_ori_n88_), .Y(ori_ori_n89_));
  NAi21      o067(.An(i_6_), .B(i_10_), .Y(ori_ori_n90_));
  NA2        o068(.A(i_6_), .B(i_9_), .Y(ori_ori_n91_));
  AOI210     o069(.A0(ori_ori_n91_), .A1(ori_ori_n90_), .B0(ori_ori_n61_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_2_), .B(i_6_), .Y(ori_ori_n93_));
  NO3        o071(.A(ori_ori_n93_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n94_), .B(ori_ori_n92_), .Y(ori_ori_n95_));
  AOI210     o073(.A0(ori_ori_n95_), .A1(ori_ori_n89_), .B0(ori_ori_n78_), .Y(ori_ori_n96_));
  AN3        o074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n97_));
  NAi21      o075(.An(i_6_), .B(i_11_), .Y(ori_ori_n98_));
  NO2        o076(.A(i_5_), .B(i_8_), .Y(ori_ori_n99_));
  NOi21      o077(.An(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  AOI220     o078(.A0(ori_ori_n100_), .A1(ori_ori_n60_), .B0(ori_ori_n97_), .B1(ori_ori_n32_), .Y(ori_ori_n101_));
  INV        o079(.A(i_7_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n46_), .B(ori_ori_n102_), .Y(ori_ori_n103_));
  NO2        o081(.A(i_0_), .B(i_5_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(ori_ori_n84_), .Y(ori_ori_n105_));
  NA2        o083(.A(i_12_), .B(i_3_), .Y(ori_ori_n106_));
  INV        o084(.A(ori_ori_n106_), .Y(ori_ori_n107_));
  NA3        o085(.A(ori_ori_n107_), .B(ori_ori_n105_), .C(ori_ori_n103_), .Y(ori_ori_n108_));
  NAi21      o086(.An(i_7_), .B(i_11_), .Y(ori_ori_n109_));
  NO3        o087(.A(ori_ori_n109_), .B(ori_ori_n90_), .C(ori_ori_n53_), .Y(ori_ori_n110_));
  AN2        o088(.A(i_2_), .B(i_10_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(i_7_), .Y(ori_ori_n112_));
  OR2        o090(.A(ori_ori_n78_), .B(ori_ori_n56_), .Y(ori_ori_n113_));
  NO2        o091(.A(i_8_), .B(ori_ori_n102_), .Y(ori_ori_n114_));
  NO3        o092(.A(ori_ori_n114_), .B(ori_ori_n113_), .C(ori_ori_n112_), .Y(ori_ori_n115_));
  NA2        o093(.A(i_12_), .B(i_7_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n61_), .B(ori_ori_n26_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n117_), .B(i_0_), .Y(ori_ori_n118_));
  NA2        o096(.A(i_11_), .B(i_12_), .Y(ori_ori_n119_));
  OAI210     o097(.A0(ori_ori_n118_), .A1(ori_ori_n116_), .B0(ori_ori_n119_), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n120_), .B(ori_ori_n115_), .Y(ori_ori_n121_));
  NAi41      o099(.An(ori_ori_n110_), .B(ori_ori_n121_), .C(ori_ori_n108_), .D(ori_ori_n101_), .Y(ori_ori_n122_));
  NOi21      o100(.An(i_1_), .B(i_5_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(i_11_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n102_), .B(ori_ori_n37_), .Y(ori_ori_n125_));
  NA2        o103(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n126_), .B(ori_ori_n125_), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n127_), .B(ori_ori_n46_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n129_));
  NAi21      o107(.An(i_3_), .B(i_8_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(ori_ori_n60_), .Y(ori_ori_n131_));
  NOi31      o109(.An(ori_ori_n131_), .B(ori_ori_n129_), .C(ori_ori_n128_), .Y(ori_ori_n132_));
  NO2        o110(.A(i_1_), .B(ori_ori_n84_), .Y(ori_ori_n133_));
  NO2        o111(.A(i_6_), .B(i_5_), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n134_), .B(i_3_), .Y(ori_ori_n135_));
  AO210      o113(.A0(ori_ori_n135_), .A1(ori_ori_n47_), .B0(ori_ori_n133_), .Y(ori_ori_n136_));
  OAI220     o114(.A0(ori_ori_n136_), .A1(ori_ori_n109_), .B0(ori_ori_n132_), .B1(ori_ori_n124_), .Y(ori_ori_n137_));
  NO3        o115(.A(ori_ori_n137_), .B(ori_ori_n122_), .C(ori_ori_n96_), .Y(ori_ori_n138_));
  NA3        o116(.A(ori_ori_n138_), .B(ori_ori_n77_), .C(ori_ori_n55_), .Y(ori2));
  NO2        o117(.A(ori_ori_n61_), .B(ori_ori_n37_), .Y(ori_ori_n140_));
  INV        o118(.A(i_6_), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n142_));
  NA4        o120(.A(ori_ori_n142_), .B(ori_ori_n75_), .C(ori_ori_n67_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o121(.A(i_8_), .B(i_7_), .Y(ori_ori_n144_));
  NA2        o122(.A(ori_ori_n144_), .B(i_6_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_12_), .B(i_13_), .Y(ori_ori_n146_));
  NAi21      o124(.An(i_5_), .B(i_11_), .Y(ori_ori_n147_));
  NOi21      o125(.An(ori_ori_n146_), .B(ori_ori_n147_), .Y(ori_ori_n148_));
  NO2        o126(.A(i_0_), .B(i_1_), .Y(ori_ori_n149_));
  NA2        o127(.A(i_2_), .B(i_3_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n150_), .B(i_4_), .Y(ori_ori_n151_));
  NA3        o129(.A(ori_ori_n151_), .B(ori_ori_n149_), .C(ori_ori_n148_), .Y(ori_ori_n152_));
  AN2        o130(.A(ori_ori_n146_), .B(ori_ori_n81_), .Y(ori_ori_n153_));
  NA2        o131(.A(i_1_), .B(i_5_), .Y(ori_ori_n154_));
  OR2        o132(.A(i_0_), .B(i_1_), .Y(ori_ori_n155_));
  NO3        o133(.A(ori_ori_n155_), .B(ori_ori_n78_), .C(i_13_), .Y(ori_ori_n156_));
  NAi32      o134(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n157_));
  NAi21      o135(.An(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  NOi21      o136(.An(i_4_), .B(i_10_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n159_), .B(ori_ori_n40_), .Y(ori_ori_n160_));
  NOi21      o138(.An(i_4_), .B(i_9_), .Y(ori_ori_n161_));
  NOi21      o139(.An(i_11_), .B(i_13_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n162_), .B(ori_ori_n161_), .Y(ori_ori_n163_));
  NO2        o141(.A(i_4_), .B(i_5_), .Y(ori_ori_n164_));
  NAi21      o142(.An(i_12_), .B(i_11_), .Y(ori_ori_n165_));
  NO2        o143(.A(ori_ori_n71_), .B(ori_ori_n61_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n166_), .B(ori_ori_n46_), .Y(ori_ori_n167_));
  NA2        o145(.A(i_3_), .B(i_5_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n71_), .B(i_5_), .Y(ori_ori_n169_));
  NO2        o147(.A(i_13_), .B(i_10_), .Y(ori_ori_n170_));
  NA3        o148(.A(ori_ori_n170_), .B(ori_ori_n169_), .C(ori_ori_n44_), .Y(ori_ori_n171_));
  NO2        o149(.A(i_2_), .B(i_1_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(i_3_), .Y(ori_ori_n173_));
  NAi21      o151(.An(i_4_), .B(i_12_), .Y(ori_ori_n174_));
  INV        o152(.A(i_8_), .Y(ori_ori_n175_));
  NO3        o153(.A(i_3_), .B(ori_ori_n84_), .C(ori_ori_n48_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(ori_ori_n114_), .Y(ori_ori_n177_));
  NO3        o155(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n178_));
  NO3        o156(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n179_));
  NO2        o157(.A(i_3_), .B(i_8_), .Y(ori_ori_n180_));
  NO3        o158(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n181_));
  NA3        o159(.A(ori_ori_n181_), .B(ori_ori_n180_), .C(ori_ori_n40_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n183_));
  INV        o161(.A(ori_ori_n183_), .Y(ori_ori_n184_));
  NO2        o162(.A(i_13_), .B(i_9_), .Y(ori_ori_n185_));
  NAi21      o163(.An(i_12_), .B(i_3_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n184_), .B(ori_ori_n182_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n188_), .B(i_7_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n189_), .B(i_4_), .Y(ori_ori_n190_));
  NAi21      o168(.An(i_12_), .B(i_7_), .Y(ori_ori_n191_));
  NA3        o169(.A(i_13_), .B(ori_ori_n175_), .C(i_10_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n192_), .B(ori_ori_n191_), .Y(ori_ori_n193_));
  NA2        o171(.A(i_0_), .B(i_5_), .Y(ori_ori_n194_));
  OAI220     o172(.A0(ori_ori_n84_), .A1(ori_ori_n173_), .B0(ori_ori_n167_), .B1(ori_ori_n135_), .Y(ori_ori_n195_));
  NAi31      o173(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n71_), .B(ori_ori_n26_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n46_), .B(ori_ori_n61_), .Y(ori_ori_n199_));
  NA3        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .C(ori_ori_n197_), .Y(ori_ori_n200_));
  INV        o178(.A(i_13_), .Y(ori_ori_n201_));
  NO2        o179(.A(i_12_), .B(ori_ori_n201_), .Y(ori_ori_n202_));
  NA3        o180(.A(ori_ori_n202_), .B(ori_ori_n178_), .C(ori_ori_n176_), .Y(ori_ori_n203_));
  OAI210     o181(.A0(ori_ori_n200_), .A1(ori_ori_n196_), .B0(ori_ori_n203_), .Y(ori_ori_n204_));
  AOI220     o182(.A0(ori_ori_n204_), .A1(ori_ori_n144_), .B0(ori_ori_n195_), .B1(ori_ori_n193_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n206_));
  OR2        o184(.A(i_8_), .B(i_7_), .Y(ori_ori_n207_));
  INV        o185(.A(i_12_), .Y(ori_ori_n208_));
  NO2        o186(.A(ori_ori_n44_), .B(ori_ori_n208_), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n210_));
  NA2        o188(.A(i_2_), .B(i_1_), .Y(ori_ori_n211_));
  NO3        o189(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n212_));
  NAi21      o190(.An(i_4_), .B(i_3_), .Y(ori_ori_n213_));
  NO2        o191(.A(i_0_), .B(i_6_), .Y(ori_ori_n214_));
  NOi41      o192(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n211_), .B(ori_ori_n168_), .Y(ori_ori_n216_));
  NO2        o194(.A(i_11_), .B(ori_ori_n201_), .Y(ori_ori_n217_));
  NOi21      o195(.An(i_1_), .B(i_6_), .Y(ori_ori_n218_));
  NAi21      o196(.An(i_3_), .B(i_7_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n208_), .B(i_9_), .Y(ori_ori_n220_));
  OR4        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .C(ori_ori_n218_), .D(ori_ori_n169_), .Y(ori_ori_n221_));
  NA2        o199(.A(ori_ori_n71_), .B(i_5_), .Y(ori_ori_n222_));
  NA2        o200(.A(i_3_), .B(i_9_), .Y(ori_ori_n223_));
  NAi21      o201(.An(i_7_), .B(i_10_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n224_), .B(ori_ori_n223_), .Y(ori_ori_n225_));
  NA3        o203(.A(ori_ori_n225_), .B(ori_ori_n222_), .C(ori_ori_n62_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n226_), .B(ori_ori_n221_), .Y(ori_ori_n227_));
  INV        o205(.A(ori_ori_n145_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n208_), .B(i_13_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n229_), .B(ori_ori_n73_), .Y(ori_ori_n230_));
  AOI220     o208(.A0(ori_ori_n230_), .A1(ori_ori_n228_), .B0(ori_ori_n227_), .B1(ori_ori_n217_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n207_), .B(ori_ori_n37_), .Y(ori_ori_n232_));
  NA2        o210(.A(i_12_), .B(i_6_), .Y(ori_ori_n233_));
  OR2        o211(.A(i_13_), .B(i_9_), .Y(ori_ori_n234_));
  NO3        o212(.A(ori_ori_n234_), .B(ori_ori_n233_), .C(ori_ori_n48_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n213_), .B(i_2_), .Y(ori_ori_n236_));
  NA3        o214(.A(ori_ori_n236_), .B(ori_ori_n235_), .C(ori_ori_n44_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n217_), .B(i_9_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n222_), .B(ori_ori_n62_), .Y(ori_ori_n239_));
  OAI210     o217(.A0(ori_ori_n239_), .A1(ori_ori_n238_), .B0(ori_ori_n237_), .Y(ori_ori_n240_));
  NO3        o218(.A(i_11_), .B(ori_ori_n201_), .C(ori_ori_n25_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n219_), .B(i_8_), .Y(ori_ori_n242_));
  NO2        o220(.A(i_6_), .B(ori_ori_n48_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n240_), .B(ori_ori_n232_), .Y(ori_ori_n244_));
  NA3        o222(.A(ori_ori_n244_), .B(ori_ori_n231_), .C(ori_ori_n205_), .Y(ori_ori_n245_));
  NO3        o223(.A(i_12_), .B(ori_ori_n201_), .C(ori_ori_n37_), .Y(ori_ori_n246_));
  INV        o224(.A(ori_ori_n246_), .Y(ori_ori_n247_));
  NO3        o225(.A(i_0_), .B(i_2_), .C(ori_ori_n61_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n211_), .B(i_0_), .Y(ori_ori_n249_));
  AOI220     o227(.A0(ori_ori_n249_), .A1(i_8_), .B0(ori_ori_n248_), .B1(ori_ori_n144_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n243_), .B(ori_ori_n26_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n251_), .B(ori_ori_n250_), .Y(ori_ori_n252_));
  INV        o230(.A(ori_ori_n252_), .Y(ori_ori_n253_));
  NO2        o231(.A(i_3_), .B(i_10_), .Y(ori_ori_n254_));
  NO2        o232(.A(i_2_), .B(ori_ori_n102_), .Y(ori_ori_n255_));
  NA2        o233(.A(i_1_), .B(ori_ori_n36_), .Y(ori_ori_n256_));
  AN2        o234(.A(i_3_), .B(i_10_), .Y(ori_ori_n257_));
  NO2        o235(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n258_));
  NO2        o236(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n253_), .B(ori_ori_n247_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n260_), .B(ori_ori_n245_), .C(ori_ori_n190_), .Y(ori_ori_n261_));
  NO3        o239(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n262_));
  NO3        o240(.A(i_6_), .B(ori_ori_n175_), .C(i_7_), .Y(ori_ori_n263_));
  NO2        o241(.A(i_2_), .B(i_3_), .Y(ori_ori_n264_));
  OR2        o242(.A(i_0_), .B(i_5_), .Y(ori_ori_n265_));
  NA2        o243(.A(ori_ori_n194_), .B(ori_ori_n265_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n155_), .B(ori_ori_n46_), .Y(ori_ori_n267_));
  NO2        o245(.A(i_12_), .B(i_10_), .Y(ori_ori_n268_));
  NOi21      o246(.An(i_5_), .B(i_0_), .Y(ori_ori_n269_));
  NO2        o247(.A(i_2_), .B(ori_ori_n102_), .Y(ori_ori_n270_));
  NO4        o248(.A(ori_ori_n270_), .B(ori_ori_n256_), .C(ori_ori_n269_), .D(ori_ori_n130_), .Y(ori_ori_n271_));
  NA4        o249(.A(ori_ori_n82_), .B(ori_ori_n36_), .C(ori_ori_n84_), .D(i_8_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n271_), .B(ori_ori_n268_), .Y(ori_ori_n273_));
  NO2        o251(.A(i_6_), .B(i_8_), .Y(ori_ori_n274_));
  NOi21      o252(.An(i_0_), .B(i_2_), .Y(ori_ori_n275_));
  AN2        o253(.A(ori_ori_n275_), .B(ori_ori_n274_), .Y(ori_ori_n276_));
  NO2        o254(.A(i_1_), .B(i_7_), .Y(ori_ori_n277_));
  NA3        o255(.A(ori_ori_n218_), .B(ori_ori_n255_), .C(ori_ori_n175_), .Y(ori_ori_n278_));
  NO2        o256(.A(ori_ori_n278_), .B(ori_ori_n266_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n279_), .B(i_3_), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n175_), .B(i_9_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n281_), .B(ori_ori_n183_), .Y(ori_ori_n282_));
  NO2        o260(.A(ori_ori_n282_), .B(ori_ori_n46_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n283_), .B(ori_ori_n252_), .Y(ori_ori_n284_));
  AOI210     o262(.A0(ori_ori_n284_), .A1(ori_ori_n280_), .B0(ori_ori_n160_), .Y(ori_ori_n285_));
  AOI210     o263(.A0(ori_ori_n871_), .A1(ori_ori_n262_), .B0(ori_ori_n285_), .Y(ori_ori_n286_));
  NOi32      o264(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n287_), .Y(ori_ori_n288_));
  NAi21      o266(.An(i_0_), .B(i_6_), .Y(ori_ori_n289_));
  NAi21      o267(.An(i_1_), .B(i_5_), .Y(ori_ori_n290_));
  NAi41      o268(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n291_));
  OAI220     o269(.A0(ori_ori_n291_), .A1(ori_ori_n290_), .B0(ori_ori_n196_), .B1(ori_ori_n157_), .Y(ori_ori_n292_));
  AOI210     o270(.A0(ori_ori_n291_), .A1(ori_ori_n157_), .B0(ori_ori_n155_), .Y(ori_ori_n293_));
  NOi32      o271(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n294_));
  NAi21      o272(.An(i_6_), .B(i_1_), .Y(ori_ori_n295_));
  NA3        o273(.A(ori_ori_n295_), .B(ori_ori_n294_), .C(ori_ori_n46_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n296_), .B(i_0_), .Y(ori_ori_n297_));
  OR3        o275(.A(ori_ori_n297_), .B(ori_ori_n293_), .C(ori_ori_n292_), .Y(ori_ori_n298_));
  NO2        o276(.A(i_1_), .B(ori_ori_n102_), .Y(ori_ori_n299_));
  NAi21      o277(.An(i_3_), .B(i_4_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n300_), .B(i_9_), .Y(ori_ori_n301_));
  AN2        o279(.A(i_6_), .B(i_7_), .Y(ori_ori_n302_));
  OAI210     o280(.A0(ori_ori_n302_), .A1(ori_ori_n299_), .B0(ori_ori_n301_), .Y(ori_ori_n303_));
  NA2        o281(.A(i_2_), .B(i_7_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n300_), .B(i_10_), .Y(ori_ori_n305_));
  NA3        o283(.A(ori_ori_n305_), .B(ori_ori_n304_), .C(ori_ori_n214_), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n306_), .A1(ori_ori_n303_), .B0(ori_ori_n169_), .Y(ori_ori_n307_));
  AOI210     o285(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n308_));
  OAI210     o286(.A0(ori_ori_n308_), .A1(ori_ori_n172_), .B0(ori_ori_n305_), .Y(ori_ori_n309_));
  AOI220     o287(.A0(ori_ori_n305_), .A1(ori_ori_n277_), .B0(ori_ori_n210_), .B1(ori_ori_n172_), .Y(ori_ori_n310_));
  AOI210     o288(.A0(ori_ori_n310_), .A1(ori_ori_n309_), .B0(i_5_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n311_), .B(ori_ori_n307_), .C(ori_ori_n298_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n312_), .B(ori_ori_n288_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n57_), .B(ori_ori_n25_), .Y(ori_ori_n314_));
  AN2        o292(.A(i_12_), .B(i_5_), .Y(ori_ori_n315_));
  NO2        o293(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n316_), .B(ori_ori_n315_), .Y(ori_ori_n317_));
  NO2        o295(.A(i_11_), .B(i_6_), .Y(ori_ori_n318_));
  NA3        o296(.A(ori_ori_n318_), .B(ori_ori_n267_), .C(ori_ori_n201_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n319_), .B(ori_ori_n317_), .Y(ori_ori_n320_));
  NO2        o298(.A(i_5_), .B(i_10_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n321_), .B(ori_ori_n236_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n146_), .B(ori_ori_n45_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n323_), .B(ori_ori_n322_), .Y(ori_ori_n324_));
  OAI210     o302(.A0(ori_ori_n324_), .A1(ori_ori_n320_), .B0(ori_ori_n314_), .Y(ori_ori_n325_));
  NO2        o303(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n326_));
  NO2        o304(.A(ori_ori_n152_), .B(ori_ori_n84_), .Y(ori_ori_n327_));
  OAI210     o305(.A0(ori_ori_n327_), .A1(ori_ori_n320_), .B0(ori_ori_n326_), .Y(ori_ori_n328_));
  NO3        o306(.A(ori_ori_n84_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n329_));
  NA3        o307(.A(ori_ori_n254_), .B(ori_ori_n91_), .C(ori_ori_n73_), .Y(ori_ori_n330_));
  NO2        o308(.A(i_11_), .B(i_12_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n331_), .B(ori_ori_n36_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n330_), .B(ori_ori_n332_), .Y(ori_ori_n333_));
  NA2        o311(.A(ori_ori_n321_), .B(ori_ori_n208_), .Y(ori_ori_n334_));
  NAi21      o312(.An(i_13_), .B(i_0_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n335_), .B(ori_ori_n211_), .Y(ori_ori_n336_));
  NA2        o314(.A(ori_ori_n333_), .B(ori_ori_n336_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n337_), .B(ori_ori_n328_), .C(ori_ori_n325_), .Y(ori_ori_n338_));
  NA2        o316(.A(ori_ori_n44_), .B(ori_ori_n201_), .Y(ori_ori_n339_));
  NO3        o317(.A(i_1_), .B(i_12_), .C(ori_ori_n84_), .Y(ori_ori_n340_));
  NO2        o318(.A(i_0_), .B(i_11_), .Y(ori_ori_n341_));
  NOi21      o319(.An(i_2_), .B(i_12_), .Y(ori_ori_n342_));
  NAi21      o320(.An(i_9_), .B(i_4_), .Y(ori_ori_n343_));
  OR2        o321(.A(i_13_), .B(i_10_), .Y(ori_ori_n344_));
  NO3        o322(.A(ori_ori_n344_), .B(ori_ori_n119_), .C(ori_ori_n343_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n163_), .B(ori_ori_n125_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n102_), .B(ori_ori_n25_), .Y(ori_ori_n347_));
  NO2        o325(.A(ori_ori_n168_), .B(ori_ori_n84_), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n175_), .B(i_10_), .Y(ori_ori_n349_));
  NA3        o327(.A(ori_ori_n222_), .B(ori_ori_n62_), .C(i_2_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n350_), .B(ori_ori_n349_), .Y(ori_ori_n351_));
  NO2        o329(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n352_));
  NA3        o330(.A(ori_ori_n277_), .B(ori_ori_n276_), .C(ori_ori_n352_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n263_), .B(ori_ori_n266_), .Y(ori_ori_n354_));
  OAI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n173_), .B0(ori_ori_n353_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n355_), .B(ori_ori_n351_), .Y(ori_ori_n356_));
  NO2        o334(.A(ori_ori_n356_), .B(ori_ori_n238_), .Y(ori_ori_n357_));
  NO3        o335(.A(ori_ori_n357_), .B(ori_ori_n338_), .C(ori_ori_n313_), .Y(ori_ori_n358_));
  NO2        o336(.A(ori_ori_n71_), .B(i_13_), .Y(ori_ori_n359_));
  NO2        o337(.A(i_10_), .B(i_9_), .Y(ori_ori_n360_));
  NAi21      o338(.An(i_12_), .B(i_8_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n361_), .B(i_3_), .Y(ori_ori_n362_));
  NO2        o340(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n363_));
  NA2        o341(.A(ori_ori_n363_), .B(ori_ori_n105_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n364_), .B(ori_ori_n182_), .Y(ori_ori_n365_));
  NA2        o343(.A(ori_ori_n259_), .B(i_0_), .Y(ori_ori_n366_));
  NO3        o344(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n367_));
  NA2        o345(.A(ori_ori_n233_), .B(ori_ori_n98_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n369_));
  NA2        o347(.A(i_8_), .B(i_9_), .Y(ori_ori_n370_));
  AOI210     o348(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n371_));
  OR2        o349(.A(ori_ori_n371_), .B(ori_ori_n370_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n246_), .B(ori_ori_n183_), .Y(ori_ori_n373_));
  OAI220     o351(.A0(ori_ori_n373_), .A1(ori_ori_n372_), .B0(ori_ori_n369_), .B1(ori_ori_n366_), .Y(ori_ori_n374_));
  NA2        o352(.A(ori_ori_n217_), .B(ori_ori_n258_), .Y(ori_ori_n375_));
  NO3        o353(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n376_));
  INV        o354(.A(ori_ori_n376_), .Y(ori_ori_n377_));
  NA3        o355(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n378_));
  NA4        o356(.A(ori_ori_n147_), .B(ori_ori_n117_), .C(ori_ori_n78_), .D(ori_ori_n23_), .Y(ori_ori_n379_));
  OAI220     o357(.A0(ori_ori_n379_), .A1(ori_ori_n378_), .B0(ori_ori_n377_), .B1(ori_ori_n375_), .Y(ori_ori_n380_));
  NO3        o358(.A(ori_ori_n380_), .B(ori_ori_n374_), .C(ori_ori_n365_), .Y(ori_ori_n381_));
  OR2        o359(.A(ori_ori_n282_), .B(ori_ori_n102_), .Y(ori_ori_n382_));
  OR2        o360(.A(ori_ori_n382_), .B(ori_ori_n160_), .Y(ori_ori_n383_));
  NA2        o361(.A(ori_ori_n97_), .B(i_13_), .Y(ori_ori_n384_));
  NA2        o362(.A(ori_ori_n348_), .B(ori_ori_n314_), .Y(ori_ori_n385_));
  NO2        o363(.A(i_2_), .B(i_13_), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n387_));
  NO3        o365(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n388_));
  NO2        o366(.A(i_6_), .B(i_7_), .Y(ori_ori_n389_));
  NO2        o367(.A(i_11_), .B(i_1_), .Y(ori_ori_n390_));
  OR2        o368(.A(i_11_), .B(i_8_), .Y(ori_ori_n391_));
  NOi21      o369(.An(i_2_), .B(i_7_), .Y(ori_ori_n392_));
  NO2        o370(.A(i_6_), .B(i_10_), .Y(ori_ori_n393_));
  NA3        o371(.A(ori_ori_n215_), .B(ori_ori_n162_), .C(ori_ori_n134_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n155_), .B(i_3_), .Y(ori_ori_n396_));
  NAi31      o374(.An(ori_ori_n395_), .B(ori_ori_n396_), .C(ori_ori_n202_), .Y(ori_ori_n397_));
  NA3        o375(.A(ori_ori_n326_), .B(ori_ori_n166_), .C(ori_ori_n151_), .Y(ori_ori_n398_));
  NA3        o376(.A(ori_ori_n398_), .B(ori_ori_n397_), .C(ori_ori_n394_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n399_), .B(ori_ori_n387_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n367_), .B(ori_ori_n315_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n376_), .B(ori_ori_n321_), .Y(ori_ori_n402_));
  NO2        o380(.A(ori_ori_n402_), .B(ori_ori_n200_), .Y(ori_ori_n403_));
  NAi21      o381(.An(ori_ori_n192_), .B(ori_ori_n331_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n277_), .B(ori_ori_n194_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n405_), .B(ori_ori_n404_), .Y(ori_ori_n406_));
  NA2        o384(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n262_), .B(ori_ori_n210_), .Y(ori_ori_n408_));
  OAI220     o386(.A0(ori_ori_n408_), .A1(ori_ori_n350_), .B0(ori_ori_n407_), .B1(ori_ori_n384_), .Y(ori_ori_n409_));
  NO3        o387(.A(ori_ori_n409_), .B(ori_ori_n406_), .C(ori_ori_n403_), .Y(ori_ori_n410_));
  NA4        o388(.A(ori_ori_n410_), .B(ori_ori_n400_), .C(ori_ori_n383_), .D(ori_ori_n381_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n124_), .B(ori_ori_n113_), .Y(ori_ori_n412_));
  AN2        o390(.A(ori_ori_n412_), .B(ori_ori_n367_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n413_), .B(ori_ori_n259_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n287_), .B(ori_ori_n71_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n302_), .B(ori_ori_n294_), .Y(ori_ori_n416_));
  NO2        o394(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n417_));
  AOI210     o395(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n345_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n222_), .B(ori_ori_n62_), .Y(ori_ori_n419_));
  OAI210     o397(.A0(i_8_), .A1(ori_ori_n419_), .B0(ori_ori_n136_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n420_), .B(ori_ori_n346_), .Y(ori_ori_n421_));
  NA3        o399(.A(ori_ori_n421_), .B(ori_ori_n418_), .C(ori_ori_n414_), .Y(ori_ori_n422_));
  NO2        o400(.A(i_12_), .B(ori_ori_n175_), .Y(ori_ori_n423_));
  NO2        o401(.A(i_8_), .B(i_7_), .Y(ori_ori_n424_));
  AOI220     o402(.A0(ori_ori_n348_), .A1(ori_ori_n267_), .B0(ori_ori_n216_), .B1(ori_ori_n214_), .Y(ori_ori_n425_));
  OAI220     o403(.A0(ori_ori_n425_), .A1(ori_ori_n229_), .B0(ori_ori_n384_), .B1(ori_ori_n135_), .Y(ori_ori_n426_));
  NA2        o404(.A(ori_ori_n426_), .B(ori_ori_n232_), .Y(ori_ori_n427_));
  NA3        o405(.A(ori_ori_n257_), .B(ori_ori_n164_), .C(ori_ori_n97_), .Y(ori_ori_n428_));
  NO2        o406(.A(ori_ori_n197_), .B(ori_ori_n44_), .Y(ori_ori_n429_));
  NO2        o407(.A(ori_ori_n155_), .B(i_5_), .Y(ori_ori_n430_));
  NA3        o408(.A(ori_ori_n430_), .B(ori_ori_n339_), .C(ori_ori_n264_), .Y(ori_ori_n431_));
  OAI210     o409(.A0(ori_ori_n431_), .A1(ori_ori_n429_), .B0(ori_ori_n428_), .Y(ori_ori_n432_));
  NA2        o410(.A(ori_ori_n432_), .B(ori_ori_n376_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n433_), .B(ori_ori_n427_), .Y(ori_ori_n434_));
  NA2        o412(.A(ori_ori_n199_), .B(ori_ori_n198_), .Y(ori_ori_n435_));
  NA2        o413(.A(ori_ori_n360_), .B(ori_ori_n197_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n435_), .B(ori_ori_n436_), .Y(ori_ori_n437_));
  AOI210     o415(.A0(ori_ori_n295_), .A1(ori_ori_n46_), .B0(ori_ori_n299_), .Y(ori_ori_n438_));
  NA2        o416(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n439_));
  NA3        o417(.A(ori_ori_n423_), .B(ori_ori_n241_), .C(ori_ori_n439_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n438_), .B(ori_ori_n440_), .Y(ori_ori_n441_));
  NO2        o419(.A(ori_ori_n441_), .B(ori_ori_n437_), .Y(ori_ori_n442_));
  NO4        o420(.A(ori_ori_n218_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n443_));
  NO3        o421(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n444_));
  NO2        o422(.A(ori_ori_n207_), .B(ori_ori_n36_), .Y(ori_ori_n445_));
  NO2        o423(.A(ori_ori_n344_), .B(i_1_), .Y(ori_ori_n446_));
  NOi31      o424(.An(ori_ori_n446_), .B(ori_ori_n368_), .C(ori_ori_n71_), .Y(ori_ori_n447_));
  NOi21      o425(.An(i_10_), .B(i_6_), .Y(ori_ori_n448_));
  NO2        o426(.A(ori_ori_n84_), .B(ori_ori_n25_), .Y(ori_ori_n449_));
  AOI220     o427(.A0(ori_ori_n246_), .A1(ori_ori_n449_), .B0(ori_ori_n241_), .B1(ori_ori_n448_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n450_), .B(ori_ori_n366_), .Y(ori_ori_n451_));
  NO2        o429(.A(ori_ori_n116_), .B(ori_ori_n23_), .Y(ori_ori_n452_));
  NO2        o430(.A(ori_ori_n178_), .B(ori_ori_n37_), .Y(ori_ori_n453_));
  NOi31      o431(.An(ori_ori_n148_), .B(ori_ori_n453_), .C(ori_ori_n272_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n454_), .B(ori_ori_n451_), .Y(ori_ori_n455_));
  NO2        o433(.A(ori_ori_n415_), .B(ori_ori_n310_), .Y(ori_ori_n456_));
  INV        o434(.A(ori_ori_n264_), .Y(ori_ori_n457_));
  NO2        o435(.A(i_12_), .B(ori_ori_n84_), .Y(ori_ori_n458_));
  NA3        o436(.A(ori_ori_n458_), .B(ori_ori_n241_), .C(ori_ori_n439_), .Y(ori_ori_n459_));
  NA3        o437(.A(ori_ori_n318_), .B(ori_ori_n246_), .C(ori_ori_n194_), .Y(ori_ori_n460_));
  AOI210     o438(.A0(ori_ori_n460_), .A1(ori_ori_n459_), .B0(ori_ori_n457_), .Y(ori_ori_n461_));
  OR2        o439(.A(i_2_), .B(i_5_), .Y(ori_ori_n462_));
  OR2        o440(.A(ori_ori_n462_), .B(i_6_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n304_), .B(ori_ori_n214_), .Y(ori_ori_n464_));
  NO2        o442(.A(ori_ori_n464_), .B(ori_ori_n404_), .Y(ori_ori_n465_));
  NO3        o443(.A(ori_ori_n465_), .B(ori_ori_n461_), .C(ori_ori_n456_), .Y(ori_ori_n466_));
  NA3        o444(.A(ori_ori_n466_), .B(ori_ori_n455_), .C(ori_ori_n442_), .Y(ori_ori_n467_));
  NO4        o445(.A(ori_ori_n467_), .B(ori_ori_n434_), .C(ori_ori_n422_), .D(ori_ori_n411_), .Y(ori_ori_n468_));
  NA4        o446(.A(ori_ori_n468_), .B(ori_ori_n358_), .C(ori_ori_n286_), .D(ori_ori_n261_), .Y(ori7));
  NO2        o447(.A(ori_ori_n93_), .B(ori_ori_n54_), .Y(ori_ori_n470_));
  NO2        o448(.A(ori_ori_n109_), .B(ori_ori_n90_), .Y(ori_ori_n471_));
  NA2        o449(.A(ori_ori_n316_), .B(ori_ori_n471_), .Y(ori_ori_n472_));
  NA2        o450(.A(ori_ori_n393_), .B(ori_ori_n82_), .Y(ori_ori_n473_));
  NA2        o451(.A(i_11_), .B(ori_ori_n175_), .Y(ori_ori_n474_));
  NA2        o452(.A(ori_ori_n146_), .B(ori_ori_n474_), .Y(ori_ori_n475_));
  OAI210     o453(.A0(ori_ori_n475_), .A1(ori_ori_n473_), .B0(ori_ori_n472_), .Y(ori_ori_n476_));
  NO2        o454(.A(ori_ori_n208_), .B(i_4_), .Y(ori_ori_n477_));
  NA2        o455(.A(ori_ori_n477_), .B(i_8_), .Y(ori_ori_n478_));
  NA2        o456(.A(i_2_), .B(ori_ori_n84_), .Y(ori_ori_n479_));
  OAI210     o457(.A0(ori_ori_n87_), .A1(ori_ori_n180_), .B0(ori_ori_n181_), .Y(ori_ori_n480_));
  NO2        o458(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n481_));
  NA2        o459(.A(i_4_), .B(i_8_), .Y(ori_ori_n482_));
  AOI210     o460(.A0(ori_ori_n482_), .A1(ori_ori_n257_), .B0(ori_ori_n481_), .Y(ori_ori_n483_));
  OAI220     o461(.A0(ori_ori_n483_), .A1(ori_ori_n479_), .B0(ori_ori_n480_), .B1(i_13_), .Y(ori_ori_n484_));
  NO3        o462(.A(ori_ori_n484_), .B(ori_ori_n476_), .C(ori_ori_n470_), .Y(ori_ori_n485_));
  AOI210     o463(.A0(ori_ori_n130_), .A1(ori_ori_n60_), .B0(i_10_), .Y(ori_ori_n486_));
  AOI210     o464(.A0(ori_ori_n486_), .A1(ori_ori_n208_), .B0(ori_ori_n159_), .Y(ori_ori_n487_));
  OR2        o465(.A(i_6_), .B(i_10_), .Y(ori_ori_n488_));
  OR3        o466(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n489_));
  INV        o467(.A(ori_ori_n179_), .Y(ori_ori_n490_));
  OR2        o468(.A(ori_ori_n487_), .B(ori_ori_n234_), .Y(ori_ori_n491_));
  AOI210     o469(.A0(ori_ori_n491_), .A1(ori_ori_n485_), .B0(ori_ori_n61_), .Y(ori_ori_n492_));
  NOi21      o470(.An(i_11_), .B(i_7_), .Y(ori_ori_n493_));
  AO210      o471(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n494_));
  NO2        o472(.A(ori_ori_n494_), .B(ori_ori_n493_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n495_), .B(ori_ori_n185_), .Y(ori_ori_n496_));
  NA3        o474(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n497_));
  NAi31      o475(.An(ori_ori_n497_), .B(ori_ori_n191_), .C(i_11_), .Y(ori_ori_n498_));
  AOI210     o476(.A0(ori_ori_n498_), .A1(ori_ori_n496_), .B0(ori_ori_n61_), .Y(ori_ori_n499_));
  NA2        o477(.A(ori_ori_n86_), .B(ori_ori_n61_), .Y(ori_ori_n500_));
  AO210      o478(.A0(ori_ori_n500_), .A1(ori_ori_n310_), .B0(ori_ori_n41_), .Y(ori_ori_n501_));
  NO3        o479(.A(ori_ori_n224_), .B(ori_ori_n186_), .C(ori_ori_n474_), .Y(ori_ori_n502_));
  OAI210     o480(.A0(ori_ori_n502_), .A1(ori_ori_n202_), .B0(ori_ori_n61_), .Y(ori_ori_n503_));
  NA2        o481(.A(ori_ori_n342_), .B(ori_ori_n31_), .Y(ori_ori_n504_));
  OR2        o482(.A(ori_ori_n186_), .B(ori_ori_n109_), .Y(ori_ori_n505_));
  NA2        o483(.A(ori_ori_n505_), .B(ori_ori_n504_), .Y(ori_ori_n506_));
  NO2        o484(.A(ori_ori_n61_), .B(i_9_), .Y(ori_ori_n507_));
  NO2        o485(.A(ori_ori_n507_), .B(i_4_), .Y(ori_ori_n508_));
  NA2        o486(.A(ori_ori_n508_), .B(ori_ori_n506_), .Y(ori_ori_n509_));
  NO2        o487(.A(i_1_), .B(i_12_), .Y(ori_ori_n510_));
  NA3        o488(.A(ori_ori_n510_), .B(ori_ori_n111_), .C(ori_ori_n24_), .Y(ori_ori_n511_));
  BUFFER     o489(.A(ori_ori_n511_), .Y(ori_ori_n512_));
  NA4        o490(.A(ori_ori_n512_), .B(ori_ori_n509_), .C(ori_ori_n503_), .D(ori_ori_n501_), .Y(ori_ori_n513_));
  OAI210     o491(.A0(ori_ori_n513_), .A1(ori_ori_n499_), .B0(i_6_), .Y(ori_ori_n514_));
  NO2        o492(.A(ori_ori_n208_), .B(ori_ori_n84_), .Y(ori_ori_n515_));
  NO2        o493(.A(ori_ori_n515_), .B(i_11_), .Y(ori_ori_n516_));
  INV        o494(.A(ori_ori_n369_), .Y(ori_ori_n517_));
  NO3        o495(.A(ori_ori_n488_), .B(ori_ori_n207_), .C(ori_ori_n23_), .Y(ori_ori_n518_));
  AOI210     o496(.A0(i_1_), .A1(ori_ori_n225_), .B0(ori_ori_n518_), .Y(ori_ori_n519_));
  NO2        o497(.A(ori_ori_n519_), .B(ori_ori_n44_), .Y(ori_ori_n520_));
  NA3        o498(.A(ori_ori_n424_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n521_));
  INV        o499(.A(i_2_), .Y(ori_ori_n522_));
  NA2        o500(.A(ori_ori_n140_), .B(i_9_), .Y(ori_ori_n523_));
  NA3        o501(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n524_));
  NO2        o502(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n525_));
  NO2        o503(.A(ori_ori_n523_), .B(ori_ori_n522_), .Y(ori_ori_n526_));
  NA3        o504(.A(ori_ori_n507_), .B(ori_ori_n264_), .C(i_6_), .Y(ori_ori_n527_));
  NO2        o505(.A(ori_ori_n527_), .B(ori_ori_n23_), .Y(ori_ori_n528_));
  AOI210     o506(.A0(ori_ori_n390_), .A1(ori_ori_n347_), .B0(ori_ori_n212_), .Y(ori_ori_n529_));
  NO2        o507(.A(ori_ori_n529_), .B(ori_ori_n479_), .Y(ori_ori_n530_));
  NAi21      o508(.An(ori_ori_n521_), .B(ori_ori_n92_), .Y(ori_ori_n531_));
  NA2        o509(.A(ori_ori_n525_), .B(ori_ori_n233_), .Y(ori_ori_n532_));
  NO2        o510(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n533_));
  NA2        o511(.A(ori_ori_n533_), .B(ori_ori_n24_), .Y(ori_ori_n534_));
  OAI210     o512(.A0(ori_ori_n534_), .A1(ori_ori_n532_), .B0(ori_ori_n531_), .Y(ori_ori_n535_));
  OR4        o513(.A(ori_ori_n535_), .B(ori_ori_n530_), .C(ori_ori_n528_), .D(ori_ori_n526_), .Y(ori_ori_n536_));
  NO3        o514(.A(ori_ori_n536_), .B(ori_ori_n520_), .C(ori_ori_n517_), .Y(ori_ori_n537_));
  NO2        o515(.A(ori_ori_n208_), .B(ori_ori_n102_), .Y(ori_ori_n538_));
  NO2        o516(.A(ori_ori_n538_), .B(ori_ori_n493_), .Y(ori_ori_n539_));
  NA2        o517(.A(ori_ori_n539_), .B(i_1_), .Y(ori_ori_n540_));
  NO2        o518(.A(ori_ori_n540_), .B(ori_ori_n489_), .Y(ori_ori_n541_));
  NO2        o519(.A(ori_ori_n343_), .B(ori_ori_n84_), .Y(ori_ori_n542_));
  NA2        o520(.A(ori_ori_n541_), .B(ori_ori_n46_), .Y(ori_ori_n543_));
  NO2        o521(.A(ori_ori_n207_), .B(ori_ori_n44_), .Y(ori_ori_n544_));
  NO3        o522(.A(ori_ori_n544_), .B(ori_ori_n259_), .C(ori_ori_n209_), .Y(ori_ori_n545_));
  NO2        o523(.A(ori_ori_n119_), .B(ori_ori_n37_), .Y(ori_ori_n546_));
  NO2        o524(.A(ori_ori_n546_), .B(i_6_), .Y(ori_ori_n547_));
  NO2        o525(.A(ori_ori_n84_), .B(i_9_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n548_), .B(ori_ori_n61_), .Y(ori_ori_n549_));
  NO2        o527(.A(ori_ori_n549_), .B(ori_ori_n510_), .Y(ori_ori_n550_));
  NO4        o528(.A(ori_ori_n550_), .B(ori_ori_n547_), .C(ori_ori_n545_), .D(i_4_), .Y(ori_ori_n551_));
  NA2        o529(.A(i_1_), .B(i_3_), .Y(ori_ori_n552_));
  INV        o530(.A(ori_ori_n551_), .Y(ori_ori_n553_));
  NA4        o531(.A(ori_ori_n553_), .B(ori_ori_n543_), .C(ori_ori_n537_), .D(ori_ori_n514_), .Y(ori_ori_n554_));
  NO3        o532(.A(ori_ori_n391_), .B(i_3_), .C(i_7_), .Y(ori_ori_n555_));
  NOi21      o533(.An(ori_ori_n555_), .B(i_10_), .Y(ori_ori_n556_));
  OA210      o534(.A0(ori_ori_n556_), .A1(ori_ori_n215_), .B0(ori_ori_n84_), .Y(ori_ori_n557_));
  NA3        o535(.A(ori_ori_n393_), .B(ori_ori_n417_), .C(ori_ori_n46_), .Y(ori_ori_n558_));
  NO3        o536(.A(ori_ori_n392_), .B(ori_ori_n482_), .C(ori_ori_n84_), .Y(ori_ori_n559_));
  NA2        o537(.A(ori_ori_n559_), .B(ori_ori_n25_), .Y(ori_ori_n560_));
  NA3        o538(.A(ori_ori_n159_), .B(ori_ori_n82_), .C(ori_ori_n84_), .Y(ori_ori_n561_));
  NA3        o539(.A(ori_ori_n561_), .B(ori_ori_n560_), .C(ori_ori_n558_), .Y(ori_ori_n562_));
  OAI210     o540(.A0(ori_ori_n562_), .A1(ori_ori_n557_), .B0(i_1_), .Y(ori_ori_n563_));
  AOI210     o541(.A0(ori_ori_n233_), .A1(ori_ori_n98_), .B0(i_1_), .Y(ori_ori_n564_));
  NO2        o542(.A(ori_ori_n300_), .B(i_2_), .Y(ori_ori_n565_));
  NA2        o543(.A(ori_ori_n565_), .B(ori_ori_n564_), .Y(ori_ori_n566_));
  OAI210     o544(.A0(ori_ori_n527_), .A1(ori_ori_n361_), .B0(ori_ori_n566_), .Y(ori_ori_n567_));
  INV        o545(.A(ori_ori_n567_), .Y(ori_ori_n568_));
  AOI210     o546(.A0(ori_ori_n568_), .A1(ori_ori_n563_), .B0(i_13_), .Y(ori_ori_n569_));
  OR2        o547(.A(i_11_), .B(i_7_), .Y(ori_ori_n570_));
  NA3        o548(.A(ori_ori_n570_), .B(ori_ori_n107_), .C(ori_ori_n140_), .Y(ori_ori_n571_));
  AOI220     o549(.A0(ori_ori_n386_), .A1(ori_ori_n159_), .B0(ori_ori_n363_), .B1(ori_ori_n140_), .Y(ori_ori_n572_));
  OAI210     o550(.A0(ori_ori_n572_), .A1(ori_ori_n44_), .B0(ori_ori_n571_), .Y(ori_ori_n573_));
  NO2        o551(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n574_));
  NO2        o552(.A(ori_ori_n392_), .B(ori_ori_n24_), .Y(ori_ori_n575_));
  NA2        o553(.A(ori_ori_n575_), .B(ori_ori_n542_), .Y(ori_ori_n576_));
  OAI220     o554(.A0(ori_ori_n576_), .A1(ori_ori_n41_), .B0(ori_ori_n870_), .B1(ori_ori_n93_), .Y(ori_ori_n577_));
  AOI210     o555(.A0(ori_ori_n573_), .A1(ori_ori_n274_), .B0(ori_ori_n577_), .Y(ori_ori_n578_));
  INV        o556(.A(ori_ori_n116_), .Y(ori_ori_n579_));
  AOI220     o557(.A0(ori_ori_n579_), .A1(ori_ori_n70_), .B0(ori_ori_n318_), .B1(ori_ori_n525_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n580_), .B(ori_ori_n213_), .Y(ori_ori_n581_));
  NA2        o559(.A(ori_ori_n129_), .B(i_13_), .Y(ori_ori_n582_));
  NO2        o560(.A(ori_ori_n524_), .B(ori_ori_n116_), .Y(ori_ori_n583_));
  INV        o561(.A(ori_ori_n583_), .Y(ori_ori_n584_));
  OAI220     o562(.A0(ori_ori_n584_), .A1(ori_ori_n69_), .B0(ori_ori_n582_), .B1(ori_ori_n564_), .Y(ori_ori_n585_));
  NO3        o563(.A(ori_ori_n69_), .B(ori_ori_n32_), .C(ori_ori_n102_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n26_), .B(ori_ori_n175_), .Y(ori_ori_n587_));
  INV        o565(.A(i_7_), .Y(ori_ori_n588_));
  AOI220     o566(.A0(ori_ori_n318_), .A1(ori_ori_n525_), .B0(ori_ori_n92_), .B1(ori_ori_n103_), .Y(ori_ori_n589_));
  OAI220     o567(.A0(ori_ori_n589_), .A1(ori_ori_n478_), .B0(ori_ori_n872_), .B1(ori_ori_n490_), .Y(ori_ori_n590_));
  NO3        o568(.A(ori_ori_n590_), .B(ori_ori_n585_), .C(ori_ori_n581_), .Y(ori_ori_n591_));
  OR2        o569(.A(i_11_), .B(i_6_), .Y(ori_ori_n592_));
  NA3        o570(.A(ori_ori_n477_), .B(ori_ori_n587_), .C(i_7_), .Y(ori_ori_n593_));
  AOI210     o571(.A0(ori_ori_n593_), .A1(ori_ori_n584_), .B0(ori_ori_n592_), .Y(ori_ori_n594_));
  NA3        o572(.A(ori_ori_n342_), .B(ori_ori_n481_), .C(ori_ori_n98_), .Y(ori_ori_n595_));
  NA2        o573(.A(ori_ori_n516_), .B(i_13_), .Y(ori_ori_n596_));
  NA2        o574(.A(ori_ori_n103_), .B(ori_ori_n587_), .Y(ori_ori_n597_));
  NAi21      o575(.An(i_11_), .B(i_12_), .Y(ori_ori_n598_));
  NOi41      o576(.An(ori_ori_n112_), .B(ori_ori_n598_), .C(i_13_), .D(ori_ori_n84_), .Y(ori_ori_n599_));
  NO3        o577(.A(ori_ori_n392_), .B(ori_ori_n458_), .C(ori_ori_n482_), .Y(ori_ori_n600_));
  AOI220     o578(.A0(ori_ori_n600_), .A1(ori_ori_n262_), .B0(ori_ori_n599_), .B1(ori_ori_n597_), .Y(ori_ori_n601_));
  NA3        o579(.A(ori_ori_n601_), .B(ori_ori_n596_), .C(ori_ori_n595_), .Y(ori_ori_n602_));
  OAI210     o580(.A0(ori_ori_n602_), .A1(ori_ori_n594_), .B0(ori_ori_n61_), .Y(ori_ori_n603_));
  NO2        o581(.A(i_2_), .B(i_12_), .Y(ori_ori_n604_));
  NA2        o582(.A(ori_ori_n299_), .B(ori_ori_n604_), .Y(ori_ori_n605_));
  INV        o583(.A(ori_ori_n605_), .Y(ori_ori_n606_));
  NA3        o584(.A(ori_ori_n606_), .B(ori_ori_n45_), .C(ori_ori_n201_), .Y(ori_ori_n607_));
  NA4        o585(.A(ori_ori_n607_), .B(ori_ori_n603_), .C(ori_ori_n591_), .D(ori_ori_n578_), .Y(ori_ori_n608_));
  OR4        o586(.A(ori_ori_n608_), .B(ori_ori_n569_), .C(ori_ori_n554_), .D(ori_ori_n492_), .Y(ori5));
  NA2        o587(.A(ori_ori_n539_), .B(ori_ori_n236_), .Y(ori_ori_n610_));
  AN2        o588(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n611_));
  NA3        o589(.A(ori_ori_n611_), .B(ori_ori_n604_), .C(ori_ori_n109_), .Y(ori_ori_n612_));
  NO2        o590(.A(ori_ori_n478_), .B(i_11_), .Y(ori_ori_n613_));
  NA2        o591(.A(ori_ori_n87_), .B(ori_ori_n613_), .Y(ori_ori_n614_));
  NA3        o592(.A(ori_ori_n614_), .B(ori_ori_n612_), .C(ori_ori_n610_), .Y(ori_ori_n615_));
  NO3        o593(.A(i_11_), .B(ori_ori_n208_), .C(i_13_), .Y(ori_ori_n616_));
  NO2        o594(.A(ori_ori_n126_), .B(ori_ori_n23_), .Y(ori_ori_n617_));
  NA2        o595(.A(i_12_), .B(i_8_), .Y(ori_ori_n618_));
  OAI210     o596(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n618_), .Y(ori_ori_n619_));
  INV        o597(.A(ori_ori_n360_), .Y(ori_ori_n620_));
  AOI220     o598(.A0(ori_ori_n264_), .A1(ori_ori_n452_), .B0(ori_ori_n619_), .B1(ori_ori_n617_), .Y(ori_ori_n621_));
  INV        o599(.A(ori_ori_n621_), .Y(ori_ori_n622_));
  NO2        o600(.A(ori_ori_n622_), .B(ori_ori_n615_), .Y(ori_ori_n623_));
  INV        o601(.A(ori_ori_n162_), .Y(ori_ori_n624_));
  INV        o602(.A(ori_ori_n215_), .Y(ori_ori_n625_));
  OAI210     o603(.A0(ori_ori_n565_), .A1(ori_ori_n362_), .B0(ori_ori_n112_), .Y(ori_ori_n626_));
  AOI210     o604(.A0(ori_ori_n626_), .A1(ori_ori_n625_), .B0(ori_ori_n624_), .Y(ori_ori_n627_));
  NO2        o605(.A(ori_ori_n370_), .B(ori_ori_n26_), .Y(ori_ori_n628_));
  NO2        o606(.A(ori_ori_n628_), .B(ori_ori_n347_), .Y(ori_ori_n629_));
  NA2        o607(.A(ori_ori_n629_), .B(i_2_), .Y(ori_ori_n630_));
  INV        o608(.A(ori_ori_n630_), .Y(ori_ori_n631_));
  AOI210     o609(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n344_), .Y(ori_ori_n632_));
  AOI210     o610(.A0(ori_ori_n632_), .A1(ori_ori_n631_), .B0(ori_ori_n627_), .Y(ori_ori_n633_));
  NO2        o611(.A(ori_ori_n174_), .B(ori_ori_n127_), .Y(ori_ori_n634_));
  OAI210     o612(.A0(ori_ori_n634_), .A1(ori_ori_n617_), .B0(i_2_), .Y(ori_ori_n635_));
  INV        o613(.A(ori_ori_n163_), .Y(ori_ori_n636_));
  NO3        o614(.A(ori_ori_n494_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n637_));
  AOI210     o615(.A0(ori_ori_n636_), .A1(ori_ori_n87_), .B0(ori_ori_n637_), .Y(ori_ori_n638_));
  AOI210     o616(.A0(ori_ori_n638_), .A1(ori_ori_n635_), .B0(ori_ori_n175_), .Y(ori_ori_n639_));
  OA210      o617(.A0(ori_ori_n495_), .A1(ori_ori_n128_), .B0(i_13_), .Y(ori_ori_n640_));
  NA2        o618(.A(ori_ori_n179_), .B(ori_ori_n180_), .Y(ori_ori_n641_));
  NA2        o619(.A(ori_ori_n153_), .B(ori_ori_n474_), .Y(ori_ori_n642_));
  AOI210     o620(.A0(ori_ori_n642_), .A1(ori_ori_n641_), .B0(ori_ori_n304_), .Y(ori_ori_n643_));
  AOI210     o621(.A0(ori_ori_n186_), .A1(ori_ori_n150_), .B0(ori_ori_n417_), .Y(ori_ori_n644_));
  NA2        o622(.A(ori_ori_n644_), .B(ori_ori_n347_), .Y(ori_ori_n645_));
  NO2        o623(.A(ori_ori_n103_), .B(ori_ori_n44_), .Y(ori_ori_n646_));
  INV        o624(.A(ori_ori_n255_), .Y(ori_ori_n647_));
  NA4        o625(.A(ori_ori_n647_), .B(ori_ori_n257_), .C(ori_ori_n126_), .D(ori_ori_n42_), .Y(ori_ori_n648_));
  OAI210     o626(.A0(ori_ori_n648_), .A1(ori_ori_n646_), .B0(ori_ori_n645_), .Y(ori_ori_n649_));
  NO4        o627(.A(ori_ori_n649_), .B(ori_ori_n643_), .C(ori_ori_n640_), .D(ori_ori_n639_), .Y(ori_ori_n650_));
  NA2        o628(.A(ori_ori_n452_), .B(ori_ori_n28_), .Y(ori_ori_n651_));
  NA2        o629(.A(ori_ori_n616_), .B(ori_ori_n242_), .Y(ori_ori_n652_));
  NA2        o630(.A(ori_ori_n652_), .B(ori_ori_n651_), .Y(ori_ori_n653_));
  NO2        o631(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n654_));
  NO2        o632(.A(ori_ori_n654_), .B(ori_ori_n128_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n655_), .B(ori_ori_n474_), .Y(ori_ori_n656_));
  AOI220     o634(.A0(ori_ori_n656_), .A1(ori_ori_n36_), .B0(ori_ori_n653_), .B1(ori_ori_n46_), .Y(ori_ori_n657_));
  NA4        o635(.A(ori_ori_n657_), .B(ori_ori_n650_), .C(ori_ori_n633_), .D(ori_ori_n623_), .Y(ori6));
  NO2        o636(.A(ori_ori_n196_), .B(ori_ori_n395_), .Y(ori_ori_n659_));
  NO2        o637(.A(i_11_), .B(i_9_), .Y(ori_ori_n660_));
  INV        o638(.A(ori_ori_n269_), .Y(ori_ori_n661_));
  OR2        o639(.A(ori_ori_n661_), .B(i_12_), .Y(ori_ori_n662_));
  NA2        o640(.A(ori_ori_n305_), .B(ori_ori_n277_), .Y(ori_ori_n663_));
  NA2        o641(.A(ori_ori_n458_), .B(ori_ori_n61_), .Y(ori_ori_n664_));
  NA2        o642(.A(ori_ori_n556_), .B(ori_ori_n69_), .Y(ori_ori_n665_));
  BUFFER     o643(.A(ori_ori_n500_), .Y(ori_ori_n666_));
  NA4        o644(.A(ori_ori_n666_), .B(ori_ori_n665_), .C(ori_ori_n664_), .D(ori_ori_n663_), .Y(ori_ori_n667_));
  INV        o645(.A(ori_ori_n177_), .Y(ori_ori_n668_));
  AOI220     o646(.A0(ori_ori_n668_), .A1(ori_ori_n660_), .B0(ori_ori_n667_), .B1(ori_ori_n71_), .Y(ori_ori_n669_));
  INV        o647(.A(ori_ori_n268_), .Y(ori_ori_n670_));
  NA2        o648(.A(ori_ori_n73_), .B(ori_ori_n133_), .Y(ori_ori_n671_));
  INV        o649(.A(ori_ori_n126_), .Y(ori_ori_n672_));
  NA2        o650(.A(ori_ori_n672_), .B(ori_ori_n46_), .Y(ori_ori_n673_));
  AOI210     o651(.A0(ori_ori_n673_), .A1(ori_ori_n671_), .B0(ori_ori_n670_), .Y(ori_ori_n674_));
  NO2        o652(.A(ori_ori_n218_), .B(i_9_), .Y(ori_ori_n675_));
  NA2        o653(.A(ori_ori_n675_), .B(ori_ori_n654_), .Y(ori_ori_n676_));
  AOI210     o654(.A0(ori_ori_n676_), .A1(ori_ori_n416_), .B0(ori_ori_n169_), .Y(ori_ori_n677_));
  NO2        o655(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n678_));
  NA3        o656(.A(ori_ori_n678_), .B(ori_ori_n389_), .C(ori_ori_n321_), .Y(ori_ori_n679_));
  NAi32      o657(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n680_));
  NO2        o658(.A(ori_ori_n592_), .B(ori_ori_n680_), .Y(ori_ori_n681_));
  OAI210     o659(.A0(ori_ori_n555_), .A1(ori_ori_n445_), .B0(ori_ori_n444_), .Y(ori_ori_n682_));
  NAi31      o660(.An(ori_ori_n681_), .B(ori_ori_n682_), .C(ori_ori_n679_), .Y(ori_ori_n683_));
  OR3        o661(.A(ori_ori_n683_), .B(ori_ori_n677_), .C(ori_ori_n674_), .Y(ori_ori_n684_));
  NO2        o662(.A(ori_ori_n570_), .B(i_2_), .Y(ori_ori_n685_));
  OR2        o663(.A(ori_ori_n495_), .B(ori_ori_n362_), .Y(ori_ori_n686_));
  NA3        o664(.A(ori_ori_n686_), .B(ori_ori_n149_), .C(ori_ori_n67_), .Y(ori_ori_n687_));
  AO210      o665(.A0(ori_ori_n402_), .A1(ori_ori_n620_), .B0(ori_ori_n36_), .Y(ori_ori_n688_));
  NA2        o666(.A(ori_ori_n688_), .B(ori_ori_n687_), .Y(ori_ori_n689_));
  OAI210     o667(.A0(ori_ori_n515_), .A1(i_11_), .B0(ori_ori_n85_), .Y(ori_ori_n690_));
  AOI220     o668(.A0(ori_ori_n690_), .A1(ori_ori_n444_), .B0(ori_ori_n659_), .B1(ori_ori_n588_), .Y(ori_ori_n691_));
  NA3        o669(.A(ori_ori_n304_), .B(ori_ori_n210_), .C(ori_ori_n149_), .Y(ori_ori_n692_));
  NA2        o670(.A(ori_ori_n329_), .B(ori_ori_n68_), .Y(ori_ori_n693_));
  NA4        o671(.A(ori_ori_n693_), .B(ori_ori_n692_), .C(ori_ori_n691_), .D(ori_ori_n480_), .Y(ori_ori_n694_));
  AO210      o672(.A0(ori_ori_n417_), .A1(ori_ori_n46_), .B0(ori_ori_n86_), .Y(ori_ori_n695_));
  NA3        o673(.A(ori_ori_n695_), .B(ori_ori_n393_), .C(ori_ori_n194_), .Y(ori_ori_n696_));
  AOI210     o674(.A0(ori_ori_n362_), .A1(ori_ori_n360_), .B0(ori_ori_n443_), .Y(ori_ori_n697_));
  NO2        o675(.A(ori_ori_n488_), .B(ori_ori_n103_), .Y(ori_ori_n698_));
  OAI210     o676(.A0(ori_ori_n698_), .A1(ori_ori_n113_), .B0(ori_ori_n341_), .Y(ori_ori_n699_));
  NA2        o677(.A(ori_ori_n214_), .B(ori_ori_n46_), .Y(ori_ori_n700_));
  INV        o678(.A(ori_ori_n463_), .Y(ori_ori_n701_));
  NA3        o679(.A(ori_ori_n701_), .B(ori_ori_n268_), .C(i_7_), .Y(ori_ori_n702_));
  NA4        o680(.A(ori_ori_n702_), .B(ori_ori_n699_), .C(ori_ori_n697_), .D(ori_ori_n696_), .Y(ori_ori_n703_));
  NO4        o681(.A(ori_ori_n703_), .B(ori_ori_n694_), .C(ori_ori_n689_), .D(ori_ori_n684_), .Y(ori_ori_n704_));
  NA4        o682(.A(ori_ori_n704_), .B(ori_ori_n669_), .C(ori_ori_n662_), .D(ori_ori_n312_), .Y(ori3));
  NA2        o683(.A(i_12_), .B(i_10_), .Y(ori_ori_n706_));
  NO2        o684(.A(i_11_), .B(ori_ori_n208_), .Y(ori_ori_n707_));
  NA3        o685(.A(ori_ori_n692_), .B(ori_ori_n480_), .C(ori_ori_n303_), .Y(ori_ori_n708_));
  NA2        o686(.A(ori_ori_n708_), .B(ori_ori_n40_), .Y(ori_ori_n709_));
  NOi21      o687(.An(ori_ori_n97_), .B(ori_ori_n629_), .Y(ori_ori_n710_));
  NO3        o688(.A(ori_ori_n505_), .B(ori_ori_n370_), .C(ori_ori_n133_), .Y(ori_ori_n711_));
  NA2        o689(.A(ori_ori_n342_), .B(ori_ori_n45_), .Y(ori_ori_n712_));
  NO2        o690(.A(ori_ori_n711_), .B(ori_ori_n710_), .Y(ori_ori_n713_));
  AOI210     o691(.A0(ori_ori_n713_), .A1(ori_ori_n709_), .B0(ori_ori_n48_), .Y(ori_ori_n714_));
  NO4        o692(.A(ori_ori_n308_), .B(ori_ori_n315_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n715_));
  NA2        o693(.A(ori_ori_n169_), .B(ori_ori_n448_), .Y(ori_ori_n716_));
  NOi21      o694(.An(ori_ori_n716_), .B(ori_ori_n715_), .Y(ori_ori_n717_));
  NO2        o695(.A(ori_ori_n717_), .B(ori_ori_n61_), .Y(ori_ori_n718_));
  NOi21      o696(.An(i_5_), .B(i_9_), .Y(ori_ori_n719_));
  NA2        o697(.A(ori_ori_n719_), .B(ori_ori_n359_), .Y(ori_ori_n720_));
  BUFFER     o698(.A(ori_ori_n233_), .Y(ori_ori_n721_));
  AOI210     o699(.A0(ori_ori_n721_), .A1(ori_ori_n390_), .B0(ori_ori_n559_), .Y(ori_ori_n722_));
  NO2        o700(.A(ori_ori_n722_), .B(ori_ori_n720_), .Y(ori_ori_n723_));
  NO3        o701(.A(ori_ori_n723_), .B(ori_ori_n718_), .C(ori_ori_n714_), .Y(ori_ori_n724_));
  NA2        o702(.A(ori_ori_n169_), .B(ori_ori_n24_), .Y(ori_ori_n725_));
  NO2        o703(.A(ori_ori_n546_), .B(ori_ori_n471_), .Y(ori_ori_n726_));
  NO2        o704(.A(ori_ori_n726_), .B(ori_ori_n725_), .Y(ori_ori_n727_));
  NA2        o705(.A(ori_ori_n262_), .B(ori_ori_n131_), .Y(ori_ori_n728_));
  NAi21      o706(.An(ori_ori_n160_), .B(ori_ori_n352_), .Y(ori_ori_n729_));
  OAI220     o707(.A0(ori_ori_n729_), .A1(ori_ori_n700_), .B0(ori_ori_n728_), .B1(ori_ori_n334_), .Y(ori_ori_n730_));
  NO2        o708(.A(ori_ori_n730_), .B(ori_ori_n727_), .Y(ori_ori_n731_));
  NA2        o709(.A(ori_ori_n449_), .B(i_0_), .Y(ori_ori_n732_));
  NO3        o710(.A(ori_ori_n732_), .B(ori_ori_n317_), .C(ori_ori_n87_), .Y(ori_ori_n733_));
  NO4        o711(.A(ori_ori_n462_), .B(ori_ori_n191_), .C(ori_ori_n344_), .D(i_6_), .Y(ori_ori_n734_));
  AOI210     o712(.A0(ori_ori_n734_), .A1(i_11_), .B0(ori_ori_n733_), .Y(ori_ori_n735_));
  INV        o713(.A(ori_ori_n389_), .Y(ori_ori_n736_));
  NA2        o714(.A(ori_ori_n616_), .B(ori_ori_n269_), .Y(ori_ori_n737_));
  AOI210     o715(.A0(ori_ori_n393_), .A1(ori_ori_n87_), .B0(ori_ori_n56_), .Y(ori_ori_n738_));
  NO2        o716(.A(ori_ori_n738_), .B(ori_ori_n737_), .Y(ori_ori_n739_));
  NO2        o717(.A(ori_ori_n220_), .B(ori_ori_n154_), .Y(ori_ori_n740_));
  NA2        o718(.A(i_0_), .B(i_10_), .Y(ori_ori_n741_));
  AN2        o719(.A(ori_ori_n740_), .B(i_6_), .Y(ori_ori_n742_));
  NO2        o720(.A(ori_ori_n742_), .B(ori_ori_n739_), .Y(ori_ori_n743_));
  NA3        o721(.A(ori_ori_n743_), .B(ori_ori_n735_), .C(ori_ori_n731_), .Y(ori_ori_n744_));
  NO2        o722(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n745_));
  NA2        o723(.A(i_11_), .B(i_9_), .Y(ori_ori_n746_));
  NO3        o724(.A(i_12_), .B(ori_ori_n746_), .C(ori_ori_n479_), .Y(ori_ori_n747_));
  AN2        o725(.A(ori_ori_n747_), .B(ori_ori_n745_), .Y(ori_ori_n748_));
  NO2        o726(.A(ori_ori_n48_), .B(i_7_), .Y(ori_ori_n749_));
  NA2        o727(.A(ori_ori_n326_), .B(ori_ori_n166_), .Y(ori_ori_n750_));
  NA2        o728(.A(ori_ori_n750_), .B(ori_ori_n158_), .Y(ori_ori_n751_));
  NO2        o729(.A(ori_ori_n746_), .B(ori_ori_n71_), .Y(ori_ori_n752_));
  NO2        o730(.A(ori_ori_n165_), .B(i_0_), .Y(ori_ori_n753_));
  INV        o731(.A(ori_ori_n340_), .Y(ori_ori_n754_));
  NO2        o732(.A(ori_ori_n754_), .B(ori_ori_n720_), .Y(ori_ori_n755_));
  NO3        o733(.A(ori_ori_n755_), .B(ori_ori_n751_), .C(ori_ori_n748_), .Y(ori_ori_n756_));
  NA2        o734(.A(ori_ori_n533_), .B(ori_ori_n123_), .Y(ori_ori_n757_));
  NO2        o735(.A(i_6_), .B(ori_ori_n757_), .Y(ori_ori_n758_));
  NA2        o736(.A(ori_ori_n162_), .B(ori_ori_n104_), .Y(ori_ori_n759_));
  NA2        o737(.A(ori_ori_n481_), .B(ori_ori_n269_), .Y(ori_ori_n760_));
  NO2        o738(.A(ori_ori_n760_), .B(ori_ori_n712_), .Y(ori_ori_n761_));
  NO2        o739(.A(ori_ori_n761_), .B(ori_ori_n758_), .Y(ori_ori_n762_));
  NOi21      o740(.An(i_7_), .B(i_5_), .Y(ori_ori_n763_));
  NOi31      o741(.An(ori_ori_n763_), .B(i_0_), .C(ori_ori_n598_), .Y(ori_ori_n764_));
  NA3        o742(.A(ori_ori_n764_), .B(ori_ori_n316_), .C(i_6_), .Y(ori_ori_n765_));
  BUFFER     o743(.A(ori_ori_n765_), .Y(ori_ori_n766_));
  INV        o744(.A(ori_ori_n265_), .Y(ori_ori_n767_));
  NA3        o745(.A(ori_ori_n766_), .B(ori_ori_n762_), .C(ori_ori_n756_), .Y(ori_ori_n768_));
  NO2        o746(.A(ori_ori_n706_), .B(ori_ori_n264_), .Y(ori_ori_n769_));
  OA210      o747(.A0(ori_ori_n389_), .A1(ori_ori_n199_), .B0(ori_ori_n388_), .Y(ori_ori_n770_));
  NA2        o748(.A(ori_ori_n769_), .B(ori_ori_n752_), .Y(ori_ori_n771_));
  NA3        o749(.A(ori_ori_n388_), .B(ori_ori_n342_), .C(ori_ori_n45_), .Y(ori_ori_n772_));
  OAI210     o750(.A0(ori_ori_n729_), .A1(ori_ori_n736_), .B0(ori_ori_n772_), .Y(ori_ori_n773_));
  NA2        o751(.A(ori_ori_n752_), .B(ori_ori_n257_), .Y(ori_ori_n774_));
  OAI210     o752(.A0(i_3_), .A1(ori_ori_n171_), .B0(ori_ori_n774_), .Y(ori_ori_n775_));
  AOI220     o753(.A0(ori_ori_n775_), .A1(ori_ori_n389_), .B0(ori_ori_n773_), .B1(ori_ori_n71_), .Y(ori_ori_n776_));
  NA3        o754(.A(i_5_), .B(ori_ori_n314_), .C(ori_ori_n515_), .Y(ori_ori_n777_));
  NA2        o755(.A(ori_ori_n93_), .B(ori_ori_n44_), .Y(ori_ori_n778_));
  NO2        o756(.A(ori_ori_n73_), .B(ori_ori_n618_), .Y(ori_ori_n779_));
  AOI220     o757(.A0(ori_ori_n779_), .A1(ori_ori_n778_), .B0(ori_ori_n164_), .B1(ori_ori_n471_), .Y(ori_ori_n780_));
  AOI210     o758(.A0(ori_ori_n780_), .A1(ori_ori_n777_), .B0(ori_ori_n47_), .Y(ori_ori_n781_));
  NO3        o759(.A(ori_ori_n462_), .B(ori_ori_n289_), .C(ori_ori_n24_), .Y(ori_ori_n782_));
  AOI210     o760(.A0(ori_ori_n575_), .A1(ori_ori_n430_), .B0(ori_ori_n782_), .Y(ori_ori_n783_));
  NAi21      o761(.An(i_9_), .B(i_5_), .Y(ori_ori_n784_));
  NO2        o762(.A(ori_ori_n784_), .B(ori_ori_n335_), .Y(ori_ori_n785_));
  NA2        o763(.A(ori_ori_n785_), .B(ori_ori_n495_), .Y(ori_ori_n786_));
  OAI220     o764(.A0(ori_ori_n786_), .A1(ori_ori_n84_), .B0(ori_ori_n783_), .B1(ori_ori_n163_), .Y(ori_ori_n787_));
  NO2        o765(.A(ori_ori_n787_), .B(ori_ori_n781_), .Y(ori_ori_n788_));
  NA3        o766(.A(ori_ori_n788_), .B(ori_ori_n776_), .C(ori_ori_n771_), .Y(ori_ori_n789_));
  NO3        o767(.A(ori_ori_n789_), .B(ori_ori_n768_), .C(ori_ori_n744_), .Y(ori_ori_n790_));
  NO2        o768(.A(i_0_), .B(ori_ori_n598_), .Y(ori_ori_n791_));
  NO2        o769(.A(ori_ori_n664_), .B(ori_ori_n759_), .Y(ori_ori_n792_));
  INV        o770(.A(ori_ori_n792_), .Y(ori_ori_n793_));
  NO2        o771(.A(ori_ori_n682_), .B(ori_ori_n335_), .Y(ori_ori_n794_));
  NA2        o772(.A(ori_ori_n214_), .B(ori_ori_n206_), .Y(ori_ori_n795_));
  AOI210     o773(.A0(ori_ori_n795_), .A1(ori_ori_n732_), .B0(ori_ori_n154_), .Y(ori_ori_n796_));
  NO2        o774(.A(ori_ori_n796_), .B(ori_ori_n794_), .Y(ori_ori_n797_));
  NA2        o775(.A(ori_ori_n797_), .B(ori_ori_n793_), .Y(ori_ori_n798_));
  NO3        o776(.A(ori_ori_n741_), .B(ori_ori_n719_), .C(ori_ori_n174_), .Y(ori_ori_n799_));
  AOI220     o777(.A0(ori_ori_n799_), .A1(i_11_), .B0(ori_ori_n447_), .B1(ori_ori_n73_), .Y(ori_ori_n800_));
  NO3        o778(.A(ori_ori_n187_), .B(ori_ori_n315_), .C(i_0_), .Y(ori_ori_n801_));
  OAI210     o779(.A0(ori_ori_n801_), .A1(ori_ori_n74_), .B0(i_13_), .Y(ori_ori_n802_));
  NA2        o780(.A(ori_ori_n802_), .B(ori_ori_n800_), .Y(ori_ori_n803_));
  NO2        o781(.A(ori_ori_n213_), .B(ori_ori_n93_), .Y(ori_ori_n804_));
  AOI210     o782(.A0(ori_ori_n804_), .A1(ori_ori_n791_), .B0(ori_ori_n110_), .Y(ori_ori_n805_));
  OR2        o783(.A(ori_ori_n805_), .B(i_5_), .Y(ori_ori_n806_));
  AOI210     o784(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n165_), .Y(ori_ori_n807_));
  NA2        o785(.A(ori_ori_n807_), .B(ori_ori_n770_), .Y(ori_ori_n808_));
  INV        o786(.A(ori_ori_n428_), .Y(ori_ori_n809_));
  NO3        o787(.A(ori_ori_n712_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n810_));
  NA2        o788(.A(ori_ori_n401_), .B(ori_ori_n394_), .Y(ori_ori_n811_));
  NO3        o789(.A(ori_ori_n811_), .B(ori_ori_n810_), .C(ori_ori_n809_), .Y(ori_ori_n812_));
  NA3        o790(.A(ori_ori_n321_), .B(ori_ori_n162_), .C(ori_ori_n161_), .Y(ori_ori_n813_));
  NA3        o791(.A(ori_ori_n749_), .B(ori_ori_n249_), .C(ori_ori_n206_), .Y(ori_ori_n814_));
  NA2        o792(.A(ori_ori_n814_), .B(ori_ori_n813_), .Y(ori_ori_n815_));
  NA3        o793(.A(ori_ori_n321_), .B(ori_ori_n276_), .C(ori_ori_n197_), .Y(ori_ori_n816_));
  INV        o794(.A(ori_ori_n816_), .Y(ori_ori_n817_));
  NO3        o795(.A(ori_ori_n746_), .B(ori_ori_n194_), .C(ori_ori_n174_), .Y(ori_ori_n818_));
  NO3        o796(.A(ori_ori_n818_), .B(ori_ori_n817_), .C(ori_ori_n815_), .Y(ori_ori_n819_));
  NA4        o797(.A(ori_ori_n819_), .B(ori_ori_n812_), .C(ori_ori_n808_), .D(ori_ori_n806_), .Y(ori_ori_n820_));
  NO2        o798(.A(ori_ori_n84_), .B(i_5_), .Y(ori_ori_n821_));
  NA3        o799(.A(ori_ori_n707_), .B(ori_ori_n111_), .C(ori_ori_n126_), .Y(ori_ori_n822_));
  INV        o800(.A(ori_ori_n822_), .Y(ori_ori_n823_));
  NA2        o801(.A(ori_ori_n823_), .B(ori_ori_n821_), .Y(ori_ori_n824_));
  NA3        o802(.A(ori_ori_n257_), .B(i_5_), .C(ori_ori_n175_), .Y(ori_ori_n825_));
  NAi31      o803(.An(ori_ori_n212_), .B(ori_ori_n825_), .C(ori_ori_n213_), .Y(ori_ori_n826_));
  NO4        o804(.A(ori_ori_n211_), .B(ori_ori_n187_), .C(i_0_), .D(i_12_), .Y(ori_ori_n827_));
  NA2        o805(.A(ori_ori_n827_), .B(ori_ori_n826_), .Y(ori_ori_n828_));
  AN2        o806(.A(ori_ori_n741_), .B(ori_ori_n154_), .Y(ori_ori_n829_));
  NO4        o807(.A(ori_ori_n829_), .B(i_12_), .C(ori_ori_n521_), .D(ori_ori_n133_), .Y(ori_ori_n830_));
  NA2        o808(.A(ori_ori_n830_), .B(ori_ori_n194_), .Y(ori_ori_n831_));
  NA2        o809(.A(ori_ori_n763_), .B(ori_ori_n386_), .Y(ori_ori_n832_));
  NA2        o810(.A(ori_ori_n62_), .B(ori_ori_n102_), .Y(ori_ori_n833_));
  OAI220     o811(.A0(ori_ori_n833_), .A1(ori_ori_n825_), .B0(ori_ori_n832_), .B1(ori_ori_n549_), .Y(ori_ori_n834_));
  NA2        o812(.A(ori_ori_n834_), .B(ori_ori_n753_), .Y(ori_ori_n835_));
  NA4        o813(.A(ori_ori_n835_), .B(ori_ori_n831_), .C(ori_ori_n828_), .D(ori_ori_n824_), .Y(ori_ori_n836_));
  NO4        o814(.A(ori_ori_n836_), .B(ori_ori_n820_), .C(ori_ori_n803_), .D(ori_ori_n798_), .Y(ori_ori_n837_));
  OAI210     o815(.A0(ori_ori_n685_), .A1(ori_ori_n678_), .B0(ori_ori_n37_), .Y(ori_ori_n838_));
  NA2        o816(.A(ori_ori_n838_), .B(ori_ori_n487_), .Y(ori_ori_n839_));
  NA2        o817(.A(ori_ori_n839_), .B(ori_ori_n185_), .Y(ori_ori_n840_));
  NAi31      o818(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n841_));
  AOI210     o819(.A0(ori_ori_n119_), .A1(ori_ori_n68_), .B0(ori_ori_n841_), .Y(ori_ori_n842_));
  NO2        o820(.A(ori_ori_n842_), .B(ori_ori_n518_), .Y(ori_ori_n843_));
  INV        o821(.A(ori_ori_n843_), .Y(ori_ori_n844_));
  AOI210     o822(.A0(ori_ori_n844_), .A1(ori_ori_n48_), .B0(ori_ori_n734_), .Y(ori_ori_n845_));
  AOI210     o823(.A0(ori_ori_n845_), .A1(ori_ori_n840_), .B0(ori_ori_n71_), .Y(ori_ori_n846_));
  INV        o824(.A(ori_ori_n311_), .Y(ori_ori_n847_));
  NO2        o825(.A(ori_ori_n847_), .B(ori_ori_n624_), .Y(ori_ori_n848_));
  OAI210     o826(.A0(ori_ori_n78_), .A1(ori_ori_n54_), .B0(ori_ori_n109_), .Y(ori_ori_n849_));
  NA2        o827(.A(ori_ori_n849_), .B(ori_ori_n74_), .Y(ori_ori_n850_));
  AOI210     o828(.A0(ori_ori_n807_), .A1(ori_ori_n749_), .B0(ori_ori_n764_), .Y(ori_ori_n851_));
  AOI210     o829(.A0(ori_ori_n851_), .A1(ori_ori_n850_), .B0(ori_ori_n552_), .Y(ori_ori_n852_));
  INV        o830(.A(ori_ori_n852_), .Y(ori_ori_n853_));
  OAI210     o831(.A0(ori_ori_n235_), .A1(ori_ori_n156_), .B0(ori_ori_n87_), .Y(ori_ori_n854_));
  NA3        o832(.A(ori_ori_n628_), .B(ori_ori_n249_), .C(ori_ori_n78_), .Y(ori_ori_n855_));
  AOI210     o833(.A0(ori_ori_n855_), .A1(ori_ori_n854_), .B0(i_11_), .Y(ori_ori_n856_));
  NO3        o834(.A(ori_ori_n57_), .B(ori_ori_n56_), .C(i_4_), .Y(ori_ori_n857_));
  OAI210     o835(.A0(ori_ori_n767_), .A1(ori_ori_n258_), .B0(ori_ori_n857_), .Y(ori_ori_n858_));
  NO2        o836(.A(ori_ori_n858_), .B(ori_ori_n598_), .Y(ori_ori_n859_));
  NO4        o837(.A(ori_ori_n784_), .B(ori_ori_n391_), .C(ori_ori_n219_), .D(ori_ori_n218_), .Y(ori_ori_n860_));
  NO2        o838(.A(ori_ori_n860_), .B(ori_ori_n443_), .Y(ori_ori_n861_));
  INV        o839(.A(ori_ori_n292_), .Y(ori_ori_n862_));
  AOI210     o840(.A0(ori_ori_n862_), .A1(ori_ori_n861_), .B0(ori_ori_n41_), .Y(ori_ori_n863_));
  NO3        o841(.A(ori_ori_n863_), .B(ori_ori_n859_), .C(ori_ori_n856_), .Y(ori_ori_n864_));
  OAI210     o842(.A0(ori_ori_n853_), .A1(i_4_), .B0(ori_ori_n864_), .Y(ori_ori_n865_));
  NO3        o843(.A(ori_ori_n865_), .B(ori_ori_n848_), .C(ori_ori_n846_), .Y(ori_ori_n866_));
  NA4        o844(.A(ori_ori_n866_), .B(ori_ori_n837_), .C(ori_ori_n790_), .D(ori_ori_n724_), .Y(ori4));
  INV        o845(.A(ori_ori_n574_), .Y(ori_ori_n870_));
  INV        o846(.A(ori_ori_n273_), .Y(ori_ori_n871_));
  INV        o847(.A(ori_ori_n586_), .Y(ori_ori_n872_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m0033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m0034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m0036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m0037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m0038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m0039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m0040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m0041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m0042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m0043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m0044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m0045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m0046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m0047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m0049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m0050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m0051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m0052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m0053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m0054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m0055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m0057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m0059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m0060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m0062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m0063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m0064(.A(i_6_), .Y(mai_mai_n87_));
  OR4        m0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n88_));
  INV        m0066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m0067(.A(i_2_), .B(i_7_), .Y(mai_mai_n90_));
  NO2        m0068(.A(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  OAI210     m0069(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NAi21      m0070(.An(i_6_), .B(i_10_), .Y(mai_mai_n93_));
  NA2        m0071(.A(i_6_), .B(i_9_), .Y(mai_mai_n94_));
  AOI210     m0072(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n64_), .Y(mai_mai_n95_));
  NA2        m0073(.A(i_2_), .B(i_6_), .Y(mai_mai_n96_));
  INV        m0074(.A(mai_mai_n95_), .Y(mai_mai_n97_));
  AOI210     m0075(.A0(mai_mai_n97_), .A1(mai_mai_n92_), .B0(mai_mai_n81_), .Y(mai_mai_n98_));
  AN3        m0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n99_));
  NAi21      m0077(.An(i_6_), .B(i_11_), .Y(mai_mai_n100_));
  NO2        m0078(.A(i_5_), .B(i_8_), .Y(mai_mai_n101_));
  NOi21      m0079(.An(mai_mai_n101_), .B(mai_mai_n100_), .Y(mai_mai_n102_));
  AOI220     m0080(.A0(mai_mai_n102_), .A1(mai_mai_n63_), .B0(mai_mai_n99_), .B1(mai_mai_n32_), .Y(mai_mai_n103_));
  INV        m0081(.A(i_7_), .Y(mai_mai_n104_));
  NA2        m0082(.A(mai_mai_n47_), .B(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m0083(.A(i_0_), .B(i_5_), .Y(mai_mai_n106_));
  NO2        m0084(.A(mai_mai_n106_), .B(mai_mai_n87_), .Y(mai_mai_n107_));
  NA2        m0085(.A(i_12_), .B(i_3_), .Y(mai_mai_n108_));
  INV        m0086(.A(mai_mai_n108_), .Y(mai_mai_n109_));
  NA3        m0087(.A(mai_mai_n109_), .B(mai_mai_n107_), .C(mai_mai_n105_), .Y(mai_mai_n110_));
  NAi21      m0088(.An(i_7_), .B(i_11_), .Y(mai_mai_n111_));
  NO3        m0089(.A(mai_mai_n111_), .B(mai_mai_n93_), .C(mai_mai_n54_), .Y(mai_mai_n112_));
  AN2        m0090(.A(i_2_), .B(i_10_), .Y(mai_mai_n113_));
  NO2        m0091(.A(mai_mai_n113_), .B(i_7_), .Y(mai_mai_n114_));
  OR2        m0092(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n115_));
  NO2        m0093(.A(i_8_), .B(mai_mai_n104_), .Y(mai_mai_n116_));
  NO3        m0094(.A(mai_mai_n116_), .B(mai_mai_n115_), .C(mai_mai_n114_), .Y(mai_mai_n117_));
  NA2        m0095(.A(i_12_), .B(i_7_), .Y(mai_mai_n118_));
  NO2        m0096(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n119_));
  NA2        m0097(.A(i_11_), .B(i_12_), .Y(mai_mai_n120_));
  INV        m0098(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NO2        m0099(.A(mai_mai_n121_), .B(mai_mai_n117_), .Y(mai_mai_n122_));
  NAi41      m0100(.An(mai_mai_n112_), .B(mai_mai_n122_), .C(mai_mai_n110_), .D(mai_mai_n103_), .Y(mai_mai_n123_));
  NOi21      m0101(.An(i_1_), .B(i_5_), .Y(mai_mai_n124_));
  NA2        m0102(.A(mai_mai_n124_), .B(i_11_), .Y(mai_mai_n125_));
  NA2        m0103(.A(mai_mai_n104_), .B(mai_mai_n37_), .Y(mai_mai_n126_));
  NA2        m0104(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n127_));
  NA2        m0105(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NO2        m0106(.A(mai_mai_n128_), .B(mai_mai_n47_), .Y(mai_mai_n129_));
  NA2        m0107(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n130_));
  NAi21      m0108(.An(i_3_), .B(i_8_), .Y(mai_mai_n131_));
  NA2        m0109(.A(mai_mai_n131_), .B(mai_mai_n63_), .Y(mai_mai_n132_));
  NOi31      m0110(.An(mai_mai_n132_), .B(mai_mai_n130_), .C(mai_mai_n129_), .Y(mai_mai_n133_));
  NO2        m0111(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n134_));
  NO2        m0112(.A(i_6_), .B(i_5_), .Y(mai_mai_n135_));
  NA2        m0113(.A(mai_mai_n135_), .B(i_3_), .Y(mai_mai_n136_));
  AO210      m0114(.A0(mai_mai_n136_), .A1(mai_mai_n48_), .B0(mai_mai_n134_), .Y(mai_mai_n137_));
  OAI220     m0115(.A0(mai_mai_n137_), .A1(mai_mai_n111_), .B0(mai_mai_n133_), .B1(mai_mai_n125_), .Y(mai_mai_n138_));
  NO3        m0116(.A(mai_mai_n138_), .B(mai_mai_n123_), .C(mai_mai_n98_), .Y(mai_mai_n139_));
  NA3        m0117(.A(mai_mai_n139_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m0118(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n141_));
  NA2        m0119(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n142_));
  NA2        m0120(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  NA4        m0121(.A(mai_mai_n143_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0122(.A(i_8_), .B(i_7_), .Y(mai_mai_n145_));
  NA2        m0123(.A(mai_mai_n145_), .B(i_6_), .Y(mai_mai_n146_));
  NO2        m0124(.A(i_12_), .B(i_13_), .Y(mai_mai_n147_));
  NAi21      m0125(.An(i_5_), .B(i_11_), .Y(mai_mai_n148_));
  NOi21      m0126(.An(mai_mai_n147_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  NO2        m0127(.A(i_0_), .B(i_1_), .Y(mai_mai_n150_));
  NA2        m0128(.A(i_2_), .B(i_3_), .Y(mai_mai_n151_));
  NO2        m0129(.A(mai_mai_n151_), .B(i_4_), .Y(mai_mai_n152_));
  NA3        m0130(.A(mai_mai_n152_), .B(mai_mai_n150_), .C(mai_mai_n149_), .Y(mai_mai_n153_));
  AN2        m0131(.A(mai_mai_n147_), .B(mai_mai_n84_), .Y(mai_mai_n154_));
  NO2        m0132(.A(mai_mai_n154_), .B(mai_mai_n27_), .Y(mai_mai_n155_));
  NA2        m0133(.A(i_1_), .B(i_5_), .Y(mai_mai_n156_));
  NO2        m0134(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n157_));
  NA2        m0135(.A(mai_mai_n157_), .B(mai_mai_n36_), .Y(mai_mai_n158_));
  NO3        m0136(.A(mai_mai_n158_), .B(mai_mai_n156_), .C(mai_mai_n155_), .Y(mai_mai_n159_));
  OR2        m0137(.A(i_0_), .B(i_1_), .Y(mai_mai_n160_));
  NO3        m0138(.A(mai_mai_n160_), .B(mai_mai_n81_), .C(i_13_), .Y(mai_mai_n161_));
  NAi32      m0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n162_));
  NAi21      m0140(.An(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  NOi21      m0141(.An(i_4_), .B(i_10_), .Y(mai_mai_n164_));
  NA2        m0142(.A(mai_mai_n164_), .B(mai_mai_n40_), .Y(mai_mai_n165_));
  NO2        m0143(.A(i_3_), .B(i_5_), .Y(mai_mai_n166_));
  NO3        m0144(.A(mai_mai_n74_), .B(i_2_), .C(i_1_), .Y(mai_mai_n167_));
  NA2        m0145(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  OAI210     m0146(.A0(mai_mai_n168_), .A1(mai_mai_n165_), .B0(mai_mai_n163_), .Y(mai_mai_n169_));
  NO2        m0147(.A(mai_mai_n169_), .B(mai_mai_n159_), .Y(mai_mai_n170_));
  AOI210     m0148(.A0(mai_mai_n170_), .A1(mai_mai_n153_), .B0(mai_mai_n146_), .Y(mai_mai_n171_));
  NA3        m0149(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n172_));
  NA2        m0150(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n173_));
  NOi21      m0151(.An(i_4_), .B(i_9_), .Y(mai_mai_n174_));
  NOi21      m0152(.An(i_11_), .B(i_13_), .Y(mai_mai_n175_));
  NA2        m0153(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  OR2        m0154(.A(mai_mai_n176_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  NO2        m0155(.A(i_4_), .B(i_5_), .Y(mai_mai_n178_));
  NAi21      m0156(.An(i_12_), .B(i_11_), .Y(mai_mai_n179_));
  NO2        m0157(.A(mai_mai_n179_), .B(i_13_), .Y(mai_mai_n180_));
  NA3        m0158(.A(mai_mai_n180_), .B(mai_mai_n178_), .C(mai_mai_n84_), .Y(mai_mai_n181_));
  AOI210     m0159(.A0(mai_mai_n181_), .A1(mai_mai_n177_), .B0(mai_mai_n172_), .Y(mai_mai_n182_));
  NO2        m0160(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n183_));
  INV        m0161(.A(mai_mai_n183_), .Y(mai_mai_n184_));
  NA2        m0162(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n185_));
  NAi31      m0163(.An(mai_mai_n185_), .B(mai_mai_n154_), .C(i_11_), .Y(mai_mai_n186_));
  NA2        m0164(.A(i_3_), .B(i_5_), .Y(mai_mai_n187_));
  OR2        m0165(.A(mai_mai_n187_), .B(mai_mai_n176_), .Y(mai_mai_n188_));
  AOI210     m0166(.A0(mai_mai_n188_), .A1(mai_mai_n186_), .B0(mai_mai_n184_), .Y(mai_mai_n189_));
  NO2        m0167(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n190_));
  NO2        m0168(.A(i_13_), .B(i_10_), .Y(mai_mai_n191_));
  NA3        m0169(.A(mai_mai_n191_), .B(mai_mai_n190_), .C(mai_mai_n45_), .Y(mai_mai_n192_));
  NO2        m0170(.A(i_2_), .B(i_1_), .Y(mai_mai_n193_));
  NA2        m0171(.A(mai_mai_n193_), .B(i_3_), .Y(mai_mai_n194_));
  NAi21      m0172(.An(i_4_), .B(i_12_), .Y(mai_mai_n195_));
  NO3        m0173(.A(mai_mai_n194_), .B(mai_mai_n192_), .C(mai_mai_n25_), .Y(mai_mai_n196_));
  NO3        m0174(.A(mai_mai_n196_), .B(mai_mai_n189_), .C(mai_mai_n182_), .Y(mai_mai_n197_));
  INV        m0175(.A(i_8_), .Y(mai_mai_n198_));
  NO2        m0176(.A(mai_mai_n198_), .B(i_7_), .Y(mai_mai_n199_));
  NA2        m0177(.A(mai_mai_n199_), .B(i_6_), .Y(mai_mai_n200_));
  NO3        m0178(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n201_));
  NA2        m0179(.A(mai_mai_n201_), .B(mai_mai_n116_), .Y(mai_mai_n202_));
  NO3        m0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n203_));
  NA3        m0181(.A(mai_mai_n203_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n204_));
  NO3        m0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n205_));
  OAI210     m0183(.A0(mai_mai_n99_), .A1(i_12_), .B0(mai_mai_n205_), .Y(mai_mai_n206_));
  AOI210     m0184(.A0(mai_mai_n206_), .A1(mai_mai_n204_), .B0(mai_mai_n202_), .Y(mai_mai_n207_));
  NO2        m0185(.A(i_3_), .B(i_8_), .Y(mai_mai_n208_));
  NO3        m0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n209_));
  NO2        m0187(.A(mai_mai_n106_), .B(mai_mai_n59_), .Y(mai_mai_n210_));
  NO2        m0188(.A(i_13_), .B(i_9_), .Y(mai_mai_n211_));
  NA3        m0189(.A(mai_mai_n211_), .B(i_6_), .C(mai_mai_n198_), .Y(mai_mai_n212_));
  NAi21      m0190(.An(i_12_), .B(i_3_), .Y(mai_mai_n213_));
  OR2        m0191(.A(mai_mai_n213_), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  NO2        m0192(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n215_));
  NO3        m0193(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n216_));
  NA2        m0194(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  NO2        m0195(.A(mai_mai_n217_), .B(mai_mai_n214_), .Y(mai_mai_n218_));
  NO2        m0196(.A(mai_mai_n218_), .B(mai_mai_n207_), .Y(mai_mai_n219_));
  OAI220     m0197(.A0(mai_mai_n219_), .A1(i_4_), .B0(mai_mai_n200_), .B1(mai_mai_n197_), .Y(mai_mai_n220_));
  NAi21      m0198(.An(i_12_), .B(i_7_), .Y(mai_mai_n221_));
  NA3        m0199(.A(i_13_), .B(mai_mai_n198_), .C(i_10_), .Y(mai_mai_n222_));
  NA2        m0200(.A(i_0_), .B(i_5_), .Y(mai_mai_n223_));
  NAi31      m0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n224_));
  NO2        m0202(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n225_));
  INV        m0203(.A(i_13_), .Y(mai_mai_n226_));
  NO2        m0204(.A(i_12_), .B(mai_mai_n226_), .Y(mai_mai_n227_));
  NO2        m0205(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n228_));
  NO2        m0206(.A(mai_mai_n187_), .B(i_4_), .Y(mai_mai_n229_));
  NA2        m0207(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  OR2        m0208(.A(i_8_), .B(i_7_), .Y(mai_mai_n231_));
  NO2        m0209(.A(mai_mai_n231_), .B(mai_mai_n87_), .Y(mai_mai_n232_));
  NO2        m0210(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n233_));
  NA2        m0211(.A(mai_mai_n233_), .B(mai_mai_n232_), .Y(mai_mai_n234_));
  INV        m0212(.A(i_12_), .Y(mai_mai_n235_));
  NO2        m0213(.A(mai_mai_n45_), .B(mai_mai_n235_), .Y(mai_mai_n236_));
  NO3        m0214(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n237_));
  NA2        m0215(.A(i_2_), .B(i_1_), .Y(mai_mai_n238_));
  NO2        m0216(.A(mai_mai_n234_), .B(mai_mai_n230_), .Y(mai_mai_n239_));
  NO3        m0217(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n240_));
  NAi21      m0218(.An(i_4_), .B(i_3_), .Y(mai_mai_n241_));
  NO2        m0219(.A(mai_mai_n241_), .B(mai_mai_n76_), .Y(mai_mai_n242_));
  NO2        m0220(.A(i_0_), .B(i_6_), .Y(mai_mai_n243_));
  NOi41      m0221(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n244_));
  NA2        m0222(.A(mai_mai_n244_), .B(mai_mai_n243_), .Y(mai_mai_n245_));
  NO2        m0223(.A(mai_mai_n238_), .B(mai_mai_n187_), .Y(mai_mai_n246_));
  NAi21      m0224(.An(mai_mai_n245_), .B(mai_mai_n246_), .Y(mai_mai_n247_));
  INV        m0225(.A(mai_mai_n247_), .Y(mai_mai_n248_));
  AOI210     m0226(.A0(mai_mai_n248_), .A1(mai_mai_n40_), .B0(mai_mai_n239_), .Y(mai_mai_n249_));
  NO2        m0227(.A(i_11_), .B(mai_mai_n226_), .Y(mai_mai_n250_));
  NOi21      m0228(.An(i_1_), .B(i_6_), .Y(mai_mai_n251_));
  NAi21      m0229(.An(i_3_), .B(i_7_), .Y(mai_mai_n252_));
  NA2        m0230(.A(mai_mai_n235_), .B(i_9_), .Y(mai_mai_n253_));
  OR4        m0231(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n251_), .D(mai_mai_n190_), .Y(mai_mai_n254_));
  NO2        m0232(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n255_));
  NO2        m0233(.A(i_12_), .B(i_3_), .Y(mai_mai_n256_));
  NA2        m0234(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n257_));
  NA2        m0235(.A(i_3_), .B(i_9_), .Y(mai_mai_n258_));
  NAi21      m0236(.An(i_7_), .B(i_10_), .Y(mai_mai_n259_));
  NO2        m0237(.A(mai_mai_n259_), .B(mai_mai_n258_), .Y(mai_mai_n260_));
  NA3        m0238(.A(mai_mai_n260_), .B(mai_mai_n257_), .C(mai_mai_n65_), .Y(mai_mai_n261_));
  NA2        m0239(.A(mai_mai_n261_), .B(mai_mai_n254_), .Y(mai_mai_n262_));
  NA3        m0240(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n263_));
  INV        m0241(.A(mai_mai_n146_), .Y(mai_mai_n264_));
  NA2        m0242(.A(mai_mai_n235_), .B(i_13_), .Y(mai_mai_n265_));
  NO2        m0243(.A(mai_mai_n265_), .B(mai_mai_n76_), .Y(mai_mai_n266_));
  AOI220     m0244(.A0(mai_mai_n266_), .A1(mai_mai_n264_), .B0(mai_mai_n262_), .B1(mai_mai_n250_), .Y(mai_mai_n267_));
  NO2        m0245(.A(mai_mai_n231_), .B(mai_mai_n37_), .Y(mai_mai_n268_));
  NA2        m0246(.A(i_12_), .B(i_6_), .Y(mai_mai_n269_));
  OR2        m0247(.A(i_13_), .B(i_9_), .Y(mai_mai_n270_));
  NO2        m0248(.A(mai_mai_n241_), .B(i_2_), .Y(mai_mai_n271_));
  NA2        m0249(.A(mai_mai_n250_), .B(i_9_), .Y(mai_mai_n272_));
  NA2        m0250(.A(mai_mai_n157_), .B(mai_mai_n64_), .Y(mai_mai_n273_));
  NO3        m0251(.A(i_11_), .B(mai_mai_n226_), .C(mai_mai_n25_), .Y(mai_mai_n274_));
  NO2        m0252(.A(mai_mai_n252_), .B(i_8_), .Y(mai_mai_n275_));
  NO2        m0253(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n276_));
  NA3        m0254(.A(mai_mai_n276_), .B(mai_mai_n275_), .C(mai_mai_n274_), .Y(mai_mai_n277_));
  NO3        m0255(.A(mai_mai_n26_), .B(mai_mai_n87_), .C(i_5_), .Y(mai_mai_n278_));
  NA3        m0256(.A(mai_mai_n278_), .B(mai_mai_n268_), .C(mai_mai_n227_), .Y(mai_mai_n279_));
  AOI210     m0257(.A0(mai_mai_n279_), .A1(mai_mai_n277_), .B0(mai_mai_n273_), .Y(mai_mai_n280_));
  INV        m0258(.A(mai_mai_n280_), .Y(mai_mai_n281_));
  NA3        m0259(.A(mai_mai_n281_), .B(mai_mai_n267_), .C(mai_mai_n249_), .Y(mai_mai_n282_));
  NO3        m0260(.A(i_12_), .B(mai_mai_n226_), .C(mai_mai_n37_), .Y(mai_mai_n283_));
  INV        m0261(.A(mai_mai_n283_), .Y(mai_mai_n284_));
  NA2        m0262(.A(i_8_), .B(mai_mai_n104_), .Y(mai_mai_n285_));
  NOi21      m0263(.An(mai_mai_n166_), .B(mai_mai_n87_), .Y(mai_mai_n286_));
  NO3        m0264(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n287_));
  AOI220     m0265(.A0(mai_mai_n287_), .A1(mai_mai_n201_), .B0(mai_mai_n286_), .B1(mai_mai_n233_), .Y(mai_mai_n288_));
  NO2        m0266(.A(mai_mai_n288_), .B(mai_mai_n285_), .Y(mai_mai_n289_));
  NO2        m0267(.A(mai_mai_n238_), .B(i_0_), .Y(mai_mai_n290_));
  NA2        m0268(.A(i_0_), .B(i_1_), .Y(mai_mai_n291_));
  NO2        m0269(.A(mai_mai_n291_), .B(i_2_), .Y(mai_mai_n292_));
  NO2        m0270(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n293_));
  NA3        m0271(.A(mai_mai_n293_), .B(mai_mai_n292_), .C(mai_mai_n166_), .Y(mai_mai_n294_));
  OAI210     m0272(.A0(mai_mai_n168_), .A1(mai_mai_n146_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  NO2        m0273(.A(mai_mai_n295_), .B(mai_mai_n289_), .Y(mai_mai_n296_));
  NO2        m0274(.A(i_3_), .B(i_10_), .Y(mai_mai_n297_));
  NA3        m0275(.A(mai_mai_n297_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n298_));
  NO2        m0276(.A(i_2_), .B(mai_mai_n104_), .Y(mai_mai_n299_));
  NA2        m0277(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n300_));
  NO2        m0278(.A(mai_mai_n300_), .B(i_8_), .Y(mai_mai_n301_));
  NOi21      m0279(.An(mai_mai_n223_), .B(mai_mai_n106_), .Y(mai_mai_n302_));
  NA3        m0280(.A(mai_mai_n302_), .B(mai_mai_n301_), .C(mai_mai_n299_), .Y(mai_mai_n303_));
  AN2        m0281(.A(i_3_), .B(i_10_), .Y(mai_mai_n304_));
  NA4        m0282(.A(mai_mai_n304_), .B(mai_mai_n203_), .C(mai_mai_n180_), .D(mai_mai_n178_), .Y(mai_mai_n305_));
  NO2        m0283(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n306_));
  NO2        m0284(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n307_));
  OR2        m0285(.A(mai_mai_n303_), .B(mai_mai_n298_), .Y(mai_mai_n308_));
  OAI220     m0286(.A0(mai_mai_n308_), .A1(i_6_), .B0(mai_mai_n296_), .B1(mai_mai_n284_), .Y(mai_mai_n309_));
  NO4        m0287(.A(mai_mai_n309_), .B(mai_mai_n282_), .C(mai_mai_n220_), .D(mai_mai_n171_), .Y(mai_mai_n310_));
  NO3        m0288(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n311_));
  NO2        m0289(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n312_));
  NA2        m0290(.A(mai_mai_n290_), .B(mai_mai_n312_), .Y(mai_mai_n313_));
  NO3        m0291(.A(i_6_), .B(mai_mai_n198_), .C(i_7_), .Y(mai_mai_n314_));
  NA2        m0292(.A(mai_mai_n314_), .B(mai_mai_n203_), .Y(mai_mai_n315_));
  AOI210     m0293(.A0(mai_mai_n315_), .A1(mai_mai_n313_), .B0(mai_mai_n173_), .Y(mai_mai_n316_));
  NO2        m0294(.A(i_2_), .B(i_3_), .Y(mai_mai_n317_));
  OR2        m0295(.A(i_0_), .B(i_5_), .Y(mai_mai_n318_));
  NA2        m0296(.A(mai_mai_n223_), .B(mai_mai_n318_), .Y(mai_mai_n319_));
  NA4        m0297(.A(mai_mai_n319_), .B(mai_mai_n232_), .C(mai_mai_n317_), .D(i_1_), .Y(mai_mai_n320_));
  NA3        m0298(.A(mai_mai_n290_), .B(mai_mai_n286_), .C(mai_mai_n116_), .Y(mai_mai_n321_));
  NAi21      m0299(.An(i_8_), .B(i_7_), .Y(mai_mai_n322_));
  NO2        m0300(.A(mai_mai_n322_), .B(i_6_), .Y(mai_mai_n323_));
  NO2        m0301(.A(mai_mai_n160_), .B(mai_mai_n47_), .Y(mai_mai_n324_));
  NA3        m0302(.A(mai_mai_n324_), .B(mai_mai_n323_), .C(mai_mai_n166_), .Y(mai_mai_n325_));
  NA3        m0303(.A(mai_mai_n325_), .B(mai_mai_n321_), .C(mai_mai_n320_), .Y(mai_mai_n326_));
  OAI210     m0304(.A0(mai_mai_n326_), .A1(mai_mai_n316_), .B0(i_4_), .Y(mai_mai_n327_));
  NO2        m0305(.A(i_12_), .B(i_10_), .Y(mai_mai_n328_));
  NOi21      m0306(.An(i_5_), .B(i_0_), .Y(mai_mai_n329_));
  NA4        m0307(.A(mai_mai_n85_), .B(mai_mai_n36_), .C(mai_mai_n87_), .D(i_8_), .Y(mai_mai_n330_));
  NO2        m0308(.A(i_6_), .B(i_8_), .Y(mai_mai_n331_));
  NOi21      m0309(.An(i_0_), .B(i_2_), .Y(mai_mai_n332_));
  AN2        m0310(.A(mai_mai_n332_), .B(mai_mai_n331_), .Y(mai_mai_n333_));
  NO2        m0311(.A(i_1_), .B(i_7_), .Y(mai_mai_n334_));
  AO220      m0312(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n323_), .B1(mai_mai_n233_), .Y(mai_mai_n335_));
  NA2        m0313(.A(mai_mai_n335_), .B(mai_mai_n42_), .Y(mai_mai_n336_));
  NA2        m0314(.A(mai_mai_n336_), .B(mai_mai_n327_), .Y(mai_mai_n337_));
  NO3        m0315(.A(mai_mai_n231_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n338_));
  NO3        m0316(.A(mai_mai_n322_), .B(i_2_), .C(i_1_), .Y(mai_mai_n339_));
  OAI210     m0317(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(i_6_), .Y(mai_mai_n340_));
  NO2        m0318(.A(mai_mai_n340_), .B(mai_mai_n319_), .Y(mai_mai_n341_));
  NOi21      m0319(.An(mai_mai_n156_), .B(mai_mai_n107_), .Y(mai_mai_n342_));
  NO2        m0320(.A(mai_mai_n342_), .B(mai_mai_n127_), .Y(mai_mai_n343_));
  OAI210     m0321(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(i_3_), .Y(mai_mai_n344_));
  INV        m0322(.A(mai_mai_n85_), .Y(mai_mai_n345_));
  NO2        m0323(.A(mai_mai_n291_), .B(mai_mai_n82_), .Y(mai_mai_n346_));
  NA2        m0324(.A(mai_mai_n346_), .B(mai_mai_n135_), .Y(mai_mai_n347_));
  NO2        m0325(.A(mai_mai_n96_), .B(mai_mai_n198_), .Y(mai_mai_n348_));
  NA3        m0326(.A(mai_mai_n302_), .B(mai_mai_n348_), .C(mai_mai_n64_), .Y(mai_mai_n349_));
  AOI210     m0327(.A0(mai_mai_n349_), .A1(mai_mai_n347_), .B0(mai_mai_n345_), .Y(mai_mai_n350_));
  NO2        m0328(.A(mai_mai_n198_), .B(i_9_), .Y(mai_mai_n351_));
  NA2        m0329(.A(mai_mai_n351_), .B(mai_mai_n210_), .Y(mai_mai_n352_));
  NO2        m0330(.A(mai_mai_n352_), .B(mai_mai_n47_), .Y(mai_mai_n353_));
  NO2        m0331(.A(mai_mai_n353_), .B(mai_mai_n350_), .Y(mai_mai_n354_));
  AOI210     m0332(.A0(mai_mai_n354_), .A1(mai_mai_n344_), .B0(mai_mai_n165_), .Y(mai_mai_n355_));
  AOI210     m0333(.A0(mai_mai_n337_), .A1(mai_mai_n311_), .B0(mai_mai_n355_), .Y(mai_mai_n356_));
  NOi32      m0334(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n357_));
  INV        m0335(.A(mai_mai_n357_), .Y(mai_mai_n358_));
  NAi21      m0336(.An(i_0_), .B(i_6_), .Y(mai_mai_n359_));
  NAi21      m0337(.An(i_1_), .B(i_5_), .Y(mai_mai_n360_));
  NA2        m0338(.A(mai_mai_n360_), .B(mai_mai_n359_), .Y(mai_mai_n361_));
  NA2        m0339(.A(mai_mai_n361_), .B(mai_mai_n25_), .Y(mai_mai_n362_));
  OAI210     m0340(.A0(mai_mai_n362_), .A1(mai_mai_n162_), .B0(mai_mai_n245_), .Y(mai_mai_n363_));
  NAi41      m0341(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n364_));
  OAI220     m0342(.A0(mai_mai_n364_), .A1(mai_mai_n360_), .B0(mai_mai_n224_), .B1(mai_mai_n162_), .Y(mai_mai_n365_));
  NO2        m0343(.A(mai_mai_n162_), .B(mai_mai_n160_), .Y(mai_mai_n366_));
  NOi32      m0344(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n367_));
  NAi21      m0345(.An(i_6_), .B(i_1_), .Y(mai_mai_n368_));
  NA3        m0346(.A(mai_mai_n368_), .B(mai_mai_n367_), .C(mai_mai_n47_), .Y(mai_mai_n369_));
  NO2        m0347(.A(mai_mai_n369_), .B(i_0_), .Y(mai_mai_n370_));
  OR3        m0348(.A(mai_mai_n370_), .B(mai_mai_n366_), .C(mai_mai_n365_), .Y(mai_mai_n371_));
  NO2        m0349(.A(i_1_), .B(mai_mai_n104_), .Y(mai_mai_n372_));
  NAi21      m0350(.An(i_3_), .B(i_4_), .Y(mai_mai_n373_));
  NO2        m0351(.A(mai_mai_n373_), .B(i_9_), .Y(mai_mai_n374_));
  AN2        m0352(.A(i_6_), .B(i_7_), .Y(mai_mai_n375_));
  OAI210     m0353(.A0(mai_mai_n375_), .A1(mai_mai_n372_), .B0(mai_mai_n374_), .Y(mai_mai_n376_));
  NA2        m0354(.A(i_2_), .B(i_7_), .Y(mai_mai_n377_));
  NO2        m0355(.A(mai_mai_n373_), .B(i_10_), .Y(mai_mai_n378_));
  NO2        m0356(.A(mai_mai_n376_), .B(mai_mai_n190_), .Y(mai_mai_n379_));
  AOI210     m0357(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n380_));
  OAI210     m0358(.A0(mai_mai_n380_), .A1(mai_mai_n193_), .B0(mai_mai_n378_), .Y(mai_mai_n381_));
  AOI220     m0359(.A0(mai_mai_n378_), .A1(mai_mai_n334_), .B0(mai_mai_n237_), .B1(mai_mai_n193_), .Y(mai_mai_n382_));
  AOI210     m0360(.A0(mai_mai_n382_), .A1(mai_mai_n381_), .B0(i_5_), .Y(mai_mai_n383_));
  NO4        m0361(.A(mai_mai_n383_), .B(mai_mai_n379_), .C(mai_mai_n371_), .D(mai_mai_n363_), .Y(mai_mai_n384_));
  NO2        m0362(.A(mai_mai_n384_), .B(mai_mai_n358_), .Y(mai_mai_n385_));
  NO2        m0363(.A(mai_mai_n60_), .B(mai_mai_n25_), .Y(mai_mai_n386_));
  AN2        m0364(.A(i_12_), .B(i_5_), .Y(mai_mai_n387_));
  NO2        m0365(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n388_));
  INV        m0366(.A(mai_mai_n387_), .Y(mai_mai_n389_));
  NO2        m0367(.A(i_11_), .B(i_6_), .Y(mai_mai_n390_));
  NO2        m0368(.A(mai_mai_n241_), .B(i_5_), .Y(mai_mai_n391_));
  NO2        m0369(.A(i_5_), .B(i_10_), .Y(mai_mai_n392_));
  AOI220     m0370(.A0(mai_mai_n392_), .A1(mai_mai_n271_), .B0(mai_mai_n391_), .B1(mai_mai_n203_), .Y(mai_mai_n393_));
  NA2        m0371(.A(mai_mai_n147_), .B(mai_mai_n46_), .Y(mai_mai_n394_));
  NO2        m0372(.A(mai_mai_n394_), .B(mai_mai_n393_), .Y(mai_mai_n395_));
  NA2        m0373(.A(mai_mai_n395_), .B(mai_mai_n386_), .Y(mai_mai_n396_));
  NO2        m0374(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n397_));
  NO3        m0375(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n398_));
  NO2        m0376(.A(i_11_), .B(i_12_), .Y(mai_mai_n399_));
  NA3        m0377(.A(mai_mai_n116_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n400_));
  NO2        m0378(.A(mai_mai_n400_), .B(mai_mai_n224_), .Y(mai_mai_n401_));
  NAi21      m0379(.An(i_13_), .B(i_0_), .Y(mai_mai_n402_));
  NO2        m0380(.A(mai_mai_n402_), .B(mai_mai_n238_), .Y(mai_mai_n403_));
  NA2        m0381(.A(mai_mai_n401_), .B(mai_mai_n403_), .Y(mai_mai_n404_));
  NA2        m0382(.A(mai_mai_n404_), .B(mai_mai_n396_), .Y(mai_mai_n405_));
  NO2        m0383(.A(i_0_), .B(i_11_), .Y(mai_mai_n406_));
  INV        m0384(.A(i_5_), .Y(mai_mai_n407_));
  AN2        m0385(.A(i_1_), .B(i_6_), .Y(mai_mai_n408_));
  NOi21      m0386(.An(i_2_), .B(i_12_), .Y(mai_mai_n409_));
  NA2        m0387(.A(mai_mai_n409_), .B(mai_mai_n408_), .Y(mai_mai_n410_));
  NO2        m0388(.A(mai_mai_n410_), .B(mai_mai_n407_), .Y(mai_mai_n411_));
  NA2        m0389(.A(mai_mai_n145_), .B(i_9_), .Y(mai_mai_n412_));
  NO2        m0390(.A(mai_mai_n412_), .B(i_4_), .Y(mai_mai_n413_));
  NA2        m0391(.A(mai_mai_n411_), .B(mai_mai_n413_), .Y(mai_mai_n414_));
  NAi21      m0392(.An(i_9_), .B(i_4_), .Y(mai_mai_n415_));
  OR2        m0393(.A(i_13_), .B(i_10_), .Y(mai_mai_n416_));
  NO3        m0394(.A(mai_mai_n416_), .B(mai_mai_n120_), .C(mai_mai_n415_), .Y(mai_mai_n417_));
  OR2        m0395(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n418_));
  NO2        m0396(.A(mai_mai_n104_), .B(mai_mai_n25_), .Y(mai_mai_n419_));
  NA2        m0397(.A(mai_mai_n283_), .B(mai_mai_n419_), .Y(mai_mai_n420_));
  NA2        m0398(.A(mai_mai_n276_), .B(mai_mai_n216_), .Y(mai_mai_n421_));
  OAI220     m0399(.A0(mai_mai_n421_), .A1(mai_mai_n418_), .B0(mai_mai_n420_), .B1(mai_mai_n342_), .Y(mai_mai_n422_));
  INV        m0400(.A(mai_mai_n422_), .Y(mai_mai_n423_));
  AOI210     m0401(.A0(mai_mai_n423_), .A1(mai_mai_n414_), .B0(mai_mai_n26_), .Y(mai_mai_n424_));
  NA2        m0402(.A(mai_mai_n321_), .B(mai_mai_n320_), .Y(mai_mai_n425_));
  AOI220     m0403(.A0(mai_mai_n293_), .A1(mai_mai_n287_), .B0(mai_mai_n290_), .B1(mai_mai_n312_), .Y(mai_mai_n426_));
  NO2        m0404(.A(mai_mai_n426_), .B(mai_mai_n173_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n187_), .B(mai_mai_n87_), .Y(mai_mai_n428_));
  AOI220     m0406(.A0(mai_mai_n428_), .A1(mai_mai_n292_), .B0(mai_mai_n278_), .B1(mai_mai_n216_), .Y(mai_mai_n429_));
  NO2        m0407(.A(mai_mai_n429_), .B(mai_mai_n285_), .Y(mai_mai_n430_));
  NO3        m0408(.A(mai_mai_n430_), .B(mai_mai_n427_), .C(mai_mai_n425_), .Y(mai_mai_n431_));
  NA2        m0409(.A(mai_mai_n201_), .B(mai_mai_n99_), .Y(mai_mai_n432_));
  NA3        m0410(.A(mai_mai_n324_), .B(mai_mai_n166_), .C(mai_mai_n87_), .Y(mai_mai_n433_));
  AOI210     m0411(.A0(mai_mai_n433_), .A1(mai_mai_n432_), .B0(mai_mai_n322_), .Y(mai_mai_n434_));
  NA2        m0412(.A(mai_mai_n198_), .B(i_10_), .Y(mai_mai_n435_));
  NA3        m0413(.A(mai_mai_n257_), .B(mai_mai_n65_), .C(i_2_), .Y(mai_mai_n436_));
  NA2        m0414(.A(mai_mai_n293_), .B(mai_mai_n233_), .Y(mai_mai_n437_));
  OAI220     m0415(.A0(mai_mai_n437_), .A1(mai_mai_n187_), .B0(mai_mai_n436_), .B1(mai_mai_n435_), .Y(mai_mai_n438_));
  NO2        m0416(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n439_));
  NA3        m0417(.A(mai_mai_n334_), .B(mai_mai_n333_), .C(mai_mai_n439_), .Y(mai_mai_n440_));
  NA2        m0418(.A(mai_mai_n314_), .B(mai_mai_n319_), .Y(mai_mai_n441_));
  OAI210     m0419(.A0(mai_mai_n441_), .A1(mai_mai_n194_), .B0(mai_mai_n440_), .Y(mai_mai_n442_));
  NO3        m0420(.A(mai_mai_n442_), .B(mai_mai_n438_), .C(mai_mai_n434_), .Y(mai_mai_n443_));
  AOI210     m0421(.A0(mai_mai_n443_), .A1(mai_mai_n431_), .B0(mai_mai_n272_), .Y(mai_mai_n444_));
  NO4        m0422(.A(mai_mai_n444_), .B(mai_mai_n424_), .C(mai_mai_n405_), .D(mai_mai_n385_), .Y(mai_mai_n445_));
  NO2        m0423(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n446_));
  NO2        m0424(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n447_));
  NA3        m0425(.A(mai_mai_n447_), .B(mai_mai_n446_), .C(i_2_), .Y(mai_mai_n448_));
  NO2        m0426(.A(i_10_), .B(i_9_), .Y(mai_mai_n449_));
  NAi21      m0427(.An(i_12_), .B(i_8_), .Y(mai_mai_n450_));
  NO2        m0428(.A(mai_mai_n450_), .B(i_3_), .Y(mai_mai_n451_));
  NA2        m0429(.A(mai_mai_n451_), .B(mai_mai_n449_), .Y(mai_mai_n452_));
  NO2        m0430(.A(mai_mai_n47_), .B(i_4_), .Y(mai_mai_n453_));
  NO2        m0431(.A(mai_mai_n452_), .B(mai_mai_n448_), .Y(mai_mai_n454_));
  NA2        m0432(.A(mai_mai_n307_), .B(i_0_), .Y(mai_mai_n455_));
  NO3        m0433(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n456_));
  NA2        m0434(.A(mai_mai_n269_), .B(mai_mai_n100_), .Y(mai_mai_n457_));
  NA2        m0435(.A(mai_mai_n457_), .B(mai_mai_n456_), .Y(mai_mai_n458_));
  NA2        m0436(.A(i_8_), .B(i_9_), .Y(mai_mai_n459_));
  NO2        m0437(.A(mai_mai_n458_), .B(mai_mai_n455_), .Y(mai_mai_n460_));
  NA2        m0438(.A(mai_mai_n250_), .B(mai_mai_n306_), .Y(mai_mai_n461_));
  NO3        m0439(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n462_));
  INV        m0440(.A(mai_mai_n462_), .Y(mai_mai_n463_));
  NA3        m0441(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n464_));
  NA4        m0442(.A(mai_mai_n148_), .B(mai_mai_n119_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n465_));
  OAI220     m0443(.A0(mai_mai_n465_), .A1(mai_mai_n464_), .B0(mai_mai_n463_), .B1(mai_mai_n461_), .Y(mai_mai_n466_));
  NO3        m0444(.A(mai_mai_n466_), .B(mai_mai_n460_), .C(mai_mai_n454_), .Y(mai_mai_n467_));
  NA2        m0445(.A(mai_mai_n292_), .B(mai_mai_n111_), .Y(mai_mai_n468_));
  OR2        m0446(.A(mai_mai_n468_), .B(mai_mai_n212_), .Y(mai_mai_n469_));
  OA210      m0447(.A0(mai_mai_n352_), .A1(mai_mai_n104_), .B0(mai_mai_n294_), .Y(mai_mai_n470_));
  OA220      m0448(.A0(mai_mai_n470_), .A1(mai_mai_n165_), .B0(mai_mai_n469_), .B1(mai_mai_n230_), .Y(mai_mai_n471_));
  NA2        m0449(.A(mai_mai_n99_), .B(i_13_), .Y(mai_mai_n472_));
  NO2        m0450(.A(i_2_), .B(i_13_), .Y(mai_mai_n473_));
  NO3        m0451(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n474_));
  NO2        m0452(.A(i_6_), .B(i_7_), .Y(mai_mai_n475_));
  NA2        m0453(.A(mai_mai_n475_), .B(mai_mai_n474_), .Y(mai_mai_n476_));
  NO2        m0454(.A(i_11_), .B(i_1_), .Y(mai_mai_n477_));
  NO2        m0455(.A(mai_mai_n74_), .B(i_3_), .Y(mai_mai_n478_));
  OR2        m0456(.A(i_11_), .B(i_8_), .Y(mai_mai_n479_));
  NOi21      m0457(.An(i_2_), .B(i_7_), .Y(mai_mai_n480_));
  NAi31      m0458(.An(mai_mai_n479_), .B(mai_mai_n480_), .C(mai_mai_n478_), .Y(mai_mai_n481_));
  NO2        m0459(.A(mai_mai_n416_), .B(i_6_), .Y(mai_mai_n482_));
  NA2        m0460(.A(mai_mai_n482_), .B(mai_mai_n446_), .Y(mai_mai_n483_));
  NO2        m0461(.A(mai_mai_n483_), .B(mai_mai_n481_), .Y(mai_mai_n484_));
  NO2        m0462(.A(i_3_), .B(mai_mai_n198_), .Y(mai_mai_n485_));
  NO2        m0463(.A(i_6_), .B(i_10_), .Y(mai_mai_n486_));
  NA4        m0464(.A(mai_mai_n486_), .B(mai_mai_n311_), .C(mai_mai_n485_), .D(mai_mai_n235_), .Y(mai_mai_n487_));
  NO2        m0465(.A(mai_mai_n487_), .B(mai_mai_n158_), .Y(mai_mai_n488_));
  NA3        m0466(.A(mai_mai_n244_), .B(mai_mai_n175_), .C(mai_mai_n135_), .Y(mai_mai_n489_));
  NA2        m0467(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n490_));
  NO2        m0468(.A(mai_mai_n160_), .B(i_3_), .Y(mai_mai_n491_));
  NAi31      m0469(.An(mai_mai_n490_), .B(mai_mai_n491_), .C(mai_mai_n227_), .Y(mai_mai_n492_));
  NA3        m0470(.A(mai_mai_n397_), .B(mai_mai_n183_), .C(mai_mai_n152_), .Y(mai_mai_n493_));
  NA3        m0471(.A(mai_mai_n493_), .B(mai_mai_n492_), .C(mai_mai_n489_), .Y(mai_mai_n494_));
  NO3        m0472(.A(mai_mai_n494_), .B(mai_mai_n488_), .C(mai_mai_n484_), .Y(mai_mai_n495_));
  NA2        m0473(.A(mai_mai_n456_), .B(mai_mai_n387_), .Y(mai_mai_n496_));
  NAi21      m0474(.An(mai_mai_n222_), .B(mai_mai_n399_), .Y(mai_mai_n497_));
  NO2        m0475(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n498_));
  NO2        m0476(.A(i_0_), .B(mai_mai_n87_), .Y(mai_mai_n499_));
  NA3        m0477(.A(mai_mai_n499_), .B(mai_mai_n498_), .C(mai_mai_n145_), .Y(mai_mai_n500_));
  OR3        m0478(.A(mai_mai_n300_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n501_));
  NO2        m0479(.A(mai_mai_n501_), .B(mai_mai_n500_), .Y(mai_mai_n502_));
  NA2        m0480(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n503_));
  NA2        m0481(.A(mai_mai_n311_), .B(mai_mai_n237_), .Y(mai_mai_n504_));
  OAI220     m0482(.A0(mai_mai_n504_), .A1(mai_mai_n436_), .B0(mai_mai_n503_), .B1(mai_mai_n472_), .Y(mai_mai_n505_));
  NA4        m0483(.A(mai_mai_n304_), .B(mai_mai_n225_), .C(mai_mai_n74_), .D(mai_mai_n235_), .Y(mai_mai_n506_));
  NO2        m0484(.A(mai_mai_n506_), .B(mai_mai_n476_), .Y(mai_mai_n507_));
  NO3        m0485(.A(mai_mai_n507_), .B(mai_mai_n505_), .C(mai_mai_n502_), .Y(mai_mai_n508_));
  NA4        m0486(.A(mai_mai_n508_), .B(mai_mai_n495_), .C(mai_mai_n471_), .D(mai_mai_n467_), .Y(mai_mai_n509_));
  NA3        m0487(.A(mai_mai_n304_), .B(mai_mai_n180_), .C(mai_mai_n178_), .Y(mai_mai_n510_));
  OAI210     m0488(.A0(mai_mai_n298_), .A1(mai_mai_n185_), .B0(mai_mai_n510_), .Y(mai_mai_n511_));
  AN2        m0489(.A(mai_mai_n287_), .B(mai_mai_n232_), .Y(mai_mai_n512_));
  NA2        m0490(.A(mai_mai_n512_), .B(mai_mai_n511_), .Y(mai_mai_n513_));
  NA2        m0491(.A(mai_mai_n311_), .B(mai_mai_n167_), .Y(mai_mai_n514_));
  OAI210     m0492(.A0(mai_mai_n514_), .A1(mai_mai_n230_), .B0(mai_mai_n305_), .Y(mai_mai_n515_));
  NA2        m0493(.A(mai_mai_n515_), .B(mai_mai_n323_), .Y(mai_mai_n516_));
  NA4        m0494(.A(mai_mai_n447_), .B(mai_mai_n446_), .C(mai_mai_n208_), .D(i_2_), .Y(mai_mai_n517_));
  INV        m0495(.A(mai_mai_n517_), .Y(mai_mai_n518_));
  NA2        m0496(.A(mai_mai_n387_), .B(mai_mai_n226_), .Y(mai_mai_n519_));
  NA2        m0497(.A(mai_mai_n357_), .B(mai_mai_n74_), .Y(mai_mai_n520_));
  NA2        m0498(.A(mai_mai_n375_), .B(mai_mai_n367_), .Y(mai_mai_n521_));
  OR2        m0499(.A(mai_mai_n519_), .B(mai_mai_n521_), .Y(mai_mai_n522_));
  NO2        m0500(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n523_));
  NAi41      m0501(.An(mai_mai_n520_), .B(mai_mai_n486_), .C(mai_mai_n523_), .D(mai_mai_n47_), .Y(mai_mai_n524_));
  AOI210     m0502(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n417_), .Y(mai_mai_n525_));
  NA3        m0503(.A(mai_mai_n525_), .B(mai_mai_n524_), .C(mai_mai_n522_), .Y(mai_mai_n526_));
  AOI210     m0504(.A0(mai_mai_n518_), .A1(mai_mai_n209_), .B0(mai_mai_n526_), .Y(mai_mai_n527_));
  AOI210     m0505(.A0(mai_mai_n199_), .A1(i_9_), .B0(mai_mai_n268_), .Y(mai_mai_n528_));
  NO2        m0506(.A(mai_mai_n528_), .B(mai_mai_n204_), .Y(mai_mai_n529_));
  NO2        m0507(.A(mai_mai_n187_), .B(mai_mai_n87_), .Y(mai_mai_n530_));
  NA2        m0508(.A(mai_mai_n530_), .B(mai_mai_n529_), .Y(mai_mai_n531_));
  NA4        m0509(.A(mai_mai_n531_), .B(mai_mai_n527_), .C(mai_mai_n516_), .D(mai_mai_n513_), .Y(mai_mai_n532_));
  NA2        m0510(.A(mai_mai_n391_), .B(mai_mai_n292_), .Y(mai_mai_n533_));
  OAI210     m0511(.A0(mai_mai_n389_), .A1(mai_mai_n172_), .B0(mai_mai_n533_), .Y(mai_mai_n534_));
  NO2        m0512(.A(i_12_), .B(mai_mai_n198_), .Y(mai_mai_n535_));
  NA2        m0513(.A(mai_mai_n535_), .B(mai_mai_n226_), .Y(mai_mai_n536_));
  NO3        m0514(.A(mai_mai_n1033_), .B(mai_mai_n536_), .C(mai_mai_n468_), .Y(mai_mai_n537_));
  NOi31      m0515(.An(mai_mai_n314_), .B(mai_mai_n416_), .C(mai_mai_n38_), .Y(mai_mai_n538_));
  OAI210     m0516(.A0(mai_mai_n538_), .A1(mai_mai_n537_), .B0(mai_mai_n534_), .Y(mai_mai_n539_));
  NO2        m0517(.A(i_8_), .B(i_7_), .Y(mai_mai_n540_));
  OAI210     m0518(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n541_));
  NA2        m0519(.A(mai_mai_n541_), .B(mai_mai_n225_), .Y(mai_mai_n542_));
  AOI220     m0520(.A0(mai_mai_n324_), .A1(mai_mai_n40_), .B0(mai_mai_n233_), .B1(mai_mai_n211_), .Y(mai_mai_n543_));
  OAI220     m0521(.A0(mai_mai_n543_), .A1(mai_mai_n187_), .B0(mai_mai_n542_), .B1(mai_mai_n241_), .Y(mai_mai_n544_));
  NA2        m0522(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n545_));
  NO2        m0523(.A(mai_mai_n545_), .B(i_6_), .Y(mai_mai_n546_));
  NA3        m0524(.A(mai_mai_n546_), .B(mai_mai_n544_), .C(mai_mai_n540_), .Y(mai_mai_n547_));
  NO2        m0525(.A(mai_mai_n472_), .B(mai_mai_n136_), .Y(mai_mai_n548_));
  NA2        m0526(.A(mai_mai_n548_), .B(mai_mai_n268_), .Y(mai_mai_n549_));
  NOi31      m0527(.An(mai_mai_n290_), .B(mai_mai_n298_), .C(mai_mai_n185_), .Y(mai_mai_n550_));
  NA2        m0528(.A(mai_mai_n550_), .B(mai_mai_n462_), .Y(mai_mai_n551_));
  NA4        m0529(.A(mai_mai_n551_), .B(mai_mai_n549_), .C(mai_mai_n547_), .D(mai_mai_n539_), .Y(mai_mai_n552_));
  NA3        m0530(.A(mai_mai_n223_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n553_));
  NA2        m0531(.A(mai_mai_n283_), .B(mai_mai_n85_), .Y(mai_mai_n554_));
  AOI210     m0532(.A0(mai_mai_n553_), .A1(mai_mai_n347_), .B0(mai_mai_n554_), .Y(mai_mai_n555_));
  NA2        m0533(.A(mai_mai_n293_), .B(mai_mai_n287_), .Y(mai_mai_n556_));
  NO2        m0534(.A(mai_mai_n556_), .B(mai_mai_n177_), .Y(mai_mai_n557_));
  AOI210     m0535(.A0(mai_mai_n368_), .A1(mai_mai_n47_), .B0(mai_mai_n372_), .Y(mai_mai_n558_));
  NA2        m0536(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n559_));
  NA3        m0537(.A(mai_mai_n535_), .B(mai_mai_n274_), .C(mai_mai_n559_), .Y(mai_mai_n560_));
  NO2        m0538(.A(mai_mai_n558_), .B(mai_mai_n560_), .Y(mai_mai_n561_));
  NO3        m0539(.A(mai_mai_n561_), .B(mai_mai_n557_), .C(mai_mai_n555_), .Y(mai_mai_n562_));
  NO4        m0540(.A(mai_mai_n251_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n563_));
  NO3        m0541(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n564_));
  NO2        m0542(.A(mai_mai_n231_), .B(mai_mai_n36_), .Y(mai_mai_n565_));
  AN2        m0543(.A(mai_mai_n565_), .B(mai_mai_n564_), .Y(mai_mai_n566_));
  OA210      m0544(.A0(mai_mai_n566_), .A1(mai_mai_n563_), .B0(mai_mai_n357_), .Y(mai_mai_n567_));
  NO2        m0545(.A(mai_mai_n416_), .B(i_1_), .Y(mai_mai_n568_));
  NOi31      m0546(.An(mai_mai_n568_), .B(mai_mai_n457_), .C(mai_mai_n74_), .Y(mai_mai_n569_));
  AN4        m0547(.A(mai_mai_n569_), .B(mai_mai_n413_), .C(mai_mai_n498_), .D(i_2_), .Y(mai_mai_n570_));
  NO2        m0548(.A(mai_mai_n426_), .B(mai_mai_n181_), .Y(mai_mai_n571_));
  NO3        m0549(.A(mai_mai_n571_), .B(mai_mai_n570_), .C(mai_mai_n567_), .Y(mai_mai_n572_));
  NOi21      m0550(.An(i_10_), .B(i_6_), .Y(mai_mai_n573_));
  NO2        m0551(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n574_));
  NO2        m0552(.A(mai_mai_n118_), .B(mai_mai_n23_), .Y(mai_mai_n575_));
  NA2        m0553(.A(mai_mai_n314_), .B(mai_mai_n167_), .Y(mai_mai_n576_));
  AOI220     m0554(.A0(mai_mai_n576_), .A1(mai_mai_n437_), .B0(mai_mai_n188_), .B1(mai_mai_n186_), .Y(mai_mai_n577_));
  NO2        m0555(.A(mai_mai_n203_), .B(mai_mai_n37_), .Y(mai_mai_n578_));
  NOi31      m0556(.An(mai_mai_n149_), .B(mai_mai_n578_), .C(mai_mai_n330_), .Y(mai_mai_n579_));
  NO2        m0557(.A(mai_mai_n579_), .B(mai_mai_n577_), .Y(mai_mai_n580_));
  INV        m0558(.A(mai_mai_n317_), .Y(mai_mai_n581_));
  NO2        m0559(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n582_));
  NA2        m0560(.A(mai_mai_n178_), .B(i_0_), .Y(mai_mai_n583_));
  NO3        m0561(.A(mai_mai_n583_), .B(mai_mai_n340_), .C(mai_mai_n298_), .Y(mai_mai_n584_));
  OR2        m0562(.A(i_2_), .B(i_5_), .Y(mai_mai_n585_));
  OR2        m0563(.A(mai_mai_n585_), .B(mai_mai_n408_), .Y(mai_mai_n586_));
  AOI210     m0564(.A0(mai_mai_n377_), .A1(mai_mai_n243_), .B0(mai_mai_n203_), .Y(mai_mai_n587_));
  AOI210     m0565(.A0(mai_mai_n587_), .A1(mai_mai_n586_), .B0(mai_mai_n497_), .Y(mai_mai_n588_));
  NO2        m0566(.A(mai_mai_n588_), .B(mai_mai_n584_), .Y(mai_mai_n589_));
  NA4        m0567(.A(mai_mai_n589_), .B(mai_mai_n580_), .C(mai_mai_n572_), .D(mai_mai_n562_), .Y(mai_mai_n590_));
  NO4        m0568(.A(mai_mai_n590_), .B(mai_mai_n552_), .C(mai_mai_n532_), .D(mai_mai_n509_), .Y(mai_mai_n591_));
  NA4        m0569(.A(mai_mai_n591_), .B(mai_mai_n445_), .C(mai_mai_n356_), .D(mai_mai_n310_), .Y(mai7));
  NO2        m0570(.A(mai_mai_n96_), .B(mai_mai_n55_), .Y(mai_mai_n593_));
  NO2        m0571(.A(mai_mai_n111_), .B(mai_mai_n93_), .Y(mai_mai_n594_));
  NA2        m0572(.A(mai_mai_n388_), .B(mai_mai_n594_), .Y(mai_mai_n595_));
  NA2        m0573(.A(mai_mai_n486_), .B(mai_mai_n85_), .Y(mai_mai_n596_));
  NA2        m0574(.A(i_11_), .B(mai_mai_n198_), .Y(mai_mai_n597_));
  NA2        m0575(.A(mai_mai_n147_), .B(mai_mai_n597_), .Y(mai_mai_n598_));
  OAI210     m0576(.A0(mai_mai_n598_), .A1(mai_mai_n596_), .B0(mai_mai_n595_), .Y(mai_mai_n599_));
  NA3        m0577(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n600_));
  NO2        m0578(.A(mai_mai_n235_), .B(i_4_), .Y(mai_mai_n601_));
  NA2        m0579(.A(mai_mai_n601_), .B(i_8_), .Y(mai_mai_n602_));
  NO2        m0580(.A(mai_mai_n108_), .B(mai_mai_n600_), .Y(mai_mai_n603_));
  NA2        m0581(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n604_));
  OAI210     m0582(.A0(mai_mai_n90_), .A1(mai_mai_n208_), .B0(mai_mai_n209_), .Y(mai_mai_n605_));
  NO2        m0583(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n606_));
  NA2        m0584(.A(i_4_), .B(i_8_), .Y(mai_mai_n607_));
  AOI210     m0585(.A0(mai_mai_n607_), .A1(mai_mai_n304_), .B0(mai_mai_n606_), .Y(mai_mai_n608_));
  OAI220     m0586(.A0(mai_mai_n608_), .A1(mai_mai_n604_), .B0(mai_mai_n605_), .B1(i_13_), .Y(mai_mai_n609_));
  NO4        m0587(.A(mai_mai_n609_), .B(mai_mai_n603_), .C(mai_mai_n599_), .D(mai_mai_n593_), .Y(mai_mai_n610_));
  AOI210     m0588(.A0(mai_mai_n131_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n611_));
  AOI210     m0589(.A0(mai_mai_n611_), .A1(mai_mai_n235_), .B0(mai_mai_n164_), .Y(mai_mai_n612_));
  OR2        m0590(.A(i_6_), .B(i_10_), .Y(mai_mai_n613_));
  NO2        m0591(.A(mai_mai_n613_), .B(mai_mai_n23_), .Y(mai_mai_n614_));
  OR3        m0592(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n615_));
  NO3        m0593(.A(mai_mai_n615_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n616_));
  INV        m0594(.A(mai_mai_n205_), .Y(mai_mai_n617_));
  NO2        m0595(.A(mai_mai_n616_), .B(mai_mai_n614_), .Y(mai_mai_n618_));
  OA220      m0596(.A0(mai_mai_n618_), .A1(mai_mai_n581_), .B0(mai_mai_n612_), .B1(mai_mai_n270_), .Y(mai_mai_n619_));
  AOI210     m0597(.A0(mai_mai_n619_), .A1(mai_mai_n610_), .B0(mai_mai_n64_), .Y(mai_mai_n620_));
  NOi21      m0598(.An(i_11_), .B(i_7_), .Y(mai_mai_n621_));
  AO210      m0599(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n622_));
  NO2        m0600(.A(mai_mai_n622_), .B(mai_mai_n621_), .Y(mai_mai_n623_));
  NA2        m0601(.A(mai_mai_n623_), .B(mai_mai_n211_), .Y(mai_mai_n624_));
  NA3        m0602(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n625_));
  NO2        m0603(.A(mai_mai_n624_), .B(mai_mai_n64_), .Y(mai_mai_n626_));
  NA2        m0604(.A(mai_mai_n89_), .B(mai_mai_n64_), .Y(mai_mai_n627_));
  AO210      m0605(.A0(mai_mai_n627_), .A1(mai_mai_n382_), .B0(mai_mai_n41_), .Y(mai_mai_n628_));
  NA2        m0606(.A(mai_mai_n227_), .B(mai_mai_n64_), .Y(mai_mai_n629_));
  NO2        m0607(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n630_));
  NO2        m0608(.A(i_1_), .B(i_12_), .Y(mai_mai_n631_));
  NA3        m0609(.A(mai_mai_n631_), .B(mai_mai_n113_), .C(mai_mai_n24_), .Y(mai_mai_n632_));
  BUFFER     m0610(.A(mai_mai_n632_), .Y(mai_mai_n633_));
  NA3        m0611(.A(mai_mai_n633_), .B(mai_mai_n629_), .C(mai_mai_n628_), .Y(mai_mai_n634_));
  OAI210     m0612(.A0(mai_mai_n634_), .A1(mai_mai_n626_), .B0(i_6_), .Y(mai_mai_n635_));
  NO2        m0613(.A(mai_mai_n625_), .B(mai_mai_n111_), .Y(mai_mai_n636_));
  NA2        m0614(.A(mai_mai_n636_), .B(mai_mai_n582_), .Y(mai_mai_n637_));
  NO2        m0615(.A(i_6_), .B(i_11_), .Y(mai_mai_n638_));
  NA2        m0616(.A(mai_mai_n637_), .B(mai_mai_n458_), .Y(mai_mai_n639_));
  NO4        m0617(.A(mai_mai_n221_), .B(mai_mai_n131_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n640_));
  NA2        m0618(.A(mai_mai_n640_), .B(mai_mai_n630_), .Y(mai_mai_n641_));
  NA2        m0619(.A(mai_mai_n235_), .B(i_6_), .Y(mai_mai_n642_));
  NA2        m0620(.A(i_1_), .B(mai_mai_n260_), .Y(mai_mai_n643_));
  OAI210     m0621(.A0(mai_mai_n643_), .A1(mai_mai_n45_), .B0(mai_mai_n641_), .Y(mai_mai_n644_));
  INV        m0622(.A(i_2_), .Y(mai_mai_n645_));
  NA2        m0623(.A(mai_mai_n141_), .B(i_9_), .Y(mai_mai_n646_));
  NA3        m0624(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n647_));
  NO2        m0625(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n648_));
  NA3        m0626(.A(mai_mai_n648_), .B(mai_mai_n269_), .C(mai_mai_n45_), .Y(mai_mai_n649_));
  OAI220     m0627(.A0(mai_mai_n649_), .A1(mai_mai_n647_), .B0(mai_mai_n646_), .B1(mai_mai_n645_), .Y(mai_mai_n650_));
  NA3        m0628(.A(mai_mai_n630_), .B(mai_mai_n317_), .C(i_6_), .Y(mai_mai_n651_));
  NO2        m0629(.A(mai_mai_n651_), .B(mai_mai_n23_), .Y(mai_mai_n652_));
  AOI210     m0630(.A0(mai_mai_n477_), .A1(mai_mai_n419_), .B0(mai_mai_n240_), .Y(mai_mai_n653_));
  NO2        m0631(.A(mai_mai_n653_), .B(mai_mai_n604_), .Y(mai_mai_n654_));
  NO2        m0632(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n655_));
  NA2        m0633(.A(mai_mai_n655_), .B(mai_mai_n24_), .Y(mai_mai_n656_));
  OR3        m0634(.A(mai_mai_n654_), .B(mai_mai_n652_), .C(mai_mai_n650_), .Y(mai_mai_n657_));
  NO3        m0635(.A(mai_mai_n657_), .B(mai_mai_n644_), .C(mai_mai_n639_), .Y(mai_mai_n658_));
  NO2        m0636(.A(mai_mai_n235_), .B(mai_mai_n104_), .Y(mai_mai_n659_));
  NO2        m0637(.A(mai_mai_n659_), .B(mai_mai_n621_), .Y(mai_mai_n660_));
  NA2        m0638(.A(mai_mai_n660_), .B(i_1_), .Y(mai_mai_n661_));
  NO2        m0639(.A(mai_mai_n661_), .B(mai_mai_n615_), .Y(mai_mai_n662_));
  NO2        m0640(.A(mai_mai_n415_), .B(mai_mai_n87_), .Y(mai_mai_n663_));
  NA2        m0641(.A(mai_mai_n662_), .B(mai_mai_n47_), .Y(mai_mai_n664_));
  NA2        m0642(.A(i_3_), .B(mai_mai_n198_), .Y(mai_mai_n665_));
  NO2        m0643(.A(mai_mai_n665_), .B(mai_mai_n118_), .Y(mai_mai_n666_));
  AN2        m0644(.A(mai_mai_n666_), .B(mai_mai_n546_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n231_), .B(mai_mai_n45_), .Y(mai_mai_n668_));
  NO3        m0646(.A(mai_mai_n668_), .B(mai_mai_n307_), .C(mai_mai_n236_), .Y(mai_mai_n669_));
  NO2        m0647(.A(mai_mai_n120_), .B(mai_mai_n37_), .Y(mai_mai_n670_));
  NO2        m0648(.A(mai_mai_n670_), .B(i_6_), .Y(mai_mai_n671_));
  NO2        m0649(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n672_));
  NO2        m0650(.A(mai_mai_n672_), .B(mai_mai_n64_), .Y(mai_mai_n673_));
  NO2        m0651(.A(mai_mai_n673_), .B(mai_mai_n631_), .Y(mai_mai_n674_));
  NO4        m0652(.A(mai_mai_n674_), .B(mai_mai_n671_), .C(mai_mai_n669_), .D(i_4_), .Y(mai_mai_n675_));
  NA2        m0653(.A(i_1_), .B(i_3_), .Y(mai_mai_n676_));
  NO2        m0654(.A(mai_mai_n459_), .B(mai_mai_n96_), .Y(mai_mai_n677_));
  AOI210     m0655(.A0(mai_mai_n668_), .A1(mai_mai_n573_), .B0(mai_mai_n677_), .Y(mai_mai_n678_));
  NO2        m0656(.A(mai_mai_n678_), .B(mai_mai_n676_), .Y(mai_mai_n679_));
  NO3        m0657(.A(mai_mai_n679_), .B(mai_mai_n675_), .C(mai_mai_n667_), .Y(mai_mai_n680_));
  NA4        m0658(.A(mai_mai_n680_), .B(mai_mai_n664_), .C(mai_mai_n658_), .D(mai_mai_n635_), .Y(mai_mai_n681_));
  AN2        m0659(.A(mai_mai_n244_), .B(mai_mai_n87_), .Y(mai_mai_n682_));
  NA2        m0660(.A(mai_mai_n375_), .B(mai_mai_n374_), .Y(mai_mai_n683_));
  INV        m0661(.A(mai_mai_n683_), .Y(mai_mai_n684_));
  OAI210     m0662(.A0(mai_mai_n684_), .A1(mai_mai_n682_), .B0(i_1_), .Y(mai_mai_n685_));
  AOI210     m0663(.A0(mai_mai_n269_), .A1(mai_mai_n100_), .B0(i_1_), .Y(mai_mai_n686_));
  NO2        m0664(.A(mai_mai_n373_), .B(i_2_), .Y(mai_mai_n687_));
  NA2        m0665(.A(mai_mai_n687_), .B(mai_mai_n686_), .Y(mai_mai_n688_));
  OAI210     m0666(.A0(mai_mai_n651_), .A1(mai_mai_n450_), .B0(mai_mai_n688_), .Y(mai_mai_n689_));
  INV        m0667(.A(mai_mai_n689_), .Y(mai_mai_n690_));
  AOI210     m0668(.A0(mai_mai_n690_), .A1(mai_mai_n685_), .B0(i_13_), .Y(mai_mai_n691_));
  OR2        m0669(.A(i_11_), .B(i_7_), .Y(mai_mai_n692_));
  NA3        m0670(.A(mai_mai_n692_), .B(mai_mai_n109_), .C(mai_mai_n141_), .Y(mai_mai_n693_));
  AOI220     m0671(.A0(mai_mai_n473_), .A1(mai_mai_n164_), .B0(mai_mai_n453_), .B1(mai_mai_n141_), .Y(mai_mai_n694_));
  OAI210     m0672(.A0(mai_mai_n694_), .A1(mai_mai_n45_), .B0(mai_mai_n693_), .Y(mai_mai_n695_));
  NO2        m0673(.A(mai_mai_n55_), .B(i_12_), .Y(mai_mai_n696_));
  INV        m0674(.A(mai_mai_n696_), .Y(mai_mai_n697_));
  NO2        m0675(.A(mai_mai_n480_), .B(mai_mai_n24_), .Y(mai_mai_n698_));
  AOI220     m0676(.A0(mai_mai_n698_), .A1(mai_mai_n663_), .B0(mai_mai_n244_), .B1(mai_mai_n134_), .Y(mai_mai_n699_));
  OAI220     m0677(.A0(mai_mai_n699_), .A1(mai_mai_n41_), .B0(mai_mai_n697_), .B1(mai_mai_n96_), .Y(mai_mai_n700_));
  AOI210     m0678(.A0(mai_mai_n695_), .A1(mai_mai_n331_), .B0(mai_mai_n700_), .Y(mai_mai_n701_));
  INV        m0679(.A(mai_mai_n118_), .Y(mai_mai_n702_));
  AOI220     m0680(.A0(mai_mai_n702_), .A1(mai_mai_n73_), .B0(mai_mai_n390_), .B1(mai_mai_n648_), .Y(mai_mai_n703_));
  NO2        m0681(.A(mai_mai_n703_), .B(mai_mai_n241_), .Y(mai_mai_n704_));
  AOI210     m0682(.A0(mai_mai_n450_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n705_));
  NOi31      m0683(.An(mai_mai_n705_), .B(mai_mai_n596_), .C(mai_mai_n45_), .Y(mai_mai_n706_));
  NA2        m0684(.A(mai_mai_n130_), .B(i_13_), .Y(mai_mai_n707_));
  NO2        m0685(.A(mai_mai_n647_), .B(mai_mai_n118_), .Y(mai_mai_n708_));
  INV        m0686(.A(mai_mai_n708_), .Y(mai_mai_n709_));
  OAI220     m0687(.A0(mai_mai_n709_), .A1(mai_mai_n72_), .B0(mai_mai_n707_), .B1(mai_mai_n686_), .Y(mai_mai_n710_));
  NO3        m0688(.A(mai_mai_n72_), .B(mai_mai_n32_), .C(mai_mai_n104_), .Y(mai_mai_n711_));
  NA2        m0689(.A(mai_mai_n26_), .B(mai_mai_n198_), .Y(mai_mai_n712_));
  NA2        m0690(.A(mai_mai_n712_), .B(i_7_), .Y(mai_mai_n713_));
  NO3        m0691(.A(mai_mai_n480_), .B(mai_mai_n235_), .C(mai_mai_n87_), .Y(mai_mai_n714_));
  AOI210     m0692(.A0(mai_mai_n714_), .A1(mai_mai_n713_), .B0(mai_mai_n711_), .Y(mai_mai_n715_));
  AOI220     m0693(.A0(mai_mai_n390_), .A1(mai_mai_n648_), .B0(mai_mai_n95_), .B1(mai_mai_n105_), .Y(mai_mai_n716_));
  OAI220     m0694(.A0(mai_mai_n716_), .A1(mai_mai_n602_), .B0(mai_mai_n715_), .B1(mai_mai_n617_), .Y(mai_mai_n717_));
  NO4        m0695(.A(mai_mai_n717_), .B(mai_mai_n710_), .C(mai_mai_n706_), .D(mai_mai_n704_), .Y(mai_mai_n718_));
  OR2        m0696(.A(i_11_), .B(i_6_), .Y(mai_mai_n719_));
  NA3        m0697(.A(mai_mai_n601_), .B(mai_mai_n712_), .C(i_7_), .Y(mai_mai_n720_));
  AOI210     m0698(.A0(mai_mai_n720_), .A1(mai_mai_n709_), .B0(mai_mai_n719_), .Y(mai_mai_n721_));
  NA3        m0699(.A(mai_mai_n409_), .B(mai_mai_n606_), .C(mai_mai_n100_), .Y(mai_mai_n722_));
  NA2        m0700(.A(mai_mai_n638_), .B(i_13_), .Y(mai_mai_n723_));
  NAi21      m0701(.An(i_11_), .B(i_12_), .Y(mai_mai_n724_));
  NOi41      m0702(.An(mai_mai_n114_), .B(mai_mai_n724_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n725_));
  NO3        m0703(.A(mai_mai_n480_), .B(mai_mai_n582_), .C(mai_mai_n607_), .Y(mai_mai_n726_));
  AOI220     m0704(.A0(mai_mai_n726_), .A1(mai_mai_n311_), .B0(mai_mai_n725_), .B1(mai_mai_n47_), .Y(mai_mai_n727_));
  NA3        m0705(.A(mai_mai_n727_), .B(mai_mai_n723_), .C(mai_mai_n722_), .Y(mai_mai_n728_));
  OAI210     m0706(.A0(mai_mai_n728_), .A1(mai_mai_n721_), .B0(mai_mai_n64_), .Y(mai_mai_n729_));
  NO2        m0707(.A(i_2_), .B(i_12_), .Y(mai_mai_n730_));
  NA2        m0708(.A(mai_mai_n372_), .B(mai_mai_n730_), .Y(mai_mai_n731_));
  NA2        m0709(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n732_));
  NO3        m0710(.A(mai_mai_n732_), .B(mai_mai_n388_), .C(mai_mai_n601_), .Y(mai_mai_n733_));
  OAI210     m0711(.A0(mai_mai_n733_), .A1(mai_mai_n374_), .B0(mai_mai_n372_), .Y(mai_mai_n734_));
  NO2        m0712(.A(mai_mai_n131_), .B(i_2_), .Y(mai_mai_n735_));
  NA2        m0713(.A(mai_mai_n735_), .B(mai_mai_n631_), .Y(mai_mai_n736_));
  NA3        m0714(.A(mai_mai_n736_), .B(mai_mai_n734_), .C(mai_mai_n731_), .Y(mai_mai_n737_));
  NA3        m0715(.A(mai_mai_n737_), .B(mai_mai_n46_), .C(mai_mai_n226_), .Y(mai_mai_n738_));
  NA4        m0716(.A(mai_mai_n738_), .B(mai_mai_n729_), .C(mai_mai_n718_), .D(mai_mai_n701_), .Y(mai_mai_n739_));
  OR4        m0717(.A(mai_mai_n739_), .B(mai_mai_n691_), .C(mai_mai_n681_), .D(mai_mai_n620_), .Y(mai5));
  NA2        m0718(.A(mai_mai_n660_), .B(mai_mai_n271_), .Y(mai_mai_n741_));
  AN2        m0719(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n742_));
  NA3        m0720(.A(mai_mai_n742_), .B(mai_mai_n730_), .C(mai_mai_n111_), .Y(mai_mai_n743_));
  NO2        m0721(.A(mai_mai_n602_), .B(i_11_), .Y(mai_mai_n744_));
  NA2        m0722(.A(mai_mai_n90_), .B(mai_mai_n744_), .Y(mai_mai_n745_));
  NA3        m0723(.A(mai_mai_n745_), .B(mai_mai_n743_), .C(mai_mai_n741_), .Y(mai_mai_n746_));
  NO3        m0724(.A(i_11_), .B(mai_mai_n235_), .C(i_13_), .Y(mai_mai_n747_));
  NO2        m0725(.A(mai_mai_n127_), .B(mai_mai_n23_), .Y(mai_mai_n748_));
  NA2        m0726(.A(i_12_), .B(i_8_), .Y(mai_mai_n749_));
  OAI210     m0727(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n749_), .Y(mai_mai_n750_));
  INV        m0728(.A(mai_mai_n449_), .Y(mai_mai_n751_));
  AOI220     m0729(.A0(mai_mai_n317_), .A1(mai_mai_n575_), .B0(mai_mai_n750_), .B1(mai_mai_n748_), .Y(mai_mai_n752_));
  INV        m0730(.A(mai_mai_n752_), .Y(mai_mai_n753_));
  NO2        m0731(.A(mai_mai_n753_), .B(mai_mai_n746_), .Y(mai_mai_n754_));
  INV        m0732(.A(mai_mai_n175_), .Y(mai_mai_n755_));
  INV        m0733(.A(mai_mai_n244_), .Y(mai_mai_n756_));
  OAI210     m0734(.A0(mai_mai_n687_), .A1(mai_mai_n451_), .B0(mai_mai_n114_), .Y(mai_mai_n757_));
  AOI210     m0735(.A0(mai_mai_n757_), .A1(mai_mai_n756_), .B0(mai_mai_n755_), .Y(mai_mai_n758_));
  NO2        m0736(.A(mai_mai_n459_), .B(mai_mai_n26_), .Y(mai_mai_n759_));
  NO2        m0737(.A(mai_mai_n759_), .B(mai_mai_n419_), .Y(mai_mai_n760_));
  NA2        m0738(.A(mai_mai_n760_), .B(i_2_), .Y(mai_mai_n761_));
  INV        m0739(.A(mai_mai_n761_), .Y(mai_mai_n762_));
  AOI210     m0740(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n416_), .Y(mai_mai_n763_));
  AOI210     m0741(.A0(mai_mai_n763_), .A1(mai_mai_n762_), .B0(mai_mai_n758_), .Y(mai_mai_n764_));
  NO2        m0742(.A(mai_mai_n195_), .B(mai_mai_n128_), .Y(mai_mai_n765_));
  OAI210     m0743(.A0(mai_mai_n765_), .A1(mai_mai_n748_), .B0(i_2_), .Y(mai_mai_n766_));
  INV        m0744(.A(mai_mai_n176_), .Y(mai_mai_n767_));
  NO3        m0745(.A(mai_mai_n622_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n768_));
  AOI210     m0746(.A0(mai_mai_n767_), .A1(mai_mai_n90_), .B0(mai_mai_n768_), .Y(mai_mai_n769_));
  AOI210     m0747(.A0(mai_mai_n769_), .A1(mai_mai_n766_), .B0(mai_mai_n198_), .Y(mai_mai_n770_));
  OA210      m0748(.A0(mai_mai_n623_), .A1(mai_mai_n129_), .B0(i_13_), .Y(mai_mai_n771_));
  NA2        m0749(.A(mai_mai_n205_), .B(mai_mai_n208_), .Y(mai_mai_n772_));
  NA2        m0750(.A(mai_mai_n154_), .B(mai_mai_n597_), .Y(mai_mai_n773_));
  AOI210     m0751(.A0(mai_mai_n773_), .A1(mai_mai_n772_), .B0(mai_mai_n377_), .Y(mai_mai_n774_));
  AOI210     m0752(.A0(mai_mai_n213_), .A1(mai_mai_n151_), .B0(mai_mai_n523_), .Y(mai_mai_n775_));
  NA2        m0753(.A(mai_mai_n775_), .B(mai_mai_n419_), .Y(mai_mai_n776_));
  NO2        m0754(.A(mai_mai_n105_), .B(mai_mai_n45_), .Y(mai_mai_n777_));
  INV        m0755(.A(mai_mai_n299_), .Y(mai_mai_n778_));
  NA4        m0756(.A(mai_mai_n778_), .B(mai_mai_n304_), .C(mai_mai_n127_), .D(mai_mai_n43_), .Y(mai_mai_n779_));
  OAI210     m0757(.A0(mai_mai_n779_), .A1(mai_mai_n777_), .B0(mai_mai_n776_), .Y(mai_mai_n780_));
  NO4        m0758(.A(mai_mai_n780_), .B(mai_mai_n774_), .C(mai_mai_n771_), .D(mai_mai_n770_), .Y(mai_mai_n781_));
  NA2        m0759(.A(mai_mai_n575_), .B(mai_mai_n28_), .Y(mai_mai_n782_));
  NA2        m0760(.A(mai_mai_n747_), .B(mai_mai_n275_), .Y(mai_mai_n783_));
  NA2        m0761(.A(mai_mai_n783_), .B(mai_mai_n782_), .Y(mai_mai_n784_));
  NO2        m0762(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n785_));
  NO2        m0763(.A(mai_mai_n785_), .B(mai_mai_n129_), .Y(mai_mai_n786_));
  NO2        m0764(.A(mai_mai_n786_), .B(mai_mai_n597_), .Y(mai_mai_n787_));
  AOI220     m0765(.A0(mai_mai_n787_), .A1(mai_mai_n36_), .B0(mai_mai_n784_), .B1(mai_mai_n47_), .Y(mai_mai_n788_));
  NA4        m0766(.A(mai_mai_n788_), .B(mai_mai_n781_), .C(mai_mai_n764_), .D(mai_mai_n754_), .Y(mai6));
  NO3        m0767(.A(mai_mai_n255_), .B(mai_mai_n306_), .C(i_1_), .Y(mai_mai_n790_));
  NO2        m0768(.A(mai_mai_n190_), .B(mai_mai_n142_), .Y(mai_mai_n791_));
  OAI210     m0769(.A0(mai_mai_n791_), .A1(mai_mai_n790_), .B0(mai_mai_n735_), .Y(mai_mai_n792_));
  NA4        m0770(.A(mai_mai_n392_), .B(mai_mai_n485_), .C(mai_mai_n72_), .D(mai_mai_n104_), .Y(mai_mai_n793_));
  INV        m0771(.A(mai_mai_n793_), .Y(mai_mai_n794_));
  NO2        m0772(.A(mai_mai_n224_), .B(mai_mai_n490_), .Y(mai_mai_n795_));
  NO2        m0773(.A(i_11_), .B(i_9_), .Y(mai_mai_n796_));
  NO2        m0774(.A(mai_mai_n794_), .B(mai_mai_n329_), .Y(mai_mai_n797_));
  AO210      m0775(.A0(mai_mai_n797_), .A1(mai_mai_n792_), .B0(i_12_), .Y(mai_mai_n798_));
  NA2        m0776(.A(mai_mai_n378_), .B(mai_mai_n334_), .Y(mai_mai_n799_));
  NA2        m0777(.A(mai_mai_n582_), .B(mai_mai_n64_), .Y(mai_mai_n800_));
  BUFFER     m0778(.A(mai_mai_n627_), .Y(mai_mai_n801_));
  NA3        m0779(.A(mai_mai_n801_), .B(mai_mai_n800_), .C(mai_mai_n799_), .Y(mai_mai_n802_));
  INV        m0780(.A(mai_mai_n202_), .Y(mai_mai_n803_));
  AOI220     m0781(.A0(mai_mai_n803_), .A1(mai_mai_n796_), .B0(mai_mai_n802_), .B1(mai_mai_n74_), .Y(mai_mai_n804_));
  INV        m0782(.A(mai_mai_n328_), .Y(mai_mai_n805_));
  NA2        m0783(.A(mai_mai_n76_), .B(mai_mai_n134_), .Y(mai_mai_n806_));
  INV        m0784(.A(mai_mai_n127_), .Y(mai_mai_n807_));
  NA2        m0785(.A(mai_mai_n807_), .B(mai_mai_n47_), .Y(mai_mai_n808_));
  AOI210     m0786(.A0(mai_mai_n808_), .A1(mai_mai_n806_), .B0(mai_mai_n805_), .Y(mai_mai_n809_));
  NO2        m0787(.A(mai_mai_n251_), .B(i_9_), .Y(mai_mai_n810_));
  NA2        m0788(.A(mai_mai_n810_), .B(mai_mai_n785_), .Y(mai_mai_n811_));
  AOI210     m0789(.A0(mai_mai_n811_), .A1(mai_mai_n521_), .B0(mai_mai_n190_), .Y(mai_mai_n812_));
  NO2        m0790(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n813_));
  NAi32      m0791(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n814_));
  NO2        m0792(.A(mai_mai_n719_), .B(mai_mai_n814_), .Y(mai_mai_n815_));
  OR3        m0793(.A(mai_mai_n815_), .B(mai_mai_n812_), .C(mai_mai_n809_), .Y(mai_mai_n816_));
  NO2        m0794(.A(mai_mai_n692_), .B(i_2_), .Y(mai_mai_n817_));
  NA2        m0795(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n818_));
  NO2        m0796(.A(mai_mai_n818_), .B(mai_mai_n408_), .Y(mai_mai_n819_));
  NA2        m0797(.A(mai_mai_n819_), .B(mai_mai_n817_), .Y(mai_mai_n820_));
  AO220      m0798(.A0(mai_mai_n361_), .A1(mai_mai_n351_), .B0(mai_mai_n398_), .B1(mai_mai_n597_), .Y(mai_mai_n821_));
  NA3        m0799(.A(mai_mai_n821_), .B(mai_mai_n256_), .C(i_7_), .Y(mai_mai_n822_));
  OR2        m0800(.A(mai_mai_n623_), .B(mai_mai_n451_), .Y(mai_mai_n823_));
  NA3        m0801(.A(mai_mai_n823_), .B(mai_mai_n150_), .C(mai_mai_n70_), .Y(mai_mai_n824_));
  OR2        m0802(.A(mai_mai_n751_), .B(mai_mai_n36_), .Y(mai_mai_n825_));
  NA4        m0803(.A(mai_mai_n825_), .B(mai_mai_n824_), .C(mai_mai_n822_), .D(mai_mai_n820_), .Y(mai_mai_n826_));
  OAI210     m0804(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n88_), .Y(mai_mai_n827_));
  AOI220     m0805(.A0(mai_mai_n827_), .A1(mai_mai_n564_), .B0(mai_mai_n795_), .B1(mai_mai_n713_), .Y(mai_mai_n828_));
  NA2        m0806(.A(mai_mai_n398_), .B(mai_mai_n71_), .Y(mai_mai_n829_));
  NA3        m0807(.A(mai_mai_n829_), .B(mai_mai_n828_), .C(mai_mai_n605_), .Y(mai_mai_n830_));
  AO210      m0808(.A0(mai_mai_n523_), .A1(mai_mai_n47_), .B0(mai_mai_n89_), .Y(mai_mai_n831_));
  NA3        m0809(.A(mai_mai_n831_), .B(mai_mai_n486_), .C(mai_mai_n223_), .Y(mai_mai_n832_));
  AOI210     m0810(.A0(mai_mai_n451_), .A1(mai_mai_n449_), .B0(mai_mai_n563_), .Y(mai_mai_n833_));
  NO2        m0811(.A(mai_mai_n613_), .B(mai_mai_n105_), .Y(mai_mai_n834_));
  OAI210     m0812(.A0(mai_mai_n834_), .A1(mai_mai_n115_), .B0(mai_mai_n406_), .Y(mai_mai_n835_));
  INV        m0813(.A(mai_mai_n586_), .Y(mai_mai_n836_));
  NA3        m0814(.A(mai_mai_n836_), .B(mai_mai_n328_), .C(i_7_), .Y(mai_mai_n837_));
  NA4        m0815(.A(mai_mai_n837_), .B(mai_mai_n835_), .C(mai_mai_n833_), .D(mai_mai_n832_), .Y(mai_mai_n838_));
  NO4        m0816(.A(mai_mai_n838_), .B(mai_mai_n830_), .C(mai_mai_n826_), .D(mai_mai_n816_), .Y(mai_mai_n839_));
  NA4        m0817(.A(mai_mai_n839_), .B(mai_mai_n804_), .C(mai_mai_n798_), .D(mai_mai_n384_), .Y(mai3));
  NA2        m0818(.A(i_6_), .B(i_7_), .Y(mai_mai_n841_));
  NO2        m0819(.A(mai_mai_n841_), .B(i_0_), .Y(mai_mai_n842_));
  NO2        m0820(.A(i_11_), .B(mai_mai_n235_), .Y(mai_mai_n843_));
  OAI210     m0821(.A0(mai_mai_n842_), .A1(mai_mai_n290_), .B0(mai_mai_n843_), .Y(mai_mai_n844_));
  NO2        m0822(.A(mai_mai_n844_), .B(mai_mai_n198_), .Y(mai_mai_n845_));
  NO3        m0823(.A(mai_mai_n455_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n846_));
  OA210      m0824(.A0(mai_mai_n846_), .A1(mai_mai_n845_), .B0(mai_mai_n178_), .Y(mai_mai_n847_));
  NOi21      m0825(.An(mai_mai_n99_), .B(mai_mai_n760_), .Y(mai_mai_n848_));
  NA2        m0826(.A(mai_mai_n409_), .B(mai_mai_n46_), .Y(mai_mai_n849_));
  AN2        m0827(.A(mai_mai_n457_), .B(mai_mai_n56_), .Y(mai_mai_n850_));
  NO2        m0828(.A(mai_mai_n850_), .B(mai_mai_n848_), .Y(mai_mai_n851_));
  NO2        m0829(.A(mai_mai_n851_), .B(mai_mai_n49_), .Y(mai_mai_n852_));
  NO4        m0830(.A(mai_mai_n380_), .B(mai_mai_n387_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n853_));
  NA2        m0831(.A(mai_mai_n190_), .B(mai_mai_n573_), .Y(mai_mai_n854_));
  NOi21      m0832(.An(mai_mai_n854_), .B(mai_mai_n853_), .Y(mai_mai_n855_));
  NA2        m0833(.A(mai_mai_n705_), .B(mai_mai_n672_), .Y(mai_mai_n856_));
  NA2        m0834(.A(mai_mai_n332_), .B(mai_mai_n439_), .Y(mai_mai_n857_));
  OAI220     m0835(.A0(mai_mai_n857_), .A1(mai_mai_n856_), .B0(mai_mai_n855_), .B1(mai_mai_n64_), .Y(mai_mai_n858_));
  NOi21      m0836(.An(i_5_), .B(i_9_), .Y(mai_mai_n859_));
  NA2        m0837(.A(mai_mai_n859_), .B(mai_mai_n447_), .Y(mai_mai_n860_));
  BUFFER     m0838(.A(mai_mai_n269_), .Y(mai_mai_n861_));
  NA2        m0839(.A(mai_mai_n861_), .B(mai_mai_n477_), .Y(mai_mai_n862_));
  NO3        m0840(.A(mai_mai_n412_), .B(mai_mai_n269_), .C(mai_mai_n74_), .Y(mai_mai_n863_));
  NO2        m0841(.A(mai_mai_n179_), .B(mai_mai_n151_), .Y(mai_mai_n864_));
  AOI210     m0842(.A0(mai_mai_n864_), .A1(mai_mai_n243_), .B0(mai_mai_n863_), .Y(mai_mai_n865_));
  OAI220     m0843(.A0(mai_mai_n865_), .A1(mai_mai_n185_), .B0(mai_mai_n862_), .B1(mai_mai_n860_), .Y(mai_mai_n866_));
  NO4        m0844(.A(mai_mai_n866_), .B(mai_mai_n858_), .C(mai_mai_n852_), .D(mai_mai_n847_), .Y(mai_mai_n867_));
  NA2        m0845(.A(mai_mai_n190_), .B(mai_mai_n24_), .Y(mai_mai_n868_));
  NO2        m0846(.A(mai_mai_n670_), .B(mai_mai_n594_), .Y(mai_mai_n869_));
  NO2        m0847(.A(mai_mai_n869_), .B(mai_mai_n868_), .Y(mai_mai_n870_));
  INV        m0848(.A(mai_mai_n870_), .Y(mai_mai_n871_));
  NO2        m0849(.A(mai_mai_n392_), .B(mai_mai_n291_), .Y(mai_mai_n872_));
  NA2        m0850(.A(mai_mai_n872_), .B(mai_mai_n708_), .Y(mai_mai_n873_));
  NA2        m0851(.A(mai_mai_n574_), .B(i_0_), .Y(mai_mai_n874_));
  NO4        m0852(.A(mai_mai_n585_), .B(mai_mai_n221_), .C(mai_mai_n416_), .D(mai_mai_n408_), .Y(mai_mai_n875_));
  NA2        m0853(.A(mai_mai_n875_), .B(i_11_), .Y(mai_mai_n876_));
  AN2        m0854(.A(mai_mai_n99_), .B(mai_mai_n242_), .Y(mai_mai_n877_));
  NA2        m0855(.A(mai_mai_n747_), .B(mai_mai_n329_), .Y(mai_mai_n878_));
  AOI210     m0856(.A0(mai_mai_n486_), .A1(mai_mai_n90_), .B0(mai_mai_n59_), .Y(mai_mai_n879_));
  OAI220     m0857(.A0(mai_mai_n879_), .A1(mai_mai_n878_), .B0(mai_mai_n656_), .B1(mai_mai_n542_), .Y(mai_mai_n880_));
  NO2        m0858(.A(mai_mai_n253_), .B(mai_mai_n156_), .Y(mai_mai_n881_));
  NA2        m0859(.A(i_0_), .B(i_10_), .Y(mai_mai_n882_));
  INV        m0860(.A(mai_mai_n545_), .Y(mai_mai_n883_));
  NO4        m0861(.A(mai_mai_n118_), .B(mai_mai_n59_), .C(mai_mai_n665_), .D(i_5_), .Y(mai_mai_n884_));
  AO220      m0862(.A0(mai_mai_n884_), .A1(mai_mai_n883_), .B0(mai_mai_n881_), .B1(i_6_), .Y(mai_mai_n885_));
  AOI220     m0863(.A0(mai_mai_n332_), .A1(mai_mai_n101_), .B0(mai_mai_n190_), .B1(mai_mai_n85_), .Y(mai_mai_n886_));
  NA2        m0864(.A(mai_mai_n568_), .B(i_4_), .Y(mai_mai_n887_));
  NA2        m0865(.A(mai_mai_n193_), .B(mai_mai_n208_), .Y(mai_mai_n888_));
  OAI220     m0866(.A0(mai_mai_n888_), .A1(mai_mai_n878_), .B0(mai_mai_n887_), .B1(mai_mai_n886_), .Y(mai_mai_n889_));
  NO4        m0867(.A(mai_mai_n889_), .B(mai_mai_n885_), .C(mai_mai_n880_), .D(mai_mai_n877_), .Y(mai_mai_n890_));
  NA4        m0868(.A(mai_mai_n890_), .B(mai_mai_n876_), .C(mai_mai_n873_), .D(mai_mai_n871_), .Y(mai_mai_n891_));
  NA2        m0869(.A(i_11_), .B(i_9_), .Y(mai_mai_n892_));
  NO2        m0870(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n893_));
  NA2        m0871(.A(mai_mai_n397_), .B(mai_mai_n183_), .Y(mai_mai_n894_));
  NA2        m0872(.A(mai_mai_n894_), .B(mai_mai_n163_), .Y(mai_mai_n895_));
  NO2        m0873(.A(mai_mai_n892_), .B(mai_mai_n74_), .Y(mai_mai_n896_));
  NO2        m0874(.A(mai_mai_n179_), .B(i_0_), .Y(mai_mai_n897_));
  INV        m0875(.A(mai_mai_n897_), .Y(mai_mai_n898_));
  NA2        m0876(.A(mai_mai_n475_), .B(mai_mai_n229_), .Y(mai_mai_n899_));
  NA2        m0877(.A(mai_mai_n375_), .B(mai_mai_n42_), .Y(mai_mai_n900_));
  OAI220     m0878(.A0(mai_mai_n900_), .A1(mai_mai_n860_), .B0(mai_mai_n899_), .B1(mai_mai_n898_), .Y(mai_mai_n901_));
  NO2        m0879(.A(mai_mai_n901_), .B(mai_mai_n895_), .Y(mai_mai_n902_));
  NA2        m0880(.A(mai_mai_n655_), .B(mai_mai_n124_), .Y(mai_mai_n903_));
  NO2        m0881(.A(i_6_), .B(mai_mai_n903_), .Y(mai_mai_n904_));
  AOI210     m0882(.A0(mai_mai_n450_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n905_));
  NA2        m0883(.A(mai_mai_n175_), .B(mai_mai_n106_), .Y(mai_mai_n906_));
  NOi32      m0884(.An(mai_mai_n905_), .Bn(mai_mai_n193_), .C(mai_mai_n906_), .Y(mai_mai_n907_));
  NA2        m0885(.A(mai_mai_n606_), .B(mai_mai_n329_), .Y(mai_mai_n908_));
  NO2        m0886(.A(mai_mai_n908_), .B(mai_mai_n849_), .Y(mai_mai_n909_));
  NO3        m0887(.A(mai_mai_n909_), .B(mai_mai_n907_), .C(mai_mai_n904_), .Y(mai_mai_n910_));
  NOi21      m0888(.An(i_7_), .B(i_5_), .Y(mai_mai_n911_));
  OR2        m0889(.A(mai_mai_n906_), .B(mai_mai_n521_), .Y(mai_mai_n912_));
  NO3        m0890(.A(mai_mai_n402_), .B(mai_mai_n364_), .C(mai_mai_n360_), .Y(mai_mai_n913_));
  NO2        m0891(.A(mai_mai_n263_), .B(mai_mai_n318_), .Y(mai_mai_n914_));
  NO2        m0892(.A(mai_mai_n724_), .B(mai_mai_n258_), .Y(mai_mai_n915_));
  AOI210     m0893(.A0(mai_mai_n915_), .A1(mai_mai_n914_), .B0(mai_mai_n913_), .Y(mai_mai_n916_));
  NA4        m0894(.A(mai_mai_n916_), .B(mai_mai_n912_), .C(mai_mai_n910_), .D(mai_mai_n902_), .Y(mai_mai_n917_));
  NO2        m0895(.A(mai_mai_n868_), .B(mai_mai_n238_), .Y(mai_mai_n918_));
  AN2        m0896(.A(mai_mai_n331_), .B(mai_mai_n329_), .Y(mai_mai_n919_));
  AN2        m0897(.A(mai_mai_n919_), .B(mai_mai_n864_), .Y(mai_mai_n920_));
  OAI210     m0898(.A0(mai_mai_n920_), .A1(mai_mai_n918_), .B0(i_10_), .Y(mai_mai_n921_));
  OA210      m0899(.A0(mai_mai_n475_), .A1(mai_mai_n225_), .B0(mai_mai_n474_), .Y(mai_mai_n922_));
  NA2        m0900(.A(mai_mai_n896_), .B(mai_mai_n304_), .Y(mai_mai_n923_));
  OAI210     m0901(.A0(i_2_), .A1(mai_mai_n192_), .B0(mai_mai_n923_), .Y(mai_mai_n924_));
  NA2        m0902(.A(mai_mai_n924_), .B(mai_mai_n475_), .Y(mai_mai_n925_));
  NO3        m0903(.A(mai_mai_n585_), .B(mai_mai_n359_), .C(mai_mai_n24_), .Y(mai_mai_n926_));
  INV        m0904(.A(mai_mai_n926_), .Y(mai_mai_n927_));
  NAi21      m0905(.An(i_9_), .B(i_5_), .Y(mai_mai_n928_));
  NO2        m0906(.A(mai_mai_n928_), .B(mai_mai_n402_), .Y(mai_mai_n929_));
  NO2        m0907(.A(mai_mai_n600_), .B(mai_mai_n108_), .Y(mai_mai_n930_));
  AOI220     m0908(.A0(mai_mai_n930_), .A1(i_0_), .B0(mai_mai_n929_), .B1(mai_mai_n623_), .Y(mai_mai_n931_));
  OAI220     m0909(.A0(mai_mai_n931_), .A1(mai_mai_n87_), .B0(mai_mai_n927_), .B1(mai_mai_n176_), .Y(mai_mai_n932_));
  NO2        m0910(.A(mai_mai_n932_), .B(mai_mai_n526_), .Y(mai_mai_n933_));
  NA3        m0911(.A(mai_mai_n933_), .B(mai_mai_n925_), .C(mai_mai_n921_), .Y(mai_mai_n934_));
  NO3        m0912(.A(mai_mai_n934_), .B(mai_mai_n917_), .C(mai_mai_n891_), .Y(mai_mai_n935_));
  NO2        m0913(.A(i_0_), .B(mai_mai_n724_), .Y(mai_mai_n936_));
  NA2        m0914(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n937_));
  INV        m0915(.A(mai_mai_n937_), .Y(mai_mai_n938_));
  NO3        m0916(.A(mai_mai_n108_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n939_));
  AO220      m0917(.A0(mai_mai_n939_), .A1(mai_mai_n938_), .B0(mai_mai_n936_), .B1(mai_mai_n178_), .Y(mai_mai_n940_));
  AOI210     m0918(.A0(mai_mai_n800_), .A1(mai_mai_n683_), .B0(mai_mai_n906_), .Y(mai_mai_n941_));
  AOI210     m0919(.A0(mai_mai_n940_), .A1(mai_mai_n348_), .B0(mai_mai_n941_), .Y(mai_mai_n942_));
  NA2        m0920(.A(mai_mai_n735_), .B(mai_mai_n149_), .Y(mai_mai_n943_));
  INV        m0921(.A(mai_mai_n943_), .Y(mai_mai_n944_));
  NA3        m0922(.A(mai_mai_n944_), .B(mai_mai_n672_), .C(mai_mai_n74_), .Y(mai_mai_n945_));
  NA3        m0923(.A(mai_mai_n842_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n946_));
  NA2        m0924(.A(mai_mai_n843_), .B(i_9_), .Y(mai_mai_n947_));
  AOI210     m0925(.A0(mai_mai_n946_), .A1(mai_mai_n500_), .B0(mai_mai_n947_), .Y(mai_mai_n948_));
  OAI210     m0926(.A0(mai_mai_n243_), .A1(i_9_), .B0(mai_mai_n228_), .Y(mai_mai_n949_));
  AOI210     m0927(.A0(mai_mai_n949_), .A1(mai_mai_n874_), .B0(mai_mai_n156_), .Y(mai_mai_n950_));
  NO2        m0928(.A(mai_mai_n950_), .B(mai_mai_n948_), .Y(mai_mai_n951_));
  NA3        m0929(.A(mai_mai_n951_), .B(mai_mai_n945_), .C(mai_mai_n942_), .Y(mai_mai_n952_));
  NA2        m0930(.A(mai_mai_n919_), .B(mai_mai_n377_), .Y(mai_mai_n953_));
  AOI210     m0931(.A0(mai_mai_n298_), .A1(mai_mai_n165_), .B0(mai_mai_n953_), .Y(mai_mai_n954_));
  NA3        m0932(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n955_));
  NA2        m0933(.A(mai_mai_n893_), .B(mai_mai_n491_), .Y(mai_mai_n956_));
  AOI210     m0934(.A0(mai_mai_n955_), .A1(mai_mai_n165_), .B0(mai_mai_n956_), .Y(mai_mai_n957_));
  NO2        m0935(.A(mai_mai_n957_), .B(mai_mai_n954_), .Y(mai_mai_n958_));
  NO3        m0936(.A(mai_mai_n882_), .B(mai_mai_n859_), .C(mai_mai_n195_), .Y(mai_mai_n959_));
  AOI220     m0937(.A0(mai_mai_n959_), .A1(i_11_), .B0(mai_mai_n569_), .B1(mai_mai_n76_), .Y(mai_mai_n960_));
  NO3        m0938(.A(mai_mai_n215_), .B(mai_mai_n387_), .C(i_0_), .Y(mai_mai_n961_));
  OAI210     m0939(.A0(mai_mai_n961_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n962_));
  INV        m0940(.A(mai_mai_n223_), .Y(mai_mai_n963_));
  OAI220     m0941(.A0(mai_mai_n536_), .A1(mai_mai_n142_), .B0(mai_mai_n642_), .B1(mai_mai_n617_), .Y(mai_mai_n964_));
  NA3        m0942(.A(mai_mai_n964_), .B(mai_mai_n1034_), .C(mai_mai_n963_), .Y(mai_mai_n965_));
  NA4        m0943(.A(mai_mai_n965_), .B(mai_mai_n962_), .C(mai_mai_n960_), .D(mai_mai_n958_), .Y(mai_mai_n966_));
  INV        m0944(.A(mai_mai_n112_), .Y(mai_mai_n967_));
  AOI220     m0945(.A0(mai_mai_n911_), .A1(mai_mai_n491_), .B0(mai_mai_n842_), .B1(mai_mai_n166_), .Y(mai_mai_n968_));
  NA2        m0946(.A(mai_mai_n351_), .B(mai_mai_n180_), .Y(mai_mai_n969_));
  OA220      m0947(.A0(mai_mai_n969_), .A1(mai_mai_n968_), .B0(mai_mai_n967_), .B1(i_5_), .Y(mai_mai_n970_));
  AOI210     m0948(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n179_), .Y(mai_mai_n971_));
  NA2        m0949(.A(mai_mai_n971_), .B(mai_mai_n922_), .Y(mai_mai_n972_));
  NA3        m0950(.A(mai_mai_n614_), .B(mai_mai_n190_), .C(mai_mai_n85_), .Y(mai_mai_n973_));
  INV        m0951(.A(mai_mai_n973_), .Y(mai_mai_n974_));
  NO3        m0952(.A(mai_mai_n849_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n975_));
  NA2        m0953(.A(mai_mai_n496_), .B(mai_mai_n489_), .Y(mai_mai_n976_));
  NO3        m0954(.A(mai_mai_n976_), .B(mai_mai_n975_), .C(mai_mai_n974_), .Y(mai_mai_n977_));
  NA3        m0955(.A(mai_mai_n893_), .B(mai_mai_n290_), .C(mai_mai_n228_), .Y(mai_mai_n978_));
  INV        m0956(.A(mai_mai_n978_), .Y(mai_mai_n979_));
  NOi31      m0957(.An(mai_mai_n391_), .B(mai_mai_n937_), .C(mai_mai_n238_), .Y(mai_mai_n980_));
  NO3        m0958(.A(mai_mai_n892_), .B(mai_mai_n223_), .C(mai_mai_n195_), .Y(mai_mai_n981_));
  NO3        m0959(.A(mai_mai_n981_), .B(mai_mai_n980_), .C(mai_mai_n979_), .Y(mai_mai_n982_));
  NA4        m0960(.A(mai_mai_n982_), .B(mai_mai_n977_), .C(mai_mai_n972_), .D(mai_mai_n970_), .Y(mai_mai_n983_));
  INV        m0961(.A(mai_mai_n616_), .Y(mai_mai_n984_));
  NO3        m0962(.A(mai_mai_n984_), .B(mai_mai_n559_), .C(mai_mai_n345_), .Y(mai_mai_n985_));
  INV        m0963(.A(mai_mai_n985_), .Y(mai_mai_n986_));
  NA2        m0964(.A(mai_mai_n794_), .B(mai_mai_n180_), .Y(mai_mai_n987_));
  NA3        m0965(.A(mai_mai_n101_), .B(mai_mai_n573_), .C(i_11_), .Y(mai_mai_n988_));
  NO2        m0966(.A(mai_mai_n988_), .B(mai_mai_n158_), .Y(mai_mai_n989_));
  INV        m0967(.A(mai_mai_n989_), .Y(mai_mai_n990_));
  NA3        m0968(.A(mai_mai_n990_), .B(mai_mai_n987_), .C(mai_mai_n986_), .Y(mai_mai_n991_));
  NO4        m0969(.A(mai_mai_n991_), .B(mai_mai_n983_), .C(mai_mai_n966_), .D(mai_mai_n952_), .Y(mai_mai_n992_));
  OAI210     m0970(.A0(mai_mai_n817_), .A1(mai_mai_n813_), .B0(mai_mai_n37_), .Y(mai_mai_n993_));
  NA3        m0971(.A(mai_mai_n905_), .B(mai_mai_n372_), .C(i_5_), .Y(mai_mai_n994_));
  NA3        m0972(.A(mai_mai_n994_), .B(mai_mai_n993_), .C(mai_mai_n612_), .Y(mai_mai_n995_));
  NA2        m0973(.A(mai_mai_n995_), .B(mai_mai_n211_), .Y(mai_mai_n996_));
  AN2        m0974(.A(mai_mai_n692_), .B(mai_mai_n373_), .Y(mai_mai_n997_));
  NA2        m0975(.A(mai_mai_n191_), .B(mai_mai_n193_), .Y(mai_mai_n998_));
  AO210      m0976(.A0(mai_mai_n997_), .A1(mai_mai_n33_), .B0(mai_mai_n998_), .Y(mai_mai_n999_));
  OAI210     m0977(.A0(mai_mai_n616_), .A1(mai_mai_n614_), .B0(mai_mai_n317_), .Y(mai_mai_n1000_));
  NAi31      m0978(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n1001_));
  NO2        m0979(.A(mai_mai_n71_), .B(mai_mai_n1001_), .Y(mai_mai_n1002_));
  INV        m0980(.A(mai_mai_n1002_), .Y(mai_mai_n1003_));
  NA3        m0981(.A(mai_mai_n1003_), .B(mai_mai_n1000_), .C(mai_mai_n999_), .Y(mai_mai_n1004_));
  NO2        m0982(.A(mai_mai_n464_), .B(mai_mai_n269_), .Y(mai_mai_n1005_));
  NO4        m0983(.A(mai_mai_n231_), .B(mai_mai_n148_), .C(mai_mai_n676_), .D(mai_mai_n37_), .Y(mai_mai_n1006_));
  NO3        m0984(.A(mai_mai_n1006_), .B(mai_mai_n1005_), .C(mai_mai_n875_), .Y(mai_mai_n1007_));
  OAI210     m0985(.A0(mai_mai_n988_), .A1(mai_mai_n151_), .B0(mai_mai_n1007_), .Y(mai_mai_n1008_));
  AOI210     m0986(.A0(mai_mai_n1004_), .A1(mai_mai_n49_), .B0(mai_mai_n1008_), .Y(mai_mai_n1009_));
  AOI210     m0987(.A0(mai_mai_n1009_), .A1(mai_mai_n996_), .B0(mai_mai_n74_), .Y(mai_mai_n1010_));
  NO2        m0988(.A(mai_mai_n566_), .B(mai_mai_n383_), .Y(mai_mai_n1011_));
  NO2        m0989(.A(mai_mai_n1011_), .B(mai_mai_n755_), .Y(mai_mai_n1012_));
  NA2        m0990(.A(mai_mai_n263_), .B(mai_mai_n58_), .Y(mai_mai_n1013_));
  AOI220     m0991(.A0(mai_mai_n1013_), .A1(mai_mai_n77_), .B0(mai_mai_n346_), .B1(mai_mai_n255_), .Y(mai_mai_n1014_));
  NO2        m0992(.A(mai_mai_n1014_), .B(mai_mai_n235_), .Y(mai_mai_n1015_));
  NA3        m0993(.A(mai_mai_n99_), .B(mai_mai_n306_), .C(mai_mai_n31_), .Y(mai_mai_n1016_));
  INV        m0994(.A(mai_mai_n1016_), .Y(mai_mai_n1017_));
  NO2        m0995(.A(mai_mai_n1017_), .B(mai_mai_n1015_), .Y(mai_mai_n1018_));
  NA2        m0996(.A(mai_mai_n607_), .B(mai_mai_n221_), .Y(mai_mai_n1019_));
  OAI210     m0997(.A0(mai_mai_n1019_), .A1(mai_mai_n905_), .B0(mai_mai_n211_), .Y(mai_mai_n1020_));
  NA2        m0998(.A(mai_mai_n167_), .B(i_5_), .Y(mai_mai_n1021_));
  NO2        m0999(.A(mai_mai_n1020_), .B(mai_mai_n1021_), .Y(mai_mai_n1022_));
  NO4        m1000(.A(mai_mai_n928_), .B(mai_mai_n479_), .C(mai_mai_n252_), .D(mai_mai_n251_), .Y(mai_mai_n1023_));
  NO2        m1001(.A(mai_mai_n1023_), .B(mai_mai_n563_), .Y(mai_mai_n1024_));
  INV        m1002(.A(mai_mai_n365_), .Y(mai_mai_n1025_));
  AOI210     m1003(.A0(mai_mai_n1025_), .A1(mai_mai_n1024_), .B0(mai_mai_n41_), .Y(mai_mai_n1026_));
  NO2        m1004(.A(mai_mai_n1026_), .B(mai_mai_n1022_), .Y(mai_mai_n1027_));
  OAI210     m1005(.A0(mai_mai_n1018_), .A1(i_4_), .B0(mai_mai_n1027_), .Y(mai_mai_n1028_));
  NO3        m1006(.A(mai_mai_n1028_), .B(mai_mai_n1012_), .C(mai_mai_n1010_), .Y(mai_mai_n1029_));
  NA4        m1007(.A(mai_mai_n1029_), .B(mai_mai_n992_), .C(mai_mai_n935_), .D(mai_mai_n867_), .Y(mai4));
  INV        m1008(.A(mai_mai_n486_), .Y(mai_mai_n1033_));
  INV        m1009(.A(i_3_), .Y(mai_mai_n1034_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  OAI210     u0028(.A0(men_men_n50_), .A1(i_3_), .B0(men_men_n48_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n50_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  NO3        u0062(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n63_), .Y(men_men_n85_));
  INV        u0063(.A(i_6_), .Y(men_men_n86_));
  NO2        u0064(.A(i_2_), .B(i_7_), .Y(men_men_n87_));
  OAI210     u0065(.A0(men_men_n85_), .A1(men_men_n82_), .B0(i_2_), .Y(men_men_n88_));
  NAi21      u0066(.An(i_6_), .B(i_10_), .Y(men_men_n89_));
  NA2        u0067(.A(i_6_), .B(i_9_), .Y(men_men_n90_));
  AOI210     u0068(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n63_), .Y(men_men_n91_));
  NA2        u0069(.A(i_2_), .B(i_6_), .Y(men_men_n92_));
  NO3        u0070(.A(men_men_n92_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n93_));
  NO2        u0071(.A(men_men_n93_), .B(men_men_n91_), .Y(men_men_n94_));
  AOI210     u0072(.A0(men_men_n94_), .A1(men_men_n88_), .B0(men_men_n80_), .Y(men_men_n95_));
  AN3        u0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n96_));
  NAi21      u0074(.An(i_6_), .B(i_11_), .Y(men_men_n97_));
  NO2        u0075(.A(i_5_), .B(i_8_), .Y(men_men_n98_));
  NOi21      u0076(.An(men_men_n98_), .B(men_men_n97_), .Y(men_men_n99_));
  AOI220     u0077(.A0(men_men_n99_), .A1(men_men_n62_), .B0(men_men_n96_), .B1(men_men_n32_), .Y(men_men_n100_));
  INV        u0078(.A(i_7_), .Y(men_men_n101_));
  NA2        u0079(.A(men_men_n46_), .B(men_men_n101_), .Y(men_men_n102_));
  NO2        u0080(.A(i_0_), .B(i_5_), .Y(men_men_n103_));
  NO2        u0081(.A(men_men_n103_), .B(men_men_n86_), .Y(men_men_n104_));
  NA2        u0082(.A(i_12_), .B(i_3_), .Y(men_men_n105_));
  INV        u0083(.A(men_men_n105_), .Y(men_men_n106_));
  NA3        u0084(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n102_), .Y(men_men_n107_));
  NAi21      u0085(.An(i_7_), .B(i_11_), .Y(men_men_n108_));
  AN2        u0086(.A(i_2_), .B(i_10_), .Y(men_men_n109_));
  NO2        u0087(.A(men_men_n109_), .B(i_7_), .Y(men_men_n110_));
  OR2        u0088(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n111_));
  NO2        u0089(.A(i_8_), .B(men_men_n101_), .Y(men_men_n112_));
  NO3        u0090(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n110_), .Y(men_men_n113_));
  NA2        u0091(.A(i_12_), .B(i_7_), .Y(men_men_n114_));
  NO2        u0092(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n115_));
  NA2        u0093(.A(men_men_n115_), .B(i_0_), .Y(men_men_n116_));
  NA2        u0094(.A(i_11_), .B(i_12_), .Y(men_men_n117_));
  OAI210     u0095(.A0(men_men_n116_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n118_), .B(men_men_n113_), .Y(men_men_n119_));
  NA3        u0097(.A(men_men_n119_), .B(men_men_n107_), .C(men_men_n100_), .Y(men_men_n120_));
  NOi21      u0098(.An(i_1_), .B(i_5_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n121_), .B(i_11_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n123_));
  NA2        u0101(.A(i_7_), .B(men_men_n25_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NO2        u0103(.A(men_men_n125_), .B(men_men_n46_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n127_));
  NAi21      u0105(.An(i_3_), .B(i_8_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(men_men_n62_), .Y(men_men_n129_));
  NOi31      u0107(.An(men_men_n129_), .B(men_men_n127_), .C(men_men_n126_), .Y(men_men_n130_));
  NO2        u0108(.A(i_1_), .B(men_men_n86_), .Y(men_men_n131_));
  NO2        u0109(.A(i_6_), .B(i_5_), .Y(men_men_n132_));
  NA2        u0110(.A(men_men_n132_), .B(i_3_), .Y(men_men_n133_));
  AO210      u0111(.A0(men_men_n133_), .A1(men_men_n47_), .B0(men_men_n131_), .Y(men_men_n134_));
  OAI220     u0112(.A0(men_men_n134_), .A1(men_men_n108_), .B0(men_men_n130_), .B1(men_men_n122_), .Y(men_men_n135_));
  NO3        u0113(.A(men_men_n135_), .B(men_men_n120_), .C(men_men_n95_), .Y(men_men_n136_));
  NA3        u0114(.A(men_men_n136_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0115(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n138_));
  NA2        u0116(.A(i_6_), .B(men_men_n25_), .Y(men_men_n139_));
  NA2        u0117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NA4        u0118(.A(men_men_n140_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0119(.A(i_8_), .B(i_7_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(i_6_), .Y(men_men_n143_));
  NO2        u0121(.A(i_12_), .B(i_13_), .Y(men_men_n144_));
  NAi21      u0122(.An(i_5_), .B(i_11_), .Y(men_men_n145_));
  NOi21      u0123(.An(men_men_n144_), .B(men_men_n145_), .Y(men_men_n146_));
  NO2        u0124(.A(i_0_), .B(i_1_), .Y(men_men_n147_));
  NA2        u0125(.A(i_2_), .B(i_3_), .Y(men_men_n148_));
  NO2        u0126(.A(men_men_n148_), .B(i_4_), .Y(men_men_n149_));
  NA3        u0127(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n150_));
  OR2        u0128(.A(men_men_n150_), .B(men_men_n25_), .Y(men_men_n151_));
  AN2        u0129(.A(men_men_n144_), .B(men_men_n83_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n152_), .B(men_men_n27_), .Y(men_men_n153_));
  NA2        u0131(.A(i_1_), .B(i_5_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n73_), .B(men_men_n46_), .Y(men_men_n155_));
  NA2        u0133(.A(men_men_n155_), .B(men_men_n36_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n156_), .B(men_men_n154_), .C(men_men_n153_), .Y(men_men_n157_));
  OR2        u0135(.A(i_0_), .B(i_1_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n159_));
  NAi32      u0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n160_));
  NAi21      u0138(.An(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0139(.An(i_4_), .B(i_10_), .Y(men_men_n162_));
  NA2        u0140(.A(men_men_n162_), .B(men_men_n40_), .Y(men_men_n163_));
  NO2        u0141(.A(i_3_), .B(i_5_), .Y(men_men_n164_));
  NO3        u0142(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  OAI210     u0144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n167_));
  NO2        u0145(.A(men_men_n167_), .B(men_men_n157_), .Y(men_men_n168_));
  AOI210     u0146(.A0(men_men_n168_), .A1(men_men_n151_), .B0(men_men_n143_), .Y(men_men_n169_));
  NA3        u0147(.A(men_men_n73_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n170_));
  NA2        u0148(.A(i_3_), .B(men_men_n48_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_4_), .B(i_9_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_11_), .B(i_13_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OR2        u0152(.A(men_men_n174_), .B(men_men_n171_), .Y(men_men_n175_));
  NO2        u0153(.A(i_4_), .B(i_5_), .Y(men_men_n176_));
  NAi21      u0154(.An(i_12_), .B(i_11_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n177_), .B(i_13_), .Y(men_men_n178_));
  NA3        u0156(.A(men_men_n178_), .B(men_men_n176_), .C(men_men_n83_), .Y(men_men_n179_));
  AOI210     u0157(.A0(men_men_n179_), .A1(men_men_n175_), .B0(men_men_n170_), .Y(men_men_n180_));
  NO2        u0158(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n181_));
  NA2        u0159(.A(men_men_n181_), .B(men_men_n46_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n36_), .B(i_5_), .Y(men_men_n183_));
  NAi31      u0161(.An(men_men_n183_), .B(men_men_n152_), .C(i_11_), .Y(men_men_n184_));
  NA2        u0162(.A(i_3_), .B(i_5_), .Y(men_men_n185_));
  OR2        u0163(.A(men_men_n185_), .B(men_men_n174_), .Y(men_men_n186_));
  AOI210     u0164(.A0(men_men_n186_), .A1(men_men_n184_), .B0(men_men_n182_), .Y(men_men_n187_));
  NO2        u0165(.A(men_men_n73_), .B(i_5_), .Y(men_men_n188_));
  NO2        u0166(.A(i_13_), .B(i_10_), .Y(men_men_n189_));
  NA3        u0167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n44_), .Y(men_men_n190_));
  NO2        u0168(.A(i_2_), .B(i_1_), .Y(men_men_n191_));
  NA2        u0169(.A(men_men_n191_), .B(i_3_), .Y(men_men_n192_));
  NAi21      u0170(.An(i_4_), .B(i_12_), .Y(men_men_n193_));
  NO4        u0171(.A(men_men_n193_), .B(men_men_n192_), .C(men_men_n190_), .D(men_men_n25_), .Y(men_men_n194_));
  NO3        u0172(.A(men_men_n194_), .B(men_men_n187_), .C(men_men_n180_), .Y(men_men_n195_));
  INV        u0173(.A(i_8_), .Y(men_men_n196_));
  NO2        u0174(.A(men_men_n196_), .B(i_7_), .Y(men_men_n197_));
  NA2        u0175(.A(men_men_n197_), .B(i_6_), .Y(men_men_n198_));
  NO3        u0176(.A(i_3_), .B(men_men_n86_), .C(men_men_n48_), .Y(men_men_n199_));
  NA2        u0177(.A(men_men_n199_), .B(men_men_n112_), .Y(men_men_n200_));
  NO3        u0178(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n201_));
  NA3        u0179(.A(men_men_n201_), .B(men_men_n40_), .C(men_men_n44_), .Y(men_men_n202_));
  NO3        u0180(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n203_));
  OAI210     u0181(.A0(men_men_n96_), .A1(i_12_), .B0(men_men_n203_), .Y(men_men_n204_));
  AOI210     u0182(.A0(men_men_n204_), .A1(men_men_n202_), .B0(men_men_n200_), .Y(men_men_n205_));
  NO2        u0183(.A(i_3_), .B(i_8_), .Y(men_men_n206_));
  NO3        u0184(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n207_));
  NA3        u0185(.A(men_men_n207_), .B(men_men_n206_), .C(men_men_n40_), .Y(men_men_n208_));
  NO2        u0186(.A(men_men_n103_), .B(men_men_n58_), .Y(men_men_n209_));
  INV        u0187(.A(men_men_n209_), .Y(men_men_n210_));
  NO2        u0188(.A(i_13_), .B(i_9_), .Y(men_men_n211_));
  NA3        u0189(.A(men_men_n211_), .B(i_6_), .C(men_men_n196_), .Y(men_men_n212_));
  NAi21      u0190(.An(i_12_), .B(i_3_), .Y(men_men_n213_));
  NO2        u0191(.A(men_men_n44_), .B(i_5_), .Y(men_men_n214_));
  NO3        u0192(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n215_));
  NA3        u0193(.A(men_men_n215_), .B(men_men_n214_), .C(i_10_), .Y(men_men_n216_));
  OAI220     u0194(.A0(men_men_n216_), .A1(men_men_n212_), .B0(men_men_n210_), .B1(men_men_n208_), .Y(men_men_n217_));
  AOI210     u0195(.A0(men_men_n217_), .A1(i_7_), .B0(men_men_n205_), .Y(men_men_n218_));
  OAI220     u0196(.A0(men_men_n218_), .A1(i_4_), .B0(men_men_n198_), .B1(men_men_n195_), .Y(men_men_n219_));
  NAi21      u0197(.An(i_12_), .B(i_7_), .Y(men_men_n220_));
  NA3        u0198(.A(i_13_), .B(men_men_n196_), .C(i_10_), .Y(men_men_n221_));
  NO2        u0199(.A(men_men_n221_), .B(men_men_n220_), .Y(men_men_n222_));
  NA2        u0200(.A(i_0_), .B(i_5_), .Y(men_men_n223_));
  NA2        u0201(.A(men_men_n223_), .B(men_men_n104_), .Y(men_men_n224_));
  OAI220     u0202(.A0(men_men_n224_), .A1(men_men_n192_), .B0(men_men_n182_), .B1(men_men_n133_), .Y(men_men_n225_));
  NAi31      u0203(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n226_));
  NO2        u0204(.A(men_men_n36_), .B(i_13_), .Y(men_men_n227_));
  NO2        u0205(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n228_));
  NO2        u0206(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n229_));
  NA3        u0207(.A(men_men_n229_), .B(men_men_n228_), .C(men_men_n227_), .Y(men_men_n230_));
  INV        u0208(.A(i_13_), .Y(men_men_n231_));
  NO2        u0209(.A(i_12_), .B(men_men_n231_), .Y(men_men_n232_));
  NA3        u0210(.A(men_men_n232_), .B(men_men_n201_), .C(men_men_n199_), .Y(men_men_n233_));
  OAI210     u0211(.A0(men_men_n230_), .A1(men_men_n226_), .B0(men_men_n233_), .Y(men_men_n234_));
  AOI220     u0212(.A0(men_men_n234_), .A1(men_men_n142_), .B0(men_men_n225_), .B1(men_men_n222_), .Y(men_men_n235_));
  NO2        u0213(.A(i_12_), .B(men_men_n37_), .Y(men_men_n236_));
  NO2        u0214(.A(men_men_n185_), .B(i_4_), .Y(men_men_n237_));
  NA2        u0215(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  OR2        u0216(.A(i_8_), .B(i_7_), .Y(men_men_n239_));
  NO2        u0217(.A(men_men_n239_), .B(men_men_n86_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n53_), .B(i_1_), .Y(men_men_n241_));
  NA2        u0219(.A(men_men_n241_), .B(men_men_n240_), .Y(men_men_n242_));
  INV        u0220(.A(i_12_), .Y(men_men_n243_));
  NO2        u0221(.A(men_men_n44_), .B(men_men_n243_), .Y(men_men_n244_));
  NO3        u0222(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n245_));
  NA2        u0223(.A(i_2_), .B(i_1_), .Y(men_men_n246_));
  NO2        u0224(.A(men_men_n242_), .B(men_men_n238_), .Y(men_men_n247_));
  NO3        u0225(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n248_));
  NAi21      u0226(.An(i_4_), .B(i_3_), .Y(men_men_n249_));
  NO2        u0227(.A(i_0_), .B(i_6_), .Y(men_men_n250_));
  NOi41      u0228(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n251_));
  NA2        u0229(.A(men_men_n251_), .B(men_men_n250_), .Y(men_men_n252_));
  NO2        u0230(.A(men_men_n246_), .B(men_men_n185_), .Y(men_men_n253_));
  NAi21      u0231(.An(men_men_n252_), .B(men_men_n253_), .Y(men_men_n254_));
  INV        u0232(.A(men_men_n254_), .Y(men_men_n255_));
  AOI220     u0233(.A0(men_men_n255_), .A1(men_men_n40_), .B0(men_men_n247_), .B1(men_men_n211_), .Y(men_men_n256_));
  NO2        u0234(.A(i_11_), .B(men_men_n231_), .Y(men_men_n257_));
  NOi21      u0235(.An(i_1_), .B(i_6_), .Y(men_men_n258_));
  NAi21      u0236(.An(i_3_), .B(i_7_), .Y(men_men_n259_));
  NA2        u0237(.A(men_men_n243_), .B(i_9_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n261_));
  NO2        u0239(.A(i_12_), .B(i_3_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n73_), .B(i_5_), .Y(men_men_n263_));
  NA2        u0241(.A(i_3_), .B(i_9_), .Y(men_men_n264_));
  NAi21      u0242(.An(i_7_), .B(i_10_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA3        u0244(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n267_));
  INV        u0245(.A(men_men_n143_), .Y(men_men_n268_));
  NA2        u0246(.A(men_men_n243_), .B(i_13_), .Y(men_men_n269_));
  NO2        u0247(.A(men_men_n269_), .B(men_men_n75_), .Y(men_men_n270_));
  NA2        u0248(.A(men_men_n270_), .B(men_men_n268_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n239_), .B(men_men_n37_), .Y(men_men_n272_));
  NA2        u0250(.A(i_12_), .B(i_6_), .Y(men_men_n273_));
  OR2        u0251(.A(i_13_), .B(i_9_), .Y(men_men_n274_));
  NO3        u0252(.A(men_men_n274_), .B(men_men_n273_), .C(men_men_n48_), .Y(men_men_n275_));
  NO2        u0253(.A(men_men_n249_), .B(i_2_), .Y(men_men_n276_));
  NA3        u0254(.A(men_men_n276_), .B(men_men_n275_), .C(men_men_n44_), .Y(men_men_n277_));
  NA2        u0255(.A(men_men_n257_), .B(i_9_), .Y(men_men_n278_));
  NA2        u0256(.A(men_men_n263_), .B(men_men_n64_), .Y(men_men_n279_));
  OAI210     u0257(.A0(men_men_n279_), .A1(men_men_n278_), .B0(men_men_n277_), .Y(men_men_n280_));
  NA2        u0258(.A(men_men_n155_), .B(men_men_n63_), .Y(men_men_n281_));
  NO3        u0259(.A(i_11_), .B(men_men_n231_), .C(men_men_n25_), .Y(men_men_n282_));
  NO2        u0260(.A(men_men_n259_), .B(i_8_), .Y(men_men_n283_));
  NO2        u0261(.A(i_6_), .B(men_men_n48_), .Y(men_men_n284_));
  NA3        u0262(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n282_), .Y(men_men_n285_));
  NO3        u0263(.A(men_men_n26_), .B(men_men_n86_), .C(i_5_), .Y(men_men_n286_));
  NA3        u0264(.A(men_men_n286_), .B(men_men_n272_), .C(men_men_n232_), .Y(men_men_n287_));
  AOI210     u0265(.A0(men_men_n287_), .A1(men_men_n285_), .B0(men_men_n281_), .Y(men_men_n288_));
  AOI210     u0266(.A0(men_men_n280_), .A1(men_men_n272_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA4        u0267(.A(men_men_n289_), .B(men_men_n271_), .C(men_men_n256_), .D(men_men_n235_), .Y(men_men_n290_));
  NO3        u0268(.A(i_12_), .B(men_men_n231_), .C(men_men_n37_), .Y(men_men_n291_));
  INV        u0269(.A(men_men_n291_), .Y(men_men_n292_));
  NA2        u0270(.A(i_8_), .B(men_men_n101_), .Y(men_men_n293_));
  NO3        u0271(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n294_));
  AOI220     u0272(.A0(men_men_n294_), .A1(men_men_n199_), .B0(men_men_n164_), .B1(men_men_n241_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n295_), .B(men_men_n293_), .Y(men_men_n296_));
  NO3        u0274(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n246_), .B(i_0_), .Y(men_men_n298_));
  AOI220     u0276(.A0(men_men_n298_), .A1(men_men_n197_), .B0(men_men_n297_), .B1(men_men_n142_), .Y(men_men_n299_));
  NA2        u0277(.A(men_men_n284_), .B(men_men_n26_), .Y(men_men_n300_));
  NO2        u0278(.A(men_men_n300_), .B(men_men_n299_), .Y(men_men_n301_));
  NA2        u0279(.A(i_0_), .B(i_1_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n302_), .B(i_2_), .Y(men_men_n303_));
  NO2        u0281(.A(men_men_n59_), .B(i_6_), .Y(men_men_n304_));
  NA3        u0282(.A(men_men_n304_), .B(men_men_n303_), .C(men_men_n164_), .Y(men_men_n305_));
  OAI210     u0283(.A0(men_men_n166_), .A1(men_men_n143_), .B0(men_men_n305_), .Y(men_men_n306_));
  NO3        u0284(.A(men_men_n306_), .B(men_men_n301_), .C(men_men_n296_), .Y(men_men_n307_));
  NO2        u0285(.A(i_3_), .B(i_10_), .Y(men_men_n308_));
  NA3        u0286(.A(men_men_n308_), .B(men_men_n40_), .C(men_men_n44_), .Y(men_men_n309_));
  NO2        u0287(.A(i_2_), .B(men_men_n101_), .Y(men_men_n310_));
  NA2        u0288(.A(i_1_), .B(men_men_n36_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n311_), .B(i_8_), .Y(men_men_n312_));
  NA2        u0290(.A(men_men_n312_), .B(men_men_n310_), .Y(men_men_n313_));
  AN2        u0291(.A(i_3_), .B(i_10_), .Y(men_men_n314_));
  NA4        u0292(.A(men_men_n314_), .B(men_men_n201_), .C(men_men_n178_), .D(men_men_n176_), .Y(men_men_n315_));
  NO2        u0293(.A(i_5_), .B(men_men_n37_), .Y(men_men_n316_));
  NO2        u0294(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n317_));
  OR2        u0295(.A(men_men_n313_), .B(men_men_n309_), .Y(men_men_n318_));
  OAI220     u0296(.A0(men_men_n318_), .A1(i_6_), .B0(men_men_n307_), .B1(men_men_n292_), .Y(men_men_n319_));
  NO4        u0297(.A(men_men_n319_), .B(men_men_n290_), .C(men_men_n219_), .D(men_men_n169_), .Y(men_men_n320_));
  NO3        u0298(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n321_));
  NO2        u0299(.A(men_men_n59_), .B(men_men_n86_), .Y(men_men_n322_));
  NA2        u0300(.A(men_men_n298_), .B(men_men_n322_), .Y(men_men_n323_));
  NO3        u0301(.A(i_6_), .B(men_men_n196_), .C(i_7_), .Y(men_men_n324_));
  NA2        u0302(.A(men_men_n324_), .B(men_men_n201_), .Y(men_men_n325_));
  AOI210     u0303(.A0(men_men_n325_), .A1(men_men_n323_), .B0(men_men_n171_), .Y(men_men_n326_));
  NO2        u0304(.A(i_2_), .B(i_3_), .Y(men_men_n327_));
  OR2        u0305(.A(i_0_), .B(i_5_), .Y(men_men_n328_));
  NA2        u0306(.A(men_men_n223_), .B(men_men_n328_), .Y(men_men_n329_));
  NA4        u0307(.A(men_men_n329_), .B(men_men_n240_), .C(men_men_n327_), .D(i_1_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n298_), .B(men_men_n164_), .C(men_men_n112_), .Y(men_men_n331_));
  NAi21      u0309(.An(i_8_), .B(i_7_), .Y(men_men_n332_));
  NO2        u0310(.A(men_men_n332_), .B(i_6_), .Y(men_men_n333_));
  NO2        u0311(.A(men_men_n158_), .B(men_men_n46_), .Y(men_men_n334_));
  NA3        u0312(.A(men_men_n334_), .B(men_men_n333_), .C(men_men_n164_), .Y(men_men_n335_));
  NA3        u0313(.A(men_men_n335_), .B(men_men_n331_), .C(men_men_n330_), .Y(men_men_n336_));
  OAI210     u0314(.A0(men_men_n336_), .A1(men_men_n326_), .B0(i_4_), .Y(men_men_n337_));
  NO2        u0315(.A(i_12_), .B(i_10_), .Y(men_men_n338_));
  NOi21      u0316(.An(i_5_), .B(i_0_), .Y(men_men_n339_));
  NO3        u0317(.A(men_men_n311_), .B(men_men_n339_), .C(men_men_n128_), .Y(men_men_n340_));
  NA4        u0318(.A(men_men_n84_), .B(men_men_n36_), .C(men_men_n86_), .D(i_8_), .Y(men_men_n341_));
  NA2        u0319(.A(men_men_n340_), .B(men_men_n338_), .Y(men_men_n342_));
  NO2        u0320(.A(i_6_), .B(i_8_), .Y(men_men_n343_));
  NOi21      u0321(.An(i_0_), .B(i_2_), .Y(men_men_n344_));
  AN2        u0322(.A(men_men_n344_), .B(men_men_n343_), .Y(men_men_n345_));
  NO2        u0323(.A(i_1_), .B(i_7_), .Y(men_men_n346_));
  AO220      u0324(.A0(men_men_n346_), .A1(men_men_n345_), .B0(men_men_n333_), .B1(men_men_n241_), .Y(men_men_n347_));
  NA3        u0325(.A(men_men_n347_), .B(i_4_), .C(i_5_), .Y(men_men_n348_));
  NA3        u0326(.A(men_men_n348_), .B(men_men_n342_), .C(men_men_n337_), .Y(men_men_n349_));
  NO3        u0327(.A(men_men_n239_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n350_));
  NO3        u0328(.A(men_men_n332_), .B(i_2_), .C(i_1_), .Y(men_men_n351_));
  OAI210     u0329(.A0(men_men_n351_), .A1(men_men_n350_), .B0(i_6_), .Y(men_men_n352_));
  NA2        u0330(.A(men_men_n258_), .B(men_men_n310_), .Y(men_men_n353_));
  AOI210     u0331(.A0(men_men_n353_), .A1(men_men_n352_), .B0(men_men_n329_), .Y(men_men_n354_));
  NOi21      u0332(.An(men_men_n154_), .B(men_men_n104_), .Y(men_men_n355_));
  NO2        u0333(.A(men_men_n355_), .B(men_men_n124_), .Y(men_men_n356_));
  OAI210     u0334(.A0(men_men_n356_), .A1(men_men_n354_), .B0(i_3_), .Y(men_men_n357_));
  INV        u0335(.A(men_men_n84_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n302_), .B(men_men_n81_), .Y(men_men_n359_));
  NA2        u0337(.A(men_men_n359_), .B(men_men_n132_), .Y(men_men_n360_));
  NO2        u0338(.A(men_men_n92_), .B(men_men_n196_), .Y(men_men_n361_));
  NA2        u0339(.A(men_men_n361_), .B(men_men_n63_), .Y(men_men_n362_));
  AOI210     u0340(.A0(men_men_n362_), .A1(men_men_n360_), .B0(men_men_n358_), .Y(men_men_n363_));
  NO2        u0341(.A(men_men_n196_), .B(i_9_), .Y(men_men_n364_));
  NO2        u0342(.A(men_men_n363_), .B(men_men_n301_), .Y(men_men_n365_));
  AOI210     u0343(.A0(men_men_n365_), .A1(men_men_n357_), .B0(men_men_n163_), .Y(men_men_n366_));
  AOI210     u0344(.A0(men_men_n349_), .A1(men_men_n321_), .B0(men_men_n366_), .Y(men_men_n367_));
  NOi32      u0345(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n368_));
  INV        u0346(.A(men_men_n368_), .Y(men_men_n369_));
  NAi21      u0347(.An(i_0_), .B(i_6_), .Y(men_men_n370_));
  NAi21      u0348(.An(i_1_), .B(i_5_), .Y(men_men_n371_));
  NA2        u0349(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  NA2        u0350(.A(men_men_n372_), .B(men_men_n25_), .Y(men_men_n373_));
  OAI210     u0351(.A0(men_men_n373_), .A1(men_men_n160_), .B0(men_men_n252_), .Y(men_men_n374_));
  NAi41      u0352(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n375_));
  AOI210     u0353(.A0(men_men_n375_), .A1(men_men_n160_), .B0(men_men_n158_), .Y(men_men_n376_));
  NOi32      u0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n377_));
  NO2        u0355(.A(i_1_), .B(men_men_n101_), .Y(men_men_n378_));
  NAi21      u0356(.An(i_3_), .B(i_4_), .Y(men_men_n379_));
  NO2        u0357(.A(men_men_n379_), .B(i_9_), .Y(men_men_n380_));
  AN2        u0358(.A(i_6_), .B(i_7_), .Y(men_men_n381_));
  OAI210     u0359(.A0(men_men_n381_), .A1(men_men_n378_), .B0(men_men_n380_), .Y(men_men_n382_));
  NA2        u0360(.A(i_2_), .B(i_7_), .Y(men_men_n383_));
  NO2        u0361(.A(men_men_n379_), .B(i_10_), .Y(men_men_n384_));
  NA3        u0362(.A(men_men_n384_), .B(men_men_n383_), .C(men_men_n250_), .Y(men_men_n385_));
  AOI210     u0363(.A0(men_men_n385_), .A1(men_men_n382_), .B0(men_men_n188_), .Y(men_men_n386_));
  AOI210     u0364(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n387_));
  OAI210     u0365(.A0(men_men_n387_), .A1(men_men_n191_), .B0(men_men_n384_), .Y(men_men_n388_));
  AOI220     u0366(.A0(men_men_n384_), .A1(men_men_n346_), .B0(men_men_n245_), .B1(men_men_n191_), .Y(men_men_n389_));
  AOI210     u0367(.A0(men_men_n389_), .A1(men_men_n388_), .B0(i_5_), .Y(men_men_n390_));
  NO4        u0368(.A(men_men_n390_), .B(men_men_n386_), .C(men_men_n376_), .D(men_men_n374_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n391_), .B(men_men_n369_), .Y(men_men_n392_));
  NO2        u0370(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n393_));
  AN2        u0371(.A(i_12_), .B(i_5_), .Y(men_men_n394_));
  NO2        u0372(.A(i_4_), .B(men_men_n26_), .Y(men_men_n395_));
  NA2        u0373(.A(men_men_n395_), .B(men_men_n394_), .Y(men_men_n396_));
  NO2        u0374(.A(i_11_), .B(i_6_), .Y(men_men_n397_));
  NA3        u0375(.A(men_men_n397_), .B(men_men_n334_), .C(men_men_n231_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n398_), .B(men_men_n396_), .Y(men_men_n399_));
  NO2        u0377(.A(men_men_n249_), .B(i_5_), .Y(men_men_n400_));
  NO2        u0378(.A(i_5_), .B(i_10_), .Y(men_men_n401_));
  NA2        u0379(.A(men_men_n400_), .B(men_men_n201_), .Y(men_men_n402_));
  NA2        u0380(.A(men_men_n144_), .B(men_men_n45_), .Y(men_men_n403_));
  NO2        u0381(.A(men_men_n403_), .B(men_men_n402_), .Y(men_men_n404_));
  OAI210     u0382(.A0(men_men_n404_), .A1(men_men_n399_), .B0(men_men_n393_), .Y(men_men_n405_));
  NO2        u0383(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n406_));
  NO2        u0384(.A(men_men_n150_), .B(men_men_n86_), .Y(men_men_n407_));
  OAI210     u0385(.A0(men_men_n407_), .A1(men_men_n399_), .B0(men_men_n406_), .Y(men_men_n408_));
  NO3        u0386(.A(men_men_n86_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n409_));
  NO2        u0387(.A(i_11_), .B(i_12_), .Y(men_men_n410_));
  NA2        u0388(.A(men_men_n401_), .B(men_men_n243_), .Y(men_men_n411_));
  NA3        u0389(.A(men_men_n112_), .B(i_4_), .C(i_11_), .Y(men_men_n412_));
  OAI220     u0390(.A0(men_men_n412_), .A1(men_men_n226_), .B0(men_men_n411_), .B1(men_men_n341_), .Y(men_men_n413_));
  NAi21      u0391(.An(i_13_), .B(i_0_), .Y(men_men_n414_));
  NO2        u0392(.A(men_men_n414_), .B(men_men_n246_), .Y(men_men_n415_));
  NA2        u0393(.A(men_men_n413_), .B(men_men_n415_), .Y(men_men_n416_));
  NA3        u0394(.A(men_men_n416_), .B(men_men_n408_), .C(men_men_n405_), .Y(men_men_n417_));
  NA2        u0395(.A(men_men_n44_), .B(men_men_n231_), .Y(men_men_n418_));
  NO3        u0396(.A(i_1_), .B(i_12_), .C(men_men_n86_), .Y(men_men_n419_));
  NO2        u0397(.A(i_0_), .B(i_11_), .Y(men_men_n420_));
  INV        u0398(.A(i_5_), .Y(men_men_n421_));
  AN2        u0399(.A(i_1_), .B(i_6_), .Y(men_men_n422_));
  NOi21      u0400(.An(i_2_), .B(i_12_), .Y(men_men_n423_));
  NA2        u0401(.A(men_men_n423_), .B(men_men_n422_), .Y(men_men_n424_));
  NO2        u0402(.A(men_men_n424_), .B(men_men_n421_), .Y(men_men_n425_));
  NA2        u0403(.A(men_men_n142_), .B(i_9_), .Y(men_men_n426_));
  NO2        u0404(.A(men_men_n426_), .B(i_4_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n425_), .B(men_men_n427_), .Y(men_men_n428_));
  NAi21      u0406(.An(i_9_), .B(i_4_), .Y(men_men_n429_));
  OR2        u0407(.A(i_13_), .B(i_10_), .Y(men_men_n430_));
  NO3        u0408(.A(men_men_n430_), .B(men_men_n117_), .C(men_men_n429_), .Y(men_men_n431_));
  NO2        u0409(.A(men_men_n174_), .B(men_men_n123_), .Y(men_men_n432_));
  OR2        u0410(.A(men_men_n221_), .B(men_men_n220_), .Y(men_men_n433_));
  NO2        u0411(.A(men_men_n101_), .B(men_men_n25_), .Y(men_men_n434_));
  NA2        u0412(.A(men_men_n291_), .B(men_men_n434_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n284_), .B(men_men_n215_), .Y(men_men_n436_));
  OAI220     u0414(.A0(men_men_n436_), .A1(men_men_n433_), .B0(men_men_n435_), .B1(men_men_n355_), .Y(men_men_n437_));
  INV        u0415(.A(men_men_n437_), .Y(men_men_n438_));
  AOI210     u0416(.A0(men_men_n438_), .A1(men_men_n428_), .B0(men_men_n26_), .Y(men_men_n439_));
  NA2        u0417(.A(men_men_n331_), .B(men_men_n330_), .Y(men_men_n440_));
  AOI220     u0418(.A0(men_men_n304_), .A1(men_men_n294_), .B0(men_men_n298_), .B1(men_men_n322_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n441_), .B(men_men_n171_), .Y(men_men_n442_));
  NO2        u0420(.A(men_men_n185_), .B(men_men_n86_), .Y(men_men_n443_));
  AOI220     u0421(.A0(men_men_n443_), .A1(men_men_n303_), .B0(men_men_n286_), .B1(men_men_n215_), .Y(men_men_n444_));
  NO2        u0422(.A(men_men_n444_), .B(men_men_n293_), .Y(men_men_n445_));
  NO3        u0423(.A(men_men_n445_), .B(men_men_n442_), .C(men_men_n440_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n199_), .B(men_men_n96_), .Y(men_men_n447_));
  NA3        u0425(.A(men_men_n334_), .B(men_men_n164_), .C(men_men_n86_), .Y(men_men_n448_));
  AOI210     u0426(.A0(men_men_n448_), .A1(men_men_n447_), .B0(men_men_n332_), .Y(men_men_n449_));
  NA2        u0427(.A(men_men_n304_), .B(men_men_n241_), .Y(men_men_n450_));
  NO2        u0428(.A(men_men_n450_), .B(men_men_n185_), .Y(men_men_n451_));
  NO2        u0429(.A(i_3_), .B(men_men_n48_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n451_), .B(men_men_n449_), .Y(men_men_n453_));
  AOI210     u0431(.A0(men_men_n453_), .A1(men_men_n446_), .B0(men_men_n278_), .Y(men_men_n454_));
  NO4        u0432(.A(men_men_n454_), .B(men_men_n439_), .C(men_men_n417_), .D(men_men_n392_), .Y(men_men_n455_));
  NO2        u0433(.A(men_men_n63_), .B(i_4_), .Y(men_men_n456_));
  NO2        u0434(.A(men_men_n73_), .B(i_13_), .Y(men_men_n457_));
  NO2        u0435(.A(i_10_), .B(i_9_), .Y(men_men_n458_));
  NAi21      u0436(.An(i_12_), .B(i_8_), .Y(men_men_n459_));
  NO2        u0437(.A(men_men_n459_), .B(i_3_), .Y(men_men_n460_));
  NO2        u0438(.A(men_men_n46_), .B(i_4_), .Y(men_men_n461_));
  NA2        u0439(.A(men_men_n461_), .B(men_men_n104_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n462_), .B(men_men_n208_), .Y(men_men_n463_));
  NA2        u0441(.A(men_men_n317_), .B(i_0_), .Y(men_men_n464_));
  NO3        u0442(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n273_), .B(men_men_n97_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n466_), .B(men_men_n465_), .Y(men_men_n467_));
  NA2        u0445(.A(i_8_), .B(i_9_), .Y(men_men_n468_));
  AOI210     u0446(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n469_));
  OR2        u0447(.A(men_men_n469_), .B(men_men_n468_), .Y(men_men_n470_));
  NA2        u0448(.A(men_men_n291_), .B(men_men_n209_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n471_), .B(men_men_n470_), .Y(men_men_n472_));
  NA2        u0450(.A(men_men_n257_), .B(men_men_n316_), .Y(men_men_n473_));
  NO3        u0451(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n474_));
  INV        u0452(.A(men_men_n474_), .Y(men_men_n475_));
  NA3        u0453(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n476_));
  NA4        u0454(.A(men_men_n145_), .B(men_men_n115_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n477_));
  OAI220     u0455(.A0(men_men_n477_), .A1(men_men_n476_), .B0(men_men_n475_), .B1(men_men_n473_), .Y(men_men_n478_));
  NO3        u0456(.A(men_men_n478_), .B(men_men_n472_), .C(men_men_n463_), .Y(men_men_n479_));
  OR2        u0457(.A(men_men_n302_), .B(men_men_n212_), .Y(men_men_n480_));
  BUFFER     u0458(.A(men_men_n305_), .Y(men_men_n481_));
  OA220      u0459(.A0(men_men_n481_), .A1(men_men_n163_), .B0(men_men_n480_), .B1(men_men_n238_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n96_), .B(i_13_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n443_), .B(men_men_n393_), .Y(men_men_n484_));
  NO2        u0462(.A(i_2_), .B(i_13_), .Y(men_men_n485_));
  NA3        u0463(.A(men_men_n485_), .B(men_men_n162_), .C(men_men_n99_), .Y(men_men_n486_));
  OAI220     u0464(.A0(men_men_n486_), .A1(men_men_n243_), .B0(men_men_n484_), .B1(men_men_n483_), .Y(men_men_n487_));
  NO3        u0465(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n488_));
  NO2        u0466(.A(i_6_), .B(i_7_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n490_));
  NO2        u0468(.A(i_11_), .B(i_1_), .Y(men_men_n491_));
  NO2        u0469(.A(men_men_n73_), .B(i_3_), .Y(men_men_n492_));
  OR2        u0470(.A(i_11_), .B(i_8_), .Y(men_men_n493_));
  NOi21      u0471(.An(i_2_), .B(i_7_), .Y(men_men_n494_));
  NAi31      u0472(.An(men_men_n493_), .B(men_men_n494_), .C(men_men_n492_), .Y(men_men_n495_));
  INV        u0473(.A(men_men_n430_), .Y(men_men_n496_));
  NA3        u0474(.A(men_men_n496_), .B(men_men_n456_), .C(men_men_n75_), .Y(men_men_n497_));
  NO2        u0475(.A(men_men_n497_), .B(men_men_n495_), .Y(men_men_n498_));
  NO2        u0476(.A(i_3_), .B(men_men_n196_), .Y(men_men_n499_));
  NO2        u0477(.A(i_6_), .B(i_10_), .Y(men_men_n500_));
  NA4        u0478(.A(men_men_n500_), .B(men_men_n321_), .C(men_men_n499_), .D(men_men_n243_), .Y(men_men_n501_));
  NO2        u0479(.A(men_men_n501_), .B(men_men_n156_), .Y(men_men_n502_));
  NA2        u0480(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n503_));
  NO2        u0481(.A(men_men_n158_), .B(i_3_), .Y(men_men_n504_));
  NAi31      u0482(.An(men_men_n503_), .B(men_men_n504_), .C(men_men_n232_), .Y(men_men_n505_));
  NA3        u0483(.A(men_men_n406_), .B(men_men_n181_), .C(men_men_n149_), .Y(men_men_n506_));
  NA2        u0484(.A(men_men_n506_), .B(men_men_n505_), .Y(men_men_n507_));
  NO4        u0485(.A(men_men_n507_), .B(men_men_n502_), .C(men_men_n498_), .D(men_men_n487_), .Y(men_men_n508_));
  NA2        u0486(.A(men_men_n474_), .B(men_men_n401_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n509_), .B(men_men_n230_), .Y(men_men_n510_));
  NAi21      u0488(.An(men_men_n221_), .B(men_men_n410_), .Y(men_men_n511_));
  NA2        u0489(.A(men_men_n346_), .B(men_men_n223_), .Y(men_men_n512_));
  NO2        u0490(.A(men_men_n26_), .B(i_5_), .Y(men_men_n513_));
  NO2        u0491(.A(i_0_), .B(men_men_n86_), .Y(men_men_n514_));
  NA3        u0492(.A(men_men_n514_), .B(men_men_n513_), .C(men_men_n142_), .Y(men_men_n515_));
  OR3        u0493(.A(men_men_n311_), .B(men_men_n38_), .C(men_men_n46_), .Y(men_men_n516_));
  OAI220     u0494(.A0(men_men_n516_), .A1(men_men_n515_), .B0(men_men_n512_), .B1(men_men_n511_), .Y(men_men_n517_));
  NA4        u0495(.A(men_men_n314_), .B(men_men_n229_), .C(men_men_n73_), .D(men_men_n243_), .Y(men_men_n518_));
  NO2        u0496(.A(men_men_n518_), .B(men_men_n490_), .Y(men_men_n519_));
  NO3        u0497(.A(men_men_n519_), .B(men_men_n517_), .C(men_men_n510_), .Y(men_men_n520_));
  NA4        u0498(.A(men_men_n520_), .B(men_men_n508_), .C(men_men_n482_), .D(men_men_n479_), .Y(men_men_n521_));
  NA3        u0499(.A(men_men_n314_), .B(men_men_n178_), .C(men_men_n176_), .Y(men_men_n522_));
  INV        u0500(.A(men_men_n522_), .Y(men_men_n523_));
  AN2        u0501(.A(men_men_n294_), .B(men_men_n240_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n524_), .B(men_men_n523_), .Y(men_men_n525_));
  NA2        u0503(.A(men_men_n122_), .B(men_men_n111_), .Y(men_men_n526_));
  AN2        u0504(.A(men_men_n526_), .B(men_men_n465_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n321_), .B(men_men_n165_), .Y(men_men_n528_));
  OAI210     u0506(.A0(men_men_n528_), .A1(men_men_n238_), .B0(men_men_n315_), .Y(men_men_n529_));
  AOI220     u0507(.A0(men_men_n529_), .A1(men_men_n333_), .B0(men_men_n527_), .B1(men_men_n317_), .Y(men_men_n530_));
  NA2        u0508(.A(men_men_n394_), .B(men_men_n231_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n368_), .B(men_men_n73_), .Y(men_men_n532_));
  NA2        u0510(.A(men_men_n381_), .B(men_men_n377_), .Y(men_men_n533_));
  AO210      u0511(.A0(men_men_n532_), .A1(men_men_n531_), .B0(men_men_n533_), .Y(men_men_n534_));
  NO2        u0512(.A(men_men_n36_), .B(i_8_), .Y(men_men_n535_));
  AOI210     u0513(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n431_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n536_), .B(men_men_n534_), .Y(men_men_n537_));
  INV        u0515(.A(men_men_n537_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n263_), .B(men_men_n64_), .Y(men_men_n539_));
  OAI210     u0517(.A0(i_8_), .A1(men_men_n539_), .B0(men_men_n134_), .Y(men_men_n540_));
  NO2        u0518(.A(i_7_), .B(men_men_n202_), .Y(men_men_n541_));
  OR2        u0519(.A(men_men_n185_), .B(i_4_), .Y(men_men_n542_));
  NO2        u0520(.A(men_men_n542_), .B(men_men_n86_), .Y(men_men_n543_));
  AOI220     u0521(.A0(men_men_n543_), .A1(men_men_n541_), .B0(men_men_n540_), .B1(men_men_n432_), .Y(men_men_n544_));
  NA4        u0522(.A(men_men_n544_), .B(men_men_n538_), .C(men_men_n530_), .D(men_men_n525_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n400_), .B(men_men_n303_), .Y(men_men_n546_));
  OAI210     u0524(.A0(men_men_n396_), .A1(men_men_n170_), .B0(men_men_n546_), .Y(men_men_n547_));
  NA2        u0525(.A(men_men_n1082_), .B(men_men_n231_), .Y(men_men_n548_));
  NA2        u0526(.A(men_men_n500_), .B(men_men_n27_), .Y(men_men_n549_));
  NO2        u0527(.A(men_men_n549_), .B(men_men_n548_), .Y(men_men_n550_));
  NOi31      u0528(.An(men_men_n324_), .B(men_men_n430_), .C(men_men_n38_), .Y(men_men_n551_));
  OAI210     u0529(.A0(men_men_n551_), .A1(men_men_n550_), .B0(men_men_n547_), .Y(men_men_n552_));
  NO2        u0530(.A(i_8_), .B(i_7_), .Y(men_men_n553_));
  OAI210     u0531(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n554_), .B(men_men_n229_), .Y(men_men_n555_));
  AOI220     u0533(.A0(men_men_n334_), .A1(men_men_n40_), .B0(men_men_n241_), .B1(men_men_n211_), .Y(men_men_n556_));
  OAI220     u0534(.A0(men_men_n556_), .A1(men_men_n542_), .B0(men_men_n555_), .B1(men_men_n249_), .Y(men_men_n557_));
  NA2        u0535(.A(men_men_n44_), .B(i_10_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n558_), .B(i_6_), .Y(men_men_n559_));
  NA3        u0537(.A(men_men_n559_), .B(men_men_n557_), .C(men_men_n553_), .Y(men_men_n560_));
  AOI220     u0538(.A0(men_men_n443_), .A1(men_men_n334_), .B0(men_men_n253_), .B1(men_men_n250_), .Y(men_men_n561_));
  NO2        u0539(.A(men_men_n561_), .B(men_men_n269_), .Y(men_men_n562_));
  NA2        u0540(.A(men_men_n562_), .B(men_men_n272_), .Y(men_men_n563_));
  NOi31      u0541(.An(men_men_n298_), .B(men_men_n309_), .C(men_men_n183_), .Y(men_men_n564_));
  NA3        u0542(.A(men_men_n314_), .B(men_men_n176_), .C(men_men_n96_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n227_), .B(men_men_n44_), .Y(men_men_n566_));
  NO2        u0544(.A(men_men_n158_), .B(i_5_), .Y(men_men_n567_));
  NA3        u0545(.A(men_men_n567_), .B(men_men_n418_), .C(men_men_n327_), .Y(men_men_n568_));
  OAI210     u0546(.A0(men_men_n568_), .A1(men_men_n566_), .B0(men_men_n565_), .Y(men_men_n569_));
  OAI210     u0547(.A0(men_men_n569_), .A1(men_men_n564_), .B0(men_men_n474_), .Y(men_men_n570_));
  NA4        u0548(.A(men_men_n570_), .B(men_men_n563_), .C(men_men_n560_), .D(men_men_n552_), .Y(men_men_n571_));
  NA3        u0549(.A(men_men_n223_), .B(men_men_n71_), .C(men_men_n44_), .Y(men_men_n572_));
  NA2        u0550(.A(men_men_n291_), .B(men_men_n84_), .Y(men_men_n573_));
  AOI210     u0551(.A0(men_men_n572_), .A1(men_men_n360_), .B0(men_men_n573_), .Y(men_men_n574_));
  NA2        u0552(.A(men_men_n304_), .B(men_men_n294_), .Y(men_men_n575_));
  NO2        u0553(.A(men_men_n575_), .B(men_men_n175_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n577_));
  NA2        u0555(.A(men_men_n458_), .B(men_men_n227_), .Y(men_men_n578_));
  NO2        u0556(.A(men_men_n577_), .B(men_men_n578_), .Y(men_men_n579_));
  NA2        u0557(.A(i_0_), .B(men_men_n48_), .Y(men_men_n580_));
  NO3        u0558(.A(men_men_n579_), .B(men_men_n576_), .C(men_men_n574_), .Y(men_men_n581_));
  NO4        u0559(.A(men_men_n258_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n582_));
  NO3        u0560(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n239_), .B(men_men_n36_), .Y(men_men_n584_));
  AN2        u0562(.A(men_men_n584_), .B(men_men_n583_), .Y(men_men_n585_));
  OA210      u0563(.A0(men_men_n585_), .A1(men_men_n582_), .B0(men_men_n368_), .Y(men_men_n586_));
  NO2        u0564(.A(men_men_n430_), .B(i_1_), .Y(men_men_n587_));
  NOi31      u0565(.An(men_men_n587_), .B(men_men_n466_), .C(men_men_n73_), .Y(men_men_n588_));
  AN4        u0566(.A(men_men_n588_), .B(men_men_n427_), .C(men_men_n513_), .D(i_2_), .Y(men_men_n589_));
  NO2        u0567(.A(men_men_n441_), .B(men_men_n179_), .Y(men_men_n590_));
  NO3        u0568(.A(men_men_n590_), .B(men_men_n589_), .C(men_men_n586_), .Y(men_men_n591_));
  NOi21      u0569(.An(i_10_), .B(i_6_), .Y(men_men_n592_));
  NO2        u0570(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n593_));
  AOI220     u0571(.A0(men_men_n291_), .A1(men_men_n593_), .B0(men_men_n282_), .B1(men_men_n592_), .Y(men_men_n594_));
  NO2        u0572(.A(men_men_n594_), .B(men_men_n464_), .Y(men_men_n595_));
  NO2        u0573(.A(men_men_n114_), .B(men_men_n23_), .Y(men_men_n596_));
  NA2        u0574(.A(men_men_n324_), .B(men_men_n165_), .Y(men_men_n597_));
  AOI220     u0575(.A0(men_men_n597_), .A1(men_men_n450_), .B0(men_men_n186_), .B1(men_men_n184_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n598_), .B(men_men_n595_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n532_), .B(men_men_n389_), .Y(men_men_n600_));
  INV        u0578(.A(men_men_n327_), .Y(men_men_n601_));
  NO2        u0579(.A(i_12_), .B(men_men_n86_), .Y(men_men_n602_));
  NA3        u0580(.A(men_men_n602_), .B(men_men_n282_), .C(men_men_n580_), .Y(men_men_n603_));
  NA3        u0581(.A(men_men_n397_), .B(men_men_n291_), .C(men_men_n223_), .Y(men_men_n604_));
  AOI210     u0582(.A0(men_men_n604_), .A1(men_men_n603_), .B0(men_men_n601_), .Y(men_men_n605_));
  NO3        u0583(.A(i_4_), .B(men_men_n352_), .C(men_men_n309_), .Y(men_men_n606_));
  OR2        u0584(.A(i_2_), .B(i_5_), .Y(men_men_n607_));
  OR2        u0585(.A(men_men_n607_), .B(men_men_n422_), .Y(men_men_n608_));
  NO2        u0586(.A(men_men_n608_), .B(men_men_n511_), .Y(men_men_n609_));
  NO4        u0587(.A(men_men_n609_), .B(men_men_n606_), .C(men_men_n605_), .D(men_men_n600_), .Y(men_men_n610_));
  NA4        u0588(.A(men_men_n610_), .B(men_men_n599_), .C(men_men_n591_), .D(men_men_n581_), .Y(men_men_n611_));
  NO4        u0589(.A(men_men_n611_), .B(men_men_n571_), .C(men_men_n545_), .D(men_men_n521_), .Y(men_men_n612_));
  NA4        u0590(.A(men_men_n612_), .B(men_men_n455_), .C(men_men_n367_), .D(men_men_n320_), .Y(men7));
  NO2        u0591(.A(men_men_n92_), .B(men_men_n54_), .Y(men_men_n614_));
  NO2        u0592(.A(men_men_n108_), .B(men_men_n89_), .Y(men_men_n615_));
  NA2        u0593(.A(men_men_n500_), .B(men_men_n84_), .Y(men_men_n616_));
  NA2        u0594(.A(i_11_), .B(men_men_n196_), .Y(men_men_n617_));
  NA3        u0595(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n618_));
  NO2        u0596(.A(men_men_n243_), .B(i_4_), .Y(men_men_n619_));
  NA2        u0597(.A(men_men_n619_), .B(i_8_), .Y(men_men_n620_));
  NO2        u0598(.A(men_men_n105_), .B(men_men_n618_), .Y(men_men_n621_));
  NA2        u0599(.A(i_2_), .B(men_men_n86_), .Y(men_men_n622_));
  OAI210     u0600(.A0(men_men_n87_), .A1(men_men_n206_), .B0(men_men_n207_), .Y(men_men_n623_));
  NO2        u0601(.A(i_7_), .B(men_men_n37_), .Y(men_men_n624_));
  NA2        u0602(.A(i_4_), .B(i_8_), .Y(men_men_n625_));
  AOI210     u0603(.A0(men_men_n625_), .A1(men_men_n314_), .B0(men_men_n624_), .Y(men_men_n626_));
  OAI220     u0604(.A0(men_men_n626_), .A1(men_men_n622_), .B0(men_men_n623_), .B1(i_13_), .Y(men_men_n627_));
  NO3        u0605(.A(men_men_n627_), .B(men_men_n621_), .C(men_men_n614_), .Y(men_men_n628_));
  AOI210     u0606(.A0(men_men_n128_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n629_));
  AOI210     u0607(.A0(men_men_n629_), .A1(men_men_n243_), .B0(men_men_n162_), .Y(men_men_n630_));
  OR2        u0608(.A(i_6_), .B(i_10_), .Y(men_men_n631_));
  NO2        u0609(.A(men_men_n631_), .B(men_men_n23_), .Y(men_men_n632_));
  OR3        u0610(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n633_));
  NO3        u0611(.A(men_men_n633_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n634_));
  INV        u0612(.A(men_men_n203_), .Y(men_men_n635_));
  NO2        u0613(.A(men_men_n634_), .B(men_men_n632_), .Y(men_men_n636_));
  OA220      u0614(.A0(men_men_n636_), .A1(men_men_n601_), .B0(men_men_n630_), .B1(men_men_n274_), .Y(men_men_n637_));
  AOI210     u0615(.A0(men_men_n637_), .A1(men_men_n628_), .B0(men_men_n63_), .Y(men_men_n638_));
  NOi21      u0616(.An(i_11_), .B(i_7_), .Y(men_men_n639_));
  AO210      u0617(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n640_));
  NO2        u0618(.A(men_men_n640_), .B(men_men_n639_), .Y(men_men_n641_));
  NA2        u0619(.A(men_men_n641_), .B(men_men_n211_), .Y(men_men_n642_));
  NA3        u0620(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n643_));
  NAi31      u0621(.An(men_men_n643_), .B(men_men_n220_), .C(i_11_), .Y(men_men_n644_));
  AOI210     u0622(.A0(men_men_n644_), .A1(men_men_n642_), .B0(men_men_n63_), .Y(men_men_n645_));
  NO3        u0623(.A(men_men_n265_), .B(men_men_n213_), .C(men_men_n617_), .Y(men_men_n646_));
  OAI210     u0624(.A0(men_men_n646_), .A1(men_men_n232_), .B0(men_men_n63_), .Y(men_men_n647_));
  NA2        u0625(.A(men_men_n423_), .B(men_men_n31_), .Y(men_men_n648_));
  OR2        u0626(.A(men_men_n213_), .B(men_men_n108_), .Y(men_men_n649_));
  NA2        u0627(.A(men_men_n649_), .B(men_men_n648_), .Y(men_men_n650_));
  NO2        u0628(.A(men_men_n63_), .B(i_9_), .Y(men_men_n651_));
  NO2        u0629(.A(men_men_n651_), .B(i_4_), .Y(men_men_n652_));
  NA2        u0630(.A(men_men_n652_), .B(men_men_n650_), .Y(men_men_n653_));
  NO2        u0631(.A(i_1_), .B(i_12_), .Y(men_men_n654_));
  NA2        u0632(.A(men_men_n653_), .B(men_men_n647_), .Y(men_men_n655_));
  OAI210     u0633(.A0(men_men_n655_), .A1(men_men_n645_), .B0(i_6_), .Y(men_men_n656_));
  NO2        u0634(.A(men_men_n643_), .B(men_men_n108_), .Y(men_men_n657_));
  NA2        u0635(.A(men_men_n657_), .B(men_men_n602_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n243_), .B(men_men_n86_), .Y(men_men_n659_));
  NO2        u0637(.A(men_men_n659_), .B(i_11_), .Y(men_men_n660_));
  NA2        u0638(.A(men_men_n658_), .B(men_men_n467_), .Y(men_men_n661_));
  NO4        u0639(.A(men_men_n220_), .B(men_men_n128_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(men_men_n651_), .Y(men_men_n663_));
  NA2        u0641(.A(men_men_n243_), .B(i_6_), .Y(men_men_n664_));
  NO3        u0642(.A(men_men_n631_), .B(men_men_n239_), .C(men_men_n23_), .Y(men_men_n665_));
  AOI210     u0643(.A0(i_1_), .A1(men_men_n266_), .B0(men_men_n665_), .Y(men_men_n666_));
  OAI210     u0644(.A0(men_men_n666_), .A1(men_men_n44_), .B0(men_men_n663_), .Y(men_men_n667_));
  NA3        u0645(.A(men_men_n553_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n668_));
  NA2        u0646(.A(men_men_n138_), .B(i_9_), .Y(men_men_n669_));
  NA3        u0647(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n670_));
  NO2        u0648(.A(men_men_n46_), .B(i_1_), .Y(men_men_n671_));
  NA3        u0649(.A(men_men_n671_), .B(men_men_n273_), .C(men_men_n44_), .Y(men_men_n672_));
  OAI220     u0650(.A0(men_men_n672_), .A1(men_men_n670_), .B0(men_men_n669_), .B1(men_men_n1080_), .Y(men_men_n673_));
  AOI210     u0651(.A0(men_men_n491_), .A1(men_men_n434_), .B0(men_men_n248_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(men_men_n622_), .Y(men_men_n675_));
  NAi21      u0653(.An(men_men_n668_), .B(men_men_n91_), .Y(men_men_n676_));
  NA2        u0654(.A(men_men_n671_), .B(men_men_n273_), .Y(men_men_n677_));
  NO2        u0655(.A(i_11_), .B(men_men_n37_), .Y(men_men_n678_));
  NA2        u0656(.A(men_men_n678_), .B(men_men_n24_), .Y(men_men_n679_));
  OAI210     u0657(.A0(men_men_n679_), .A1(men_men_n677_), .B0(men_men_n676_), .Y(men_men_n680_));
  OR3        u0658(.A(men_men_n680_), .B(men_men_n675_), .C(men_men_n673_), .Y(men_men_n681_));
  NO3        u0659(.A(men_men_n681_), .B(men_men_n667_), .C(men_men_n661_), .Y(men_men_n682_));
  NO2        u0660(.A(men_men_n243_), .B(men_men_n101_), .Y(men_men_n683_));
  NO2        u0661(.A(men_men_n683_), .B(men_men_n639_), .Y(men_men_n684_));
  NA2        u0662(.A(men_men_n684_), .B(i_1_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n685_), .B(men_men_n633_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n429_), .B(men_men_n86_), .Y(men_men_n687_));
  NA2        u0665(.A(men_men_n686_), .B(men_men_n46_), .Y(men_men_n688_));
  NA2        u0666(.A(i_3_), .B(men_men_n196_), .Y(men_men_n689_));
  NO2        u0667(.A(men_men_n689_), .B(men_men_n114_), .Y(men_men_n690_));
  AN2        u0668(.A(men_men_n690_), .B(men_men_n559_), .Y(men_men_n691_));
  NO2        u0669(.A(men_men_n239_), .B(men_men_n44_), .Y(men_men_n692_));
  NO3        u0670(.A(men_men_n692_), .B(men_men_n317_), .C(men_men_n244_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n117_), .B(men_men_n37_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n694_), .B(i_6_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n86_), .B(i_9_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n696_), .B(men_men_n63_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n697_), .B(men_men_n654_), .Y(men_men_n698_));
  NO4        u0676(.A(men_men_n698_), .B(men_men_n695_), .C(men_men_n693_), .D(i_4_), .Y(men_men_n699_));
  NA2        u0677(.A(i_1_), .B(i_3_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n468_), .B(men_men_n92_), .Y(men_men_n701_));
  AOI210     u0679(.A0(men_men_n692_), .A1(men_men_n592_), .B0(men_men_n701_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n702_), .B(men_men_n700_), .Y(men_men_n703_));
  NO3        u0681(.A(men_men_n703_), .B(men_men_n699_), .C(men_men_n691_), .Y(men_men_n704_));
  NA4        u0682(.A(men_men_n704_), .B(men_men_n688_), .C(men_men_n682_), .D(men_men_n656_), .Y(men_men_n705_));
  NO3        u0683(.A(men_men_n493_), .B(i_3_), .C(i_7_), .Y(men_men_n706_));
  NOi21      u0684(.An(men_men_n706_), .B(i_10_), .Y(men_men_n707_));
  OA210      u0685(.A0(men_men_n707_), .A1(men_men_n251_), .B0(men_men_n86_), .Y(men_men_n708_));
  NA2        u0686(.A(men_men_n381_), .B(men_men_n380_), .Y(men_men_n709_));
  NA3        u0687(.A(men_men_n500_), .B(men_men_n535_), .C(men_men_n46_), .Y(men_men_n710_));
  NO3        u0688(.A(men_men_n494_), .B(men_men_n625_), .C(men_men_n86_), .Y(men_men_n711_));
  NA2        u0689(.A(men_men_n711_), .B(men_men_n25_), .Y(men_men_n712_));
  NA3        u0690(.A(men_men_n162_), .B(men_men_n84_), .C(men_men_n86_), .Y(men_men_n713_));
  NA4        u0691(.A(men_men_n713_), .B(men_men_n712_), .C(men_men_n710_), .D(men_men_n709_), .Y(men_men_n714_));
  OAI210     u0692(.A0(men_men_n714_), .A1(men_men_n708_), .B0(i_1_), .Y(men_men_n715_));
  AOI210     u0693(.A0(men_men_n273_), .A1(men_men_n97_), .B0(i_1_), .Y(men_men_n716_));
  NO2        u0694(.A(men_men_n379_), .B(i_2_), .Y(men_men_n717_));
  NA2        u0695(.A(men_men_n717_), .B(men_men_n716_), .Y(men_men_n718_));
  AOI210     u0696(.A0(men_men_n718_), .A1(men_men_n715_), .B0(i_13_), .Y(men_men_n719_));
  OR2        u0697(.A(i_11_), .B(i_7_), .Y(men_men_n720_));
  NO2        u0698(.A(men_men_n54_), .B(i_12_), .Y(men_men_n721_));
  INV        u0699(.A(men_men_n721_), .Y(men_men_n722_));
  NO2        u0700(.A(men_men_n494_), .B(men_men_n24_), .Y(men_men_n723_));
  AOI220     u0701(.A0(men_men_n723_), .A1(men_men_n687_), .B0(men_men_n251_), .B1(men_men_n131_), .Y(men_men_n724_));
  OAI220     u0702(.A0(men_men_n724_), .A1(men_men_n41_), .B0(men_men_n722_), .B1(men_men_n92_), .Y(men_men_n725_));
  INV        u0703(.A(men_men_n725_), .Y(men_men_n726_));
  NA2        u0704(.A(men_men_n397_), .B(men_men_n671_), .Y(men_men_n727_));
  NO2        u0705(.A(men_men_n727_), .B(men_men_n249_), .Y(men_men_n728_));
  AOI210     u0706(.A0(men_men_n459_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n729_));
  NOi31      u0707(.An(men_men_n729_), .B(men_men_n616_), .C(men_men_n44_), .Y(men_men_n730_));
  NA2        u0708(.A(men_men_n127_), .B(i_13_), .Y(men_men_n731_));
  NO2        u0709(.A(men_men_n670_), .B(men_men_n114_), .Y(men_men_n732_));
  INV        u0710(.A(men_men_n732_), .Y(men_men_n733_));
  NO2        u0711(.A(men_men_n731_), .B(men_men_n716_), .Y(men_men_n734_));
  NA2        u0712(.A(men_men_n26_), .B(men_men_n196_), .Y(men_men_n735_));
  NA2        u0713(.A(men_men_n735_), .B(i_7_), .Y(men_men_n736_));
  NO3        u0714(.A(men_men_n494_), .B(men_men_n243_), .C(men_men_n86_), .Y(men_men_n737_));
  NA2        u0715(.A(men_men_n737_), .B(men_men_n736_), .Y(men_men_n738_));
  AOI220     u0716(.A0(men_men_n397_), .A1(men_men_n671_), .B0(men_men_n91_), .B1(men_men_n102_), .Y(men_men_n739_));
  OAI220     u0717(.A0(men_men_n739_), .A1(men_men_n620_), .B0(men_men_n738_), .B1(men_men_n635_), .Y(men_men_n740_));
  NO4        u0718(.A(men_men_n740_), .B(men_men_n734_), .C(men_men_n730_), .D(men_men_n728_), .Y(men_men_n741_));
  OR2        u0719(.A(i_11_), .B(i_6_), .Y(men_men_n742_));
  NA3        u0720(.A(men_men_n619_), .B(men_men_n735_), .C(i_7_), .Y(men_men_n743_));
  AOI210     u0721(.A0(men_men_n743_), .A1(men_men_n733_), .B0(men_men_n742_), .Y(men_men_n744_));
  NA3        u0722(.A(men_men_n423_), .B(men_men_n624_), .C(men_men_n97_), .Y(men_men_n745_));
  NA2        u0723(.A(men_men_n660_), .B(i_13_), .Y(men_men_n746_));
  NA2        u0724(.A(men_men_n102_), .B(men_men_n735_), .Y(men_men_n747_));
  NAi21      u0725(.An(i_11_), .B(i_12_), .Y(men_men_n748_));
  NOi41      u0726(.An(men_men_n110_), .B(men_men_n748_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n749_));
  NA2        u0727(.A(men_men_n749_), .B(men_men_n747_), .Y(men_men_n750_));
  NA3        u0728(.A(men_men_n750_), .B(men_men_n746_), .C(men_men_n745_), .Y(men_men_n751_));
  OAI210     u0729(.A0(men_men_n751_), .A1(men_men_n744_), .B0(men_men_n63_), .Y(men_men_n752_));
  NO2        u0730(.A(i_2_), .B(i_12_), .Y(men_men_n753_));
  NA2        u0731(.A(men_men_n378_), .B(men_men_n753_), .Y(men_men_n754_));
  NA2        u0732(.A(i_8_), .B(men_men_n25_), .Y(men_men_n755_));
  NO3        u0733(.A(men_men_n755_), .B(men_men_n395_), .C(men_men_n619_), .Y(men_men_n756_));
  OAI210     u0734(.A0(men_men_n756_), .A1(men_men_n380_), .B0(men_men_n378_), .Y(men_men_n757_));
  NO2        u0735(.A(men_men_n128_), .B(i_2_), .Y(men_men_n758_));
  NA2        u0736(.A(men_men_n758_), .B(men_men_n654_), .Y(men_men_n759_));
  NA3        u0737(.A(men_men_n759_), .B(men_men_n757_), .C(men_men_n754_), .Y(men_men_n760_));
  NA3        u0738(.A(men_men_n760_), .B(men_men_n45_), .C(men_men_n231_), .Y(men_men_n761_));
  NA4        u0739(.A(men_men_n761_), .B(men_men_n752_), .C(men_men_n741_), .D(men_men_n726_), .Y(men_men_n762_));
  OR4        u0740(.A(men_men_n762_), .B(men_men_n719_), .C(men_men_n705_), .D(men_men_n638_), .Y(men5));
  AOI210     u0741(.A0(men_men_n684_), .A1(men_men_n276_), .B0(men_men_n432_), .Y(men_men_n764_));
  AN2        u0742(.A(men_men_n24_), .B(i_10_), .Y(men_men_n765_));
  NA3        u0743(.A(men_men_n765_), .B(men_men_n753_), .C(men_men_n108_), .Y(men_men_n766_));
  NO2        u0744(.A(men_men_n620_), .B(i_11_), .Y(men_men_n767_));
  NA2        u0745(.A(men_men_n87_), .B(men_men_n767_), .Y(men_men_n768_));
  NA3        u0746(.A(men_men_n768_), .B(men_men_n766_), .C(men_men_n764_), .Y(men_men_n769_));
  NO3        u0747(.A(i_11_), .B(men_men_n243_), .C(i_13_), .Y(men_men_n770_));
  NO2        u0748(.A(men_men_n124_), .B(men_men_n23_), .Y(men_men_n771_));
  NA2        u0749(.A(i_12_), .B(i_8_), .Y(men_men_n772_));
  OAI210     u0750(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n772_), .Y(men_men_n773_));
  INV        u0751(.A(men_men_n458_), .Y(men_men_n774_));
  AOI220     u0752(.A0(men_men_n327_), .A1(men_men_n596_), .B0(men_men_n773_), .B1(men_men_n771_), .Y(men_men_n775_));
  INV        u0753(.A(men_men_n775_), .Y(men_men_n776_));
  NO2        u0754(.A(men_men_n776_), .B(men_men_n769_), .Y(men_men_n777_));
  INV        u0755(.A(men_men_n173_), .Y(men_men_n778_));
  INV        u0756(.A(men_men_n251_), .Y(men_men_n779_));
  OAI210     u0757(.A0(men_men_n717_), .A1(men_men_n460_), .B0(men_men_n110_), .Y(men_men_n780_));
  AOI210     u0758(.A0(men_men_n780_), .A1(men_men_n779_), .B0(men_men_n778_), .Y(men_men_n781_));
  NO2        u0759(.A(men_men_n468_), .B(men_men_n26_), .Y(men_men_n782_));
  NO2        u0760(.A(men_men_n782_), .B(men_men_n434_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(i_2_), .Y(men_men_n784_));
  INV        u0762(.A(men_men_n784_), .Y(men_men_n785_));
  AOI210     u0763(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n430_), .Y(men_men_n786_));
  AOI210     u0764(.A0(men_men_n786_), .A1(men_men_n785_), .B0(men_men_n781_), .Y(men_men_n787_));
  NO2        u0765(.A(men_men_n193_), .B(men_men_n125_), .Y(men_men_n788_));
  OAI210     u0766(.A0(men_men_n788_), .A1(men_men_n771_), .B0(i_2_), .Y(men_men_n789_));
  INV        u0767(.A(men_men_n174_), .Y(men_men_n790_));
  NO3        u0768(.A(men_men_n640_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n791_));
  AOI210     u0769(.A0(men_men_n790_), .A1(men_men_n87_), .B0(men_men_n791_), .Y(men_men_n792_));
  AOI210     u0770(.A0(men_men_n792_), .A1(men_men_n789_), .B0(men_men_n196_), .Y(men_men_n793_));
  OA210      u0771(.A0(men_men_n641_), .A1(men_men_n126_), .B0(i_13_), .Y(men_men_n794_));
  NA2        u0772(.A(men_men_n203_), .B(men_men_n206_), .Y(men_men_n795_));
  NA2        u0773(.A(men_men_n152_), .B(men_men_n617_), .Y(men_men_n796_));
  AOI210     u0774(.A0(men_men_n796_), .A1(men_men_n795_), .B0(men_men_n383_), .Y(men_men_n797_));
  AOI210     u0775(.A0(men_men_n213_), .A1(men_men_n148_), .B0(men_men_n535_), .Y(men_men_n798_));
  NA2        u0776(.A(men_men_n798_), .B(men_men_n434_), .Y(men_men_n799_));
  NO2        u0777(.A(men_men_n102_), .B(men_men_n44_), .Y(men_men_n800_));
  INV        u0778(.A(men_men_n310_), .Y(men_men_n801_));
  NA4        u0779(.A(men_men_n801_), .B(men_men_n314_), .C(men_men_n124_), .D(men_men_n42_), .Y(men_men_n802_));
  OAI210     u0780(.A0(men_men_n802_), .A1(men_men_n800_), .B0(men_men_n799_), .Y(men_men_n803_));
  NO4        u0781(.A(men_men_n803_), .B(men_men_n797_), .C(men_men_n794_), .D(men_men_n793_), .Y(men_men_n804_));
  NA2        u0782(.A(men_men_n596_), .B(men_men_n28_), .Y(men_men_n805_));
  NA2        u0783(.A(men_men_n770_), .B(men_men_n283_), .Y(men_men_n806_));
  NA2        u0784(.A(men_men_n806_), .B(men_men_n805_), .Y(men_men_n807_));
  NO2        u0785(.A(men_men_n62_), .B(i_12_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n808_), .B(men_men_n126_), .Y(men_men_n809_));
  NO2        u0787(.A(men_men_n809_), .B(men_men_n617_), .Y(men_men_n810_));
  AOI220     u0788(.A0(men_men_n810_), .A1(men_men_n36_), .B0(men_men_n807_), .B1(men_men_n46_), .Y(men_men_n811_));
  NA4        u0789(.A(men_men_n811_), .B(men_men_n804_), .C(men_men_n787_), .D(men_men_n777_), .Y(men6));
  NO3        u0790(.A(men_men_n261_), .B(men_men_n316_), .C(i_1_), .Y(men_men_n813_));
  NO2        u0791(.A(men_men_n188_), .B(men_men_n139_), .Y(men_men_n814_));
  OAI210     u0792(.A0(men_men_n814_), .A1(men_men_n813_), .B0(men_men_n758_), .Y(men_men_n815_));
  NA4        u0793(.A(men_men_n401_), .B(men_men_n499_), .C(men_men_n71_), .D(men_men_n101_), .Y(men_men_n816_));
  INV        u0794(.A(men_men_n816_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n226_), .B(men_men_n503_), .Y(men_men_n818_));
  NO2        u0796(.A(men_men_n817_), .B(men_men_n339_), .Y(men_men_n819_));
  AO210      u0797(.A0(men_men_n819_), .A1(men_men_n815_), .B0(i_12_), .Y(men_men_n820_));
  NA2        u0798(.A(men_men_n602_), .B(men_men_n63_), .Y(men_men_n821_));
  NA2        u0799(.A(men_men_n707_), .B(men_men_n71_), .Y(men_men_n822_));
  NA2        u0800(.A(men_men_n822_), .B(men_men_n821_), .Y(men_men_n823_));
  NA2        u0801(.A(men_men_n823_), .B(men_men_n73_), .Y(men_men_n824_));
  INV        u0802(.A(men_men_n338_), .Y(men_men_n825_));
  NA2        u0803(.A(men_men_n75_), .B(men_men_n131_), .Y(men_men_n826_));
  INV        u0804(.A(men_men_n124_), .Y(men_men_n827_));
  NA2        u0805(.A(men_men_n827_), .B(men_men_n46_), .Y(men_men_n828_));
  AOI210     u0806(.A0(men_men_n828_), .A1(men_men_n826_), .B0(men_men_n825_), .Y(men_men_n829_));
  NO2        u0807(.A(men_men_n258_), .B(i_9_), .Y(men_men_n830_));
  NA2        u0808(.A(men_men_n830_), .B(men_men_n808_), .Y(men_men_n831_));
  AOI210     u0809(.A0(men_men_n831_), .A1(men_men_n533_), .B0(men_men_n188_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n32_), .B(i_11_), .Y(men_men_n833_));
  NA3        u0811(.A(men_men_n833_), .B(men_men_n489_), .C(men_men_n401_), .Y(men_men_n834_));
  NAi32      u0812(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n835_));
  NO2        u0813(.A(men_men_n742_), .B(men_men_n835_), .Y(men_men_n836_));
  OAI210     u0814(.A0(men_men_n706_), .A1(men_men_n584_), .B0(men_men_n583_), .Y(men_men_n837_));
  NAi31      u0815(.An(men_men_n836_), .B(men_men_n837_), .C(men_men_n834_), .Y(men_men_n838_));
  OR3        u0816(.A(men_men_n838_), .B(men_men_n832_), .C(men_men_n829_), .Y(men_men_n839_));
  NO2        u0817(.A(men_men_n720_), .B(i_2_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n841_));
  NO2        u0819(.A(men_men_n841_), .B(men_men_n422_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n842_), .B(men_men_n840_), .Y(men_men_n843_));
  AO210      u0821(.A0(men_men_n372_), .A1(men_men_n364_), .B0(men_men_n409_), .Y(men_men_n844_));
  NA3        u0822(.A(men_men_n844_), .B(men_men_n262_), .C(i_7_), .Y(men_men_n845_));
  BUFFER     u0823(.A(men_men_n641_), .Y(men_men_n846_));
  NA3        u0824(.A(men_men_n846_), .B(men_men_n147_), .C(men_men_n69_), .Y(men_men_n847_));
  AO210      u0825(.A0(men_men_n509_), .A1(men_men_n774_), .B0(men_men_n36_), .Y(men_men_n848_));
  NA4        u0826(.A(men_men_n848_), .B(men_men_n847_), .C(men_men_n845_), .D(men_men_n843_), .Y(men_men_n849_));
  NO2        u0827(.A(men_men_n659_), .B(i_11_), .Y(men_men_n850_));
  AOI220     u0828(.A0(men_men_n850_), .A1(men_men_n583_), .B0(men_men_n818_), .B1(men_men_n736_), .Y(men_men_n851_));
  NA3        u0829(.A(men_men_n383_), .B(men_men_n245_), .C(men_men_n147_), .Y(men_men_n852_));
  NA2        u0830(.A(men_men_n409_), .B(men_men_n70_), .Y(men_men_n853_));
  NA4        u0831(.A(men_men_n853_), .B(men_men_n852_), .C(men_men_n851_), .D(men_men_n623_), .Y(men_men_n854_));
  AOI210     u0832(.A0(men_men_n460_), .A1(men_men_n458_), .B0(men_men_n582_), .Y(men_men_n855_));
  NA2        u0833(.A(men_men_n111_), .B(men_men_n420_), .Y(men_men_n856_));
  NA2        u0834(.A(men_men_n250_), .B(men_men_n46_), .Y(men_men_n857_));
  INV        u0835(.A(men_men_n608_), .Y(men_men_n858_));
  NA3        u0836(.A(men_men_n858_), .B(men_men_n338_), .C(i_7_), .Y(men_men_n859_));
  NA3        u0837(.A(men_men_n859_), .B(men_men_n856_), .C(men_men_n855_), .Y(men_men_n860_));
  NO4        u0838(.A(men_men_n860_), .B(men_men_n854_), .C(men_men_n849_), .D(men_men_n839_), .Y(men_men_n861_));
  NA4        u0839(.A(men_men_n861_), .B(men_men_n824_), .C(men_men_n820_), .D(men_men_n391_), .Y(men3));
  NA2        u0840(.A(i_12_), .B(i_10_), .Y(men_men_n863_));
  NA2        u0841(.A(i_6_), .B(i_7_), .Y(men_men_n864_));
  NO2        u0842(.A(men_men_n864_), .B(i_0_), .Y(men_men_n865_));
  NO2        u0843(.A(i_11_), .B(men_men_n243_), .Y(men_men_n866_));
  OAI210     u0844(.A0(men_men_n865_), .A1(men_men_n298_), .B0(men_men_n866_), .Y(men_men_n867_));
  NO2        u0845(.A(men_men_n867_), .B(men_men_n196_), .Y(men_men_n868_));
  NO3        u0846(.A(men_men_n464_), .B(men_men_n89_), .C(men_men_n44_), .Y(men_men_n869_));
  OA210      u0847(.A0(men_men_n869_), .A1(men_men_n868_), .B0(men_men_n176_), .Y(men_men_n870_));
  NA3        u0848(.A(men_men_n852_), .B(men_men_n623_), .C(men_men_n382_), .Y(men_men_n871_));
  NA2        u0849(.A(men_men_n871_), .B(men_men_n40_), .Y(men_men_n872_));
  NO3        u0850(.A(men_men_n649_), .B(men_men_n468_), .C(men_men_n131_), .Y(men_men_n873_));
  AN2        u0851(.A(men_men_n466_), .B(men_men_n55_), .Y(men_men_n874_));
  NO2        u0852(.A(men_men_n874_), .B(men_men_n873_), .Y(men_men_n875_));
  AOI210     u0853(.A0(men_men_n875_), .A1(men_men_n872_), .B0(men_men_n48_), .Y(men_men_n876_));
  NO4        u0854(.A(men_men_n387_), .B(men_men_n394_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n877_));
  NA2        u0855(.A(men_men_n188_), .B(men_men_n592_), .Y(men_men_n878_));
  NOi21      u0856(.An(men_men_n878_), .B(men_men_n877_), .Y(men_men_n879_));
  NA2        u0857(.A(men_men_n729_), .B(men_men_n696_), .Y(men_men_n880_));
  NA2        u0858(.A(men_men_n344_), .B(men_men_n452_), .Y(men_men_n881_));
  OAI220     u0859(.A0(men_men_n881_), .A1(men_men_n880_), .B0(men_men_n879_), .B1(men_men_n63_), .Y(men_men_n882_));
  NOi21      u0860(.An(i_5_), .B(i_9_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n883_), .B(men_men_n457_), .Y(men_men_n884_));
  AOI210     u0862(.A0(men_men_n273_), .A1(men_men_n491_), .B0(men_men_n711_), .Y(men_men_n885_));
  NO3        u0863(.A(men_men_n426_), .B(men_men_n273_), .C(men_men_n73_), .Y(men_men_n886_));
  NO2        u0864(.A(men_men_n177_), .B(men_men_n148_), .Y(men_men_n887_));
  AOI210     u0865(.A0(men_men_n887_), .A1(men_men_n250_), .B0(men_men_n886_), .Y(men_men_n888_));
  OAI220     u0866(.A0(men_men_n888_), .A1(men_men_n183_), .B0(men_men_n885_), .B1(men_men_n884_), .Y(men_men_n889_));
  NO4        u0867(.A(men_men_n889_), .B(men_men_n882_), .C(men_men_n876_), .D(men_men_n870_), .Y(men_men_n890_));
  NA2        u0868(.A(men_men_n188_), .B(men_men_n24_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n321_), .B(men_men_n129_), .Y(men_men_n892_));
  NAi21      u0870(.An(men_men_n163_), .B(men_men_n452_), .Y(men_men_n893_));
  OAI220     u0871(.A0(men_men_n893_), .A1(men_men_n857_), .B0(men_men_n892_), .B1(men_men_n411_), .Y(men_men_n894_));
  INV        u0872(.A(men_men_n894_), .Y(men_men_n895_));
  NO2        u0873(.A(men_men_n401_), .B(men_men_n302_), .Y(men_men_n896_));
  NA2        u0874(.A(men_men_n896_), .B(men_men_n732_), .Y(men_men_n897_));
  NA2        u0875(.A(men_men_n593_), .B(i_0_), .Y(men_men_n898_));
  NO3        u0876(.A(men_men_n898_), .B(men_men_n396_), .C(men_men_n87_), .Y(men_men_n899_));
  INV        u0877(.A(men_men_n899_), .Y(men_men_n900_));
  INV        u0878(.A(men_men_n489_), .Y(men_men_n901_));
  NA2        u0879(.A(men_men_n770_), .B(men_men_n339_), .Y(men_men_n902_));
  INV        u0880(.A(men_men_n58_), .Y(men_men_n903_));
  OAI220     u0881(.A0(men_men_n903_), .A1(men_men_n902_), .B0(men_men_n679_), .B1(men_men_n555_), .Y(men_men_n904_));
  NO2        u0882(.A(men_men_n260_), .B(men_men_n154_), .Y(men_men_n905_));
  NA2        u0883(.A(i_0_), .B(i_10_), .Y(men_men_n906_));
  OAI210     u0884(.A0(men_men_n906_), .A1(men_men_n86_), .B0(men_men_n558_), .Y(men_men_n907_));
  NO4        u0885(.A(men_men_n114_), .B(men_men_n58_), .C(men_men_n689_), .D(i_5_), .Y(men_men_n908_));
  AO220      u0886(.A0(men_men_n908_), .A1(men_men_n907_), .B0(men_men_n905_), .B1(i_6_), .Y(men_men_n909_));
  AOI220     u0887(.A0(men_men_n344_), .A1(men_men_n98_), .B0(men_men_n188_), .B1(men_men_n84_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n587_), .B(i_4_), .Y(men_men_n911_));
  NA2        u0889(.A(men_men_n191_), .B(men_men_n206_), .Y(men_men_n912_));
  OAI220     u0890(.A0(men_men_n912_), .A1(men_men_n902_), .B0(men_men_n911_), .B1(men_men_n910_), .Y(men_men_n913_));
  NO3        u0891(.A(men_men_n913_), .B(men_men_n909_), .C(men_men_n904_), .Y(men_men_n914_));
  NA4        u0892(.A(men_men_n914_), .B(men_men_n900_), .C(men_men_n897_), .D(men_men_n895_), .Y(men_men_n915_));
  NO2        u0893(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n916_));
  NA2        u0894(.A(i_11_), .B(i_9_), .Y(men_men_n917_));
  NO3        u0895(.A(i_12_), .B(men_men_n917_), .C(men_men_n622_), .Y(men_men_n918_));
  AN2        u0896(.A(men_men_n918_), .B(men_men_n916_), .Y(men_men_n919_));
  NO2        u0897(.A(men_men_n48_), .B(i_7_), .Y(men_men_n920_));
  NA2        u0898(.A(men_men_n406_), .B(men_men_n181_), .Y(men_men_n921_));
  NA2        u0899(.A(men_men_n921_), .B(men_men_n161_), .Y(men_men_n922_));
  NO2        u0900(.A(men_men_n917_), .B(men_men_n73_), .Y(men_men_n923_));
  NO2        u0901(.A(men_men_n177_), .B(i_0_), .Y(men_men_n924_));
  INV        u0902(.A(men_men_n924_), .Y(men_men_n925_));
  NA2        u0903(.A(men_men_n489_), .B(men_men_n237_), .Y(men_men_n926_));
  INV        u0904(.A(men_men_n419_), .Y(men_men_n927_));
  OAI220     u0905(.A0(men_men_n927_), .A1(men_men_n884_), .B0(men_men_n926_), .B1(men_men_n925_), .Y(men_men_n928_));
  NO3        u0906(.A(men_men_n928_), .B(men_men_n922_), .C(men_men_n919_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n678_), .B(men_men_n121_), .Y(men_men_n930_));
  NO2        u0908(.A(i_6_), .B(men_men_n930_), .Y(men_men_n931_));
  AOI210     u0909(.A0(men_men_n459_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n932_));
  NA2        u0910(.A(men_men_n173_), .B(men_men_n103_), .Y(men_men_n933_));
  NOi32      u0911(.An(men_men_n932_), .Bn(men_men_n191_), .C(men_men_n933_), .Y(men_men_n934_));
  NO2        u0912(.A(men_men_n934_), .B(men_men_n931_), .Y(men_men_n935_));
  NOi21      u0913(.An(i_7_), .B(i_5_), .Y(men_men_n936_));
  NOi31      u0914(.An(men_men_n936_), .B(i_0_), .C(men_men_n748_), .Y(men_men_n937_));
  NA3        u0915(.A(men_men_n937_), .B(men_men_n395_), .C(i_6_), .Y(men_men_n938_));
  OA210      u0916(.A0(men_men_n933_), .A1(men_men_n533_), .B0(men_men_n938_), .Y(men_men_n939_));
  NO3        u0917(.A(men_men_n414_), .B(men_men_n375_), .C(men_men_n371_), .Y(men_men_n940_));
  NO2        u0918(.A(men_men_n267_), .B(men_men_n328_), .Y(men_men_n941_));
  NO2        u0919(.A(men_men_n748_), .B(men_men_n264_), .Y(men_men_n942_));
  AOI210     u0920(.A0(men_men_n942_), .A1(men_men_n941_), .B0(men_men_n940_), .Y(men_men_n943_));
  NA4        u0921(.A(men_men_n943_), .B(men_men_n939_), .C(men_men_n935_), .D(men_men_n929_), .Y(men_men_n944_));
  NO2        u0922(.A(men_men_n891_), .B(men_men_n246_), .Y(men_men_n945_));
  AN2        u0923(.A(men_men_n343_), .B(men_men_n339_), .Y(men_men_n946_));
  AN2        u0924(.A(men_men_n946_), .B(men_men_n887_), .Y(men_men_n947_));
  OAI210     u0925(.A0(men_men_n947_), .A1(men_men_n945_), .B0(i_10_), .Y(men_men_n948_));
  NO2        u0926(.A(men_men_n863_), .B(men_men_n327_), .Y(men_men_n949_));
  NA2        u0927(.A(men_men_n949_), .B(men_men_n923_), .Y(men_men_n950_));
  NA3        u0928(.A(men_men_n488_), .B(men_men_n423_), .C(men_men_n45_), .Y(men_men_n951_));
  OAI210     u0929(.A0(men_men_n893_), .A1(men_men_n901_), .B0(men_men_n951_), .Y(men_men_n952_));
  NO2        u0930(.A(men_men_n262_), .B(men_men_n46_), .Y(men_men_n953_));
  NO2        u0931(.A(men_men_n953_), .B(men_men_n190_), .Y(men_men_n954_));
  AOI220     u0932(.A0(men_men_n954_), .A1(men_men_n489_), .B0(men_men_n952_), .B1(men_men_n73_), .Y(men_men_n955_));
  NA3        u0933(.A(men_men_n841_), .B(men_men_n393_), .C(men_men_n659_), .Y(men_men_n956_));
  NA2        u0934(.A(men_men_n92_), .B(men_men_n44_), .Y(men_men_n957_));
  NO2        u0935(.A(men_men_n75_), .B(men_men_n772_), .Y(men_men_n958_));
  AOI220     u0936(.A0(men_men_n958_), .A1(men_men_n957_), .B0(men_men_n176_), .B1(men_men_n615_), .Y(men_men_n959_));
  AOI210     u0937(.A0(men_men_n959_), .A1(men_men_n956_), .B0(men_men_n47_), .Y(men_men_n960_));
  NA2        u0938(.A(men_men_n723_), .B(men_men_n567_), .Y(men_men_n961_));
  NO2        u0939(.A(men_men_n618_), .B(men_men_n105_), .Y(men_men_n962_));
  NA2        u0940(.A(men_men_n962_), .B(i_0_), .Y(men_men_n963_));
  OAI220     u0941(.A0(men_men_n963_), .A1(men_men_n86_), .B0(men_men_n961_), .B1(men_men_n174_), .Y(men_men_n964_));
  NO3        u0942(.A(men_men_n964_), .B(men_men_n960_), .C(men_men_n537_), .Y(men_men_n965_));
  NA4        u0943(.A(men_men_n965_), .B(men_men_n955_), .C(men_men_n950_), .D(men_men_n948_), .Y(men_men_n966_));
  NO3        u0944(.A(men_men_n966_), .B(men_men_n944_), .C(men_men_n915_), .Y(men_men_n967_));
  NO2        u0945(.A(i_0_), .B(men_men_n748_), .Y(men_men_n968_));
  NA2        u0946(.A(men_men_n73_), .B(men_men_n44_), .Y(men_men_n969_));
  NA2        u0947(.A(men_men_n906_), .B(men_men_n969_), .Y(men_men_n970_));
  NO3        u0948(.A(men_men_n105_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n971_));
  AO220      u0949(.A0(men_men_n971_), .A1(men_men_n970_), .B0(men_men_n968_), .B1(men_men_n176_), .Y(men_men_n972_));
  AOI210     u0950(.A0(men_men_n821_), .A1(men_men_n709_), .B0(men_men_n933_), .Y(men_men_n973_));
  AOI210     u0951(.A0(men_men_n972_), .A1(men_men_n361_), .B0(men_men_n973_), .Y(men_men_n974_));
  NA2        u0952(.A(men_men_n758_), .B(men_men_n146_), .Y(men_men_n975_));
  INV        u0953(.A(men_men_n975_), .Y(men_men_n976_));
  NA3        u0954(.A(men_men_n976_), .B(men_men_n696_), .C(men_men_n73_), .Y(men_men_n977_));
  NO2        u0955(.A(men_men_n837_), .B(men_men_n414_), .Y(men_men_n978_));
  NA3        u0956(.A(men_men_n865_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n866_), .B(i_9_), .Y(men_men_n980_));
  AOI210     u0958(.A0(men_men_n979_), .A1(men_men_n515_), .B0(men_men_n980_), .Y(men_men_n981_));
  NA2        u0959(.A(men_men_n250_), .B(men_men_n236_), .Y(men_men_n982_));
  AOI210     u0960(.A0(men_men_n982_), .A1(men_men_n898_), .B0(men_men_n154_), .Y(men_men_n983_));
  NO3        u0961(.A(men_men_n983_), .B(men_men_n981_), .C(men_men_n978_), .Y(men_men_n984_));
  NA3        u0962(.A(men_men_n984_), .B(men_men_n977_), .C(men_men_n974_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n946_), .B(men_men_n383_), .Y(men_men_n986_));
  AOI210     u0964(.A0(men_men_n309_), .A1(men_men_n163_), .B0(men_men_n986_), .Y(men_men_n987_));
  NA3        u0965(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n988_));
  NA2        u0966(.A(men_men_n920_), .B(men_men_n504_), .Y(men_men_n989_));
  AOI210     u0967(.A0(men_men_n988_), .A1(men_men_n163_), .B0(men_men_n989_), .Y(men_men_n990_));
  NO2        u0968(.A(men_men_n990_), .B(men_men_n987_), .Y(men_men_n991_));
  NO3        u0969(.A(men_men_n906_), .B(men_men_n883_), .C(men_men_n193_), .Y(men_men_n992_));
  AOI220     u0970(.A0(men_men_n992_), .A1(i_11_), .B0(men_men_n588_), .B1(men_men_n75_), .Y(men_men_n993_));
  NO3        u0971(.A(men_men_n214_), .B(men_men_n394_), .C(i_0_), .Y(men_men_n994_));
  OAI210     u0972(.A0(men_men_n994_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n995_));
  INV        u0973(.A(men_men_n223_), .Y(men_men_n996_));
  OAI220     u0974(.A0(men_men_n548_), .A1(men_men_n139_), .B0(men_men_n664_), .B1(men_men_n635_), .Y(men_men_n997_));
  NA3        u0975(.A(men_men_n997_), .B(i_7_), .C(men_men_n996_), .Y(men_men_n998_));
  NA4        u0976(.A(men_men_n998_), .B(men_men_n995_), .C(men_men_n993_), .D(men_men_n991_), .Y(men_men_n999_));
  NO2        u0977(.A(men_men_n249_), .B(men_men_n92_), .Y(men_men_n1000_));
  NA2        u0978(.A(men_men_n1000_), .B(men_men_n968_), .Y(men_men_n1001_));
  AOI220     u0979(.A0(men_men_n936_), .A1(men_men_n504_), .B0(men_men_n865_), .B1(men_men_n164_), .Y(men_men_n1002_));
  NA2        u0980(.A(men_men_n364_), .B(men_men_n178_), .Y(men_men_n1003_));
  OA220      u0981(.A0(men_men_n1003_), .A1(men_men_n1002_), .B0(men_men_n1001_), .B1(i_5_), .Y(men_men_n1004_));
  AOI210     u0982(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n177_), .Y(men_men_n1005_));
  NA3        u0983(.A(men_men_n632_), .B(men_men_n188_), .C(men_men_n84_), .Y(men_men_n1006_));
  NA2        u0984(.A(men_men_n1006_), .B(men_men_n565_), .Y(men_men_n1007_));
  INV        u0985(.A(men_men_n486_), .Y(men_men_n1008_));
  NO2        u0986(.A(men_men_n1008_), .B(men_men_n1007_), .Y(men_men_n1009_));
  NA3        u0987(.A(men_men_n401_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n1010_));
  NA3        u0988(.A(men_men_n401_), .B(men_men_n345_), .C(men_men_n227_), .Y(men_men_n1011_));
  INV        u0989(.A(men_men_n1011_), .Y(men_men_n1012_));
  NOi31      u0990(.An(men_men_n400_), .B(men_men_n969_), .C(men_men_n246_), .Y(men_men_n1013_));
  NO3        u0991(.A(men_men_n917_), .B(men_men_n223_), .C(men_men_n193_), .Y(men_men_n1014_));
  NO4        u0992(.A(men_men_n1014_), .B(men_men_n1013_), .C(men_men_n1012_), .D(men_men_n1081_), .Y(men_men_n1015_));
  NA3        u0993(.A(men_men_n1015_), .B(men_men_n1009_), .C(men_men_n1004_), .Y(men_men_n1016_));
  INV        u0994(.A(men_men_n634_), .Y(men_men_n1017_));
  NO3        u0995(.A(men_men_n1017_), .B(men_men_n580_), .C(men_men_n358_), .Y(men_men_n1018_));
  NO2        u0996(.A(men_men_n86_), .B(i_5_), .Y(men_men_n1019_));
  NA3        u0997(.A(men_men_n866_), .B(men_men_n109_), .C(men_men_n124_), .Y(men_men_n1020_));
  INV        u0998(.A(men_men_n1020_), .Y(men_men_n1021_));
  AOI210     u0999(.A0(men_men_n1021_), .A1(men_men_n1019_), .B0(men_men_n1018_), .Y(men_men_n1022_));
  NA3        u1000(.A(men_men_n314_), .B(i_5_), .C(men_men_n196_), .Y(men_men_n1023_));
  NAi31      u1001(.An(men_men_n248_), .B(men_men_n1023_), .C(men_men_n249_), .Y(men_men_n1024_));
  NO4        u1002(.A(men_men_n246_), .B(men_men_n214_), .C(i_0_), .D(i_12_), .Y(men_men_n1025_));
  AOI220     u1003(.A0(men_men_n1025_), .A1(men_men_n1024_), .B0(men_men_n817_), .B1(men_men_n178_), .Y(men_men_n1026_));
  AN2        u1004(.A(men_men_n906_), .B(men_men_n154_), .Y(men_men_n1027_));
  NO4        u1005(.A(men_men_n1027_), .B(i_12_), .C(men_men_n668_), .D(men_men_n131_), .Y(men_men_n1028_));
  NA2        u1006(.A(men_men_n1028_), .B(men_men_n223_), .Y(men_men_n1029_));
  NA3        u1007(.A(men_men_n98_), .B(men_men_n592_), .C(i_11_), .Y(men_men_n1030_));
  NO2        u1008(.A(men_men_n1030_), .B(men_men_n156_), .Y(men_men_n1031_));
  NA2        u1009(.A(men_men_n936_), .B(men_men_n485_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n64_), .B(men_men_n101_), .Y(men_men_n1033_));
  OAI220     u1011(.A0(men_men_n1033_), .A1(men_men_n1023_), .B0(men_men_n1032_), .B1(men_men_n697_), .Y(men_men_n1034_));
  AOI210     u1012(.A0(men_men_n1034_), .A1(men_men_n924_), .B0(men_men_n1031_), .Y(men_men_n1035_));
  NA4        u1013(.A(men_men_n1035_), .B(men_men_n1029_), .C(men_men_n1026_), .D(men_men_n1022_), .Y(men_men_n1036_));
  NO4        u1014(.A(men_men_n1036_), .B(men_men_n1016_), .C(men_men_n999_), .D(men_men_n985_), .Y(men_men_n1037_));
  OAI210     u1015(.A0(men_men_n840_), .A1(men_men_n833_), .B0(men_men_n37_), .Y(men_men_n1038_));
  NA3        u1016(.A(men_men_n932_), .B(men_men_n378_), .C(i_5_), .Y(men_men_n1039_));
  NA3        u1017(.A(men_men_n1039_), .B(men_men_n1038_), .C(men_men_n630_), .Y(men_men_n1040_));
  NA2        u1018(.A(men_men_n1040_), .B(men_men_n211_), .Y(men_men_n1041_));
  NA2        u1019(.A(men_men_n189_), .B(men_men_n191_), .Y(men_men_n1042_));
  AO210      u1020(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n1042_), .Y(men_men_n1043_));
  OAI210     u1021(.A0(men_men_n634_), .A1(men_men_n632_), .B0(men_men_n327_), .Y(men_men_n1044_));
  INV        u1022(.A(men_men_n665_), .Y(men_men_n1045_));
  NA3        u1023(.A(men_men_n1045_), .B(men_men_n1044_), .C(men_men_n1043_), .Y(men_men_n1046_));
  NO2        u1024(.A(men_men_n476_), .B(men_men_n273_), .Y(men_men_n1047_));
  NO4        u1025(.A(men_men_n239_), .B(men_men_n145_), .C(men_men_n700_), .D(men_men_n37_), .Y(men_men_n1048_));
  NO2        u1026(.A(men_men_n1048_), .B(men_men_n1047_), .Y(men_men_n1049_));
  OAI210     u1027(.A0(men_men_n1030_), .A1(men_men_n148_), .B0(men_men_n1049_), .Y(men_men_n1050_));
  AOI210     u1028(.A0(men_men_n1046_), .A1(men_men_n48_), .B0(men_men_n1050_), .Y(men_men_n1051_));
  AOI210     u1029(.A0(men_men_n1051_), .A1(men_men_n1041_), .B0(men_men_n73_), .Y(men_men_n1052_));
  NO2        u1030(.A(men_men_n585_), .B(men_men_n390_), .Y(men_men_n1053_));
  NO2        u1031(.A(men_men_n1053_), .B(men_men_n778_), .Y(men_men_n1054_));
  INV        u1032(.A(men_men_n76_), .Y(men_men_n1055_));
  AOI210     u1033(.A0(men_men_n1005_), .A1(men_men_n920_), .B0(men_men_n937_), .Y(men_men_n1056_));
  AOI210     u1034(.A0(men_men_n1056_), .A1(men_men_n1055_), .B0(men_men_n700_), .Y(men_men_n1057_));
  NA2        u1035(.A(men_men_n267_), .B(men_men_n57_), .Y(men_men_n1058_));
  AOI220     u1036(.A0(men_men_n1058_), .A1(men_men_n76_), .B0(men_men_n359_), .B1(men_men_n261_), .Y(men_men_n1059_));
  NO2        u1037(.A(men_men_n1059_), .B(men_men_n243_), .Y(men_men_n1060_));
  NA3        u1038(.A(men_men_n96_), .B(men_men_n316_), .C(men_men_n31_), .Y(men_men_n1061_));
  INV        u1039(.A(men_men_n1061_), .Y(men_men_n1062_));
  NO3        u1040(.A(men_men_n1062_), .B(men_men_n1060_), .C(men_men_n1057_), .Y(men_men_n1063_));
  OAI210     u1041(.A0(men_men_n275_), .A1(men_men_n159_), .B0(men_men_n87_), .Y(men_men_n1064_));
  NA3        u1042(.A(men_men_n782_), .B(men_men_n298_), .C(men_men_n80_), .Y(men_men_n1065_));
  AOI210     u1043(.A0(men_men_n1065_), .A1(men_men_n1064_), .B0(i_11_), .Y(men_men_n1066_));
  NA2        u1044(.A(men_men_n625_), .B(men_men_n220_), .Y(men_men_n1067_));
  OAI210     u1045(.A0(men_men_n1067_), .A1(men_men_n932_), .B0(men_men_n211_), .Y(men_men_n1068_));
  NA2        u1046(.A(men_men_n165_), .B(i_5_), .Y(men_men_n1069_));
  NO2        u1047(.A(men_men_n1068_), .B(men_men_n1069_), .Y(men_men_n1070_));
  NO3        u1048(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1071_));
  OAI210     u1049(.A0(men_men_n941_), .A1(men_men_n316_), .B0(men_men_n1071_), .Y(men_men_n1072_));
  NO2        u1050(.A(men_men_n1072_), .B(men_men_n748_), .Y(men_men_n1073_));
  NO3        u1051(.A(men_men_n1073_), .B(men_men_n1070_), .C(men_men_n1066_), .Y(men_men_n1074_));
  OAI210     u1052(.A0(men_men_n1063_), .A1(i_4_), .B0(men_men_n1074_), .Y(men_men_n1075_));
  NO3        u1053(.A(men_men_n1075_), .B(men_men_n1054_), .C(men_men_n1052_), .Y(men_men_n1076_));
  NA4        u1054(.A(men_men_n1076_), .B(men_men_n1037_), .C(men_men_n967_), .D(men_men_n890_), .Y(men4));
  INV        u1055(.A(i_2_), .Y(men_men_n1080_));
  INV        u1056(.A(men_men_n1010_), .Y(men_men_n1081_));
  INV        u1057(.A(i_12_), .Y(men_men_n1082_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule