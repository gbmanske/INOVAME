//Benchmark atmr_max1024_476_0.125

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n426_, mai_mai_n427_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n439_, men_men_n440_, men_men_n441_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n60_));
  INV        o044(.A(x9), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n60_), .B(x5), .Y(ori_ori_n62_));
  OAI210     o046(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n63_));
  OAI210     o047(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n63_), .Y(ori_ori_n64_));
  INV        o048(.A(ori_ori_n64_), .Y(ori_ori_n65_));
  NA2        o049(.A(ori_ori_n65_), .B(x4), .Y(ori_ori_n66_));
  NA2        o050(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n67_));
  OAI210     o051(.A0(ori_ori_n67_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n68_));
  NA2        o052(.A(x5), .B(x3), .Y(ori_ori_n69_));
  NO2        o053(.A(x8), .B(x6), .Y(ori_ori_n70_));
  NO3        o054(.A(ori_ori_n70_), .B(ori_ori_n69_), .C(ori_ori_n54_), .Y(ori_ori_n71_));
  NAi21      o055(.An(x4), .B(x3), .Y(ori_ori_n72_));
  INV        o056(.A(ori_ori_n72_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n22_), .Y(ori_ori_n74_));
  NO2        o058(.A(x4), .B(x2), .Y(ori_ori_n75_));
  NO2        o059(.A(ori_ori_n75_), .B(x3), .Y(ori_ori_n76_));
  NO3        o060(.A(ori_ori_n76_), .B(ori_ori_n74_), .C(ori_ori_n18_), .Y(ori_ori_n77_));
  NO3        o061(.A(ori_ori_n77_), .B(ori_ori_n71_), .C(ori_ori_n68_), .Y(ori_ori_n78_));
  NA2        o062(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n25_), .Y(ori_ori_n80_));
  INV        o064(.A(x8), .Y(ori_ori_n81_));
  NA2        o065(.A(x2), .B(x1), .Y(ori_ori_n82_));
  INV        o066(.A(ori_ori_n80_), .Y(ori_ori_n83_));
  NO2        o067(.A(ori_ori_n83_), .B(ori_ori_n26_), .Y(ori_ori_n84_));
  AOI210     o068(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n85_));
  OAI210     o069(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n86_));
  NO3        o070(.A(ori_ori_n86_), .B(ori_ori_n85_), .C(ori_ori_n84_), .Y(ori_ori_n87_));
  NA2        o071(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n89_));
  OAI210     o073(.A0(ori_ori_n89_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n88_), .A1(ori_ori_n52_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NO2        o075(.A(x3), .B(x2), .Y(ori_ori_n92_));
  NA3        o076(.A(ori_ori_n92_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n93_));
  AOI210     o077(.A0(x8), .A1(x6), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NA2        o078(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n95_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n96_));
  NO4        o080(.A(ori_ori_n96_), .B(ori_ori_n94_), .C(ori_ori_n91_), .D(ori_ori_n87_), .Y(ori_ori_n97_));
  AO210      o081(.A0(ori_ori_n78_), .A1(ori_ori_n66_), .B0(ori_ori_n97_), .Y(ori02));
  NO2        o082(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n99_));
  NO2        o083(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n101_));
  OR2        o085(.A(x8), .B(x0), .Y(ori_ori_n102_));
  INV        o086(.A(ori_ori_n102_), .Y(ori_ori_n103_));
  NAi21      o087(.An(x2), .B(x8), .Y(ori_ori_n104_));
  INV        o088(.A(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o089(.A(x4), .B(x1), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n106_), .B(x2), .Y(ori_ori_n107_));
  NOi21      o091(.An(x0), .B(x4), .Y(ori_ori_n108_));
  NO2        o092(.A(ori_ori_n107_), .B(ori_ori_n69_), .Y(ori_ori_n109_));
  NO2        o093(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n110_));
  NA2        o094(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n111_));
  AOI210     o095(.A0(ori_ori_n111_), .A1(ori_ori_n95_), .B0(ori_ori_n101_), .Y(ori_ori_n112_));
  OAI210     o096(.A0(ori_ori_n112_), .A1(ori_ori_n35_), .B0(ori_ori_n110_), .Y(ori_ori_n113_));
  NO2        o097(.A(x7), .B(x0), .Y(ori_ori_n114_));
  NO2        o098(.A(ori_ori_n75_), .B(ori_ori_n89_), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n115_), .B(x3), .Y(ori_ori_n116_));
  NA2        o100(.A(ori_ori_n114_), .B(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o101(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n118_));
  NA2        o102(.A(x5), .B(x0), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n120_));
  NA3        o104(.A(ori_ori_n120_), .B(ori_ori_n119_), .C(ori_ori_n118_), .Y(ori_ori_n121_));
  NA4        o105(.A(ori_ori_n121_), .B(ori_ori_n117_), .C(ori_ori_n113_), .D(ori_ori_n36_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n122_), .B(ori_ori_n109_), .Y(ori_ori_n123_));
  NO3        o107(.A(ori_ori_n69_), .B(ori_ori_n67_), .C(ori_ori_n24_), .Y(ori_ori_n124_));
  NO2        o108(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n125_));
  NA2        o109(.A(x7), .B(x3), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n88_), .B(x5), .Y(ori_ori_n127_));
  INV        o111(.A(x7), .Y(ori_ori_n128_));
  NOi21      o112(.An(x8), .B(x0), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n130_));
  INV        o114(.A(x7), .Y(ori_ori_n131_));
  NA2        o115(.A(ori_ori_n131_), .B(ori_ori_n18_), .Y(ori_ori_n132_));
  AOI220     o116(.A0(ori_ori_n132_), .A1(ori_ori_n130_), .B0(ori_ori_n99_), .B1(ori_ori_n38_), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n134_), .B(ori_ori_n108_), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n135_), .B(ori_ori_n133_), .Y(ori_ori_n136_));
  AOI210     o120(.A0(ori_ori_n129_), .A1(ori_ori_n127_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  OAI210     o121(.A0(ori_ori_n126_), .A1(ori_ori_n50_), .B0(ori_ori_n137_), .Y(ori_ori_n138_));
  NA2        o122(.A(x5), .B(x1), .Y(ori_ori_n139_));
  INV        o123(.A(ori_ori_n139_), .Y(ori_ori_n140_));
  AOI210     o124(.A0(ori_ori_n140_), .A1(ori_ori_n108_), .B0(ori_ori_n36_), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n61_), .B(ori_ori_n81_), .Y(ori_ori_n142_));
  NAi21      o126(.An(x2), .B(x7), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n143_), .B(ori_ori_n48_), .Y(ori_ori_n144_));
  NA2        o128(.A(ori_ori_n144_), .B(ori_ori_n62_), .Y(ori_ori_n145_));
  NAi31      o129(.An(ori_ori_n69_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n146_));
  NA3        o130(.A(ori_ori_n146_), .B(ori_ori_n145_), .C(ori_ori_n141_), .Y(ori_ori_n147_));
  NO3        o131(.A(ori_ori_n147_), .B(ori_ori_n138_), .C(ori_ori_n124_), .Y(ori_ori_n148_));
  NO2        o132(.A(ori_ori_n148_), .B(ori_ori_n123_), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n119_), .B(ori_ori_n115_), .Y(ori_ori_n150_));
  NA2        o134(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n151_));
  NA2        o135(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n152_));
  NA3        o136(.A(ori_ori_n152_), .B(ori_ori_n151_), .C(ori_ori_n24_), .Y(ori_ori_n153_));
  AN2        o137(.A(ori_ori_n153_), .B(ori_ori_n120_), .Y(ori_ori_n154_));
  NA2        o138(.A(x8), .B(x0), .Y(ori_ori_n155_));
  NO2        o139(.A(ori_ori_n131_), .B(ori_ori_n25_), .Y(ori_ori_n156_));
  NA2        o140(.A(x2), .B(x0), .Y(ori_ori_n157_));
  NA2        o141(.A(x4), .B(x1), .Y(ori_ori_n158_));
  NAi21      o142(.An(ori_ori_n106_), .B(ori_ori_n158_), .Y(ori_ori_n159_));
  NOi31      o143(.An(ori_ori_n159_), .B(ori_ori_n134_), .C(ori_ori_n157_), .Y(ori_ori_n160_));
  NO3        o144(.A(ori_ori_n160_), .B(ori_ori_n154_), .C(ori_ori_n150_), .Y(ori_ori_n161_));
  NO2        o145(.A(ori_ori_n161_), .B(ori_ori_n43_), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n153_), .B(ori_ori_n67_), .Y(ori_ori_n163_));
  INV        o147(.A(ori_ori_n110_), .Y(ori_ori_n164_));
  NO2        o148(.A(ori_ori_n95_), .B(ori_ori_n17_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n35_), .B(ori_ori_n165_), .Y(ori_ori_n166_));
  NO3        o150(.A(ori_ori_n166_), .B(ori_ori_n164_), .C(x7), .Y(ori_ori_n167_));
  NA3        o151(.A(ori_ori_n159_), .B(ori_ori_n164_), .C(ori_ori_n42_), .Y(ori_ori_n168_));
  OAI210     o152(.A0(ori_ori_n152_), .A1(ori_ori_n115_), .B0(ori_ori_n168_), .Y(ori_ori_n169_));
  NO3        o153(.A(ori_ori_n169_), .B(ori_ori_n167_), .C(ori_ori_n163_), .Y(ori_ori_n170_));
  NO2        o154(.A(ori_ori_n170_), .B(x3), .Y(ori_ori_n171_));
  NO3        o155(.A(ori_ori_n171_), .B(ori_ori_n162_), .C(ori_ori_n149_), .Y(ori03));
  NO2        o156(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n69_), .B(x6), .Y(ori_ori_n175_));
  NA2        o159(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n176_));
  NO2        o160(.A(ori_ori_n176_), .B(x4), .Y(ori_ori_n177_));
  NO2        o161(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n178_));
  AN2        o162(.A(ori_ori_n175_), .B(ori_ori_n55_), .Y(ori_ori_n179_));
  INV        o163(.A(ori_ori_n179_), .Y(ori_ori_n180_));
  NA2        o164(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n181_), .B(ori_ori_n176_), .Y(ori_ori_n182_));
  NA2        o166(.A(x2), .B(x4), .Y(ori_ori_n183_));
  NA2        o167(.A(ori_ori_n183_), .B(ori_ori_n182_), .Y(ori_ori_n184_));
  NO3        o168(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n185_));
  NO2        o169(.A(x5), .B(x1), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n181_), .B(ori_ori_n151_), .Y(ori_ori_n187_));
  NO3        o171(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n188_));
  NO2        o172(.A(ori_ori_n188_), .B(ori_ori_n187_), .Y(ori_ori_n189_));
  INV        o173(.A(ori_ori_n189_), .Y(ori_ori_n190_));
  AOI220     o174(.A0(ori_ori_n190_), .A1(ori_ori_n48_), .B0(ori_ori_n185_), .B1(ori_ori_n110_), .Y(ori_ori_n191_));
  NA3        o175(.A(ori_ori_n191_), .B(ori_ori_n184_), .C(ori_ori_n180_), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n193_));
  NA2        o177(.A(ori_ori_n193_), .B(ori_ori_n19_), .Y(ori_ori_n194_));
  NO2        o178(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n195_), .B(x6), .Y(ori_ori_n196_));
  NOi21      o180(.An(ori_ori_n75_), .B(ori_ori_n196_), .Y(ori_ori_n197_));
  NA2        o181(.A(ori_ori_n195_), .B(x6), .Y(ori_ori_n198_));
  AOI210     o182(.A0(ori_ori_n198_), .A1(ori_ori_n197_), .B0(ori_ori_n131_), .Y(ori_ori_n199_));
  AO210      o183(.A0(ori_ori_n199_), .A1(ori_ori_n194_), .B0(ori_ori_n156_), .Y(ori_ori_n200_));
  NA2        o184(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n120_), .B(ori_ori_n80_), .Y(ori_ori_n202_));
  NA2        o186(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n203_));
  OAI210     o187(.A0(ori_ori_n103_), .A1(ori_ori_n70_), .B0(x4), .Y(ori_ori_n204_));
  AOI210     o188(.A0(ori_ori_n204_), .A1(ori_ori_n203_), .B0(ori_ori_n69_), .Y(ori_ori_n205_));
  NA3        o189(.A(ori_ori_n181_), .B(ori_ori_n110_), .C(x6), .Y(ori_ori_n206_));
  INV        o190(.A(ori_ori_n62_), .Y(ori_ori_n207_));
  NA2        o191(.A(ori_ori_n207_), .B(ori_ori_n206_), .Y(ori_ori_n208_));
  OAI210     o192(.A0(ori_ori_n208_), .A1(ori_ori_n205_), .B0(x2), .Y(ori_ori_n209_));
  NA3        o193(.A(ori_ori_n209_), .B(ori_ori_n202_), .C(ori_ori_n200_), .Y(ori_ori_n210_));
  AOI210     o194(.A0(ori_ori_n192_), .A1(x8), .B0(ori_ori_n210_), .Y(ori_ori_n211_));
  NO2        o195(.A(ori_ori_n79_), .B(ori_ori_n25_), .Y(ori_ori_n212_));
  AOI210     o196(.A0(ori_ori_n196_), .A1(ori_ori_n134_), .B0(ori_ori_n212_), .Y(ori_ori_n213_));
  NO2        o197(.A(ori_ori_n213_), .B(x2), .Y(ori_ori_n214_));
  AOI220     o198(.A0(ori_ori_n177_), .A1(ori_ori_n165_), .B0(x2), .B1(ori_ori_n62_), .Y(ori_ori_n215_));
  NA2        o199(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n216_));
  NA2        o200(.A(ori_ori_n181_), .B(x6), .Y(ori_ori_n217_));
  NO2        o201(.A(ori_ori_n181_), .B(x6), .Y(ori_ori_n218_));
  NAi21      o202(.An(ori_ori_n142_), .B(ori_ori_n218_), .Y(ori_ori_n219_));
  NA3        o203(.A(ori_ori_n219_), .B(ori_ori_n217_), .C(ori_ori_n125_), .Y(ori_ori_n220_));
  NA3        o204(.A(ori_ori_n220_), .B(ori_ori_n215_), .C(ori_ori_n131_), .Y(ori_ori_n221_));
  AOI210     o205(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n222_));
  OAI210     o206(.A0(ori_ori_n119_), .A1(x3), .B0(ori_ori_n222_), .Y(ori_ori_n223_));
  NA2        o207(.A(ori_ori_n223_), .B(x1), .Y(ori_ori_n224_));
  INV        o208(.A(ori_ori_n224_), .Y(ori_ori_n225_));
  NA2        o209(.A(x6), .B(x2), .Y(ori_ori_n226_));
  NA2        o210(.A(x4), .B(ori_ori_n225_), .Y(ori_ori_n227_));
  OR2        o211(.A(ori_ori_n175_), .B(ori_ori_n127_), .Y(ori_ori_n228_));
  NA2        o212(.A(x4), .B(x0), .Y(ori_ori_n229_));
  NA2        o213(.A(ori_ori_n228_), .B(ori_ori_n42_), .Y(ori_ori_n230_));
  AOI210     o214(.A0(ori_ori_n230_), .A1(ori_ori_n227_), .B0(x8), .Y(ori_ori_n231_));
  NA2        o215(.A(ori_ori_n186_), .B(x6), .Y(ori_ori_n232_));
  INV        o216(.A(ori_ori_n155_), .Y(ori_ori_n233_));
  OAI210     o217(.A0(ori_ori_n233_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n234_));
  AOI210     o218(.A0(ori_ori_n234_), .A1(ori_ori_n232_), .B0(ori_ori_n201_), .Y(ori_ori_n235_));
  NO4        o219(.A(ori_ori_n235_), .B(ori_ori_n231_), .C(ori_ori_n221_), .D(ori_ori_n214_), .Y(ori_ori_n236_));
  NA2        o220(.A(ori_ori_n218_), .B(x2), .Y(ori_ori_n237_));
  OAI210     o221(.A0(ori_ori_n233_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n238_));
  AOI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n237_), .B0(ori_ori_n164_), .Y(ori_ori_n239_));
  NOi21      o223(.An(ori_ori_n226_), .B(ori_ori_n17_), .Y(ori_ori_n240_));
  NA3        o224(.A(ori_ori_n240_), .B(ori_ori_n186_), .C(ori_ori_n40_), .Y(ori_ori_n241_));
  AOI210     o225(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n242_));
  NA3        o226(.A(ori_ori_n242_), .B(ori_ori_n140_), .C(ori_ori_n32_), .Y(ori_ori_n243_));
  NA2        o227(.A(x3), .B(x2), .Y(ori_ori_n244_));
  AOI220     o228(.A0(ori_ori_n244_), .A1(ori_ori_n201_), .B0(ori_ori_n243_), .B1(ori_ori_n241_), .Y(ori_ori_n245_));
  NAi21      o229(.An(x4), .B(x0), .Y(ori_ori_n246_));
  NO3        o230(.A(ori_ori_n246_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n247_));
  OAI210     o231(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n247_), .Y(ori_ori_n248_));
  NO2        o232(.A(ori_ori_n242_), .B(ori_ori_n240_), .Y(ori_ori_n249_));
  AOI220     o233(.A0(ori_ori_n249_), .A1(ori_ori_n73_), .B0(ori_ori_n18_), .B1(ori_ori_n31_), .Y(ori_ori_n250_));
  AOI210     o234(.A0(ori_ori_n250_), .A1(ori_ori_n248_), .B0(ori_ori_n25_), .Y(ori_ori_n251_));
  NA3        o235(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n252_));
  NO2        o236(.A(ori_ori_n242_), .B(ori_ori_n240_), .Y(ori_ori_n253_));
  INV        o237(.A(ori_ori_n187_), .Y(ori_ori_n254_));
  NA2        o238(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n255_));
  OR2        o239(.A(ori_ori_n255_), .B(ori_ori_n229_), .Y(ori_ori_n256_));
  OAI220     o240(.A0(ori_ori_n256_), .A1(ori_ori_n139_), .B0(ori_ori_n203_), .B1(ori_ori_n254_), .Y(ori_ori_n257_));
  AO210      o241(.A0(ori_ori_n253_), .A1(ori_ori_n127_), .B0(ori_ori_n257_), .Y(ori_ori_n258_));
  NO4        o242(.A(ori_ori_n258_), .B(ori_ori_n251_), .C(ori_ori_n245_), .D(ori_ori_n239_), .Y(ori_ori_n259_));
  OAI210     o243(.A0(ori_ori_n236_), .A1(ori_ori_n211_), .B0(ori_ori_n259_), .Y(ori04));
  NO2        o244(.A(x2), .B(x1), .Y(ori_ori_n261_));
  OAI210     o245(.A0(ori_ori_n216_), .A1(ori_ori_n261_), .B0(ori_ori_n36_), .Y(ori_ori_n262_));
  NO2        o246(.A(ori_ori_n244_), .B(ori_ori_n178_), .Y(ori_ori_n263_));
  NA2        o247(.A(ori_ori_n263_), .B(ori_ori_n81_), .Y(ori_ori_n264_));
  NA2        o248(.A(ori_ori_n264_), .B(x6), .Y(ori_ori_n265_));
  NA2        o249(.A(ori_ori_n265_), .B(ori_ori_n262_), .Y(ori_ori_n266_));
  NO2        o250(.A(x2), .B(ori_ori_n101_), .Y(ori_ori_n267_));
  NO3        o251(.A(ori_ori_n374_), .B(ori_ori_n104_), .C(ori_ori_n18_), .Y(ori_ori_n268_));
  NO2        o252(.A(ori_ori_n268_), .B(ori_ori_n267_), .Y(ori_ori_n269_));
  OAI210     o253(.A0(ori_ori_n102_), .A1(ori_ori_n95_), .B0(ori_ori_n155_), .Y(ori_ori_n270_));
  NA3        o254(.A(ori_ori_n270_), .B(x6), .C(x3), .Y(ori_ori_n271_));
  NOi21      o255(.An(ori_ori_n129_), .B(ori_ori_n111_), .Y(ori_ori_n272_));
  NO2        o256(.A(ori_ori_n377_), .B(ori_ori_n252_), .Y(ori_ori_n273_));
  AOI210     o257(.A0(ori_ori_n272_), .A1(x6), .B0(ori_ori_n273_), .Y(ori_ori_n274_));
  NA2        o258(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n275_));
  OAI210     o259(.A0(ori_ori_n95_), .A1(ori_ori_n17_), .B0(ori_ori_n275_), .Y(ori_ori_n276_));
  NA2        o260(.A(ori_ori_n276_), .B(ori_ori_n70_), .Y(ori_ori_n277_));
  NA4        o261(.A(ori_ori_n277_), .B(ori_ori_n274_), .C(ori_ori_n271_), .D(ori_ori_n269_), .Y(ori_ori_n278_));
  OAI210     o262(.A0(ori_ori_n100_), .A1(x3), .B0(ori_ori_n247_), .Y(ori_ori_n279_));
  NA2        o263(.A(ori_ori_n185_), .B(ori_ori_n75_), .Y(ori_ori_n280_));
  NA3        o264(.A(ori_ori_n280_), .B(ori_ori_n279_), .C(ori_ori_n131_), .Y(ori_ori_n281_));
  AOI210     o265(.A0(ori_ori_n278_), .A1(x4), .B0(ori_ori_n281_), .Y(ori_ori_n282_));
  XO2        o266(.A(x4), .B(x0), .Y(ori_ori_n283_));
  NA2        o267(.A(x4), .B(ori_ori_n82_), .Y(ori_ori_n284_));
  NO2        o268(.A(ori_ori_n284_), .B(x3), .Y(ori_ori_n285_));
  INV        o269(.A(ori_ori_n82_), .Y(ori_ori_n286_));
  NO2        o270(.A(ori_ori_n81_), .B(x4), .Y(ori_ori_n287_));
  AOI220     o271(.A0(ori_ori_n287_), .A1(ori_ori_n44_), .B0(ori_ori_n108_), .B1(ori_ori_n286_), .Y(ori_ori_n288_));
  NO3        o272(.A(ori_ori_n283_), .B(ori_ori_n142_), .C(x2), .Y(ori_ori_n289_));
  INV        o273(.A(ori_ori_n289_), .Y(ori_ori_n290_));
  NA4        o274(.A(ori_ori_n290_), .B(ori_ori_n288_), .C(ori_ori_n194_), .D(x6), .Y(ori_ori_n291_));
  OAI220     o275(.A0(ori_ori_n246_), .A1(ori_ori_n79_), .B0(ori_ori_n157_), .B1(ori_ori_n81_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n292_), .B(ori_ori_n60_), .Y(ori_ori_n293_));
  NO2        o277(.A(ori_ori_n129_), .B(ori_ori_n72_), .Y(ori_ori_n294_));
  NO2        o278(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n295_));
  NOi21      o279(.An(ori_ori_n106_), .B(ori_ori_n27_), .Y(ori_ori_n296_));
  AOI210     o280(.A0(ori_ori_n295_), .A1(ori_ori_n294_), .B0(ori_ori_n296_), .Y(ori_ori_n297_));
  OAI210     o281(.A0(ori_ori_n293_), .A1(ori_ori_n61_), .B0(ori_ori_n297_), .Y(ori_ori_n298_));
  OAI220     o282(.A0(ori_ori_n298_), .A1(x6), .B0(ori_ori_n291_), .B1(ori_ori_n285_), .Y(ori_ori_n299_));
  OAI210     o283(.A0(x6), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n300_));
  OAI210     o284(.A0(ori_ori_n300_), .A1(ori_ori_n81_), .B0(ori_ori_n256_), .Y(ori_ori_n301_));
  AOI210     o285(.A0(ori_ori_n301_), .A1(ori_ori_n18_), .B0(ori_ori_n131_), .Y(ori_ori_n302_));
  AO220      o286(.A0(ori_ori_n302_), .A1(ori_ori_n299_), .B0(ori_ori_n282_), .B1(ori_ori_n266_), .Y(ori_ori_n303_));
  NA2        o287(.A(ori_ori_n295_), .B(x6), .Y(ori_ori_n304_));
  AOI210     o288(.A0(x6), .A1(x1), .B0(ori_ori_n130_), .Y(ori_ori_n305_));
  NA2        o289(.A(ori_ori_n287_), .B(x0), .Y(ori_ori_n306_));
  NA2        o290(.A(ori_ori_n75_), .B(x6), .Y(ori_ori_n307_));
  OAI210     o291(.A0(ori_ori_n306_), .A1(ori_ori_n305_), .B0(ori_ori_n307_), .Y(ori_ori_n308_));
  NA2        o292(.A(ori_ori_n308_), .B(ori_ori_n304_), .Y(ori_ori_n309_));
  NA2        o293(.A(ori_ori_n309_), .B(ori_ori_n303_), .Y(ori_ori_n310_));
  AOI210     o294(.A0(ori_ori_n174_), .A1(x8), .B0(ori_ori_n100_), .Y(ori_ori_n311_));
  NA2        o295(.A(ori_ori_n311_), .B(ori_ori_n275_), .Y(ori_ori_n312_));
  NA3        o296(.A(ori_ori_n312_), .B(ori_ori_n173_), .C(ori_ori_n131_), .Y(ori_ori_n313_));
  OAI210     o297(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n201_), .Y(ori_ori_n314_));
  AO220      o298(.A0(ori_ori_n314_), .A1(ori_ori_n128_), .B0(ori_ori_n99_), .B1(x4), .Y(ori_ori_n315_));
  NA3        o299(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n316_));
  NA2        o300(.A(ori_ori_n193_), .B(x0), .Y(ori_ori_n317_));
  OAI220     o301(.A0(ori_ori_n317_), .A1(x2), .B0(ori_ori_n316_), .B1(ori_ori_n286_), .Y(ori_ori_n318_));
  AOI210     o302(.A0(ori_ori_n315_), .A1(ori_ori_n103_), .B0(ori_ori_n318_), .Y(ori_ori_n319_));
  AOI210     o303(.A0(ori_ori_n319_), .A1(ori_ori_n313_), .B0(ori_ori_n25_), .Y(ori_ori_n320_));
  NA3        o304(.A(ori_ori_n105_), .B(ori_ori_n193_), .C(x0), .Y(ori_ori_n321_));
  NAi31      o305(.An(ori_ori_n50_), .B(ori_ori_n375_), .C(ori_ori_n156_), .Y(ori_ori_n322_));
  NA2        o306(.A(ori_ori_n322_), .B(ori_ori_n321_), .Y(ori_ori_n323_));
  OAI210     o307(.A0(ori_ori_n323_), .A1(ori_ori_n320_), .B0(x6), .Y(ori_ori_n324_));
  OAI210     o308(.A0(ori_ori_n142_), .A1(ori_ori_n48_), .B0(ori_ori_n114_), .Y(ori_ori_n325_));
  NA2        o309(.A(ori_ori_n55_), .B(ori_ori_n38_), .Y(ori_ori_n326_));
  AOI220     o310(.A0(ori_ori_n326_), .A1(ori_ori_n325_), .B0(ori_ori_n40_), .B1(ori_ori_n32_), .Y(ori_ori_n327_));
  NO2        o311(.A(ori_ori_n131_), .B(x0), .Y(ori_ori_n328_));
  AOI220     o312(.A0(ori_ori_n328_), .A1(ori_ori_n193_), .B0(ori_ori_n173_), .B1(ori_ori_n131_), .Y(ori_ori_n329_));
  OAI210     o313(.A0(ori_ori_n329_), .A1(x8), .B0(ori_ori_n373_), .Y(ori_ori_n330_));
  NAi31      o314(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n331_));
  OAI210     o315(.A0(ori_ori_n331_), .A1(x4), .B0(ori_ori_n143_), .Y(ori_ori_n332_));
  NA2        o316(.A(ori_ori_n332_), .B(ori_ori_n126_), .Y(ori_ori_n333_));
  NO2        o317(.A(ori_ori_n131_), .B(x0), .Y(ori_ori_n334_));
  AOI220     o318(.A0(ori_ori_n334_), .A1(ori_ori_n376_), .B0(ori_ori_n294_), .B1(ori_ori_n131_), .Y(ori_ori_n335_));
  NA4        o319(.A(ori_ori_n335_), .B(x1), .C(ori_ori_n333_), .D(ori_ori_n50_), .Y(ori_ori_n336_));
  OAI210     o320(.A0(ori_ori_n330_), .A1(ori_ori_n327_), .B0(ori_ori_n336_), .Y(ori_ori_n337_));
  NO2        o321(.A(x1), .B(x0), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n338_), .B(x3), .Y(ori_ori_n339_));
  NO3        o323(.A(ori_ori_n339_), .B(x3), .C(x2), .Y(ori_ori_n340_));
  OAI210     o324(.A0(ori_ori_n246_), .A1(ori_ori_n43_), .B0(ori_ori_n283_), .Y(ori_ori_n341_));
  INV        o325(.A(ori_ori_n316_), .Y(ori_ori_n342_));
  AOI220     o326(.A0(ori_ori_n342_), .A1(ori_ori_n81_), .B0(ori_ori_n341_), .B1(ori_ori_n131_), .Y(ori_ori_n343_));
  NO2        o327(.A(ori_ori_n343_), .B(ori_ori_n54_), .Y(ori_ori_n344_));
  NO2        o328(.A(ori_ori_n344_), .B(ori_ori_n340_), .Y(ori_ori_n345_));
  AOI210     o329(.A0(ori_ori_n345_), .A1(ori_ori_n337_), .B0(ori_ori_n25_), .Y(ori_ori_n346_));
  NA4        o330(.A(ori_ori_n31_), .B(ori_ori_n81_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n347_));
  NO2        o331(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n348_));
  NA2        o332(.A(ori_ori_n348_), .B(ori_ori_n222_), .Y(ori_ori_n349_));
  NO2        o333(.A(ori_ori_n349_), .B(ori_ori_n92_), .Y(ori_ori_n350_));
  NA2        o334(.A(ori_ori_n350_), .B(x7), .Y(ori_ori_n351_));
  NA2        o335(.A(ori_ori_n351_), .B(ori_ori_n347_), .Y(ori_ori_n352_));
  OAI210     o336(.A0(ori_ori_n352_), .A1(ori_ori_n346_), .B0(ori_ori_n36_), .Y(ori_ori_n353_));
  INV        o337(.A(ori_ori_n334_), .Y(ori_ori_n354_));
  NO4        o338(.A(ori_ori_n354_), .B(ori_ori_n69_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n355_));
  NA2        o339(.A(ori_ori_n216_), .B(ori_ori_n21_), .Y(ori_ori_n356_));
  NO2        o340(.A(ori_ori_n139_), .B(ori_ori_n114_), .Y(ori_ori_n357_));
  NA2        o341(.A(ori_ori_n357_), .B(ori_ori_n356_), .Y(ori_ori_n358_));
  AOI210     o342(.A0(ori_ori_n358_), .A1(ori_ori_n146_), .B0(ori_ori_n28_), .Y(ori_ori_n359_));
  NA2        o343(.A(ori_ori_n129_), .B(ori_ori_n174_), .Y(ori_ori_n360_));
  NA3        o344(.A(ori_ori_n360_), .B(ori_ori_n331_), .C(ori_ori_n79_), .Y(ori_ori_n361_));
  NA2        o345(.A(ori_ori_n361_), .B(ori_ori_n156_), .Y(ori_ori_n362_));
  NO2        o346(.A(ori_ori_n139_), .B(ori_ori_n43_), .Y(ori_ori_n363_));
  NA2        o347(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n364_));
  NO2        o348(.A(ori_ori_n132_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  AOI220     o349(.A0(ori_ori_n365_), .A1(x0), .B0(ori_ori_n363_), .B1(ori_ori_n114_), .Y(ori_ori_n366_));
  AOI210     o350(.A0(ori_ori_n366_), .A1(ori_ori_n362_), .B0(ori_ori_n203_), .Y(ori_ori_n367_));
  NO3        o351(.A(ori_ori_n367_), .B(ori_ori_n359_), .C(ori_ori_n355_), .Y(ori_ori_n368_));
  NA3        o352(.A(ori_ori_n368_), .B(ori_ori_n353_), .C(ori_ori_n324_), .Y(ori_ori_n369_));
  AOI210     o353(.A0(ori_ori_n310_), .A1(ori_ori_n25_), .B0(ori_ori_n369_), .Y(ori05));
  INV        o354(.A(x1), .Y(ori_ori_n373_));
  INV        o355(.A(x6), .Y(ori_ori_n374_));
  INV        o356(.A(x1), .Y(ori_ori_n375_));
  INV        o357(.A(x3), .Y(ori_ori_n376_));
  INV        o358(.A(x2), .Y(ori_ori_n377_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  INV        m005(.A(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x7), .B(x6), .Y(mai_mai_n25_));
  NA2        m009(.A(x8), .B(x3), .Y(mai_mai_n26_));
  NA2        m010(.A(x4), .B(x2), .Y(mai_mai_n27_));
  INV        m011(.A(mai_mai_n23_), .Y(mai_mai_n28_));
  NO2        m012(.A(x4), .B(x3), .Y(mai_mai_n29_));
  INV        m013(.A(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m014(.An(mai_mai_n22_), .B(mai_mai_n28_), .Y(mai00));
  NO2        m015(.A(x1), .B(x0), .Y(mai_mai_n32_));
  INV        m016(.A(x6), .Y(mai_mai_n33_));
  NO2        m017(.A(mai_mai_n33_), .B(mai_mai_n24_), .Y(mai_mai_n34_));
  NA2        m018(.A(x4), .B(x3), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n22_), .B(mai_mai_n35_), .Y(mai_mai_n36_));
  NO2        m020(.A(x2), .B(x0), .Y(mai_mai_n37_));
  INV        m021(.A(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n39_));
  INV        m023(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n34_), .B(x4), .Y(mai_mai_n41_));
  OAI210     m025(.A0(mai_mai_n41_), .A1(mai_mai_n40_), .B0(mai_mai_n37_), .Y(mai_mai_n42_));
  INV        m026(.A(x4), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n44_));
  NA2        m028(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n45_));
  OAI210     m029(.A0(mai_mai_n45_), .A1(mai_mai_n20_), .B0(mai_mai_n42_), .Y(mai_mai_n46_));
  INV        m030(.A(mai_mai_n32_), .Y(mai_mai_n47_));
  INV        m031(.A(x2), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n51_));
  OAI210     m035(.A0(mai_mai_n47_), .A1(mai_mai_n30_), .B0(mai_mai_n51_), .Y(mai_mai_n52_));
  NO3        m036(.A(mai_mai_n52_), .B(mai_mai_n46_), .C(mai_mai_n36_), .Y(mai01));
  NA2        m037(.A(x8), .B(x7), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n38_), .B(x1), .Y(mai_mai_n55_));
  INV        m039(.A(x9), .Y(mai_mai_n56_));
  NO2        m040(.A(mai_mai_n56_), .B(mai_mai_n33_), .Y(mai_mai_n57_));
  INV        m041(.A(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n55_), .C(mai_mai_n54_), .Y(mai_mai_n59_));
  NO2        m043(.A(x7), .B(x6), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n61_));
  NO2        m045(.A(x8), .B(x2), .Y(mai_mai_n62_));
  INV        m046(.A(mai_mai_n62_), .Y(mai_mai_n63_));
  NO2        m047(.A(mai_mai_n63_), .B(x1), .Y(mai_mai_n64_));
  OA210      m048(.A0(mai_mai_n64_), .A1(mai_mai_n61_), .B0(mai_mai_n60_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n39_), .A1(mai_mai_n24_), .B0(mai_mai_n48_), .Y(mai_mai_n66_));
  OAI210     m050(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  NAi31      m051(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n67_), .B(mai_mai_n65_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n69_), .A1(mai_mai_n59_), .B0(x4), .Y(mai_mai_n70_));
  NA2        m054(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n71_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n72_));
  NA2        m056(.A(x5), .B(x3), .Y(mai_mai_n73_));
  NO2        m057(.A(x8), .B(x6), .Y(mai_mai_n74_));
  NO4        m058(.A(mai_mai_n74_), .B(mai_mai_n73_), .C(mai_mai_n60_), .D(mai_mai_n48_), .Y(mai_mai_n75_));
  NAi21      m059(.An(x4), .B(x3), .Y(mai_mai_n76_));
  INV        m060(.A(mai_mai_n76_), .Y(mai_mai_n77_));
  NO2        m061(.A(x4), .B(x2), .Y(mai_mai_n78_));
  NO2        m062(.A(mai_mai_n78_), .B(x3), .Y(mai_mai_n79_));
  NO2        m063(.A(mai_mai_n76_), .B(mai_mai_n18_), .Y(mai_mai_n80_));
  NO3        m064(.A(mai_mai_n80_), .B(mai_mai_n75_), .C(mai_mai_n72_), .Y(mai_mai_n81_));
  NO3        m065(.A(mai_mai_n21_), .B(mai_mai_n38_), .C(x1), .Y(mai_mai_n82_));
  INV        m066(.A(x4), .Y(mai_mai_n83_));
  NA2        m067(.A(mai_mai_n82_), .B(mai_mai_n83_), .Y(mai_mai_n84_));
  NA2        m068(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n85_));
  NO2        m069(.A(mai_mai_n85_), .B(mai_mai_n24_), .Y(mai_mai_n86_));
  INV        m070(.A(x8), .Y(mai_mai_n87_));
  NA2        m071(.A(x2), .B(x1), .Y(mai_mai_n88_));
  NO2        m072(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n89_), .B(mai_mai_n86_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n25_), .Y(mai_mai_n91_));
  AOI210     m075(.A0(mai_mai_n50_), .A1(mai_mai_n24_), .B0(mai_mai_n48_), .Y(mai_mai_n92_));
  OAI210     m076(.A0(mai_mai_n40_), .A1(mai_mai_n34_), .B0(mai_mai_n43_), .Y(mai_mai_n93_));
  NO3        m077(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n94_));
  NA2        m078(.A(x4), .B(mai_mai_n38_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n43_), .B(mai_mai_n48_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n95_), .B(x1), .Y(mai_mai_n97_));
  NO2        m081(.A(x3), .B(x2), .Y(mai_mai_n98_));
  NA3        m082(.A(mai_mai_n98_), .B(mai_mai_n25_), .C(mai_mai_n24_), .Y(mai_mai_n99_));
  INV        m083(.A(mai_mai_n99_), .Y(mai_mai_n100_));
  NA2        m084(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n101_));
  OAI210     m085(.A0(mai_mai_n101_), .A1(mai_mai_n35_), .B0(mai_mai_n17_), .Y(mai_mai_n102_));
  NO4        m086(.A(mai_mai_n102_), .B(mai_mai_n100_), .C(mai_mai_n97_), .D(mai_mai_n94_), .Y(mai_mai_n103_));
  AO220      m087(.A0(mai_mai_n103_), .A1(mai_mai_n84_), .B0(mai_mai_n81_), .B1(mai_mai_n70_), .Y(mai02));
  NO2        m088(.A(x3), .B(mai_mai_n48_), .Y(mai_mai_n105_));
  NO2        m089(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n106_));
  NA2        m090(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n107_));
  NA2        m091(.A(mai_mai_n38_), .B(x0), .Y(mai_mai_n108_));
  OAI210     m092(.A0(x4), .A1(mai_mai_n107_), .B0(mai_mai_n108_), .Y(mai_mai_n109_));
  AOI220     m093(.A0(mai_mai_n109_), .A1(mai_mai_n106_), .B0(mai_mai_n105_), .B1(x4), .Y(mai_mai_n110_));
  NO3        m094(.A(mai_mai_n110_), .B(x7), .C(x5), .Y(mai_mai_n111_));
  NA2        m095(.A(x9), .B(x2), .Y(mai_mai_n112_));
  OR2        m096(.A(x8), .B(x0), .Y(mai_mai_n113_));
  INV        m097(.A(mai_mai_n113_), .Y(mai_mai_n114_));
  NAi21      m098(.An(x2), .B(x8), .Y(mai_mai_n115_));
  INV        m099(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  OAI220     m100(.A0(mai_mai_n116_), .A1(mai_mai_n114_), .B0(mai_mai_n112_), .B1(x7), .Y(mai_mai_n117_));
  NO2        m101(.A(x4), .B(x1), .Y(mai_mai_n118_));
  NA3        m102(.A(mai_mai_n118_), .B(mai_mai_n117_), .C(mai_mai_n54_), .Y(mai_mai_n119_));
  NOi21      m103(.An(x0), .B(x1), .Y(mai_mai_n120_));
  NO3        m104(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n121_));
  NOi21      m105(.An(x0), .B(x4), .Y(mai_mai_n122_));
  NO2        m106(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n123_));
  AOI220     m107(.A0(mai_mai_n123_), .A1(mai_mai_n122_), .B0(mai_mai_n121_), .B1(mai_mai_n120_), .Y(mai_mai_n124_));
  AOI210     m108(.A0(mai_mai_n124_), .A1(mai_mai_n119_), .B0(mai_mai_n73_), .Y(mai_mai_n125_));
  NO2        m109(.A(x5), .B(mai_mai_n43_), .Y(mai_mai_n126_));
  NA2        m110(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n127_));
  AOI210     m111(.A0(mai_mai_n127_), .A1(mai_mai_n101_), .B0(mai_mai_n108_), .Y(mai_mai_n128_));
  OAI210     m112(.A0(mai_mai_n128_), .A1(mai_mai_n32_), .B0(mai_mai_n126_), .Y(mai_mai_n129_));
  NAi21      m113(.An(x0), .B(x4), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n130_), .B(x1), .Y(mai_mai_n131_));
  NO2        m115(.A(x7), .B(x0), .Y(mai_mai_n132_));
  NO2        m116(.A(mai_mai_n78_), .B(mai_mai_n96_), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n133_), .B(x3), .Y(mai_mai_n134_));
  OAI210     m118(.A0(mai_mai_n132_), .A1(mai_mai_n131_), .B0(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n21_), .B(mai_mai_n38_), .Y(mai_mai_n136_));
  NA2        m120(.A(x5), .B(x0), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n138_));
  NA3        m122(.A(mai_mai_n138_), .B(mai_mai_n137_), .C(mai_mai_n136_), .Y(mai_mai_n139_));
  NA4        m123(.A(mai_mai_n139_), .B(mai_mai_n135_), .C(mai_mai_n129_), .D(mai_mai_n33_), .Y(mai_mai_n140_));
  NO3        m124(.A(mai_mai_n140_), .B(mai_mai_n125_), .C(mai_mai_n111_), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n27_), .B(mai_mai_n24_), .Y(mai_mai_n142_));
  AOI220     m126(.A0(mai_mai_n120_), .A1(mai_mai_n142_), .B0(mai_mai_n61_), .B1(mai_mai_n17_), .Y(mai_mai_n143_));
  NO3        m127(.A(mai_mai_n143_), .B(mai_mai_n54_), .C(mai_mai_n56_), .Y(mai_mai_n144_));
  NO2        m128(.A(x9), .B(x7), .Y(mai_mai_n145_));
  NO2        m129(.A(mai_mai_n38_), .B(x2), .Y(mai_mai_n146_));
  INV        m130(.A(x7), .Y(mai_mai_n147_));
  NA2        m131(.A(mai_mai_n147_), .B(mai_mai_n18_), .Y(mai_mai_n148_));
  NA2        m132(.A(mai_mai_n148_), .B(mai_mai_n146_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n24_), .B(x4), .Y(mai_mai_n150_));
  NO2        m134(.A(mai_mai_n150_), .B(mai_mai_n122_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n151_), .B(mai_mai_n149_), .Y(mai_mai_n152_));
  NA2        m136(.A(x5), .B(x1), .Y(mai_mai_n153_));
  INV        m137(.A(mai_mai_n153_), .Y(mai_mai_n154_));
  AOI210     m138(.A0(mai_mai_n154_), .A1(mai_mai_n122_), .B0(mai_mai_n33_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n56_), .B(mai_mai_n87_), .Y(mai_mai_n156_));
  NO3        m140(.A(x2), .B(mai_mai_n156_), .C(mai_mai_n43_), .Y(mai_mai_n157_));
  NA2        m141(.A(mai_mai_n157_), .B(mai_mai_n61_), .Y(mai_mai_n158_));
  NA2        m142(.A(mai_mai_n158_), .B(mai_mai_n155_), .Y(mai_mai_n159_));
  NO3        m143(.A(mai_mai_n159_), .B(mai_mai_n152_), .C(mai_mai_n144_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n141_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n137_), .B(mai_mai_n133_), .Y(mai_mai_n162_));
  NA2        m146(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n163_));
  NA2        m147(.A(mai_mai_n24_), .B(mai_mai_n17_), .Y(mai_mai_n164_));
  NA3        m148(.A(mai_mai_n164_), .B(mai_mai_n163_), .C(mai_mai_n23_), .Y(mai_mai_n165_));
  AN2        m149(.A(mai_mai_n165_), .B(mai_mai_n138_), .Y(mai_mai_n166_));
  NA2        m150(.A(x8), .B(x0), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n147_), .B(mai_mai_n24_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n120_), .B(x4), .Y(mai_mai_n169_));
  NA2        m153(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  AOI210     m154(.A0(mai_mai_n167_), .A1(mai_mai_n127_), .B0(mai_mai_n170_), .Y(mai_mai_n171_));
  NA2        m155(.A(x2), .B(x0), .Y(mai_mai_n172_));
  NA2        m156(.A(x4), .B(x1), .Y(mai_mai_n173_));
  NAi21      m157(.An(mai_mai_n118_), .B(mai_mai_n173_), .Y(mai_mai_n174_));
  NOi31      m158(.An(mai_mai_n174_), .B(mai_mai_n150_), .C(mai_mai_n172_), .Y(mai_mai_n175_));
  NO4        m159(.A(mai_mai_n175_), .B(mai_mai_n171_), .C(mai_mai_n166_), .D(mai_mai_n162_), .Y(mai_mai_n176_));
  NO2        m160(.A(mai_mai_n176_), .B(mai_mai_n38_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n165_), .B(mai_mai_n71_), .Y(mai_mai_n178_));
  INV        m162(.A(mai_mai_n126_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n101_), .B(mai_mai_n17_), .Y(mai_mai_n180_));
  NA3        m164(.A(mai_mai_n174_), .B(mai_mai_n179_), .C(mai_mai_n37_), .Y(mai_mai_n181_));
  OAI210     m165(.A0(mai_mai_n164_), .A1(mai_mai_n133_), .B0(mai_mai_n181_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n182_), .B(mai_mai_n178_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n183_), .B(x3), .Y(mai_mai_n184_));
  NO3        m168(.A(mai_mai_n184_), .B(mai_mai_n177_), .C(mai_mai_n161_), .Y(mai03));
  NO2        m169(.A(mai_mai_n43_), .B(x3), .Y(mai_mai_n186_));
  NO2        m170(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n187_));
  NO2        m171(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n188_));
  OAI210     m172(.A0(mai_mai_n188_), .A1(mai_mai_n24_), .B0(mai_mai_n57_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n189_), .B(mai_mai_n17_), .Y(mai_mai_n190_));
  NA2        m174(.A(mai_mai_n190_), .B(mai_mai_n186_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n73_), .B(x6), .Y(mai_mai_n192_));
  NA2        m176(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n193_), .B(x4), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n195_));
  NA2        m179(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n196_));
  NA2        m180(.A(mai_mai_n193_), .B(mai_mai_n76_), .Y(mai_mai_n197_));
  AOI210     m181(.A0(mai_mai_n24_), .A1(x3), .B0(mai_mai_n172_), .Y(mai_mai_n198_));
  NA2        m182(.A(mai_mai_n198_), .B(mai_mai_n197_), .Y(mai_mai_n199_));
  NO2        m183(.A(x5), .B(x1), .Y(mai_mai_n200_));
  AOI220     m184(.A0(mai_mai_n200_), .A1(mai_mai_n17_), .B0(mai_mai_n98_), .B1(x5), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n196_), .B(mai_mai_n163_), .Y(mai_mai_n202_));
  NO3        m186(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  OAI210     m188(.A0(mai_mai_n201_), .A1(mai_mai_n58_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  NA2        m189(.A(mai_mai_n205_), .B(mai_mai_n43_), .Y(mai_mai_n206_));
  NA3        m190(.A(mai_mai_n206_), .B(mai_mai_n199_), .C(mai_mai_n191_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n43_), .B(mai_mai_n38_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n19_), .Y(mai_mai_n209_));
  NO2        m193(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n210_));
  NO2        m194(.A(mai_mai_n210_), .B(x6), .Y(mai_mai_n211_));
  NOi21      m195(.An(mai_mai_n78_), .B(mai_mai_n211_), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n212_), .B(mai_mai_n147_), .Y(mai_mai_n213_));
  OR2        m197(.A(mai_mai_n213_), .B(mai_mai_n168_), .Y(mai_mai_n214_));
  NA2        m198(.A(mai_mai_n38_), .B(mai_mai_n48_), .Y(mai_mai_n215_));
  OAI210     m199(.A0(mai_mai_n215_), .A1(mai_mai_n24_), .B0(mai_mai_n164_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n173_), .B(x6), .Y(mai_mai_n217_));
  AOI220     m201(.A0(mai_mai_n217_), .A1(mai_mai_n216_), .B0(mai_mai_n138_), .B1(mai_mai_n86_), .Y(mai_mai_n218_));
  NA2        m202(.A(x6), .B(mai_mai_n43_), .Y(mai_mai_n219_));
  OAI210     m203(.A0(mai_mai_n114_), .A1(mai_mai_n74_), .B0(x4), .Y(mai_mai_n220_));
  AOI210     m204(.A0(mai_mai_n220_), .A1(mai_mai_n219_), .B0(mai_mai_n73_), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n153_), .B(mai_mai_n38_), .Y(mai_mai_n222_));
  OAI210     m206(.A0(mai_mai_n222_), .A1(mai_mai_n202_), .B0(mai_mai_n426_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n187_), .B(mai_mai_n131_), .Y(mai_mai_n224_));
  OAI210     m208(.A0(mai_mai_n87_), .A1(mai_mai_n33_), .B0(mai_mai_n61_), .Y(mai_mai_n225_));
  NA3        m209(.A(mai_mai_n225_), .B(mai_mai_n224_), .C(mai_mai_n223_), .Y(mai_mai_n226_));
  OAI210     m210(.A0(mai_mai_n226_), .A1(mai_mai_n221_), .B0(x2), .Y(mai_mai_n227_));
  NA3        m211(.A(mai_mai_n227_), .B(mai_mai_n218_), .C(mai_mai_n214_), .Y(mai_mai_n228_));
  AOI210     m212(.A0(mai_mai_n207_), .A1(x8), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  NO2        m213(.A(mai_mai_n87_), .B(x3), .Y(mai_mai_n230_));
  NA2        m214(.A(mai_mai_n230_), .B(mai_mai_n194_), .Y(mai_mai_n231_));
  NO3        m215(.A(mai_mai_n85_), .B(mai_mai_n74_), .C(mai_mai_n24_), .Y(mai_mai_n232_));
  AOI210     m216(.A0(mai_mai_n211_), .A1(mai_mai_n150_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  AOI210     m217(.A0(mai_mai_n233_), .A1(mai_mai_n231_), .B0(x2), .Y(mai_mai_n234_));
  NO2        m218(.A(x4), .B(mai_mai_n48_), .Y(mai_mai_n235_));
  AOI220     m219(.A0(mai_mai_n194_), .A1(mai_mai_n180_), .B0(mai_mai_n235_), .B1(mai_mai_n61_), .Y(mai_mai_n236_));
  NA2        m220(.A(mai_mai_n56_), .B(x6), .Y(mai_mai_n237_));
  NA3        m221(.A(mai_mai_n24_), .B(x3), .C(x2), .Y(mai_mai_n238_));
  AOI210     m222(.A0(mai_mai_n238_), .A1(mai_mai_n137_), .B0(mai_mai_n237_), .Y(mai_mai_n239_));
  NA2        m223(.A(mai_mai_n38_), .B(mai_mai_n17_), .Y(mai_mai_n240_));
  NO2        m224(.A(mai_mai_n240_), .B(mai_mai_n24_), .Y(mai_mai_n241_));
  OAI210     m225(.A0(mai_mai_n241_), .A1(mai_mai_n239_), .B0(mai_mai_n118_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n196_), .B(x6), .Y(mai_mai_n243_));
  NO2        m227(.A(mai_mai_n196_), .B(x6), .Y(mai_mai_n244_));
  NA2        m228(.A(mai_mai_n243_), .B(mai_mai_n142_), .Y(mai_mai_n245_));
  NA4        m229(.A(mai_mai_n245_), .B(mai_mai_n242_), .C(mai_mai_n236_), .D(mai_mai_n147_), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n187_), .B(mai_mai_n210_), .Y(mai_mai_n247_));
  NO2        m231(.A(x9), .B(x6), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n137_), .B(mai_mai_n18_), .Y(mai_mai_n249_));
  NAi21      m233(.An(mai_mai_n249_), .B(mai_mai_n238_), .Y(mai_mai_n250_));
  NAi21      m234(.An(x1), .B(x4), .Y(mai_mai_n251_));
  AOI210     m235(.A0(x3), .A1(x2), .B0(mai_mai_n43_), .Y(mai_mai_n252_));
  AOI220     m236(.A0(mai_mai_n43_), .A1(mai_mai_n251_), .B0(mai_mai_n250_), .B1(mai_mai_n248_), .Y(mai_mai_n253_));
  NA2        m237(.A(mai_mai_n253_), .B(mai_mai_n247_), .Y(mai_mai_n254_));
  NA2        m238(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n255_));
  NO2        m239(.A(mai_mai_n255_), .B(mai_mai_n247_), .Y(mai_mai_n256_));
  NO3        m240(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n257_));
  NA2        m241(.A(mai_mai_n101_), .B(mai_mai_n24_), .Y(mai_mai_n258_));
  NA2        m242(.A(x6), .B(x2), .Y(mai_mai_n259_));
  NO2        m243(.A(mai_mai_n259_), .B(mai_mai_n163_), .Y(mai_mai_n260_));
  AOI210     m244(.A0(mai_mai_n258_), .A1(mai_mai_n257_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  OAI220     m245(.A0(mai_mai_n261_), .A1(mai_mai_n38_), .B0(mai_mai_n169_), .B1(mai_mai_n41_), .Y(mai_mai_n262_));
  OAI210     m246(.A0(mai_mai_n262_), .A1(mai_mai_n256_), .B0(mai_mai_n254_), .Y(mai_mai_n263_));
  NA2        m247(.A(x9), .B(mai_mai_n38_), .Y(mai_mai_n264_));
  NO2        m248(.A(mai_mai_n264_), .B(mai_mai_n193_), .Y(mai_mai_n265_));
  OR2        m249(.A(mai_mai_n265_), .B(mai_mai_n192_), .Y(mai_mai_n266_));
  NA2        m250(.A(mai_mai_n266_), .B(mai_mai_n37_), .Y(mai_mai_n267_));
  AOI210     m251(.A0(mai_mai_n267_), .A1(mai_mai_n263_), .B0(x8), .Y(mai_mai_n268_));
  OAI210     m252(.A0(x0), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n269_));
  AOI210     m253(.A0(mai_mai_n269_), .A1(mai_mai_n427_), .B0(mai_mai_n215_), .Y(mai_mai_n270_));
  NO4        m254(.A(mai_mai_n270_), .B(mai_mai_n268_), .C(mai_mai_n246_), .D(mai_mai_n234_), .Y(mai_mai_n271_));
  NO2        m255(.A(mai_mai_n156_), .B(x1), .Y(mai_mai_n272_));
  NO2        m256(.A(x3), .B(mai_mai_n33_), .Y(mai_mai_n273_));
  OAI210     m257(.A0(mai_mai_n273_), .A1(mai_mai_n244_), .B0(x2), .Y(mai_mai_n274_));
  OAI210     m258(.A0(x0), .A1(x6), .B0(mai_mai_n39_), .Y(mai_mai_n275_));
  AOI210     m259(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n179_), .Y(mai_mai_n276_));
  NOi21      m260(.An(mai_mai_n259_), .B(mai_mai_n17_), .Y(mai_mai_n277_));
  NA3        m261(.A(mai_mai_n277_), .B(mai_mai_n200_), .C(mai_mai_n35_), .Y(mai_mai_n278_));
  AOI210     m262(.A0(mai_mai_n33_), .A1(mai_mai_n48_), .B0(x0), .Y(mai_mai_n279_));
  NA3        m263(.A(mai_mai_n279_), .B(mai_mai_n154_), .C(mai_mai_n30_), .Y(mai_mai_n280_));
  NA2        m264(.A(x3), .B(x2), .Y(mai_mai_n281_));
  AOI220     m265(.A0(mai_mai_n281_), .A1(mai_mai_n215_), .B0(mai_mai_n280_), .B1(mai_mai_n278_), .Y(mai_mai_n282_));
  NAi21      m266(.An(x4), .B(x0), .Y(mai_mai_n283_));
  NO3        m267(.A(mai_mai_n283_), .B(mai_mai_n39_), .C(x2), .Y(mai_mai_n284_));
  OAI210     m268(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  OAI220     m269(.A0(mai_mai_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n286_));
  NO2        m270(.A(x9), .B(x8), .Y(mai_mai_n287_));
  NA3        m271(.A(mai_mai_n287_), .B(mai_mai_n33_), .C(mai_mai_n48_), .Y(mai_mai_n288_));
  OAI210     m272(.A0(mai_mai_n279_), .A1(mai_mai_n277_), .B0(mai_mai_n288_), .Y(mai_mai_n289_));
  AOI220     m273(.A0(mai_mai_n289_), .A1(mai_mai_n77_), .B0(mai_mai_n286_), .B1(mai_mai_n29_), .Y(mai_mai_n290_));
  AOI210     m274(.A0(mai_mai_n290_), .A1(mai_mai_n285_), .B0(mai_mai_n24_), .Y(mai_mai_n291_));
  NA3        m275(.A(mai_mai_n33_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n292_));
  INV        m276(.A(mai_mai_n202_), .Y(mai_mai_n293_));
  NA2        m277(.A(mai_mai_n33_), .B(mai_mai_n38_), .Y(mai_mai_n294_));
  NO2        m278(.A(mai_mai_n219_), .B(mai_mai_n293_), .Y(mai_mai_n295_));
  NO4        m279(.A(mai_mai_n295_), .B(mai_mai_n291_), .C(mai_mai_n282_), .D(mai_mai_n276_), .Y(mai_mai_n296_));
  OAI210     m280(.A0(mai_mai_n271_), .A1(mai_mai_n229_), .B0(mai_mai_n296_), .Y(mai04));
  OAI210     m281(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n298_), .B(mai_mai_n257_), .C(mai_mai_n79_), .Y(mai_mai_n299_));
  NO2        m283(.A(x2), .B(x1), .Y(mai_mai_n300_));
  OAI210     m284(.A0(mai_mai_n240_), .A1(mai_mai_n300_), .B0(mai_mai_n33_), .Y(mai_mai_n301_));
  NO2        m285(.A(mai_mai_n300_), .B(mai_mai_n283_), .Y(mai_mai_n302_));
  INV        m286(.A(mai_mai_n107_), .Y(mai_mai_n303_));
  OAI210     m287(.A0(mai_mai_n303_), .A1(mai_mai_n302_), .B0(mai_mai_n230_), .Y(mai_mai_n304_));
  NO2        m288(.A(mai_mai_n255_), .B(mai_mai_n85_), .Y(mai_mai_n305_));
  NO2        m289(.A(mai_mai_n305_), .B(mai_mai_n33_), .Y(mai_mai_n306_));
  NO2        m290(.A(mai_mai_n281_), .B(mai_mai_n195_), .Y(mai_mai_n307_));
  NA2        m291(.A(x9), .B(x0), .Y(mai_mai_n308_));
  AOI210     m292(.A0(mai_mai_n85_), .A1(mai_mai_n71_), .B0(mai_mai_n308_), .Y(mai_mai_n309_));
  OAI210     m293(.A0(mai_mai_n309_), .A1(mai_mai_n307_), .B0(mai_mai_n87_), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n306_), .C(mai_mai_n304_), .Y(mai_mai_n311_));
  NA2        m295(.A(mai_mai_n311_), .B(mai_mai_n301_), .Y(mai_mai_n312_));
  AOI210     m296(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n313_));
  OAI220     m297(.A0(mai_mai_n313_), .A1(mai_mai_n294_), .B0(mai_mai_n255_), .B1(mai_mai_n292_), .Y(mai_mai_n314_));
  INV        m298(.A(mai_mai_n314_), .Y(mai_mai_n315_));
  NA2        m299(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n316_));
  OAI210     m300(.A0(mai_mai_n101_), .A1(mai_mai_n17_), .B0(mai_mai_n316_), .Y(mai_mai_n317_));
  AOI220     m301(.A0(mai_mai_n317_), .A1(mai_mai_n74_), .B0(mai_mai_n305_), .B1(mai_mai_n87_), .Y(mai_mai_n318_));
  NA2        m302(.A(mai_mai_n318_), .B(mai_mai_n315_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n106_), .A1(x3), .B0(mai_mai_n284_), .Y(mai_mai_n320_));
  NA2        m304(.A(mai_mai_n320_), .B(mai_mai_n147_), .Y(mai_mai_n321_));
  AOI210     m305(.A0(mai_mai_n319_), .A1(x4), .B0(mai_mai_n321_), .Y(mai_mai_n322_));
  NA2        m306(.A(mai_mai_n302_), .B(mai_mai_n87_), .Y(mai_mai_n323_));
  NOi21      m307(.An(x4), .B(x0), .Y(mai_mai_n324_));
  XO2        m308(.A(x4), .B(x0), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n325_), .A1(mai_mai_n112_), .B0(mai_mai_n251_), .Y(mai_mai_n326_));
  AOI220     m310(.A0(mai_mai_n326_), .A1(x8), .B0(mai_mai_n324_), .B1(mai_mai_n88_), .Y(mai_mai_n327_));
  AOI210     m311(.A0(mai_mai_n327_), .A1(mai_mai_n323_), .B0(x3), .Y(mai_mai_n328_));
  INV        m312(.A(mai_mai_n88_), .Y(mai_mai_n329_));
  NO2        m313(.A(mai_mai_n87_), .B(x4), .Y(mai_mai_n330_));
  NO3        m314(.A(mai_mai_n325_), .B(mai_mai_n156_), .C(x2), .Y(mai_mai_n331_));
  NO2        m315(.A(mai_mai_n27_), .B(mai_mai_n23_), .Y(mai_mai_n332_));
  NO2        m316(.A(mai_mai_n332_), .B(mai_mai_n331_), .Y(mai_mai_n333_));
  NA3        m317(.A(mai_mai_n333_), .B(mai_mai_n209_), .C(x6), .Y(mai_mai_n334_));
  OAI220     m318(.A0(mai_mai_n283_), .A1(mai_mai_n85_), .B0(mai_mai_n172_), .B1(mai_mai_n87_), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n38_), .B(x0), .Y(mai_mai_n336_));
  OR2        m320(.A(mai_mai_n330_), .B(mai_mai_n336_), .Y(mai_mai_n337_));
  INV        m321(.A(mai_mai_n101_), .Y(mai_mai_n338_));
  AOI220     m322(.A0(mai_mai_n338_), .A1(mai_mai_n337_), .B0(mai_mai_n335_), .B1(mai_mai_n55_), .Y(mai_mai_n339_));
  INV        m323(.A(mai_mai_n76_), .Y(mai_mai_n340_));
  NO2        m324(.A(mai_mai_n32_), .B(x2), .Y(mai_mai_n341_));
  NOi21      m325(.An(mai_mai_n118_), .B(mai_mai_n26_), .Y(mai_mai_n342_));
  AOI210     m326(.A0(mai_mai_n341_), .A1(mai_mai_n340_), .B0(mai_mai_n342_), .Y(mai_mai_n343_));
  OAI210     m327(.A0(mai_mai_n339_), .A1(mai_mai_n56_), .B0(mai_mai_n343_), .Y(mai_mai_n344_));
  OAI220     m328(.A0(mai_mai_n344_), .A1(x6), .B0(mai_mai_n334_), .B1(mai_mai_n328_), .Y(mai_mai_n345_));
  AO220      m329(.A0(x7), .A1(mai_mai_n345_), .B0(mai_mai_n322_), .B1(mai_mai_n312_), .Y(mai_mai_n346_));
  NA2        m330(.A(mai_mai_n341_), .B(x6), .Y(mai_mai_n347_));
  AOI210     m331(.A0(x6), .A1(x1), .B0(mai_mai_n146_), .Y(mai_mai_n348_));
  NA2        m332(.A(mai_mai_n330_), .B(x0), .Y(mai_mai_n349_));
  NA2        m333(.A(mai_mai_n78_), .B(x6), .Y(mai_mai_n350_));
  OAI210     m334(.A0(mai_mai_n349_), .A1(mai_mai_n348_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  AOI220     m335(.A0(mai_mai_n351_), .A1(mai_mai_n347_), .B0(mai_mai_n203_), .B1(mai_mai_n44_), .Y(mai_mai_n352_));
  NA3        m336(.A(mai_mai_n352_), .B(mai_mai_n346_), .C(mai_mai_n299_), .Y(mai_mai_n353_));
  AOI210     m337(.A0(mai_mai_n188_), .A1(x8), .B0(mai_mai_n106_), .Y(mai_mai_n354_));
  NA2        m338(.A(mai_mai_n354_), .B(mai_mai_n316_), .Y(mai_mai_n355_));
  NA3        m339(.A(mai_mai_n355_), .B(mai_mai_n186_), .C(mai_mai_n147_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n27_), .A1(x1), .B0(mai_mai_n215_), .Y(mai_mai_n357_));
  AO220      m341(.A0(mai_mai_n357_), .A1(mai_mai_n145_), .B0(mai_mai_n105_), .B1(x4), .Y(mai_mai_n358_));
  NA3        m342(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n359_));
  NO2        m343(.A(mai_mai_n359_), .B(mai_mai_n329_), .Y(mai_mai_n360_));
  AOI210     m344(.A0(mai_mai_n358_), .A1(mai_mai_n114_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  AOI210     m345(.A0(mai_mai_n361_), .A1(mai_mai_n356_), .B0(mai_mai_n24_), .Y(mai_mai_n362_));
  NA3        m346(.A(mai_mai_n116_), .B(mai_mai_n208_), .C(x0), .Y(mai_mai_n363_));
  OAI210     m347(.A0(mai_mai_n186_), .A1(mai_mai_n62_), .B0(mai_mai_n195_), .Y(mai_mai_n364_));
  NA3        m348(.A(mai_mai_n188_), .B(mai_mai_n210_), .C(x8), .Y(mai_mai_n365_));
  AOI210     m349(.A0(mai_mai_n365_), .A1(mai_mai_n364_), .B0(mai_mai_n24_), .Y(mai_mai_n366_));
  AOI210     m350(.A0(mai_mai_n115_), .A1(mai_mai_n113_), .B0(mai_mai_n37_), .Y(mai_mai_n367_));
  NOi31      m351(.An(mai_mai_n367_), .B(mai_mai_n336_), .C(mai_mai_n173_), .Y(mai_mai_n368_));
  OAI210     m352(.A0(mai_mai_n368_), .A1(mai_mai_n366_), .B0(mai_mai_n145_), .Y(mai_mai_n369_));
  NAi31      m353(.An(mai_mai_n45_), .B(mai_mai_n272_), .C(mai_mai_n168_), .Y(mai_mai_n370_));
  NA3        m354(.A(mai_mai_n370_), .B(mai_mai_n369_), .C(mai_mai_n363_), .Y(mai_mai_n371_));
  OAI210     m355(.A0(mai_mai_n371_), .A1(mai_mai_n362_), .B0(x6), .Y(mai_mai_n372_));
  INV        m356(.A(mai_mai_n132_), .Y(mai_mai_n373_));
  AOI210     m357(.A0(mai_mai_n35_), .A1(mai_mai_n30_), .B0(mai_mai_n373_), .Y(mai_mai_n374_));
  NO2        m358(.A(mai_mai_n147_), .B(x0), .Y(mai_mai_n375_));
  AOI220     m359(.A0(mai_mai_n375_), .A1(mai_mai_n208_), .B0(mai_mai_n186_), .B1(mai_mai_n147_), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n123_), .A1(mai_mai_n235_), .B0(x1), .Y(mai_mai_n377_));
  OAI210     m361(.A0(mai_mai_n376_), .A1(x8), .B0(mai_mai_n377_), .Y(mai_mai_n378_));
  NO4        m362(.A(x8), .B(mai_mai_n283_), .C(x9), .D(x2), .Y(mai_mai_n379_));
  NOi21      m363(.An(mai_mai_n121_), .B(mai_mai_n172_), .Y(mai_mai_n380_));
  NO3        m364(.A(mai_mai_n380_), .B(mai_mai_n379_), .C(mai_mai_n18_), .Y(mai_mai_n381_));
  NO3        m365(.A(x9), .B(mai_mai_n147_), .C(x0), .Y(mai_mai_n382_));
  AOI220     m366(.A0(mai_mai_n382_), .A1(mai_mai_n230_), .B0(mai_mai_n340_), .B1(mai_mai_n147_), .Y(mai_mai_n383_));
  NA3        m367(.A(mai_mai_n383_), .B(mai_mai_n381_), .C(mai_mai_n45_), .Y(mai_mai_n384_));
  OAI210     m368(.A0(mai_mai_n378_), .A1(mai_mai_n374_), .B0(mai_mai_n384_), .Y(mai_mai_n385_));
  NOi31      m369(.An(mai_mai_n375_), .B(mai_mai_n30_), .C(x8), .Y(mai_mai_n386_));
  INV        m370(.A(mai_mai_n130_), .Y(mai_mai_n387_));
  NO3        m371(.A(mai_mai_n387_), .B(mai_mai_n121_), .C(mai_mai_n38_), .Y(mai_mai_n388_));
  NOi31      m372(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n389_));
  AOI220     m373(.A0(mai_mai_n389_), .A1(mai_mai_n324_), .B0(mai_mai_n122_), .B1(x3), .Y(mai_mai_n390_));
  AOI210     m374(.A0(mai_mai_n251_), .A1(mai_mai_n54_), .B0(mai_mai_n120_), .Y(mai_mai_n391_));
  OAI210     m375(.A0(mai_mai_n391_), .A1(x3), .B0(mai_mai_n390_), .Y(mai_mai_n392_));
  NO3        m376(.A(mai_mai_n392_), .B(mai_mai_n388_), .C(x2), .Y(mai_mai_n393_));
  OAI220     m377(.A0(mai_mai_n325_), .A1(mai_mai_n287_), .B0(mai_mai_n283_), .B1(mai_mai_n38_), .Y(mai_mai_n394_));
  NA2        m378(.A(mai_mai_n394_), .B(mai_mai_n147_), .Y(mai_mai_n395_));
  NO2        m379(.A(mai_mai_n395_), .B(mai_mai_n48_), .Y(mai_mai_n396_));
  NO3        m380(.A(mai_mai_n396_), .B(mai_mai_n393_), .C(mai_mai_n386_), .Y(mai_mai_n397_));
  AOI210     m381(.A0(mai_mai_n397_), .A1(mai_mai_n385_), .B0(mai_mai_n24_), .Y(mai_mai_n398_));
  NO3        m382(.A(mai_mai_n56_), .B(x4), .C(x1), .Y(mai_mai_n399_));
  NO3        m383(.A(mai_mai_n62_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n400_));
  AOI220     m384(.A0(mai_mai_n400_), .A1(mai_mai_n252_), .B0(mai_mai_n399_), .B1(mai_mai_n367_), .Y(mai_mai_n401_));
  NO2        m385(.A(mai_mai_n401_), .B(mai_mai_n98_), .Y(mai_mai_n402_));
  NO3        m386(.A(mai_mai_n255_), .B(mai_mai_n167_), .C(mai_mai_n35_), .Y(mai_mai_n403_));
  OAI210     m387(.A0(mai_mai_n403_), .A1(mai_mai_n402_), .B0(x7), .Y(mai_mai_n404_));
  NA2        m388(.A(mai_mai_n146_), .B(mai_mai_n131_), .Y(mai_mai_n405_));
  NA2        m389(.A(mai_mai_n405_), .B(mai_mai_n404_), .Y(mai_mai_n406_));
  OAI210     m390(.A0(mai_mai_n406_), .A1(mai_mai_n398_), .B0(mai_mai_n33_), .Y(mai_mai_n407_));
  NO2        m391(.A(mai_mai_n382_), .B(mai_mai_n195_), .Y(mai_mai_n408_));
  NO4        m392(.A(mai_mai_n408_), .B(mai_mai_n73_), .C(x4), .D(mai_mai_n48_), .Y(mai_mai_n409_));
  NA2        m393(.A(mai_mai_n336_), .B(mai_mai_n168_), .Y(mai_mai_n410_));
  OAI220     m394(.A0(mai_mai_n264_), .A1(mai_mai_n63_), .B0(mai_mai_n153_), .B1(mai_mai_n38_), .Y(mai_mai_n411_));
  AOI210     m395(.A0(x2), .A1(mai_mai_n26_), .B0(mai_mai_n68_), .Y(mai_mai_n412_));
  OAI210     m396(.A0(mai_mai_n145_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n413_));
  NO3        m397(.A(mai_mai_n389_), .B(x3), .C(mai_mai_n48_), .Y(mai_mai_n414_));
  AOI210     m398(.A0(mai_mai_n414_), .A1(mai_mai_n413_), .B0(mai_mai_n412_), .Y(mai_mai_n415_));
  INV        m399(.A(mai_mai_n415_), .Y(mai_mai_n416_));
  AOI220     m400(.A0(mai_mai_n416_), .A1(x0), .B0(mai_mai_n411_), .B1(mai_mai_n132_), .Y(mai_mai_n417_));
  AOI210     m401(.A0(mai_mai_n417_), .A1(mai_mai_n410_), .B0(mai_mai_n219_), .Y(mai_mai_n418_));
  INV        m402(.A(x5), .Y(mai_mai_n419_));
  NO4        m403(.A(mai_mai_n101_), .B(mai_mai_n419_), .C(mai_mai_n54_), .D(mai_mai_n30_), .Y(mai_mai_n420_));
  NO3        m404(.A(mai_mai_n420_), .B(mai_mai_n418_), .C(mai_mai_n409_), .Y(mai_mai_n421_));
  NA3        m405(.A(mai_mai_n421_), .B(mai_mai_n407_), .C(mai_mai_n372_), .Y(mai_mai_n422_));
  AOI210     m406(.A0(mai_mai_n353_), .A1(mai_mai_n24_), .B0(mai_mai_n422_), .Y(mai05));
  INV        m407(.A(x6), .Y(mai_mai_n426_));
  INV        m408(.A(mai_mai_n249_), .Y(mai_mai_n427_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n63_));
  NO3        u047(.A(men_men_n36_), .B(men_men_n61_), .C(men_men_n60_), .Y(men_men_n64_));
  NO2        u048(.A(x7), .B(x6), .Y(men_men_n65_));
  NO2        u049(.A(men_men_n61_), .B(x5), .Y(men_men_n66_));
  NO2        u050(.A(x8), .B(x2), .Y(men_men_n67_));
  INV        u051(.A(men_men_n67_), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n67_), .A1(men_men_n66_), .B0(men_men_n65_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n43_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n64_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n48_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO3        u062(.A(men_men_n77_), .B(men_men_n65_), .C(men_men_n54_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(men_men_n22_), .Y(men_men_n82_));
  NO2        u066(.A(x4), .B(x2), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(x3), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n82_), .C(men_men_n18_), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n86_));
  NO3        u070(.A(x6), .B(men_men_n43_), .C(x1), .Y(men_men_n87_));
  NA2        u071(.A(men_men_n62_), .B(men_men_n48_), .Y(men_men_n88_));
  INV        u072(.A(men_men_n88_), .Y(men_men_n89_));
  OAI210     u073(.A0(men_men_n87_), .A1(men_men_n66_), .B0(men_men_n89_), .Y(men_men_n90_));
  NA2        u074(.A(x3), .B(men_men_n18_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n25_), .Y(men_men_n92_));
  INV        u076(.A(x8), .Y(men_men_n93_));
  NA2        u077(.A(x2), .B(x1), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n92_), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n26_), .Y(men_men_n97_));
  AOI210     u081(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n98_));
  OAI210     u082(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n99_));
  NO3        u083(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n100_));
  NA2        u084(.A(x4), .B(men_men_n43_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n102_));
  OAI210     u086(.A0(men_men_n102_), .A1(men_men_n43_), .B0(men_men_n18_), .Y(men_men_n103_));
  AOI210     u087(.A0(men_men_n101_), .A1(men_men_n52_), .B0(men_men_n103_), .Y(men_men_n104_));
  NO2        u088(.A(x3), .B(x2), .Y(men_men_n105_));
  NA2        u089(.A(men_men_n105_), .B(men_men_n25_), .Y(men_men_n106_));
  AOI210     u090(.A0(x8), .A1(x6), .B0(men_men_n106_), .Y(men_men_n107_));
  NA2        u091(.A(men_men_n54_), .B(x1), .Y(men_men_n108_));
  OAI210     u092(.A0(men_men_n108_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n109_));
  NO4        u093(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n104_), .D(men_men_n100_), .Y(men_men_n110_));
  AO220      u094(.A0(men_men_n110_), .A1(men_men_n90_), .B0(men_men_n86_), .B1(men_men_n74_), .Y(men02));
  NO2        u095(.A(x3), .B(men_men_n54_), .Y(men_men_n112_));
  NO2        u096(.A(x8), .B(men_men_n18_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n114_));
  NA2        u098(.A(men_men_n43_), .B(x0), .Y(men_men_n115_));
  OAI210     u099(.A0(men_men_n88_), .A1(men_men_n114_), .B0(men_men_n115_), .Y(men_men_n116_));
  AOI220     u100(.A0(men_men_n116_), .A1(men_men_n113_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n117_));
  NO3        u101(.A(men_men_n117_), .B(x7), .C(x5), .Y(men_men_n118_));
  NA2        u102(.A(x9), .B(x2), .Y(men_men_n119_));
  OR2        u103(.A(x8), .B(x0), .Y(men_men_n120_));
  NAi21      u104(.An(x2), .B(x8), .Y(men_men_n121_));
  NO2        u105(.A(x4), .B(x1), .Y(men_men_n122_));
  NOi21      u106(.An(x0), .B(x1), .Y(men_men_n123_));
  NO3        u107(.A(x9), .B(x8), .C(x7), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x4), .Y(men_men_n125_));
  NAi21      u109(.An(x8), .B(x7), .Y(men_men_n126_));
  NO2        u110(.A(men_men_n126_), .B(men_men_n62_), .Y(men_men_n127_));
  AOI220     u111(.A0(men_men_n127_), .A1(men_men_n125_), .B0(men_men_n124_), .B1(men_men_n123_), .Y(men_men_n128_));
  NO2        u112(.A(men_men_n128_), .B(men_men_n77_), .Y(men_men_n129_));
  NO2        u113(.A(x5), .B(men_men_n48_), .Y(men_men_n130_));
  NA2        u114(.A(x2), .B(men_men_n18_), .Y(men_men_n131_));
  AOI210     u115(.A0(men_men_n131_), .A1(men_men_n108_), .B0(men_men_n115_), .Y(men_men_n132_));
  OAI210     u116(.A0(men_men_n132_), .A1(men_men_n35_), .B0(men_men_n130_), .Y(men_men_n133_));
  NAi21      u117(.An(x0), .B(x4), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x1), .Y(men_men_n135_));
  NO2        u119(.A(x7), .B(x0), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n83_), .B(men_men_n102_), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x3), .Y(men_men_n138_));
  OAI210     u122(.A0(men_men_n136_), .A1(men_men_n135_), .B0(men_men_n138_), .Y(men_men_n139_));
  NA2        u123(.A(x5), .B(x0), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n48_), .B(x2), .Y(men_men_n141_));
  NA3        u125(.A(men_men_n139_), .B(men_men_n133_), .C(men_men_n36_), .Y(men_men_n142_));
  NO3        u126(.A(men_men_n142_), .B(men_men_n129_), .C(men_men_n118_), .Y(men_men_n143_));
  NO3        u127(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n24_), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n145_));
  AOI220     u129(.A0(men_men_n123_), .A1(men_men_n145_), .B0(men_men_n66_), .B1(men_men_n17_), .Y(men_men_n146_));
  NO2        u130(.A(men_men_n146_), .B(men_men_n60_), .Y(men_men_n147_));
  NA2        u131(.A(x7), .B(x3), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n101_), .B(x5), .Y(men_men_n149_));
  NO2        u133(.A(x9), .B(x7), .Y(men_men_n150_));
  NOi21      u134(.An(x8), .B(x0), .Y(men_men_n151_));
  OA210      u135(.A0(men_men_n150_), .A1(x1), .B0(men_men_n151_), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n43_), .B(x2), .Y(men_men_n153_));
  INV        u137(.A(x7), .Y(men_men_n154_));
  NA2        u138(.A(men_men_n154_), .B(men_men_n18_), .Y(men_men_n155_));
  AOI220     u139(.A0(men_men_n155_), .A1(men_men_n153_), .B0(men_men_n112_), .B1(men_men_n38_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n25_), .B(x4), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n157_), .B(men_men_n125_), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n158_), .B(men_men_n156_), .Y(men_men_n159_));
  AOI210     u143(.A0(men_men_n152_), .A1(men_men_n149_), .B0(men_men_n159_), .Y(men_men_n160_));
  OAI210     u144(.A0(men_men_n148_), .A1(men_men_n50_), .B0(men_men_n160_), .Y(men_men_n161_));
  NA2        u145(.A(x5), .B(x1), .Y(men_men_n162_));
  INV        u146(.A(men_men_n162_), .Y(men_men_n163_));
  AOI210     u147(.A0(men_men_n163_), .A1(men_men_n125_), .B0(men_men_n36_), .Y(men_men_n164_));
  NO2        u148(.A(men_men_n62_), .B(men_men_n93_), .Y(men_men_n165_));
  NAi21      u149(.An(x2), .B(x7), .Y(men_men_n166_));
  NAi31      u150(.An(men_men_n77_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n167_));
  NA2        u151(.A(men_men_n167_), .B(men_men_n164_), .Y(men_men_n168_));
  NO4        u152(.A(men_men_n168_), .B(men_men_n161_), .C(men_men_n147_), .D(men_men_n144_), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n169_), .B(men_men_n143_), .Y(men_men_n170_));
  NO2        u154(.A(men_men_n140_), .B(men_men_n137_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n172_));
  NA2        u156(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n173_));
  NA3        u157(.A(men_men_n173_), .B(men_men_n172_), .C(men_men_n24_), .Y(men_men_n174_));
  AN2        u158(.A(men_men_n174_), .B(men_men_n141_), .Y(men_men_n175_));
  NA2        u159(.A(x8), .B(x0), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n154_), .B(men_men_n25_), .Y(men_men_n177_));
  NO2        u161(.A(men_men_n123_), .B(x4), .Y(men_men_n178_));
  NA2        u162(.A(men_men_n178_), .B(men_men_n177_), .Y(men_men_n179_));
  AOI210     u163(.A0(men_men_n176_), .A1(men_men_n131_), .B0(men_men_n179_), .Y(men_men_n180_));
  NA2        u164(.A(x2), .B(x0), .Y(men_men_n181_));
  NA2        u165(.A(x4), .B(x1), .Y(men_men_n182_));
  NAi21      u166(.An(men_men_n122_), .B(men_men_n182_), .Y(men_men_n183_));
  NOi31      u167(.An(men_men_n183_), .B(men_men_n157_), .C(men_men_n181_), .Y(men_men_n184_));
  NO4        u168(.A(men_men_n184_), .B(men_men_n180_), .C(men_men_n175_), .D(men_men_n171_), .Y(men_men_n185_));
  NO2        u169(.A(men_men_n185_), .B(men_men_n43_), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n174_), .B(men_men_n75_), .Y(men_men_n187_));
  INV        u171(.A(men_men_n130_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n108_), .B(men_men_n17_), .Y(men_men_n189_));
  AOI210     u173(.A0(men_men_n35_), .A1(men_men_n93_), .B0(men_men_n189_), .Y(men_men_n190_));
  NO3        u174(.A(men_men_n190_), .B(men_men_n188_), .C(x7), .Y(men_men_n191_));
  NA3        u175(.A(men_men_n183_), .B(men_men_n188_), .C(men_men_n42_), .Y(men_men_n192_));
  OAI210     u176(.A0(men_men_n173_), .A1(men_men_n137_), .B0(men_men_n192_), .Y(men_men_n193_));
  NO3        u177(.A(men_men_n193_), .B(men_men_n191_), .C(men_men_n187_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n194_), .B(x3), .Y(men_men_n195_));
  NO3        u179(.A(men_men_n195_), .B(men_men_n186_), .C(men_men_n170_), .Y(men03));
  NO2        u180(.A(men_men_n48_), .B(x3), .Y(men_men_n197_));
  NO2        u181(.A(x6), .B(men_men_n25_), .Y(men_men_n198_));
  INV        u182(.A(men_men_n198_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n54_), .B(x1), .Y(men_men_n200_));
  OAI210     u184(.A0(men_men_n200_), .A1(men_men_n25_), .B0(men_men_n63_), .Y(men_men_n201_));
  OAI220     u185(.A0(men_men_n201_), .A1(men_men_n17_), .B0(men_men_n199_), .B1(men_men_n108_), .Y(men_men_n202_));
  NA2        u186(.A(men_men_n202_), .B(men_men_n197_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n77_), .B(x6), .Y(men_men_n204_));
  NA2        u188(.A(x6), .B(men_men_n25_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n205_), .B(x4), .Y(men_men_n206_));
  AO220      u190(.A0(men_men_n440_), .A1(men_men_n206_), .B0(men_men_n204_), .B1(men_men_n55_), .Y(men_men_n207_));
  NA2        u191(.A(men_men_n207_), .B(men_men_n62_), .Y(men_men_n208_));
  NA2        u192(.A(x3), .B(men_men_n17_), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n209_), .B(men_men_n205_), .Y(men_men_n210_));
  NA2        u194(.A(x9), .B(men_men_n54_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n205_), .B(men_men_n80_), .Y(men_men_n212_));
  AOI210     u196(.A0(men_men_n25_), .A1(x3), .B0(men_men_n181_), .Y(men_men_n213_));
  AOI220     u197(.A0(men_men_n213_), .A1(men_men_n212_), .B0(x9), .B1(men_men_n210_), .Y(men_men_n214_));
  NO3        u198(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n215_));
  NO2        u199(.A(x5), .B(x1), .Y(men_men_n216_));
  AOI220     u200(.A0(men_men_n216_), .A1(men_men_n17_), .B0(men_men_n105_), .B1(x5), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n209_), .B(men_men_n172_), .Y(men_men_n218_));
  NO2        u202(.A(men_men_n217_), .B(men_men_n36_), .Y(men_men_n219_));
  AOI220     u203(.A0(men_men_n219_), .A1(men_men_n48_), .B0(men_men_n215_), .B1(men_men_n130_), .Y(men_men_n220_));
  NA4        u204(.A(men_men_n220_), .B(men_men_n214_), .C(men_men_n208_), .D(men_men_n203_), .Y(men_men_n221_));
  NO2        u205(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n222_), .B(men_men_n19_), .Y(men_men_n223_));
  NO2        u207(.A(x3), .B(men_men_n17_), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n224_), .B(x6), .Y(men_men_n225_));
  NOi21      u209(.An(men_men_n83_), .B(men_men_n225_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n62_), .B(men_men_n93_), .Y(men_men_n227_));
  NA3        u211(.A(men_men_n227_), .B(men_men_n224_), .C(x6), .Y(men_men_n228_));
  AOI210     u212(.A0(men_men_n228_), .A1(men_men_n226_), .B0(men_men_n154_), .Y(men_men_n229_));
  AO210      u213(.A0(men_men_n229_), .A1(men_men_n223_), .B0(men_men_n177_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n25_), .B0(men_men_n173_), .Y(men_men_n232_));
  NO3        u216(.A(men_men_n182_), .B(men_men_n62_), .C(x6), .Y(men_men_n233_));
  AOI220     u217(.A0(men_men_n233_), .A1(men_men_n232_), .B0(men_men_n141_), .B1(men_men_n92_), .Y(men_men_n234_));
  NA2        u218(.A(x6), .B(men_men_n48_), .Y(men_men_n235_));
  NO2        u219(.A(men_men_n235_), .B(men_men_n77_), .Y(men_men_n236_));
  NO2        u220(.A(men_men_n62_), .B(x6), .Y(men_men_n237_));
  NO2        u221(.A(men_men_n162_), .B(men_men_n43_), .Y(men_men_n238_));
  OAI210     u222(.A0(men_men_n238_), .A1(men_men_n218_), .B0(men_men_n237_), .Y(men_men_n239_));
  NA2        u223(.A(men_men_n198_), .B(men_men_n135_), .Y(men_men_n240_));
  NA3        u224(.A(men_men_n209_), .B(men_men_n130_), .C(x6), .Y(men_men_n241_));
  OAI210     u225(.A0(men_men_n93_), .A1(men_men_n36_), .B0(men_men_n66_), .Y(men_men_n242_));
  NA4        u226(.A(men_men_n242_), .B(men_men_n241_), .C(men_men_n240_), .D(men_men_n239_), .Y(men_men_n243_));
  OAI210     u227(.A0(men_men_n243_), .A1(men_men_n236_), .B0(x2), .Y(men_men_n244_));
  NA3        u228(.A(men_men_n244_), .B(men_men_n234_), .C(men_men_n230_), .Y(men_men_n245_));
  AOI210     u229(.A0(men_men_n221_), .A1(x8), .B0(men_men_n245_), .Y(men_men_n246_));
  NO2        u230(.A(men_men_n93_), .B(x3), .Y(men_men_n247_));
  NA2        u231(.A(men_men_n247_), .B(men_men_n206_), .Y(men_men_n248_));
  NO3        u232(.A(men_men_n91_), .B(men_men_n78_), .C(men_men_n25_), .Y(men_men_n249_));
  AOI210     u233(.A0(men_men_n225_), .A1(men_men_n157_), .B0(men_men_n249_), .Y(men_men_n250_));
  AOI210     u234(.A0(men_men_n250_), .A1(men_men_n248_), .B0(x2), .Y(men_men_n251_));
  NO2        u235(.A(x4), .B(men_men_n54_), .Y(men_men_n252_));
  AOI220     u236(.A0(men_men_n206_), .A1(men_men_n189_), .B0(men_men_n252_), .B1(men_men_n66_), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n62_), .B(x6), .Y(men_men_n254_));
  NA3        u238(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n255_), .A1(men_men_n140_), .B0(men_men_n254_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n257_));
  NO2        u241(.A(men_men_n257_), .B(men_men_n25_), .Y(men_men_n258_));
  OAI210     u242(.A0(men_men_n258_), .A1(men_men_n256_), .B0(men_men_n122_), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n209_), .B(x6), .Y(men_men_n260_));
  NO2        u244(.A(men_men_n209_), .B(x6), .Y(men_men_n261_));
  INV        u245(.A(men_men_n261_), .Y(men_men_n262_));
  NA3        u246(.A(men_men_n262_), .B(men_men_n260_), .C(men_men_n145_), .Y(men_men_n263_));
  NA4        u247(.A(men_men_n263_), .B(men_men_n259_), .C(men_men_n253_), .D(men_men_n154_), .Y(men_men_n264_));
  NA2        u248(.A(men_men_n198_), .B(men_men_n224_), .Y(men_men_n265_));
  NO2        u249(.A(x9), .B(x6), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n140_), .B(men_men_n18_), .Y(men_men_n267_));
  NAi21      u251(.An(men_men_n267_), .B(men_men_n255_), .Y(men_men_n268_));
  NAi21      u252(.An(x1), .B(x4), .Y(men_men_n269_));
  AOI210     u253(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n270_));
  OAI210     u254(.A0(men_men_n140_), .A1(x3), .B0(men_men_n270_), .Y(men_men_n271_));
  AOI220     u255(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n268_), .B1(men_men_n266_), .Y(men_men_n272_));
  NA2        u256(.A(men_men_n272_), .B(men_men_n265_), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n62_), .B(x2), .Y(men_men_n274_));
  NO2        u258(.A(men_men_n274_), .B(men_men_n265_), .Y(men_men_n275_));
  NO3        u259(.A(x9), .B(x6), .C(x0), .Y(men_men_n276_));
  NA2        u260(.A(x6), .B(x2), .Y(men_men_n277_));
  NO2        u261(.A(men_men_n277_), .B(men_men_n172_), .Y(men_men_n278_));
  NO2        u262(.A(men_men_n276_), .B(men_men_n278_), .Y(men_men_n279_));
  OAI220     u263(.A0(men_men_n279_), .A1(men_men_n43_), .B0(men_men_n178_), .B1(men_men_n46_), .Y(men_men_n280_));
  OAI210     u264(.A0(men_men_n280_), .A1(men_men_n275_), .B0(men_men_n273_), .Y(men_men_n281_));
  NO2        u265(.A(x3), .B(men_men_n205_), .Y(men_men_n282_));
  NA2        u266(.A(x4), .B(x0), .Y(men_men_n283_));
  NO3        u267(.A(men_men_n72_), .B(men_men_n283_), .C(x6), .Y(men_men_n284_));
  AOI210     u268(.A0(men_men_n282_), .A1(men_men_n42_), .B0(men_men_n284_), .Y(men_men_n285_));
  AOI210     u269(.A0(men_men_n285_), .A1(men_men_n281_), .B0(x8), .Y(men_men_n286_));
  INV        u270(.A(men_men_n254_), .Y(men_men_n287_));
  OAI210     u271(.A0(men_men_n267_), .A1(men_men_n216_), .B0(men_men_n287_), .Y(men_men_n288_));
  INV        u272(.A(men_men_n176_), .Y(men_men_n289_));
  OAI210     u273(.A0(men_men_n289_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n290_), .A1(men_men_n288_), .B0(men_men_n231_), .Y(men_men_n291_));
  NO4        u275(.A(men_men_n291_), .B(men_men_n286_), .C(men_men_n264_), .D(men_men_n251_), .Y(men_men_n292_));
  NO2        u276(.A(men_men_n165_), .B(x1), .Y(men_men_n293_));
  NO3        u277(.A(men_men_n293_), .B(x3), .C(men_men_n36_), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n294_), .A1(men_men_n261_), .B0(x2), .Y(men_men_n295_));
  OAI210     u279(.A0(men_men_n289_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n296_));
  AOI210     u280(.A0(men_men_n296_), .A1(men_men_n295_), .B0(men_men_n188_), .Y(men_men_n297_));
  NOi21      u281(.An(men_men_n277_), .B(men_men_n17_), .Y(men_men_n298_));
  NA3        u282(.A(men_men_n298_), .B(men_men_n216_), .C(men_men_n40_), .Y(men_men_n299_));
  AOI210     u283(.A0(men_men_n36_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n300_));
  NA3        u284(.A(men_men_n300_), .B(men_men_n163_), .C(men_men_n32_), .Y(men_men_n301_));
  NA2        u285(.A(x3), .B(x2), .Y(men_men_n302_));
  AOI220     u286(.A0(men_men_n302_), .A1(men_men_n231_), .B0(men_men_n301_), .B1(men_men_n299_), .Y(men_men_n303_));
  NAi21      u287(.An(x4), .B(x0), .Y(men_men_n304_));
  NO3        u288(.A(men_men_n304_), .B(men_men_n44_), .C(x2), .Y(men_men_n305_));
  OAI210     u289(.A0(x6), .A1(men_men_n18_), .B0(men_men_n305_), .Y(men_men_n306_));
  OAI220     u290(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n307_));
  NO2        u291(.A(x9), .B(x8), .Y(men_men_n308_));
  NA2        u292(.A(men_men_n36_), .B(men_men_n54_), .Y(men_men_n309_));
  OAI210     u293(.A0(men_men_n300_), .A1(men_men_n298_), .B0(men_men_n309_), .Y(men_men_n310_));
  AOI220     u294(.A0(men_men_n310_), .A1(men_men_n81_), .B0(men_men_n307_), .B1(men_men_n31_), .Y(men_men_n311_));
  AOI210     u295(.A0(men_men_n311_), .A1(men_men_n306_), .B0(men_men_n25_), .Y(men_men_n312_));
  NA3        u296(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n313_));
  OAI210     u297(.A0(men_men_n300_), .A1(men_men_n298_), .B0(men_men_n313_), .Y(men_men_n314_));
  INV        u298(.A(men_men_n218_), .Y(men_men_n315_));
  NA2        u299(.A(men_men_n36_), .B(men_men_n43_), .Y(men_men_n316_));
  OR2        u300(.A(men_men_n316_), .B(men_men_n283_), .Y(men_men_n317_));
  OAI220     u301(.A0(men_men_n317_), .A1(men_men_n162_), .B0(men_men_n235_), .B1(men_men_n315_), .Y(men_men_n318_));
  AO210      u302(.A0(men_men_n314_), .A1(men_men_n149_), .B0(men_men_n318_), .Y(men_men_n319_));
  NO4        u303(.A(men_men_n319_), .B(men_men_n312_), .C(men_men_n303_), .D(men_men_n297_), .Y(men_men_n320_));
  OAI210     u304(.A0(men_men_n292_), .A1(men_men_n246_), .B0(men_men_n320_), .Y(men04));
  OAI210     u305(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n322_));
  NA3        u306(.A(men_men_n322_), .B(men_men_n276_), .C(men_men_n84_), .Y(men_men_n323_));
  NO2        u307(.A(x2), .B(x1), .Y(men_men_n324_));
  OAI210     u308(.A0(men_men_n257_), .A1(men_men_n324_), .B0(men_men_n36_), .Y(men_men_n325_));
  NO2        u309(.A(men_men_n324_), .B(men_men_n304_), .Y(men_men_n326_));
  AOI210     u310(.A0(men_men_n62_), .A1(x4), .B0(men_men_n114_), .Y(men_men_n327_));
  OAI210     u311(.A0(men_men_n327_), .A1(men_men_n326_), .B0(men_men_n247_), .Y(men_men_n328_));
  NO2        u312(.A(men_men_n274_), .B(men_men_n91_), .Y(men_men_n329_));
  NA3        u313(.A(men_men_n91_), .B(x6), .C(men_men_n328_), .Y(men_men_n330_));
  NA2        u314(.A(men_men_n330_), .B(men_men_n325_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n211_), .B(men_men_n115_), .Y(men_men_n332_));
  NO3        u316(.A(men_men_n254_), .B(men_men_n121_), .C(men_men_n18_), .Y(men_men_n333_));
  NO2        u317(.A(men_men_n333_), .B(men_men_n332_), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n120_), .A1(men_men_n108_), .B0(men_men_n176_), .Y(men_men_n335_));
  NA3        u319(.A(men_men_n335_), .B(x6), .C(x3), .Y(men_men_n336_));
  NOi21      u320(.An(men_men_n151_), .B(men_men_n131_), .Y(men_men_n337_));
  AOI210     u321(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n338_), .B(men_men_n316_), .Y(men_men_n339_));
  AOI210     u323(.A0(men_men_n337_), .A1(men_men_n63_), .B0(men_men_n339_), .Y(men_men_n340_));
  NA2        u324(.A(men_men_n329_), .B(men_men_n93_), .Y(men_men_n341_));
  NA4        u325(.A(men_men_n341_), .B(men_men_n340_), .C(men_men_n336_), .D(men_men_n334_), .Y(men_men_n342_));
  OAI210     u326(.A0(men_men_n113_), .A1(x3), .B0(men_men_n305_), .Y(men_men_n343_));
  NA3        u327(.A(men_men_n227_), .B(men_men_n215_), .C(men_men_n83_), .Y(men_men_n344_));
  NA3        u328(.A(men_men_n344_), .B(men_men_n343_), .C(men_men_n154_), .Y(men_men_n345_));
  AOI210     u329(.A0(men_men_n342_), .A1(x4), .B0(men_men_n345_), .Y(men_men_n346_));
  NA3        u330(.A(men_men_n326_), .B(men_men_n211_), .C(men_men_n93_), .Y(men_men_n347_));
  XO2        u331(.A(x4), .B(x0), .Y(men_men_n348_));
  OAI210     u332(.A0(men_men_n348_), .A1(men_men_n119_), .B0(men_men_n269_), .Y(men_men_n349_));
  NA2        u333(.A(men_men_n349_), .B(x8), .Y(men_men_n350_));
  AOI210     u334(.A0(men_men_n350_), .A1(men_men_n347_), .B0(x3), .Y(men_men_n351_));
  INV        u335(.A(men_men_n94_), .Y(men_men_n352_));
  NO2        u336(.A(men_men_n93_), .B(x4), .Y(men_men_n353_));
  AOI220     u337(.A0(men_men_n353_), .A1(men_men_n44_), .B0(men_men_n125_), .B1(men_men_n352_), .Y(men_men_n354_));
  NO3        u338(.A(men_men_n348_), .B(men_men_n165_), .C(x2), .Y(men_men_n355_));
  NO3        u339(.A(men_men_n227_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n356_));
  NO2        u340(.A(men_men_n356_), .B(men_men_n355_), .Y(men_men_n357_));
  NA4        u341(.A(men_men_n357_), .B(men_men_n354_), .C(men_men_n223_), .D(x6), .Y(men_men_n358_));
  NO2        u342(.A(men_men_n181_), .B(men_men_n93_), .Y(men_men_n359_));
  NO2        u343(.A(men_men_n43_), .B(x0), .Y(men_men_n360_));
  OR2        u344(.A(men_men_n353_), .B(men_men_n360_), .Y(men_men_n361_));
  NO2        u345(.A(men_men_n151_), .B(men_men_n108_), .Y(men_men_n362_));
  AOI220     u346(.A0(men_men_n362_), .A1(men_men_n361_), .B0(men_men_n359_), .B1(men_men_n61_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n363_), .B(men_men_n62_), .Y(men_men_n364_));
  OAI220     u348(.A0(men_men_n364_), .A1(x6), .B0(men_men_n358_), .B1(men_men_n351_), .Y(men_men_n365_));
  OAI210     u349(.A0(men_men_n63_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n366_));
  OAI210     u350(.A0(men_men_n366_), .A1(men_men_n93_), .B0(men_men_n317_), .Y(men_men_n367_));
  AOI210     u351(.A0(men_men_n367_), .A1(men_men_n18_), .B0(men_men_n154_), .Y(men_men_n368_));
  AO220      u352(.A0(men_men_n368_), .A1(men_men_n365_), .B0(men_men_n346_), .B1(men_men_n331_), .Y(men_men_n369_));
  NA2        u353(.A(men_men_n369_), .B(men_men_n323_), .Y(men_men_n370_));
  NA3        u354(.A(x7), .B(x3), .C(x0), .Y(men_men_n371_));
  NA2        u355(.A(men_men_n222_), .B(x0), .Y(men_men_n372_));
  OAI220     u356(.A0(men_men_n372_), .A1(men_men_n211_), .B0(men_men_n371_), .B1(men_men_n352_), .Y(men_men_n373_));
  INV        u357(.A(men_men_n373_), .Y(men_men_n374_));
  NO2        u358(.A(men_men_n374_), .B(men_men_n25_), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n197_), .A1(men_men_n67_), .B0(men_men_n440_), .Y(men_men_n376_));
  NA3        u360(.A(men_men_n200_), .B(men_men_n224_), .C(x8), .Y(men_men_n377_));
  AOI210     u361(.A0(men_men_n377_), .A1(men_men_n376_), .B0(men_men_n25_), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n121_), .A1(men_men_n120_), .B0(men_men_n42_), .Y(men_men_n379_));
  NOi31      u363(.An(men_men_n379_), .B(men_men_n360_), .C(men_men_n182_), .Y(men_men_n380_));
  OAI210     u364(.A0(men_men_n380_), .A1(men_men_n378_), .B0(men_men_n150_), .Y(men_men_n381_));
  INV        u365(.A(men_men_n381_), .Y(men_men_n382_));
  OAI210     u366(.A0(men_men_n382_), .A1(men_men_n375_), .B0(x6), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n439_), .A1(x0), .B0(men_men_n32_), .Y(men_men_n384_));
  AOI210     u368(.A0(men_men_n127_), .A1(men_men_n252_), .B0(x1), .Y(men_men_n385_));
  INV        u369(.A(men_men_n385_), .Y(men_men_n386_));
  NAi31      u370(.An(x2), .B(x8), .C(x0), .Y(men_men_n387_));
  OAI210     u371(.A0(men_men_n387_), .A1(x4), .B0(men_men_n166_), .Y(men_men_n388_));
  NA3        u372(.A(men_men_n388_), .B(men_men_n148_), .C(x9), .Y(men_men_n389_));
  NO4        u373(.A(men_men_n126_), .B(men_men_n304_), .C(x9), .D(x2), .Y(men_men_n390_));
  NOi21      u374(.An(men_men_n124_), .B(men_men_n181_), .Y(men_men_n391_));
  NO3        u375(.A(men_men_n391_), .B(men_men_n390_), .C(men_men_n18_), .Y(men_men_n392_));
  NA3        u376(.A(men_men_n392_), .B(men_men_n389_), .C(men_men_n50_), .Y(men_men_n393_));
  OAI210     u377(.A0(men_men_n386_), .A1(men_men_n384_), .B0(men_men_n393_), .Y(men_men_n394_));
  AOI210     u378(.A0(men_men_n38_), .A1(x9), .B0(men_men_n134_), .Y(men_men_n395_));
  NO3        u379(.A(men_men_n395_), .B(men_men_n124_), .C(men_men_n43_), .Y(men_men_n396_));
  AOI210     u380(.A0(men_men_n269_), .A1(men_men_n60_), .B0(men_men_n123_), .Y(men_men_n397_));
  NO2        u381(.A(men_men_n397_), .B(x3), .Y(men_men_n398_));
  NO3        u382(.A(men_men_n398_), .B(men_men_n396_), .C(x2), .Y(men_men_n399_));
  OAI220     u383(.A0(men_men_n348_), .A1(men_men_n308_), .B0(men_men_n304_), .B1(men_men_n43_), .Y(men_men_n400_));
  AOI210     u384(.A0(x9), .A1(men_men_n48_), .B0(men_men_n371_), .Y(men_men_n401_));
  AOI220     u385(.A0(men_men_n401_), .A1(men_men_n93_), .B0(men_men_n400_), .B1(men_men_n154_), .Y(men_men_n402_));
  NO2        u386(.A(men_men_n402_), .B(men_men_n54_), .Y(men_men_n403_));
  NO2        u387(.A(men_men_n403_), .B(men_men_n399_), .Y(men_men_n404_));
  AOI210     u388(.A0(men_men_n404_), .A1(men_men_n394_), .B0(men_men_n25_), .Y(men_men_n405_));
  NA4        u389(.A(men_men_n31_), .B(men_men_n93_), .C(x2), .D(men_men_n17_), .Y(men_men_n406_));
  NO3        u390(.A(men_men_n67_), .B(men_men_n18_), .C(x0), .Y(men_men_n407_));
  AOI220     u391(.A0(men_men_n407_), .A1(men_men_n270_), .B0(men_men_n441_), .B1(men_men_n379_), .Y(men_men_n408_));
  NO2        u392(.A(men_men_n408_), .B(men_men_n105_), .Y(men_men_n409_));
  NO3        u393(.A(men_men_n274_), .B(men_men_n176_), .C(men_men_n40_), .Y(men_men_n410_));
  OAI210     u394(.A0(men_men_n410_), .A1(men_men_n409_), .B0(x7), .Y(men_men_n411_));
  NA2        u395(.A(men_men_n227_), .B(x7), .Y(men_men_n412_));
  NA3        u396(.A(men_men_n412_), .B(men_men_n153_), .C(men_men_n135_), .Y(men_men_n413_));
  NA3        u397(.A(men_men_n413_), .B(men_men_n411_), .C(men_men_n406_), .Y(men_men_n414_));
  OAI210     u398(.A0(men_men_n414_), .A1(men_men_n405_), .B0(men_men_n36_), .Y(men_men_n415_));
  NA2        u399(.A(men_men_n257_), .B(men_men_n21_), .Y(men_men_n416_));
  NO2        u400(.A(men_men_n162_), .B(men_men_n136_), .Y(men_men_n417_));
  NA2        u401(.A(men_men_n417_), .B(men_men_n416_), .Y(men_men_n418_));
  AOI210     u402(.A0(men_men_n418_), .A1(men_men_n167_), .B0(men_men_n28_), .Y(men_men_n419_));
  AOI220     u403(.A0(men_men_n360_), .A1(men_men_n93_), .B0(men_men_n151_), .B1(men_men_n200_), .Y(men_men_n420_));
  NA3        u404(.A(men_men_n420_), .B(men_men_n387_), .C(men_men_n91_), .Y(men_men_n421_));
  NA2        u405(.A(men_men_n421_), .B(men_men_n177_), .Y(men_men_n422_));
  OAI220     u406(.A0(x3), .A1(men_men_n68_), .B0(men_men_n162_), .B1(men_men_n43_), .Y(men_men_n423_));
  NA2        u407(.A(x3), .B(men_men_n54_), .Y(men_men_n424_));
  AOI210     u408(.A0(men_men_n166_), .A1(men_men_n27_), .B0(men_men_n72_), .Y(men_men_n425_));
  OAI210     u409(.A0(men_men_n150_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n426_));
  NO2        u410(.A(x3), .B(men_men_n54_), .Y(men_men_n427_));
  AOI210     u411(.A0(men_men_n427_), .A1(men_men_n426_), .B0(men_men_n425_), .Y(men_men_n428_));
  OAI210     u412(.A0(men_men_n155_), .A1(men_men_n424_), .B0(men_men_n428_), .Y(men_men_n429_));
  AOI220     u413(.A0(men_men_n429_), .A1(x0), .B0(men_men_n423_), .B1(men_men_n136_), .Y(men_men_n430_));
  AOI210     u414(.A0(men_men_n430_), .A1(men_men_n422_), .B0(men_men_n235_), .Y(men_men_n431_));
  NA2        u415(.A(x9), .B(x5), .Y(men_men_n432_));
  NO4        u416(.A(men_men_n108_), .B(men_men_n432_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n433_));
  NO3        u417(.A(men_men_n433_), .B(men_men_n431_), .C(men_men_n419_), .Y(men_men_n434_));
  NA3        u418(.A(men_men_n434_), .B(men_men_n415_), .C(men_men_n383_), .Y(men_men_n435_));
  AOI210     u419(.A0(men_men_n370_), .A1(men_men_n25_), .B0(men_men_n435_), .Y(men05));
  INV        u420(.A(men_men_n38_), .Y(men_men_n439_));
  INV        u421(.A(x0), .Y(men_men_n440_));
  INV        u422(.A(x4), .Y(men_men_n441_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule