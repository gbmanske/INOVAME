// Benchmark "top" written by ABC on Thu Jun 20 14:00:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n143_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n781_,
    new_new_n782_, new_new_n783_, new_new_n784_, new_new_n785_,
    new_new_n786_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n827_, new_new_n828_, new_new_n829_, new_new_n830_,
    new_new_n831_, new_new_n832_, new_new_n833_, new_new_n834_,
    new_new_n835_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n881_, new_new_n882_, new_new_n883_,
    new_new_n884_, new_new_n885_, new_new_n886_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1107_, new_new_n1108_,
    new_new_n1109_, new_new_n1110_, new_new_n1114_, new_new_n1115_,
    new_new_n1116_, new_new_n1117_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(zz01));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  OR4        g0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g0066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  AOI210     g0067(.A0(new_new_n88_), .A1(new_new_n86_), .B0(new_new_n89_), .Y(new_new_n90_));
  OAI210     g0068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g0069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g0070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g0072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g0073(.A(new_new_n95_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g0074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g0075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n98_));
  AN3        g0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g0077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g0078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g0079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g0080(.A0(new_new_n102_), .A1(new_new_n62_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g0081(.A(i_7_), .Y(new_new_n104_));
  NA2        g0082(.A(new_new_n47_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g0083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g0084(.A(new_new_n106_), .B(new_new_n86_), .Y(new_new_n107_));
  NA2        g0085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g0086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g0087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g0088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  NO3        g0089(.A(new_new_n111_), .B(new_new_n92_), .C(new_new_n54_), .Y(new_new_n112_));
  AN2        g0090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g0092(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n115_));
  NO2        g0093(.A(i_8_), .B(new_new_n104_), .Y(new_new_n116_));
  NO3        g0094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g0095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g0097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  INV        g0098(.A(new_new_n120_), .Y(new_new_n121_));
  NO2        g0099(.A(new_new_n121_), .B(new_new_n117_), .Y(new_new_n122_));
  NAi41      g0100(.An(new_new_n112_), .B(new_new_n122_), .C(new_new_n110_), .D(new_new_n103_), .Y(new_new_n123_));
  NOi21      g0101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g0104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g0106(.A(new_new_n128_), .B(new_new_n47_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n130_));
  NAi21      g0108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(new_new_n62_), .Y(new_new_n132_));
  NOi31      g0110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g0111(.A(i_1_), .B(new_new_n86_), .Y(new_new_n134_));
  NO2        g0112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g0113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g0114(.A0(new_new_n136_), .A1(new_new_n48_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g0115(.A0(new_new_n137_), .A1(new_new_n111_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g0116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n98_), .Y(new_new_n139_));
  NA3        g0117(.A(new_new_n139_), .B(new_new_n79_), .C(new_new_n56_), .Y(zz02));
  NO2        g0118(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g0119(.A(i_6_), .B(new_new_n25_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(new_new_n141_), .Y(new_new_n143_));
  NA4        g0121(.A(new_new_n143_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(zz00));
  AN2        g0122(.A(i_8_), .B(i_7_), .Y(new_new_n145_));
  NA2        g0123(.A(new_new_n145_), .B(i_6_), .Y(new_new_n146_));
  NO2        g0124(.A(i_12_), .B(i_13_), .Y(new_new_n147_));
  NAi21      g0125(.An(i_5_), .B(i_11_), .Y(new_new_n148_));
  NOi21      g0126(.An(new_new_n147_), .B(new_new_n148_), .Y(new_new_n149_));
  NO2        g0127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NA2        g0128(.A(i_2_), .B(i_3_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(i_4_), .Y(new_new_n152_));
  NA3        g0130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  OR2        g0131(.A(new_new_n153_), .B(new_new_n25_), .Y(new_new_n154_));
  AN2        g0132(.A(new_new_n147_), .B(new_new_n83_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n155_), .B(new_new_n27_), .Y(new_new_n156_));
  NA2        g0134(.A(i_1_), .B(i_5_), .Y(new_new_n157_));
  NO2        g0135(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n158_));
  NA2        g0136(.A(new_new_n158_), .B(new_new_n36_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n157_), .C(new_new_n156_), .Y(new_new_n160_));
  OR2        g0138(.A(i_0_), .B(i_1_), .Y(new_new_n161_));
  NO3        g0139(.A(new_new_n161_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n162_));
  NAi32      g0140(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n163_));
  NAi21      g0141(.An(new_new_n163_), .B(new_new_n162_), .Y(new_new_n164_));
  NOi21      g0142(.An(i_4_), .B(i_10_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n40_), .Y(new_new_n166_));
  NO2        g0144(.A(i_3_), .B(i_5_), .Y(new_new_n167_));
  NO3        g0145(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n168_));
  NA2        g0146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  OAI210     g0147(.A0(new_new_n169_), .A1(new_new_n166_), .B0(new_new_n164_), .Y(new_new_n170_));
  NO2        g0148(.A(new_new_n170_), .B(new_new_n160_), .Y(new_new_n171_));
  AOI210     g0149(.A0(new_new_n171_), .A1(new_new_n154_), .B0(new_new_n146_), .Y(new_new_n172_));
  NA3        g0150(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n173_));
  NA2        g0151(.A(i_3_), .B(new_new_n49_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_4_), .B(i_9_), .Y(new_new_n175_));
  NOi21      g0153(.An(i_11_), .B(i_13_), .Y(new_new_n176_));
  NA2        g0154(.A(new_new_n176_), .B(new_new_n175_), .Y(new_new_n177_));
  OR2        g0155(.A(new_new_n177_), .B(new_new_n174_), .Y(new_new_n178_));
  NO2        g0156(.A(i_4_), .B(i_5_), .Y(new_new_n179_));
  NAi21      g0157(.An(i_12_), .B(i_11_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n180_), .B(i_13_), .Y(new_new_n181_));
  NA3        g0159(.A(new_new_n181_), .B(new_new_n179_), .C(new_new_n83_), .Y(new_new_n182_));
  AOI210     g0160(.A0(new_new_n182_), .A1(new_new_n178_), .B0(new_new_n173_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n184_), .B(new_new_n47_), .Y(new_new_n185_));
  NA2        g0163(.A(new_new_n36_), .B(i_5_), .Y(new_new_n186_));
  NAi31      g0164(.An(new_new_n186_), .B(new_new_n155_), .C(i_11_), .Y(new_new_n187_));
  NA2        g0165(.A(i_3_), .B(i_5_), .Y(new_new_n188_));
  OR2        g0166(.A(new_new_n188_), .B(new_new_n177_), .Y(new_new_n189_));
  AOI210     g0167(.A0(new_new_n189_), .A1(new_new_n187_), .B0(new_new_n185_), .Y(new_new_n190_));
  NO2        g0168(.A(new_new_n73_), .B(i_5_), .Y(new_new_n191_));
  NO2        g0169(.A(i_13_), .B(i_10_), .Y(new_new_n192_));
  NA3        g0170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n45_), .Y(new_new_n193_));
  NO2        g0171(.A(i_2_), .B(i_1_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(i_3_), .Y(new_new_n195_));
  NAi21      g0173(.An(i_4_), .B(i_12_), .Y(new_new_n196_));
  NO4        g0174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n193_), .D(new_new_n25_), .Y(new_new_n197_));
  NO3        g0175(.A(new_new_n197_), .B(new_new_n190_), .C(new_new_n183_), .Y(new_new_n198_));
  INV        g0176(.A(i_8_), .Y(new_new_n199_));
  NO2        g0177(.A(new_new_n199_), .B(i_7_), .Y(new_new_n200_));
  NA2        g0178(.A(new_new_n200_), .B(i_6_), .Y(new_new_n201_));
  NO3        g0179(.A(i_3_), .B(new_new_n86_), .C(new_new_n49_), .Y(new_new_n202_));
  NA2        g0180(.A(new_new_n202_), .B(new_new_n116_), .Y(new_new_n203_));
  NO3        g0181(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n206_));
  OAI210     g0184(.A0(new_new_n99_), .A1(i_12_), .B0(new_new_n206_), .Y(new_new_n207_));
  AOI210     g0185(.A0(new_new_n207_), .A1(new_new_n205_), .B0(new_new_n203_), .Y(new_new_n208_));
  NO2        g0186(.A(i_3_), .B(i_8_), .Y(new_new_n209_));
  NO3        g0187(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n210_));
  NA3        g0188(.A(new_new_n210_), .B(new_new_n209_), .C(new_new_n40_), .Y(new_new_n211_));
  NO2        g0189(.A(new_new_n106_), .B(new_new_n58_), .Y(new_new_n212_));
  NA2        g0190(.A(new_new_n212_), .B(new_new_n161_), .Y(new_new_n213_));
  NO2        g0191(.A(i_13_), .B(i_9_), .Y(new_new_n214_));
  NA3        g0192(.A(new_new_n214_), .B(i_6_), .C(new_new_n199_), .Y(new_new_n215_));
  NAi21      g0193(.An(i_12_), .B(i_3_), .Y(new_new_n216_));
  OR2        g0194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n45_), .B(i_5_), .Y(new_new_n218_));
  NO3        g0196(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n219_));
  NA3        g0197(.A(new_new_n219_), .B(new_new_n218_), .C(i_10_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n220_), .A1(new_new_n217_), .B0(new_new_n213_), .B1(new_new_n211_), .Y(new_new_n221_));
  AOI210     g0199(.A0(new_new_n221_), .A1(i_7_), .B0(new_new_n208_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(i_4_), .B0(new_new_n201_), .B1(new_new_n198_), .Y(new_new_n223_));
  NAi21      g0201(.An(i_12_), .B(i_7_), .Y(new_new_n224_));
  NA3        g0202(.A(i_13_), .B(new_new_n199_), .C(i_10_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  NA2        g0204(.A(i_0_), .B(i_5_), .Y(new_new_n227_));
  NA2        g0205(.A(new_new_n227_), .B(new_new_n107_), .Y(new_new_n228_));
  OAI220     g0206(.A0(new_new_n228_), .A1(new_new_n195_), .B0(new_new_n185_), .B1(new_new_n136_), .Y(new_new_n229_));
  NAi31      g0207(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n36_), .B(i_13_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n233_));
  NA3        g0211(.A(new_new_n233_), .B(new_new_n232_), .C(new_new_n231_), .Y(new_new_n234_));
  INV        g0212(.A(i_13_), .Y(new_new_n235_));
  NO2        g0213(.A(i_12_), .B(new_new_n235_), .Y(new_new_n236_));
  NA3        g0214(.A(new_new_n236_), .B(new_new_n204_), .C(new_new_n202_), .Y(new_new_n237_));
  OAI210     g0215(.A0(new_new_n234_), .A1(new_new_n230_), .B0(new_new_n237_), .Y(new_new_n238_));
  AOI220     g0216(.A0(new_new_n238_), .A1(new_new_n145_), .B0(new_new_n229_), .B1(new_new_n226_), .Y(new_new_n239_));
  NO2        g0217(.A(i_12_), .B(new_new_n37_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n188_), .B(i_4_), .Y(new_new_n241_));
  NA2        g0219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  OR2        g0220(.A(i_8_), .B(i_7_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n243_), .B(new_new_n86_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n54_), .B(i_1_), .Y(new_new_n245_));
  NA2        g0223(.A(new_new_n245_), .B(new_new_n244_), .Y(new_new_n246_));
  INV        g0224(.A(i_12_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n45_), .B(new_new_n247_), .Y(new_new_n248_));
  NO3        g0226(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n249_));
  NA2        g0227(.A(i_2_), .B(i_1_), .Y(new_new_n250_));
  NO2        g0228(.A(new_new_n246_), .B(new_new_n242_), .Y(new_new_n251_));
  NO3        g0229(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n252_));
  NAi21      g0230(.An(i_4_), .B(i_3_), .Y(new_new_n253_));
  NO2        g0231(.A(new_new_n253_), .B(new_new_n75_), .Y(new_new_n254_));
  NO2        g0232(.A(i_0_), .B(i_6_), .Y(new_new_n255_));
  NOi41      g0233(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n256_), .B(new_new_n255_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n250_), .B(new_new_n188_), .Y(new_new_n258_));
  NAi21      g0236(.An(new_new_n257_), .B(new_new_n258_), .Y(new_new_n259_));
  INV        g0237(.A(new_new_n259_), .Y(new_new_n260_));
  AOI220     g0238(.A0(new_new_n260_), .A1(new_new_n40_), .B0(new_new_n251_), .B1(new_new_n214_), .Y(new_new_n261_));
  NO2        g0239(.A(i_11_), .B(new_new_n235_), .Y(new_new_n262_));
  NOi21      g0240(.An(i_1_), .B(i_6_), .Y(new_new_n263_));
  NAi21      g0241(.An(i_3_), .B(i_7_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n247_), .B(i_9_), .Y(new_new_n265_));
  OR4        g0243(.A(new_new_n265_), .B(new_new_n264_), .C(new_new_n263_), .D(new_new_n191_), .Y(new_new_n266_));
  NO2        g0244(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n267_));
  NO2        g0245(.A(i_12_), .B(i_3_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n73_), .B(i_5_), .Y(new_new_n269_));
  NA2        g0247(.A(i_3_), .B(i_9_), .Y(new_new_n270_));
  NAi21      g0248(.An(i_7_), .B(i_10_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n270_), .Y(new_new_n272_));
  NA3        g0250(.A(new_new_n272_), .B(new_new_n269_), .C(new_new_n64_), .Y(new_new_n273_));
  NA2        g0251(.A(new_new_n273_), .B(new_new_n266_), .Y(new_new_n274_));
  NA3        g0252(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n275_));
  INV        g0253(.A(new_new_n146_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n247_), .B(i_13_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n277_), .B(new_new_n75_), .Y(new_new_n278_));
  AOI220     g0256(.A0(new_new_n278_), .A1(new_new_n276_), .B0(new_new_n274_), .B1(new_new_n262_), .Y(new_new_n279_));
  NO2        g0257(.A(new_new_n243_), .B(new_new_n37_), .Y(new_new_n280_));
  NA2        g0258(.A(i_12_), .B(i_6_), .Y(new_new_n281_));
  OR2        g0259(.A(i_13_), .B(i_9_), .Y(new_new_n282_));
  NO3        g0260(.A(new_new_n282_), .B(new_new_n281_), .C(new_new_n49_), .Y(new_new_n283_));
  NO2        g0261(.A(new_new_n253_), .B(i_2_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(new_new_n283_), .C(new_new_n45_), .Y(new_new_n285_));
  NA2        g0263(.A(new_new_n262_), .B(i_9_), .Y(new_new_n286_));
  NA3        g0264(.A(new_new_n269_), .B(new_new_n161_), .C(new_new_n64_), .Y(new_new_n287_));
  OAI210     g0265(.A0(new_new_n287_), .A1(new_new_n286_), .B0(new_new_n285_), .Y(new_new_n288_));
  NA2        g0266(.A(new_new_n158_), .B(new_new_n63_), .Y(new_new_n289_));
  NO3        g0267(.A(i_11_), .B(new_new_n235_), .C(new_new_n25_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n264_), .B(i_8_), .Y(new_new_n291_));
  NO2        g0269(.A(i_6_), .B(new_new_n49_), .Y(new_new_n292_));
  NA3        g0270(.A(new_new_n292_), .B(new_new_n291_), .C(new_new_n290_), .Y(new_new_n293_));
  NO3        g0271(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n294_));
  NA3        g0272(.A(new_new_n294_), .B(new_new_n280_), .C(new_new_n236_), .Y(new_new_n295_));
  AOI210     g0273(.A0(new_new_n295_), .A1(new_new_n293_), .B0(new_new_n289_), .Y(new_new_n296_));
  AOI210     g0274(.A0(new_new_n288_), .A1(new_new_n280_), .B0(new_new_n296_), .Y(new_new_n297_));
  NA4        g0275(.A(new_new_n297_), .B(new_new_n279_), .C(new_new_n261_), .D(new_new_n239_), .Y(new_new_n298_));
  NO3        g0276(.A(i_12_), .B(new_new_n235_), .C(new_new_n37_), .Y(new_new_n299_));
  INV        g0277(.A(new_new_n299_), .Y(new_new_n300_));
  NA2        g0278(.A(i_8_), .B(new_new_n104_), .Y(new_new_n301_));
  NOi21      g0279(.An(new_new_n167_), .B(new_new_n86_), .Y(new_new_n302_));
  NO3        g0280(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n303_));
  AOI220     g0281(.A0(new_new_n303_), .A1(new_new_n202_), .B0(new_new_n302_), .B1(new_new_n245_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n304_), .B(new_new_n301_), .Y(new_new_n305_));
  NO3        g0283(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n306_));
  NO2        g0284(.A(new_new_n250_), .B(i_0_), .Y(new_new_n307_));
  AOI220     g0285(.A0(new_new_n307_), .A1(new_new_n200_), .B0(new_new_n306_), .B1(new_new_n145_), .Y(new_new_n308_));
  NA2        g0286(.A(new_new_n292_), .B(new_new_n26_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n309_), .B(new_new_n308_), .Y(new_new_n310_));
  NA2        g0288(.A(i_0_), .B(i_1_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n311_), .B(i_2_), .Y(new_new_n312_));
  NO2        g0290(.A(new_new_n59_), .B(i_6_), .Y(new_new_n313_));
  NA3        g0291(.A(new_new_n313_), .B(new_new_n312_), .C(new_new_n167_), .Y(new_new_n314_));
  OAI210     g0292(.A0(new_new_n169_), .A1(new_new_n146_), .B0(new_new_n314_), .Y(new_new_n315_));
  NO3        g0293(.A(new_new_n315_), .B(new_new_n310_), .C(new_new_n305_), .Y(new_new_n316_));
  NO2        g0294(.A(i_3_), .B(i_10_), .Y(new_new_n317_));
  NA3        g0295(.A(new_new_n317_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n318_));
  NO2        g0296(.A(i_2_), .B(new_new_n104_), .Y(new_new_n319_));
  NA2        g0297(.A(i_1_), .B(new_new_n36_), .Y(new_new_n320_));
  NO2        g0298(.A(new_new_n320_), .B(i_8_), .Y(new_new_n321_));
  NOi21      g0299(.An(new_new_n227_), .B(new_new_n106_), .Y(new_new_n322_));
  NA3        g0300(.A(new_new_n322_), .B(new_new_n321_), .C(new_new_n319_), .Y(new_new_n323_));
  AN2        g0301(.A(i_3_), .B(i_10_), .Y(new_new_n324_));
  NA4        g0302(.A(new_new_n324_), .B(new_new_n204_), .C(new_new_n181_), .D(new_new_n179_), .Y(new_new_n325_));
  NO2        g0303(.A(i_5_), .B(new_new_n37_), .Y(new_new_n326_));
  NO2        g0304(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n327_));
  OR2        g0305(.A(new_new_n323_), .B(new_new_n318_), .Y(new_new_n328_));
  OAI220     g0306(.A0(new_new_n328_), .A1(i_6_), .B0(new_new_n316_), .B1(new_new_n300_), .Y(new_new_n329_));
  NO4        g0307(.A(new_new_n329_), .B(new_new_n298_), .C(new_new_n223_), .D(new_new_n172_), .Y(new_new_n330_));
  NO3        g0308(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n332_));
  NA2        g0310(.A(new_new_n307_), .B(new_new_n332_), .Y(new_new_n333_));
  NO3        g0311(.A(i_6_), .B(new_new_n199_), .C(i_7_), .Y(new_new_n334_));
  NA2        g0312(.A(new_new_n334_), .B(new_new_n204_), .Y(new_new_n335_));
  AOI210     g0313(.A0(new_new_n335_), .A1(new_new_n333_), .B0(new_new_n174_), .Y(new_new_n336_));
  NO2        g0314(.A(i_2_), .B(i_3_), .Y(new_new_n337_));
  OR2        g0315(.A(i_0_), .B(i_5_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n227_), .B(new_new_n338_), .Y(new_new_n339_));
  NA4        g0317(.A(new_new_n339_), .B(new_new_n244_), .C(new_new_n337_), .D(i_1_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n307_), .B(new_new_n302_), .C(new_new_n116_), .Y(new_new_n341_));
  NAi21      g0319(.An(i_8_), .B(i_7_), .Y(new_new_n342_));
  NO2        g0320(.A(new_new_n342_), .B(i_6_), .Y(new_new_n343_));
  NO2        g0321(.A(new_new_n161_), .B(new_new_n47_), .Y(new_new_n344_));
  NA3        g0322(.A(new_new_n344_), .B(new_new_n343_), .C(new_new_n167_), .Y(new_new_n345_));
  NA3        g0323(.A(new_new_n345_), .B(new_new_n341_), .C(new_new_n340_), .Y(new_new_n346_));
  OAI210     g0324(.A0(new_new_n346_), .A1(new_new_n336_), .B0(i_4_), .Y(new_new_n347_));
  NO2        g0325(.A(i_12_), .B(i_10_), .Y(new_new_n348_));
  NOi21      g0326(.An(i_5_), .B(i_0_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n320_), .B(new_new_n349_), .C(new_new_n131_), .Y(new_new_n350_));
  NA4        g0328(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n351_));
  NA2        g0329(.A(new_new_n350_), .B(new_new_n348_), .Y(new_new_n352_));
  NO2        g0330(.A(i_6_), .B(i_8_), .Y(new_new_n353_));
  NOi21      g0331(.An(i_0_), .B(i_2_), .Y(new_new_n354_));
  AN2        g0332(.A(new_new_n354_), .B(new_new_n353_), .Y(new_new_n355_));
  NO2        g0333(.A(i_1_), .B(i_7_), .Y(new_new_n356_));
  AO220      g0334(.A0(new_new_n356_), .A1(new_new_n355_), .B0(new_new_n343_), .B1(new_new_n245_), .Y(new_new_n357_));
  NA3        g0335(.A(new_new_n357_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n358_));
  NA3        g0336(.A(new_new_n358_), .B(new_new_n352_), .C(new_new_n347_), .Y(new_new_n359_));
  NO3        g0337(.A(new_new_n243_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n360_));
  NO3        g0338(.A(new_new_n342_), .B(i_2_), .C(i_1_), .Y(new_new_n361_));
  OAI210     g0339(.A0(new_new_n361_), .A1(new_new_n360_), .B0(i_6_), .Y(new_new_n362_));
  NA3        g0340(.A(new_new_n263_), .B(new_new_n319_), .C(new_new_n199_), .Y(new_new_n363_));
  AOI210     g0341(.A0(new_new_n363_), .A1(new_new_n362_), .B0(new_new_n339_), .Y(new_new_n364_));
  NOi21      g0342(.An(new_new_n157_), .B(new_new_n107_), .Y(new_new_n365_));
  NA2        g0343(.A(new_new_n364_), .B(i_3_), .Y(new_new_n366_));
  INV        g0344(.A(new_new_n84_), .Y(new_new_n367_));
  NO2        g0345(.A(new_new_n311_), .B(new_new_n81_), .Y(new_new_n368_));
  NA2        g0346(.A(new_new_n368_), .B(new_new_n135_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n95_), .B(new_new_n199_), .Y(new_new_n370_));
  NA3        g0348(.A(new_new_n322_), .B(new_new_n370_), .C(new_new_n63_), .Y(new_new_n371_));
  AOI210     g0349(.A0(new_new_n371_), .A1(new_new_n369_), .B0(new_new_n367_), .Y(new_new_n372_));
  NO2        g0350(.A(new_new_n199_), .B(i_9_), .Y(new_new_n373_));
  NA3        g0351(.A(new_new_n373_), .B(new_new_n212_), .C(new_new_n161_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n372_), .B(new_new_n310_), .Y(new_new_n375_));
  AOI210     g0353(.A0(new_new_n375_), .A1(new_new_n366_), .B0(new_new_n166_), .Y(new_new_n376_));
  AOI210     g0354(.A0(new_new_n359_), .A1(new_new_n331_), .B0(new_new_n376_), .Y(new_new_n377_));
  NOi32      g0355(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n378_));
  INV        g0356(.A(new_new_n378_), .Y(new_new_n379_));
  NAi21      g0357(.An(i_0_), .B(i_6_), .Y(new_new_n380_));
  NAi21      g0358(.An(i_1_), .B(i_5_), .Y(new_new_n381_));
  NA2        g0359(.A(new_new_n381_), .B(new_new_n380_), .Y(new_new_n382_));
  NA2        g0360(.A(new_new_n382_), .B(new_new_n25_), .Y(new_new_n383_));
  OAI210     g0361(.A0(new_new_n383_), .A1(new_new_n163_), .B0(new_new_n257_), .Y(new_new_n384_));
  NAi41      g0362(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n385_));
  OAI220     g0363(.A0(new_new_n385_), .A1(new_new_n381_), .B0(new_new_n230_), .B1(new_new_n163_), .Y(new_new_n386_));
  AOI210     g0364(.A0(new_new_n385_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n387_));
  NOi32      g0365(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n388_));
  OR2        g0366(.A(new_new_n387_), .B(new_new_n386_), .Y(new_new_n389_));
  NO2        g0367(.A(i_1_), .B(new_new_n104_), .Y(new_new_n390_));
  NAi21      g0368(.An(i_3_), .B(i_4_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(i_9_), .Y(new_new_n392_));
  AN2        g0370(.A(i_6_), .B(i_7_), .Y(new_new_n393_));
  OAI210     g0371(.A0(new_new_n393_), .A1(new_new_n390_), .B0(new_new_n392_), .Y(new_new_n394_));
  NA2        g0372(.A(i_2_), .B(i_7_), .Y(new_new_n395_));
  NO2        g0373(.A(new_new_n391_), .B(i_10_), .Y(new_new_n396_));
  NA3        g0374(.A(new_new_n396_), .B(new_new_n395_), .C(new_new_n255_), .Y(new_new_n397_));
  AOI210     g0375(.A0(new_new_n397_), .A1(new_new_n394_), .B0(new_new_n191_), .Y(new_new_n398_));
  AOI210     g0376(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n399_));
  OAI210     g0377(.A0(new_new_n399_), .A1(new_new_n194_), .B0(new_new_n396_), .Y(new_new_n400_));
  AOI220     g0378(.A0(new_new_n396_), .A1(new_new_n356_), .B0(new_new_n249_), .B1(new_new_n194_), .Y(new_new_n401_));
  AOI210     g0379(.A0(new_new_n401_), .A1(new_new_n400_), .B0(i_5_), .Y(new_new_n402_));
  NO4        g0380(.A(new_new_n402_), .B(new_new_n398_), .C(new_new_n389_), .D(new_new_n384_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n379_), .Y(new_new_n404_));
  NO2        g0382(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n405_));
  AN2        g0383(.A(i_12_), .B(i_5_), .Y(new_new_n406_));
  NO2        g0384(.A(i_4_), .B(new_new_n26_), .Y(new_new_n407_));
  NA2        g0385(.A(new_new_n407_), .B(new_new_n406_), .Y(new_new_n408_));
  NO2        g0386(.A(i_11_), .B(i_6_), .Y(new_new_n409_));
  NA3        g0387(.A(new_new_n409_), .B(new_new_n344_), .C(new_new_n235_), .Y(new_new_n410_));
  NO2        g0388(.A(new_new_n410_), .B(new_new_n408_), .Y(new_new_n411_));
  NO2        g0389(.A(new_new_n253_), .B(i_5_), .Y(new_new_n412_));
  NO2        g0390(.A(i_5_), .B(i_10_), .Y(new_new_n413_));
  AOI220     g0391(.A0(new_new_n413_), .A1(new_new_n284_), .B0(new_new_n412_), .B1(new_new_n204_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n147_), .B(new_new_n46_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n415_), .B(new_new_n414_), .Y(new_new_n416_));
  OAI210     g0394(.A0(new_new_n416_), .A1(new_new_n411_), .B0(new_new_n405_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n153_), .B(new_new_n86_), .Y(new_new_n419_));
  OAI210     g0397(.A0(new_new_n419_), .A1(new_new_n411_), .B0(new_new_n418_), .Y(new_new_n420_));
  NO3        g0398(.A(new_new_n86_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n421_));
  NO2        g0399(.A(i_11_), .B(i_12_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n413_), .B(new_new_n247_), .Y(new_new_n423_));
  NA3        g0401(.A(new_new_n116_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n424_));
  OAI220     g0402(.A0(new_new_n424_), .A1(new_new_n230_), .B0(new_new_n423_), .B1(new_new_n351_), .Y(new_new_n425_));
  NAi21      g0403(.An(i_13_), .B(i_0_), .Y(new_new_n426_));
  NO2        g0404(.A(new_new_n426_), .B(new_new_n250_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n425_), .B(new_new_n427_), .Y(new_new_n428_));
  NA3        g0406(.A(new_new_n428_), .B(new_new_n420_), .C(new_new_n417_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n45_), .B(new_new_n235_), .Y(new_new_n430_));
  NO3        g0408(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n431_));
  NO2        g0409(.A(i_0_), .B(i_11_), .Y(new_new_n432_));
  INV        g0410(.A(i_5_), .Y(new_new_n433_));
  AN2        g0411(.A(i_1_), .B(i_6_), .Y(new_new_n434_));
  NOi21      g0412(.An(i_2_), .B(i_12_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n435_), .B(new_new_n434_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(new_new_n433_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n145_), .B(i_9_), .Y(new_new_n438_));
  NO2        g0416(.A(new_new_n438_), .B(i_4_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n437_), .B(new_new_n439_), .Y(new_new_n440_));
  NAi21      g0418(.An(i_9_), .B(i_4_), .Y(new_new_n441_));
  OR2        g0419(.A(i_13_), .B(i_10_), .Y(new_new_n442_));
  NO3        g0420(.A(new_new_n442_), .B(new_new_n120_), .C(new_new_n441_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n177_), .B(new_new_n126_), .Y(new_new_n444_));
  OR2        g0422(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n299_), .B(new_new_n446_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n292_), .B(new_new_n219_), .Y(new_new_n448_));
  OAI220     g0426(.A0(new_new_n448_), .A1(new_new_n445_), .B0(new_new_n447_), .B1(new_new_n365_), .Y(new_new_n449_));
  INV        g0427(.A(new_new_n449_), .Y(new_new_n450_));
  AOI210     g0428(.A0(new_new_n450_), .A1(new_new_n440_), .B0(new_new_n26_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n452_));
  AOI220     g0430(.A0(new_new_n313_), .A1(new_new_n303_), .B0(new_new_n307_), .B1(new_new_n332_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n453_), .B(new_new_n174_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n188_), .B(new_new_n86_), .Y(new_new_n455_));
  AOI220     g0433(.A0(new_new_n455_), .A1(new_new_n312_), .B0(new_new_n294_), .B1(new_new_n219_), .Y(new_new_n456_));
  NO2        g0434(.A(new_new_n456_), .B(new_new_n301_), .Y(new_new_n457_));
  NO3        g0435(.A(new_new_n457_), .B(new_new_n454_), .C(new_new_n452_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n202_), .B(new_new_n99_), .Y(new_new_n459_));
  NA3        g0437(.A(new_new_n344_), .B(new_new_n167_), .C(new_new_n86_), .Y(new_new_n460_));
  AOI210     g0438(.A0(new_new_n460_), .A1(new_new_n459_), .B0(new_new_n342_), .Y(new_new_n461_));
  NA2        g0439(.A(new_new_n313_), .B(new_new_n245_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n462_), .B(new_new_n188_), .Y(new_new_n463_));
  NO2        g0441(.A(i_3_), .B(new_new_n49_), .Y(new_new_n464_));
  NA3        g0442(.A(new_new_n356_), .B(new_new_n355_), .C(new_new_n464_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n334_), .B(new_new_n339_), .Y(new_new_n466_));
  OAI210     g0444(.A0(new_new_n466_), .A1(new_new_n195_), .B0(new_new_n465_), .Y(new_new_n467_));
  NO3        g0445(.A(new_new_n467_), .B(new_new_n463_), .C(new_new_n461_), .Y(new_new_n468_));
  AOI210     g0446(.A0(new_new_n468_), .A1(new_new_n458_), .B0(new_new_n286_), .Y(new_new_n469_));
  NO4        g0447(.A(new_new_n469_), .B(new_new_n451_), .C(new_new_n429_), .D(new_new_n404_), .Y(new_new_n470_));
  NO2        g0448(.A(new_new_n63_), .B(i_4_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n73_), .B(i_13_), .Y(new_new_n472_));
  NA3        g0450(.A(new_new_n472_), .B(new_new_n471_), .C(i_2_), .Y(new_new_n473_));
  NO2        g0451(.A(i_10_), .B(i_9_), .Y(new_new_n474_));
  NAi21      g0452(.An(i_12_), .B(i_8_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n475_), .B(i_3_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n476_), .B(new_new_n474_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n47_), .B(i_4_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n478_), .B(new_new_n107_), .Y(new_new_n479_));
  OAI220     g0457(.A0(new_new_n479_), .A1(new_new_n211_), .B0(new_new_n477_), .B1(new_new_n473_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n327_), .B(i_0_), .Y(new_new_n481_));
  NO3        g0459(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n281_), .B(new_new_n100_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n483_), .B(new_new_n482_), .Y(new_new_n484_));
  NA2        g0462(.A(i_8_), .B(i_9_), .Y(new_new_n485_));
  AOI210     g0463(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n486_));
  OR2        g0464(.A(new_new_n486_), .B(new_new_n485_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n299_), .B(new_new_n212_), .Y(new_new_n488_));
  OAI220     g0466(.A0(new_new_n488_), .A1(new_new_n487_), .B0(new_new_n484_), .B1(new_new_n481_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n262_), .B(new_new_n326_), .Y(new_new_n490_));
  NO3        g0468(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n491_));
  INV        g0469(.A(new_new_n491_), .Y(new_new_n492_));
  NA3        g0470(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n493_));
  NA4        g0471(.A(new_new_n148_), .B(new_new_n119_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n494_));
  OAI220     g0472(.A0(new_new_n494_), .A1(new_new_n493_), .B0(new_new_n492_), .B1(new_new_n490_), .Y(new_new_n495_));
  NO3        g0473(.A(new_new_n495_), .B(new_new_n489_), .C(new_new_n480_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n312_), .B(new_new_n111_), .Y(new_new_n497_));
  OR2        g0475(.A(new_new_n497_), .B(new_new_n215_), .Y(new_new_n498_));
  OA210      g0476(.A0(new_new_n374_), .A1(new_new_n104_), .B0(new_new_n314_), .Y(new_new_n499_));
  OA220      g0477(.A0(new_new_n499_), .A1(new_new_n166_), .B0(new_new_n498_), .B1(new_new_n242_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n99_), .B(i_13_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n455_), .B(new_new_n405_), .Y(new_new_n502_));
  NO2        g0480(.A(i_2_), .B(i_13_), .Y(new_new_n503_));
  NA3        g0481(.A(new_new_n503_), .B(new_new_n165_), .C(new_new_n102_), .Y(new_new_n504_));
  OAI220     g0482(.A0(new_new_n504_), .A1(new_new_n247_), .B0(new_new_n502_), .B1(new_new_n501_), .Y(new_new_n505_));
  NO3        g0483(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n506_));
  NO2        g0484(.A(i_6_), .B(i_7_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n507_), .B(new_new_n506_), .Y(new_new_n508_));
  NO2        g0486(.A(i_11_), .B(i_1_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n73_), .B(i_3_), .Y(new_new_n510_));
  OR2        g0488(.A(i_11_), .B(i_8_), .Y(new_new_n511_));
  NOi21      g0489(.An(i_2_), .B(i_7_), .Y(new_new_n512_));
  NAi31      g0490(.An(new_new_n511_), .B(new_new_n512_), .C(new_new_n510_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n442_), .B(i_6_), .Y(new_new_n514_));
  NA3        g0492(.A(new_new_n514_), .B(new_new_n471_), .C(new_new_n75_), .Y(new_new_n515_));
  NO2        g0493(.A(new_new_n515_), .B(new_new_n513_), .Y(new_new_n516_));
  NO2        g0494(.A(i_3_), .B(new_new_n199_), .Y(new_new_n517_));
  NO2        g0495(.A(i_6_), .B(i_10_), .Y(new_new_n518_));
  NA4        g0496(.A(new_new_n518_), .B(new_new_n331_), .C(new_new_n517_), .D(new_new_n247_), .Y(new_new_n519_));
  NO2        g0497(.A(new_new_n519_), .B(new_new_n159_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n256_), .B(new_new_n176_), .C(new_new_n135_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n161_), .B(i_3_), .Y(new_new_n523_));
  NAi31      g0501(.An(new_new_n522_), .B(new_new_n523_), .C(new_new_n236_), .Y(new_new_n524_));
  NA3        g0502(.A(new_new_n418_), .B(new_new_n184_), .C(new_new_n152_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n525_), .B(new_new_n524_), .C(new_new_n521_), .Y(new_new_n526_));
  NO4        g0504(.A(new_new_n526_), .B(new_new_n520_), .C(new_new_n516_), .D(new_new_n505_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n482_), .B(new_new_n406_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n491_), .B(new_new_n413_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n529_), .B(new_new_n234_), .Y(new_new_n530_));
  NAi21      g0508(.An(new_new_n225_), .B(new_new_n422_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n356_), .B(new_new_n227_), .Y(new_new_n532_));
  NO2        g0510(.A(new_new_n26_), .B(i_5_), .Y(new_new_n533_));
  NO2        g0511(.A(i_0_), .B(new_new_n86_), .Y(new_new_n534_));
  NA3        g0512(.A(new_new_n534_), .B(new_new_n533_), .C(new_new_n145_), .Y(new_new_n535_));
  OR3        g0513(.A(new_new_n320_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n536_));
  OAI220     g0514(.A0(new_new_n536_), .A1(new_new_n535_), .B0(new_new_n532_), .B1(new_new_n531_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n27_), .B(i_10_), .Y(new_new_n538_));
  NO2        g0516(.A(new_new_n538_), .B(new_new_n501_), .Y(new_new_n539_));
  NA4        g0517(.A(new_new_n324_), .B(new_new_n233_), .C(new_new_n73_), .D(new_new_n247_), .Y(new_new_n540_));
  NO2        g0518(.A(new_new_n540_), .B(new_new_n508_), .Y(new_new_n541_));
  NO4        g0519(.A(new_new_n541_), .B(new_new_n539_), .C(new_new_n537_), .D(new_new_n530_), .Y(new_new_n542_));
  NA4        g0520(.A(new_new_n542_), .B(new_new_n527_), .C(new_new_n500_), .D(new_new_n496_), .Y(new_new_n543_));
  NA3        g0521(.A(new_new_n324_), .B(new_new_n181_), .C(new_new_n179_), .Y(new_new_n544_));
  OAI210     g0522(.A0(new_new_n318_), .A1(new_new_n186_), .B0(new_new_n544_), .Y(new_new_n545_));
  AN2        g0523(.A(new_new_n303_), .B(new_new_n244_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n546_), .B(new_new_n545_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n125_), .B(new_new_n115_), .Y(new_new_n548_));
  AO220      g0526(.A0(new_new_n548_), .A1(new_new_n482_), .B0(new_new_n443_), .B1(i_6_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n331_), .B(new_new_n168_), .Y(new_new_n550_));
  OAI210     g0528(.A0(new_new_n550_), .A1(new_new_n242_), .B0(new_new_n325_), .Y(new_new_n551_));
  AOI220     g0529(.A0(new_new_n551_), .A1(new_new_n343_), .B0(new_new_n549_), .B1(new_new_n327_), .Y(new_new_n552_));
  NA2        g0530(.A(new_new_n406_), .B(new_new_n235_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n378_), .B(new_new_n73_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n393_), .B(new_new_n388_), .Y(new_new_n555_));
  AO210      g0533(.A0(new_new_n554_), .A1(new_new_n553_), .B0(new_new_n555_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n36_), .B(i_8_), .Y(new_new_n557_));
  AOI210     g0535(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n443_), .Y(new_new_n558_));
  NA2        g0536(.A(new_new_n558_), .B(new_new_n556_), .Y(new_new_n559_));
  INV        g0537(.A(new_new_n559_), .Y(new_new_n560_));
  NA2        g0538(.A(new_new_n269_), .B(new_new_n64_), .Y(new_new_n561_));
  OAI210     g0539(.A0(i_8_), .A1(new_new_n561_), .B0(new_new_n137_), .Y(new_new_n562_));
  NO2        g0540(.A(i_7_), .B(new_new_n205_), .Y(new_new_n563_));
  OR2        g0541(.A(new_new_n188_), .B(i_4_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n564_), .B(new_new_n86_), .Y(new_new_n565_));
  AOI220     g0543(.A0(new_new_n565_), .A1(new_new_n563_), .B0(new_new_n562_), .B1(new_new_n444_), .Y(new_new_n566_));
  NA4        g0544(.A(new_new_n566_), .B(new_new_n560_), .C(new_new_n552_), .D(new_new_n547_), .Y(new_new_n567_));
  NA2        g0545(.A(new_new_n412_), .B(new_new_n312_), .Y(new_new_n568_));
  OAI210     g0546(.A0(new_new_n408_), .A1(new_new_n173_), .B0(new_new_n568_), .Y(new_new_n569_));
  NO2        g0547(.A(i_12_), .B(new_new_n199_), .Y(new_new_n570_));
  NA2        g0548(.A(new_new_n570_), .B(new_new_n235_), .Y(new_new_n571_));
  NO3        g0549(.A(new_new_n1116_), .B(new_new_n571_), .C(new_new_n497_), .Y(new_new_n572_));
  NOi31      g0550(.An(new_new_n334_), .B(new_new_n442_), .C(new_new_n38_), .Y(new_new_n573_));
  OAI210     g0551(.A0(new_new_n573_), .A1(new_new_n572_), .B0(new_new_n569_), .Y(new_new_n574_));
  NO2        g0552(.A(i_8_), .B(i_7_), .Y(new_new_n575_));
  OAI210     g0553(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n576_), .B(new_new_n233_), .Y(new_new_n577_));
  AOI220     g0555(.A0(new_new_n344_), .A1(new_new_n40_), .B0(new_new_n245_), .B1(new_new_n214_), .Y(new_new_n578_));
  OAI220     g0556(.A0(new_new_n578_), .A1(new_new_n564_), .B0(new_new_n577_), .B1(new_new_n253_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n45_), .B(i_10_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n580_), .B(i_6_), .Y(new_new_n581_));
  NA3        g0559(.A(new_new_n581_), .B(new_new_n579_), .C(new_new_n575_), .Y(new_new_n582_));
  AOI220     g0560(.A0(new_new_n455_), .A1(new_new_n344_), .B0(new_new_n258_), .B1(new_new_n255_), .Y(new_new_n583_));
  OAI220     g0561(.A0(new_new_n583_), .A1(new_new_n277_), .B0(new_new_n501_), .B1(new_new_n136_), .Y(new_new_n584_));
  NA2        g0562(.A(new_new_n584_), .B(new_new_n280_), .Y(new_new_n585_));
  NOi31      g0563(.An(new_new_n307_), .B(new_new_n318_), .C(new_new_n186_), .Y(new_new_n586_));
  NA3        g0564(.A(new_new_n324_), .B(new_new_n179_), .C(new_new_n99_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n231_), .B(new_new_n45_), .Y(new_new_n588_));
  NO2        g0566(.A(new_new_n161_), .B(i_5_), .Y(new_new_n589_));
  NA3        g0567(.A(new_new_n589_), .B(new_new_n430_), .C(new_new_n337_), .Y(new_new_n590_));
  OAI210     g0568(.A0(new_new_n590_), .A1(new_new_n588_), .B0(new_new_n587_), .Y(new_new_n591_));
  OAI210     g0569(.A0(new_new_n591_), .A1(new_new_n586_), .B0(new_new_n491_), .Y(new_new_n592_));
  NA4        g0570(.A(new_new_n592_), .B(new_new_n585_), .C(new_new_n582_), .D(new_new_n574_), .Y(new_new_n593_));
  NA3        g0571(.A(new_new_n227_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n594_));
  NA2        g0572(.A(new_new_n299_), .B(new_new_n84_), .Y(new_new_n595_));
  AOI210     g0573(.A0(new_new_n594_), .A1(new_new_n369_), .B0(new_new_n595_), .Y(new_new_n596_));
  NA2        g0574(.A(new_new_n313_), .B(new_new_n303_), .Y(new_new_n597_));
  NO2        g0575(.A(new_new_n597_), .B(new_new_n178_), .Y(new_new_n598_));
  NA2        g0576(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n599_));
  NA2        g0577(.A(new_new_n474_), .B(new_new_n231_), .Y(new_new_n600_));
  NO2        g0578(.A(new_new_n599_), .B(new_new_n600_), .Y(new_new_n601_));
  AOI210     g0579(.A0(i_6_), .A1(new_new_n47_), .B0(new_new_n390_), .Y(new_new_n602_));
  NA2        g0580(.A(i_0_), .B(new_new_n49_), .Y(new_new_n603_));
  NA3        g0581(.A(new_new_n570_), .B(new_new_n290_), .C(new_new_n603_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n602_), .B(new_new_n604_), .Y(new_new_n605_));
  NO4        g0583(.A(new_new_n605_), .B(new_new_n601_), .C(new_new_n598_), .D(new_new_n596_), .Y(new_new_n606_));
  NO4        g0584(.A(new_new_n263_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n607_));
  NO3        g0585(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n608_));
  NO2        g0586(.A(new_new_n243_), .B(new_new_n36_), .Y(new_new_n609_));
  AN2        g0587(.A(new_new_n609_), .B(new_new_n608_), .Y(new_new_n610_));
  OA210      g0588(.A0(new_new_n610_), .A1(new_new_n607_), .B0(new_new_n378_), .Y(new_new_n611_));
  NO2        g0589(.A(new_new_n442_), .B(i_1_), .Y(new_new_n612_));
  NOi31      g0590(.An(new_new_n612_), .B(new_new_n483_), .C(new_new_n73_), .Y(new_new_n613_));
  AN4        g0591(.A(new_new_n613_), .B(new_new_n439_), .C(new_new_n533_), .D(i_2_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n453_), .B(new_new_n182_), .Y(new_new_n615_));
  NO3        g0593(.A(new_new_n615_), .B(new_new_n614_), .C(new_new_n611_), .Y(new_new_n616_));
  NOi21      g0594(.An(i_10_), .B(i_6_), .Y(new_new_n617_));
  NO2        g0595(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n618_));
  AOI220     g0596(.A0(new_new_n299_), .A1(new_new_n618_), .B0(new_new_n290_), .B1(new_new_n617_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n619_), .B(new_new_n481_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n334_), .B(new_new_n168_), .Y(new_new_n622_));
  AOI220     g0600(.A0(new_new_n622_), .A1(new_new_n462_), .B0(new_new_n189_), .B1(new_new_n187_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n204_), .B(new_new_n37_), .Y(new_new_n624_));
  NOi31      g0602(.An(new_new_n149_), .B(new_new_n624_), .C(new_new_n351_), .Y(new_new_n625_));
  NO3        g0603(.A(new_new_n625_), .B(new_new_n623_), .C(new_new_n620_), .Y(new_new_n626_));
  NO2        g0604(.A(new_new_n554_), .B(new_new_n401_), .Y(new_new_n627_));
  INV        g0605(.A(new_new_n337_), .Y(new_new_n628_));
  NO2        g0606(.A(i_12_), .B(new_new_n86_), .Y(new_new_n629_));
  NA3        g0607(.A(new_new_n629_), .B(new_new_n290_), .C(new_new_n603_), .Y(new_new_n630_));
  NA3        g0608(.A(new_new_n409_), .B(new_new_n299_), .C(new_new_n227_), .Y(new_new_n631_));
  AOI210     g0609(.A0(new_new_n631_), .A1(new_new_n630_), .B0(new_new_n628_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n179_), .B(i_0_), .Y(new_new_n633_));
  NO3        g0611(.A(new_new_n633_), .B(new_new_n362_), .C(new_new_n318_), .Y(new_new_n634_));
  OR2        g0612(.A(i_2_), .B(i_5_), .Y(new_new_n635_));
  OR2        g0613(.A(new_new_n635_), .B(new_new_n434_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n636_), .B(new_new_n531_), .Y(new_new_n637_));
  NO4        g0615(.A(new_new_n637_), .B(new_new_n634_), .C(new_new_n632_), .D(new_new_n627_), .Y(new_new_n638_));
  NA4        g0616(.A(new_new_n638_), .B(new_new_n626_), .C(new_new_n616_), .D(new_new_n606_), .Y(new_new_n639_));
  NO4        g0617(.A(new_new_n639_), .B(new_new_n593_), .C(new_new_n567_), .D(new_new_n543_), .Y(new_new_n640_));
  NA4        g0618(.A(new_new_n640_), .B(new_new_n470_), .C(new_new_n377_), .D(new_new_n330_), .Y(zz07));
  NO2        g0619(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n642_));
  NO2        g0620(.A(new_new_n111_), .B(new_new_n92_), .Y(new_new_n643_));
  NA2        g0621(.A(new_new_n407_), .B(new_new_n643_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n518_), .B(new_new_n84_), .Y(new_new_n645_));
  NA2        g0623(.A(i_11_), .B(new_new_n199_), .Y(new_new_n646_));
  INV        g0624(.A(new_new_n644_), .Y(new_new_n647_));
  NA3        g0625(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n247_), .B(i_4_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n649_), .B(i_8_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n108_), .B(new_new_n648_), .Y(new_new_n651_));
  NA2        g0629(.A(i_2_), .B(new_new_n86_), .Y(new_new_n652_));
  OAI210     g0630(.A0(new_new_n89_), .A1(new_new_n209_), .B0(new_new_n210_), .Y(new_new_n653_));
  NO2        g0631(.A(i_7_), .B(new_new_n37_), .Y(new_new_n654_));
  NA2        g0632(.A(i_4_), .B(i_8_), .Y(new_new_n655_));
  AOI210     g0633(.A0(new_new_n655_), .A1(new_new_n324_), .B0(new_new_n654_), .Y(new_new_n656_));
  OAI220     g0634(.A0(new_new_n656_), .A1(new_new_n652_), .B0(new_new_n653_), .B1(i_13_), .Y(new_new_n657_));
  NO4        g0635(.A(new_new_n657_), .B(new_new_n651_), .C(new_new_n647_), .D(new_new_n642_), .Y(new_new_n658_));
  AOI210     g0636(.A0(new_new_n131_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n659_));
  AOI210     g0637(.A0(new_new_n659_), .A1(new_new_n247_), .B0(new_new_n165_), .Y(new_new_n660_));
  OR2        g0638(.A(i_6_), .B(i_10_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n23_), .Y(new_new_n662_));
  OR3        g0640(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n663_));
  NO3        g0641(.A(new_new_n663_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n664_));
  INV        g0642(.A(new_new_n206_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n664_), .B(new_new_n662_), .Y(new_new_n666_));
  OA220      g0644(.A0(new_new_n666_), .A1(new_new_n628_), .B0(new_new_n660_), .B1(new_new_n282_), .Y(new_new_n667_));
  AOI210     g0645(.A0(new_new_n667_), .A1(new_new_n658_), .B0(new_new_n63_), .Y(new_new_n668_));
  NOi21      g0646(.An(i_11_), .B(i_7_), .Y(new_new_n669_));
  AO210      g0647(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n670_), .B(new_new_n669_), .Y(new_new_n671_));
  NA2        g0649(.A(new_new_n671_), .B(new_new_n214_), .Y(new_new_n672_));
  NA3        g0650(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n673_));
  NAi31      g0651(.An(new_new_n673_), .B(new_new_n224_), .C(i_11_), .Y(new_new_n674_));
  AOI210     g0652(.A0(new_new_n674_), .A1(new_new_n672_), .B0(new_new_n63_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n676_));
  AO210      g0654(.A0(new_new_n676_), .A1(new_new_n401_), .B0(new_new_n41_), .Y(new_new_n677_));
  NO3        g0655(.A(new_new_n271_), .B(new_new_n216_), .C(new_new_n646_), .Y(new_new_n678_));
  OAI210     g0656(.A0(new_new_n678_), .A1(new_new_n236_), .B0(new_new_n63_), .Y(new_new_n679_));
  NA2        g0657(.A(new_new_n435_), .B(new_new_n31_), .Y(new_new_n680_));
  OR2        g0658(.A(new_new_n216_), .B(new_new_n111_), .Y(new_new_n681_));
  NA2        g0659(.A(new_new_n681_), .B(new_new_n680_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n63_), .B(i_9_), .Y(new_new_n683_));
  NO2        g0661(.A(new_new_n683_), .B(i_4_), .Y(new_new_n684_));
  NA2        g0662(.A(new_new_n684_), .B(new_new_n682_), .Y(new_new_n685_));
  NO2        g0663(.A(i_1_), .B(i_12_), .Y(new_new_n686_));
  NA3        g0664(.A(new_new_n686_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n687_));
  NA4        g0665(.A(new_new_n687_), .B(new_new_n685_), .C(new_new_n679_), .D(new_new_n677_), .Y(new_new_n688_));
  OAI210     g0666(.A0(new_new_n688_), .A1(new_new_n675_), .B0(i_6_), .Y(new_new_n689_));
  NO2        g0667(.A(new_new_n247_), .B(new_new_n86_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n690_), .B(i_11_), .Y(new_new_n691_));
  INV        g0669(.A(new_new_n484_), .Y(new_new_n692_));
  NO4        g0670(.A(new_new_n224_), .B(new_new_n131_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n693_), .B(new_new_n683_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n247_), .B(i_6_), .Y(new_new_n695_));
  NO3        g0673(.A(new_new_n661_), .B(new_new_n243_), .C(new_new_n23_), .Y(new_new_n696_));
  AOI210     g0674(.A0(i_1_), .A1(new_new_n272_), .B0(new_new_n696_), .Y(new_new_n697_));
  OAI210     g0675(.A0(new_new_n697_), .A1(new_new_n45_), .B0(new_new_n694_), .Y(new_new_n698_));
  NA3        g0676(.A(new_new_n575_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n699_));
  NA2        g0677(.A(new_new_n141_), .B(i_9_), .Y(new_new_n700_));
  NA3        g0678(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n47_), .B(i_1_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n700_), .B(new_new_n1114_), .Y(new_new_n703_));
  NA3        g0681(.A(new_new_n683_), .B(new_new_n337_), .C(i_6_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n704_), .B(new_new_n23_), .Y(new_new_n705_));
  AOI210     g0683(.A0(new_new_n509_), .A1(new_new_n446_), .B0(new_new_n252_), .Y(new_new_n706_));
  NO2        g0684(.A(new_new_n706_), .B(new_new_n652_), .Y(new_new_n707_));
  NO2        g0685(.A(i_11_), .B(new_new_n37_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n708_), .B(new_new_n24_), .Y(new_new_n709_));
  OR3        g0687(.A(new_new_n707_), .B(new_new_n705_), .C(new_new_n703_), .Y(new_new_n710_));
  NO3        g0688(.A(new_new_n710_), .B(new_new_n698_), .C(new_new_n692_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n247_), .B(new_new_n104_), .Y(new_new_n712_));
  NO2        g0690(.A(new_new_n712_), .B(new_new_n669_), .Y(new_new_n713_));
  NA2        g0691(.A(new_new_n713_), .B(i_1_), .Y(new_new_n714_));
  NO2        g0692(.A(new_new_n714_), .B(new_new_n663_), .Y(new_new_n715_));
  NO2        g0693(.A(new_new_n441_), .B(new_new_n86_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n715_), .B(new_new_n47_), .Y(new_new_n717_));
  NO2        g0695(.A(new_new_n243_), .B(new_new_n45_), .Y(new_new_n718_));
  NO3        g0696(.A(new_new_n718_), .B(new_new_n327_), .C(new_new_n248_), .Y(new_new_n719_));
  NO2        g0697(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n720_));
  NO2        g0698(.A(new_new_n720_), .B(i_6_), .Y(new_new_n721_));
  NO2        g0699(.A(new_new_n86_), .B(i_9_), .Y(new_new_n722_));
  NO2        g0700(.A(new_new_n722_), .B(new_new_n63_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n723_), .B(new_new_n686_), .Y(new_new_n724_));
  NO4        g0702(.A(new_new_n724_), .B(new_new_n721_), .C(new_new_n719_), .D(i_4_), .Y(new_new_n725_));
  NA2        g0703(.A(i_1_), .B(i_3_), .Y(new_new_n726_));
  INV        g0704(.A(new_new_n725_), .Y(new_new_n727_));
  NA4        g0705(.A(new_new_n727_), .B(new_new_n717_), .C(new_new_n711_), .D(new_new_n689_), .Y(new_new_n728_));
  NO3        g0706(.A(new_new_n511_), .B(i_3_), .C(i_7_), .Y(new_new_n729_));
  NOi21      g0707(.An(new_new_n729_), .B(i_10_), .Y(new_new_n730_));
  OA210      g0708(.A0(new_new_n730_), .A1(new_new_n256_), .B0(new_new_n86_), .Y(new_new_n731_));
  NO3        g0709(.A(new_new_n512_), .B(new_new_n655_), .C(new_new_n86_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n732_), .B(new_new_n25_), .Y(new_new_n733_));
  NA3        g0711(.A(new_new_n165_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n734_), .B(new_new_n733_), .Y(new_new_n735_));
  OAI210     g0713(.A0(new_new_n735_), .A1(new_new_n731_), .B0(i_1_), .Y(new_new_n736_));
  AOI210     g0714(.A0(new_new_n281_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n737_));
  NO2        g0715(.A(new_new_n391_), .B(i_2_), .Y(new_new_n738_));
  NA2        g0716(.A(new_new_n738_), .B(new_new_n737_), .Y(new_new_n739_));
  OAI210     g0717(.A0(new_new_n704_), .A1(new_new_n475_), .B0(new_new_n739_), .Y(new_new_n740_));
  INV        g0718(.A(new_new_n740_), .Y(new_new_n741_));
  AOI210     g0719(.A0(new_new_n741_), .A1(new_new_n736_), .B0(i_13_), .Y(new_new_n742_));
  OR2        g0720(.A(i_11_), .B(i_7_), .Y(new_new_n743_));
  NA3        g0721(.A(new_new_n743_), .B(new_new_n109_), .C(new_new_n141_), .Y(new_new_n744_));
  AOI220     g0722(.A0(new_new_n503_), .A1(new_new_n165_), .B0(new_new_n478_), .B1(new_new_n141_), .Y(new_new_n745_));
  OAI210     g0723(.A0(new_new_n745_), .A1(new_new_n45_), .B0(new_new_n744_), .Y(new_new_n746_));
  AOI210     g0724(.A0(new_new_n701_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n747_));
  INV        g0725(.A(new_new_n747_), .Y(new_new_n748_));
  NO2        g0726(.A(new_new_n512_), .B(new_new_n24_), .Y(new_new_n749_));
  AOI220     g0727(.A0(new_new_n749_), .A1(new_new_n716_), .B0(new_new_n256_), .B1(new_new_n134_), .Y(new_new_n750_));
  OAI220     g0728(.A0(new_new_n750_), .A1(new_new_n41_), .B0(new_new_n748_), .B1(new_new_n95_), .Y(new_new_n751_));
  AOI210     g0729(.A0(new_new_n746_), .A1(new_new_n353_), .B0(new_new_n751_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n409_), .B(new_new_n702_), .Y(new_new_n753_));
  NO2        g0731(.A(new_new_n753_), .B(new_new_n253_), .Y(new_new_n754_));
  AOI210     g0732(.A0(new_new_n475_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n755_));
  NOi31      g0733(.An(new_new_n755_), .B(new_new_n645_), .C(new_new_n45_), .Y(new_new_n756_));
  NA2        g0734(.A(new_new_n130_), .B(i_13_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n701_), .B(new_new_n118_), .Y(new_new_n758_));
  INV        g0736(.A(new_new_n758_), .Y(new_new_n759_));
  OAI220     g0737(.A0(new_new_n759_), .A1(new_new_n71_), .B0(new_new_n757_), .B1(new_new_n737_), .Y(new_new_n760_));
  NO3        g0738(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n761_));
  NA2        g0739(.A(new_new_n26_), .B(new_new_n199_), .Y(new_new_n762_));
  AOI220     g0740(.A0(new_new_n409_), .A1(new_new_n702_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n763_));
  OAI220     g0741(.A0(new_new_n763_), .A1(new_new_n650_), .B0(new_new_n1115_), .B1(new_new_n665_), .Y(new_new_n764_));
  NO4        g0742(.A(new_new_n764_), .B(new_new_n760_), .C(new_new_n756_), .D(new_new_n754_), .Y(new_new_n765_));
  OR2        g0743(.A(i_11_), .B(i_6_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n649_), .B(new_new_n762_), .C(i_7_), .Y(new_new_n767_));
  AOI210     g0745(.A0(new_new_n767_), .A1(new_new_n759_), .B0(new_new_n766_), .Y(new_new_n768_));
  NA3        g0746(.A(new_new_n435_), .B(new_new_n654_), .C(new_new_n100_), .Y(new_new_n769_));
  NA2        g0747(.A(new_new_n691_), .B(i_13_), .Y(new_new_n770_));
  NA2        g0748(.A(new_new_n105_), .B(new_new_n762_), .Y(new_new_n771_));
  NAi21      g0749(.An(i_11_), .B(i_12_), .Y(new_new_n772_));
  NOi41      g0750(.An(new_new_n114_), .B(new_new_n772_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n773_), .B(new_new_n771_), .Y(new_new_n774_));
  NA3        g0752(.A(new_new_n774_), .B(new_new_n770_), .C(new_new_n769_), .Y(new_new_n775_));
  OAI210     g0753(.A0(new_new_n775_), .A1(new_new_n768_), .B0(new_new_n63_), .Y(new_new_n776_));
  NO2        g0754(.A(i_2_), .B(i_12_), .Y(new_new_n777_));
  NA2        g0755(.A(new_new_n390_), .B(new_new_n777_), .Y(new_new_n778_));
  NA2        g0756(.A(i_8_), .B(new_new_n25_), .Y(new_new_n779_));
  NO3        g0757(.A(new_new_n779_), .B(new_new_n407_), .C(new_new_n649_), .Y(new_new_n780_));
  OAI210     g0758(.A0(new_new_n780_), .A1(new_new_n392_), .B0(new_new_n390_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n131_), .B(i_2_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n782_), .B(new_new_n686_), .Y(new_new_n783_));
  NA3        g0761(.A(new_new_n783_), .B(new_new_n781_), .C(new_new_n778_), .Y(new_new_n784_));
  NA3        g0762(.A(new_new_n784_), .B(new_new_n46_), .C(new_new_n235_), .Y(new_new_n785_));
  NA4        g0763(.A(new_new_n785_), .B(new_new_n776_), .C(new_new_n765_), .D(new_new_n752_), .Y(new_new_n786_));
  OR4        g0764(.A(new_new_n786_), .B(new_new_n742_), .C(new_new_n728_), .D(new_new_n668_), .Y(zz05));
  AOI210     g0765(.A0(new_new_n713_), .A1(new_new_n284_), .B0(new_new_n444_), .Y(new_new_n788_));
  AN2        g0766(.A(new_new_n24_), .B(i_10_), .Y(new_new_n789_));
  NA3        g0767(.A(new_new_n789_), .B(new_new_n777_), .C(new_new_n111_), .Y(new_new_n790_));
  NO2        g0768(.A(new_new_n650_), .B(i_11_), .Y(new_new_n791_));
  OAI210     g0769(.A0(new_new_n654_), .A1(new_new_n89_), .B0(new_new_n791_), .Y(new_new_n792_));
  NA3        g0770(.A(new_new_n792_), .B(new_new_n790_), .C(new_new_n788_), .Y(new_new_n793_));
  NO3        g0771(.A(i_11_), .B(new_new_n247_), .C(i_13_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n795_));
  NA2        g0773(.A(i_12_), .B(i_8_), .Y(new_new_n796_));
  OAI210     g0774(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n796_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n474_), .Y(new_new_n798_));
  AOI220     g0776(.A0(new_new_n337_), .A1(new_new_n621_), .B0(new_new_n797_), .B1(new_new_n795_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n799_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n800_), .B(new_new_n793_), .Y(new_new_n801_));
  INV        g0779(.A(new_new_n176_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n256_), .Y(new_new_n803_));
  OAI210     g0781(.A0(new_new_n738_), .A1(new_new_n476_), .B0(new_new_n114_), .Y(new_new_n804_));
  AOI210     g0782(.A0(new_new_n804_), .A1(new_new_n803_), .B0(new_new_n802_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n485_), .B(new_new_n26_), .Y(new_new_n806_));
  NO2        g0784(.A(new_new_n806_), .B(new_new_n446_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n807_), .B(i_2_), .Y(new_new_n808_));
  INV        g0786(.A(new_new_n808_), .Y(new_new_n809_));
  AOI210     g0787(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n442_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n810_), .A1(new_new_n809_), .B0(new_new_n805_), .Y(new_new_n811_));
  NO2        g0789(.A(new_new_n196_), .B(new_new_n128_), .Y(new_new_n812_));
  OAI210     g0790(.A0(new_new_n812_), .A1(new_new_n795_), .B0(i_2_), .Y(new_new_n813_));
  INV        g0791(.A(new_new_n177_), .Y(new_new_n814_));
  NO3        g0792(.A(new_new_n670_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n815_));
  AOI210     g0793(.A0(new_new_n814_), .A1(new_new_n89_), .B0(new_new_n815_), .Y(new_new_n816_));
  AOI210     g0794(.A0(new_new_n816_), .A1(new_new_n813_), .B0(new_new_n199_), .Y(new_new_n817_));
  OA210      g0795(.A0(new_new_n671_), .A1(new_new_n129_), .B0(i_13_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n206_), .B(new_new_n209_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n155_), .B(new_new_n646_), .Y(new_new_n820_));
  AOI210     g0798(.A0(new_new_n820_), .A1(new_new_n819_), .B0(new_new_n395_), .Y(new_new_n821_));
  AOI210     g0799(.A0(new_new_n216_), .A1(new_new_n151_), .B0(new_new_n557_), .Y(new_new_n822_));
  OAI210     g0800(.A0(new_new_n822_), .A1(new_new_n236_), .B0(new_new_n446_), .Y(new_new_n823_));
  NO2        g0801(.A(new_new_n105_), .B(new_new_n45_), .Y(new_new_n824_));
  INV        g0802(.A(new_new_n319_), .Y(new_new_n825_));
  NA4        g0803(.A(new_new_n825_), .B(new_new_n324_), .C(new_new_n127_), .D(new_new_n43_), .Y(new_new_n826_));
  OAI210     g0804(.A0(new_new_n826_), .A1(new_new_n824_), .B0(new_new_n823_), .Y(new_new_n827_));
  NO4        g0805(.A(new_new_n827_), .B(new_new_n821_), .C(new_new_n818_), .D(new_new_n817_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n621_), .B(new_new_n28_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n794_), .B(new_new_n291_), .Y(new_new_n830_));
  NA2        g0808(.A(new_new_n830_), .B(new_new_n829_), .Y(new_new_n831_));
  NO2        g0809(.A(new_new_n62_), .B(i_12_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n832_), .B(new_new_n129_), .Y(new_new_n833_));
  NO2        g0811(.A(new_new_n833_), .B(new_new_n646_), .Y(new_new_n834_));
  AOI220     g0812(.A0(new_new_n834_), .A1(new_new_n36_), .B0(new_new_n831_), .B1(new_new_n47_), .Y(new_new_n835_));
  NA4        g0813(.A(new_new_n835_), .B(new_new_n828_), .C(new_new_n811_), .D(new_new_n801_), .Y(zz06));
  NO3        g0814(.A(new_new_n267_), .B(new_new_n326_), .C(i_1_), .Y(new_new_n837_));
  NO2        g0815(.A(new_new_n191_), .B(new_new_n142_), .Y(new_new_n838_));
  OAI210     g0816(.A0(new_new_n838_), .A1(new_new_n837_), .B0(new_new_n782_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n230_), .B(new_new_n522_), .Y(new_new_n840_));
  INV        g0818(.A(new_new_n349_), .Y(new_new_n841_));
  AO210      g0819(.A0(new_new_n841_), .A1(new_new_n839_), .B0(i_12_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n629_), .B(new_new_n63_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n730_), .B(new_new_n71_), .Y(new_new_n844_));
  BUFFER     g0822(.A(new_new_n676_), .Y(new_new_n845_));
  NA3        g0823(.A(new_new_n845_), .B(new_new_n844_), .C(new_new_n843_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n846_), .B(new_new_n73_), .Y(new_new_n847_));
  INV        g0825(.A(new_new_n348_), .Y(new_new_n848_));
  NA2        g0826(.A(new_new_n75_), .B(new_new_n134_), .Y(new_new_n849_));
  INV        g0827(.A(new_new_n127_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n850_), .B(new_new_n47_), .Y(new_new_n851_));
  AOI210     g0829(.A0(new_new_n851_), .A1(new_new_n849_), .B0(new_new_n848_), .Y(new_new_n852_));
  NO3        g0830(.A(new_new_n263_), .B(new_new_n135_), .C(i_9_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n853_), .B(new_new_n832_), .Y(new_new_n854_));
  AOI210     g0832(.A0(new_new_n854_), .A1(new_new_n555_), .B0(new_new_n191_), .Y(new_new_n855_));
  NO2        g0833(.A(new_new_n32_), .B(i_11_), .Y(new_new_n856_));
  NA3        g0834(.A(new_new_n856_), .B(new_new_n507_), .C(new_new_n413_), .Y(new_new_n857_));
  NAi32      g0835(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n858_));
  AOI210     g0836(.A0(new_new_n766_), .A1(new_new_n87_), .B0(new_new_n858_), .Y(new_new_n859_));
  OAI210     g0837(.A0(new_new_n729_), .A1(new_new_n609_), .B0(new_new_n608_), .Y(new_new_n860_));
  NAi31      g0838(.An(new_new_n859_), .B(new_new_n860_), .C(new_new_n857_), .Y(new_new_n861_));
  OR3        g0839(.A(new_new_n861_), .B(new_new_n855_), .C(new_new_n852_), .Y(new_new_n862_));
  NO2        g0840(.A(new_new_n743_), .B(i_2_), .Y(new_new_n863_));
  NA2        g0841(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n864_));
  OAI210     g0842(.A0(new_new_n864_), .A1(new_new_n434_), .B0(new_new_n383_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n865_), .B(new_new_n863_), .Y(new_new_n866_));
  AO220      g0844(.A0(new_new_n382_), .A1(new_new_n373_), .B0(new_new_n421_), .B1(new_new_n646_), .Y(new_new_n867_));
  NA3        g0845(.A(new_new_n867_), .B(new_new_n268_), .C(i_7_), .Y(new_new_n868_));
  OR2        g0846(.A(new_new_n671_), .B(new_new_n476_), .Y(new_new_n869_));
  NA3        g0847(.A(new_new_n869_), .B(new_new_n150_), .C(new_new_n69_), .Y(new_new_n870_));
  AO210      g0848(.A0(new_new_n529_), .A1(new_new_n798_), .B0(new_new_n36_), .Y(new_new_n871_));
  NA4        g0849(.A(new_new_n871_), .B(new_new_n870_), .C(new_new_n868_), .D(new_new_n866_), .Y(new_new_n872_));
  OAI210     g0850(.A0(new_new_n690_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n873_));
  AOI220     g0851(.A0(new_new_n873_), .A1(new_new_n608_), .B0(new_new_n840_), .B1(new_new_n1117_), .Y(new_new_n874_));
  NA3        g0852(.A(new_new_n395_), .B(new_new_n249_), .C(new_new_n150_), .Y(new_new_n875_));
  OAI210     g0853(.A0(new_new_n421_), .A1(new_new_n210_), .B0(new_new_n70_), .Y(new_new_n876_));
  NA4        g0854(.A(new_new_n876_), .B(new_new_n875_), .C(new_new_n874_), .D(new_new_n653_), .Y(new_new_n877_));
  NA3        g0855(.A(new_new_n88_), .B(new_new_n518_), .C(new_new_n227_), .Y(new_new_n878_));
  AOI210     g0856(.A0(new_new_n476_), .A1(new_new_n474_), .B0(new_new_n607_), .Y(new_new_n879_));
  NO2        g0857(.A(new_new_n661_), .B(new_new_n105_), .Y(new_new_n880_));
  OAI210     g0858(.A0(new_new_n880_), .A1(new_new_n115_), .B0(new_new_n432_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n255_), .B(new_new_n47_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n882_), .B(new_new_n636_), .Y(new_new_n883_));
  NA3        g0861(.A(new_new_n883_), .B(new_new_n348_), .C(i_7_), .Y(new_new_n884_));
  NA4        g0862(.A(new_new_n884_), .B(new_new_n881_), .C(new_new_n879_), .D(new_new_n878_), .Y(new_new_n885_));
  NO4        g0863(.A(new_new_n885_), .B(new_new_n877_), .C(new_new_n872_), .D(new_new_n862_), .Y(new_new_n886_));
  NA4        g0864(.A(new_new_n886_), .B(new_new_n847_), .C(new_new_n842_), .D(new_new_n403_), .Y(zz03));
  NA2        g0865(.A(i_6_), .B(i_7_), .Y(new_new_n888_));
  NO2        g0866(.A(new_new_n888_), .B(i_0_), .Y(new_new_n889_));
  NO2        g0867(.A(i_11_), .B(new_new_n247_), .Y(new_new_n890_));
  OAI210     g0868(.A0(new_new_n889_), .A1(new_new_n307_), .B0(new_new_n890_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n891_), .B(new_new_n199_), .Y(new_new_n892_));
  NO3        g0870(.A(new_new_n481_), .B(new_new_n92_), .C(new_new_n45_), .Y(new_new_n893_));
  OA210      g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n179_), .Y(new_new_n894_));
  NA3        g0872(.A(new_new_n875_), .B(new_new_n653_), .C(new_new_n394_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n895_), .B(new_new_n40_), .Y(new_new_n896_));
  NOi21      g0874(.An(new_new_n99_), .B(new_new_n807_), .Y(new_new_n897_));
  NO3        g0875(.A(new_new_n681_), .B(new_new_n485_), .C(new_new_n134_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n435_), .B(new_new_n46_), .Y(new_new_n899_));
  NO2        g0877(.A(new_new_n898_), .B(new_new_n897_), .Y(new_new_n900_));
  AOI210     g0878(.A0(new_new_n900_), .A1(new_new_n896_), .B0(new_new_n49_), .Y(new_new_n901_));
  NO4        g0879(.A(new_new_n399_), .B(new_new_n406_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n191_), .B(new_new_n617_), .Y(new_new_n903_));
  NOi31      g0881(.An(new_new_n903_), .B(new_new_n902_), .C(new_new_n39_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n755_), .B(new_new_n722_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n354_), .B(new_new_n464_), .Y(new_new_n906_));
  OAI220     g0884(.A0(new_new_n906_), .A1(new_new_n905_), .B0(new_new_n904_), .B1(new_new_n63_), .Y(new_new_n907_));
  NOi21      g0885(.An(i_5_), .B(i_9_), .Y(new_new_n908_));
  NA2        g0886(.A(new_new_n908_), .B(new_new_n472_), .Y(new_new_n909_));
  AOI210     g0887(.A0(new_new_n281_), .A1(new_new_n509_), .B0(new_new_n732_), .Y(new_new_n910_));
  NO3        g0888(.A(new_new_n438_), .B(new_new_n281_), .C(new_new_n73_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n180_), .B(new_new_n151_), .Y(new_new_n912_));
  AOI210     g0890(.A0(new_new_n912_), .A1(new_new_n255_), .B0(new_new_n911_), .Y(new_new_n913_));
  OAI220     g0891(.A0(new_new_n913_), .A1(new_new_n186_), .B0(new_new_n910_), .B1(new_new_n909_), .Y(new_new_n914_));
  NO4        g0892(.A(new_new_n914_), .B(new_new_n907_), .C(new_new_n901_), .D(new_new_n894_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n191_), .B(new_new_n24_), .Y(new_new_n916_));
  NO2        g0894(.A(new_new_n720_), .B(new_new_n643_), .Y(new_new_n917_));
  NO2        g0895(.A(new_new_n917_), .B(new_new_n916_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n331_), .B(new_new_n132_), .Y(new_new_n919_));
  NAi21      g0897(.An(new_new_n166_), .B(new_new_n464_), .Y(new_new_n920_));
  OAI220     g0898(.A0(new_new_n920_), .A1(new_new_n882_), .B0(new_new_n919_), .B1(new_new_n423_), .Y(new_new_n921_));
  NO2        g0899(.A(new_new_n921_), .B(new_new_n918_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n413_), .B(new_new_n311_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n923_), .B(new_new_n758_), .Y(new_new_n924_));
  NA2        g0902(.A(new_new_n618_), .B(i_0_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n925_), .B(new_new_n408_), .C(new_new_n89_), .Y(new_new_n926_));
  NO4        g0904(.A(new_new_n635_), .B(new_new_n224_), .C(new_new_n442_), .D(new_new_n434_), .Y(new_new_n927_));
  AOI210     g0905(.A0(new_new_n927_), .A1(i_11_), .B0(new_new_n926_), .Y(new_new_n928_));
  INV        g0906(.A(new_new_n507_), .Y(new_new_n929_));
  AN2        g0907(.A(new_new_n99_), .B(new_new_n254_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n794_), .B(new_new_n349_), .Y(new_new_n931_));
  AOI210     g0909(.A0(new_new_n518_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n932_));
  OAI220     g0910(.A0(new_new_n932_), .A1(new_new_n931_), .B0(new_new_n709_), .B1(new_new_n577_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n265_), .B(new_new_n157_), .Y(new_new_n934_));
  NA2        g0912(.A(i_0_), .B(i_10_), .Y(new_new_n935_));
  AN2        g0913(.A(new_new_n934_), .B(i_6_), .Y(new_new_n936_));
  AOI220     g0914(.A0(new_new_n354_), .A1(new_new_n101_), .B0(new_new_n191_), .B1(new_new_n84_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n612_), .B(i_4_), .Y(new_new_n938_));
  NA2        g0916(.A(new_new_n194_), .B(new_new_n209_), .Y(new_new_n939_));
  OAI220     g0917(.A0(new_new_n939_), .A1(new_new_n931_), .B0(new_new_n938_), .B1(new_new_n937_), .Y(new_new_n940_));
  NO4        g0918(.A(new_new_n940_), .B(new_new_n936_), .C(new_new_n933_), .D(new_new_n930_), .Y(new_new_n941_));
  NA4        g0919(.A(new_new_n941_), .B(new_new_n928_), .C(new_new_n924_), .D(new_new_n922_), .Y(new_new_n942_));
  NA2        g0920(.A(i_11_), .B(i_9_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n49_), .B(i_7_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n418_), .B(new_new_n184_), .Y(new_new_n945_));
  NA3        g0923(.A(new_new_n945_), .B(new_new_n490_), .C(new_new_n164_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n943_), .B(new_new_n73_), .Y(new_new_n947_));
  NO2        g0925(.A(new_new_n180_), .B(i_0_), .Y(new_new_n948_));
  INV        g0926(.A(new_new_n948_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n507_), .B(new_new_n241_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n393_), .A1(new_new_n42_), .B0(new_new_n431_), .Y(new_new_n951_));
  OAI220     g0929(.A0(new_new_n951_), .A1(new_new_n909_), .B0(new_new_n950_), .B1(new_new_n949_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n952_), .B(new_new_n946_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n708_), .B(new_new_n124_), .Y(new_new_n954_));
  NO2        g0932(.A(i_6_), .B(new_new_n954_), .Y(new_new_n955_));
  AOI210     g0933(.A0(new_new_n475_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n176_), .B(new_new_n106_), .Y(new_new_n957_));
  NOi32      g0935(.An(new_new_n956_), .Bn(new_new_n194_), .C(new_new_n957_), .Y(new_new_n958_));
  AOI210     g0936(.A0(new_new_n654_), .A1(new_new_n349_), .B0(new_new_n254_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n959_), .B(new_new_n899_), .Y(new_new_n960_));
  NO3        g0938(.A(new_new_n960_), .B(new_new_n958_), .C(new_new_n955_), .Y(new_new_n961_));
  NOi21      g0939(.An(i_7_), .B(i_5_), .Y(new_new_n962_));
  NOi31      g0940(.An(new_new_n962_), .B(i_0_), .C(new_new_n772_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n963_), .B(new_new_n407_), .C(i_6_), .Y(new_new_n964_));
  OA210      g0942(.A0(new_new_n957_), .A1(new_new_n555_), .B0(new_new_n964_), .Y(new_new_n965_));
  NO3        g0943(.A(new_new_n426_), .B(new_new_n385_), .C(new_new_n381_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n275_), .B(new_new_n338_), .Y(new_new_n967_));
  NO2        g0945(.A(new_new_n772_), .B(new_new_n270_), .Y(new_new_n968_));
  AOI210     g0946(.A0(new_new_n968_), .A1(new_new_n967_), .B0(new_new_n966_), .Y(new_new_n969_));
  NA4        g0947(.A(new_new_n969_), .B(new_new_n965_), .C(new_new_n961_), .D(new_new_n953_), .Y(new_new_n970_));
  NO2        g0948(.A(new_new_n916_), .B(new_new_n250_), .Y(new_new_n971_));
  AN2        g0949(.A(new_new_n353_), .B(new_new_n349_), .Y(new_new_n972_));
  AO220      g0950(.A0(new_new_n972_), .A1(new_new_n912_), .B0(new_new_n368_), .B1(new_new_n27_), .Y(new_new_n973_));
  OAI210     g0951(.A0(new_new_n973_), .A1(new_new_n971_), .B0(i_10_), .Y(new_new_n974_));
  OA210      g0952(.A0(new_new_n507_), .A1(new_new_n233_), .B0(new_new_n506_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n506_), .B(new_new_n435_), .C(new_new_n46_), .Y(new_new_n976_));
  OAI210     g0954(.A0(new_new_n920_), .A1(new_new_n929_), .B0(new_new_n976_), .Y(new_new_n977_));
  NO2        g0955(.A(new_new_n268_), .B(new_new_n47_), .Y(new_new_n978_));
  NA2        g0956(.A(new_new_n947_), .B(new_new_n324_), .Y(new_new_n979_));
  OAI210     g0957(.A0(new_new_n978_), .A1(new_new_n193_), .B0(new_new_n979_), .Y(new_new_n980_));
  AOI220     g0958(.A0(new_new_n980_), .A1(new_new_n507_), .B0(new_new_n977_), .B1(new_new_n73_), .Y(new_new_n981_));
  NA3        g0959(.A(new_new_n864_), .B(new_new_n405_), .C(new_new_n690_), .Y(new_new_n982_));
  NA2        g0960(.A(new_new_n95_), .B(new_new_n45_), .Y(new_new_n983_));
  NO2        g0961(.A(new_new_n75_), .B(new_new_n796_), .Y(new_new_n984_));
  AOI220     g0962(.A0(new_new_n984_), .A1(new_new_n983_), .B0(new_new_n179_), .B1(new_new_n643_), .Y(new_new_n985_));
  AOI210     g0963(.A0(new_new_n985_), .A1(new_new_n982_), .B0(new_new_n48_), .Y(new_new_n986_));
  NO3        g0964(.A(new_new_n635_), .B(new_new_n380_), .C(new_new_n24_), .Y(new_new_n987_));
  AOI210     g0965(.A0(new_new_n749_), .A1(new_new_n589_), .B0(new_new_n987_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n648_), .B(new_new_n108_), .Y(new_new_n989_));
  NA2        g0967(.A(new_new_n989_), .B(i_0_), .Y(new_new_n990_));
  OAI220     g0968(.A0(new_new_n990_), .A1(new_new_n86_), .B0(new_new_n988_), .B1(new_new_n177_), .Y(new_new_n991_));
  NO3        g0969(.A(new_new_n991_), .B(new_new_n986_), .C(new_new_n559_), .Y(new_new_n992_));
  NA3        g0970(.A(new_new_n992_), .B(new_new_n981_), .C(new_new_n974_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n993_), .B(new_new_n970_), .C(new_new_n942_), .Y(new_new_n994_));
  NO2        g0972(.A(i_0_), .B(new_new_n772_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n935_), .B(new_new_n996_), .Y(new_new_n997_));
  NO3        g0975(.A(new_new_n108_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n998_));
  AO220      g0976(.A0(new_new_n998_), .A1(new_new_n997_), .B0(new_new_n995_), .B1(new_new_n179_), .Y(new_new_n999_));
  NO2        g0977(.A(new_new_n843_), .B(new_new_n957_), .Y(new_new_n1000_));
  AOI210     g0978(.A0(new_new_n999_), .A1(new_new_n370_), .B0(new_new_n1000_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n782_), .B(new_new_n149_), .Y(new_new_n1002_));
  INV        g0980(.A(new_new_n1002_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n1003_), .B(new_new_n722_), .C(new_new_n73_), .Y(new_new_n1004_));
  NO2        g0982(.A(new_new_n860_), .B(new_new_n426_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n889_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n1006_));
  NA2        g0984(.A(new_new_n890_), .B(i_9_), .Y(new_new_n1007_));
  AOI210     g0985(.A0(new_new_n1006_), .A1(new_new_n535_), .B0(new_new_n1007_), .Y(new_new_n1008_));
  OAI210     g0986(.A0(new_new_n255_), .A1(i_9_), .B0(new_new_n240_), .Y(new_new_n1009_));
  AOI210     g0987(.A0(new_new_n1009_), .A1(new_new_n925_), .B0(new_new_n157_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n1010_), .B(new_new_n1008_), .C(new_new_n1005_), .Y(new_new_n1011_));
  NA3        g0989(.A(new_new_n1011_), .B(new_new_n1004_), .C(new_new_n1001_), .Y(new_new_n1012_));
  NA2        g0990(.A(new_new_n972_), .B(new_new_n395_), .Y(new_new_n1013_));
  AOI210     g0991(.A0(new_new_n318_), .A1(new_new_n166_), .B0(new_new_n1013_), .Y(new_new_n1014_));
  NA3        g0992(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n1015_));
  NA2        g0993(.A(new_new_n944_), .B(new_new_n523_), .Y(new_new_n1016_));
  AOI210     g0994(.A0(new_new_n1015_), .A1(new_new_n166_), .B0(new_new_n1016_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n1017_), .B(new_new_n1014_), .Y(new_new_n1018_));
  NO3        g0996(.A(new_new_n935_), .B(new_new_n908_), .C(new_new_n196_), .Y(new_new_n1019_));
  AOI220     g0997(.A0(new_new_n1019_), .A1(i_11_), .B0(new_new_n613_), .B1(new_new_n75_), .Y(new_new_n1020_));
  NO3        g0998(.A(new_new_n218_), .B(new_new_n406_), .C(i_0_), .Y(new_new_n1021_));
  OAI210     g0999(.A0(new_new_n1021_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n1022_));
  INV        g1000(.A(new_new_n227_), .Y(new_new_n1023_));
  OAI220     g1001(.A0(new_new_n571_), .A1(new_new_n142_), .B0(new_new_n695_), .B1(new_new_n665_), .Y(new_new_n1024_));
  NA3        g1002(.A(new_new_n1024_), .B(i_7_), .C(new_new_n1023_), .Y(new_new_n1025_));
  NA4        g1003(.A(new_new_n1025_), .B(new_new_n1022_), .C(new_new_n1020_), .D(new_new_n1018_), .Y(new_new_n1026_));
  NO2        g1004(.A(new_new_n253_), .B(new_new_n95_), .Y(new_new_n1027_));
  AOI210     g1005(.A0(new_new_n1027_), .A1(new_new_n995_), .B0(new_new_n112_), .Y(new_new_n1028_));
  AOI220     g1006(.A0(new_new_n962_), .A1(new_new_n523_), .B0(new_new_n889_), .B1(new_new_n167_), .Y(new_new_n1029_));
  NA2        g1007(.A(new_new_n373_), .B(new_new_n181_), .Y(new_new_n1030_));
  OA220      g1008(.A0(new_new_n1030_), .A1(new_new_n1029_), .B0(new_new_n1028_), .B1(i_5_), .Y(new_new_n1031_));
  AOI210     g1009(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n180_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n1032_), .B(new_new_n975_), .Y(new_new_n1033_));
  NA3        g1011(.A(new_new_n662_), .B(new_new_n191_), .C(new_new_n84_), .Y(new_new_n1034_));
  NA2        g1012(.A(new_new_n1034_), .B(new_new_n587_), .Y(new_new_n1035_));
  NO3        g1013(.A(new_new_n899_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n528_), .B(new_new_n521_), .C(new_new_n504_), .Y(new_new_n1037_));
  NO3        g1015(.A(new_new_n1037_), .B(new_new_n1036_), .C(new_new_n1035_), .Y(new_new_n1038_));
  NA3        g1016(.A(new_new_n413_), .B(new_new_n176_), .C(new_new_n175_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n944_), .B(new_new_n307_), .C(new_new_n240_), .Y(new_new_n1040_));
  NA2        g1018(.A(new_new_n1040_), .B(new_new_n1039_), .Y(new_new_n1041_));
  NA3        g1019(.A(new_new_n413_), .B(new_new_n355_), .C(new_new_n231_), .Y(new_new_n1042_));
  OAI210     g1020(.A0(new_new_n903_), .A1(new_new_n699_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  NOi31      g1021(.An(new_new_n412_), .B(new_new_n996_), .C(new_new_n250_), .Y(new_new_n1044_));
  NO3        g1022(.A(new_new_n943_), .B(new_new_n227_), .C(new_new_n196_), .Y(new_new_n1045_));
  NO4        g1023(.A(new_new_n1045_), .B(new_new_n1044_), .C(new_new_n1043_), .D(new_new_n1041_), .Y(new_new_n1046_));
  NA4        g1024(.A(new_new_n1046_), .B(new_new_n1038_), .C(new_new_n1033_), .D(new_new_n1031_), .Y(new_new_n1047_));
  INV        g1025(.A(new_new_n664_), .Y(new_new_n1048_));
  NO3        g1026(.A(new_new_n1048_), .B(new_new_n603_), .C(new_new_n367_), .Y(new_new_n1049_));
  INV        g1027(.A(new_new_n1049_), .Y(new_new_n1050_));
  NA3        g1028(.A(new_new_n324_), .B(i_5_), .C(new_new_n199_), .Y(new_new_n1051_));
  NAi31      g1029(.An(new_new_n252_), .B(new_new_n1051_), .C(new_new_n253_), .Y(new_new_n1052_));
  NO4        g1030(.A(new_new_n250_), .B(new_new_n218_), .C(i_0_), .D(i_12_), .Y(new_new_n1053_));
  NA2        g1031(.A(new_new_n1053_), .B(new_new_n1052_), .Y(new_new_n1054_));
  AN2        g1032(.A(new_new_n935_), .B(new_new_n157_), .Y(new_new_n1055_));
  NO4        g1033(.A(new_new_n1055_), .B(i_12_), .C(new_new_n699_), .D(new_new_n134_), .Y(new_new_n1056_));
  NA2        g1034(.A(new_new_n1056_), .B(new_new_n227_), .Y(new_new_n1057_));
  NA3        g1035(.A(new_new_n101_), .B(new_new_n617_), .C(i_11_), .Y(new_new_n1058_));
  NO2        g1036(.A(new_new_n1058_), .B(new_new_n159_), .Y(new_new_n1059_));
  NA2        g1037(.A(new_new_n962_), .B(new_new_n503_), .Y(new_new_n1060_));
  NA2        g1038(.A(new_new_n64_), .B(new_new_n104_), .Y(new_new_n1061_));
  OAI220     g1039(.A0(new_new_n1061_), .A1(new_new_n1051_), .B0(new_new_n1060_), .B1(new_new_n723_), .Y(new_new_n1062_));
  AOI210     g1040(.A0(new_new_n1062_), .A1(new_new_n948_), .B0(new_new_n1059_), .Y(new_new_n1063_));
  NA4        g1041(.A(new_new_n1063_), .B(new_new_n1057_), .C(new_new_n1054_), .D(new_new_n1050_), .Y(new_new_n1064_));
  NO4        g1042(.A(new_new_n1064_), .B(new_new_n1047_), .C(new_new_n1026_), .D(new_new_n1012_), .Y(new_new_n1065_));
  OAI210     g1043(.A0(new_new_n863_), .A1(new_new_n856_), .B0(new_new_n37_), .Y(new_new_n1066_));
  NA3        g1044(.A(new_new_n956_), .B(new_new_n390_), .C(i_5_), .Y(new_new_n1067_));
  NA3        g1045(.A(new_new_n1067_), .B(new_new_n1066_), .C(new_new_n660_), .Y(new_new_n1068_));
  NA2        g1046(.A(new_new_n1068_), .B(new_new_n214_), .Y(new_new_n1069_));
  BUFFER     g1047(.A(new_new_n391_), .Y(new_new_n1070_));
  NA2        g1048(.A(new_new_n192_), .B(new_new_n194_), .Y(new_new_n1071_));
  AO210      g1049(.A0(new_new_n1070_), .A1(new_new_n33_), .B0(new_new_n1071_), .Y(new_new_n1072_));
  OAI210     g1050(.A0(new_new_n664_), .A1(new_new_n662_), .B0(new_new_n337_), .Y(new_new_n1073_));
  NAi31      g1051(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1074_));
  AOI210     g1052(.A0(new_new_n120_), .A1(new_new_n70_), .B0(new_new_n1074_), .Y(new_new_n1075_));
  NO2        g1053(.A(new_new_n1075_), .B(new_new_n696_), .Y(new_new_n1076_));
  NA3        g1054(.A(new_new_n1076_), .B(new_new_n1073_), .C(new_new_n1072_), .Y(new_new_n1077_));
  NO2        g1055(.A(new_new_n493_), .B(new_new_n281_), .Y(new_new_n1078_));
  NO4        g1056(.A(new_new_n243_), .B(new_new_n148_), .C(new_new_n726_), .D(new_new_n37_), .Y(new_new_n1079_));
  NO3        g1057(.A(new_new_n1079_), .B(new_new_n1078_), .C(new_new_n927_), .Y(new_new_n1080_));
  OAI210     g1058(.A0(new_new_n1058_), .A1(new_new_n151_), .B0(new_new_n1080_), .Y(new_new_n1081_));
  AOI210     g1059(.A0(new_new_n1077_), .A1(new_new_n49_), .B0(new_new_n1081_), .Y(new_new_n1082_));
  AOI210     g1060(.A0(new_new_n1082_), .A1(new_new_n1069_), .B0(new_new_n73_), .Y(new_new_n1083_));
  NO2        g1061(.A(new_new_n610_), .B(new_new_n402_), .Y(new_new_n1084_));
  NO2        g1062(.A(new_new_n1084_), .B(new_new_n802_), .Y(new_new_n1085_));
  OAI210     g1063(.A0(new_new_n80_), .A1(new_new_n55_), .B0(new_new_n111_), .Y(new_new_n1086_));
  NA2        g1064(.A(new_new_n1086_), .B(new_new_n76_), .Y(new_new_n1087_));
  AOI210     g1065(.A0(new_new_n1032_), .A1(new_new_n944_), .B0(new_new_n963_), .Y(new_new_n1088_));
  AOI210     g1066(.A0(new_new_n1088_), .A1(new_new_n1087_), .B0(new_new_n726_), .Y(new_new_n1089_));
  NA2        g1067(.A(new_new_n275_), .B(new_new_n57_), .Y(new_new_n1090_));
  AOI220     g1068(.A0(new_new_n1090_), .A1(new_new_n76_), .B0(new_new_n368_), .B1(new_new_n267_), .Y(new_new_n1091_));
  NO2        g1069(.A(new_new_n1091_), .B(new_new_n247_), .Y(new_new_n1092_));
  NA3        g1070(.A(new_new_n99_), .B(new_new_n326_), .C(new_new_n31_), .Y(new_new_n1093_));
  INV        g1071(.A(new_new_n1093_), .Y(new_new_n1094_));
  NO3        g1072(.A(new_new_n1094_), .B(new_new_n1092_), .C(new_new_n1089_), .Y(new_new_n1095_));
  OAI210     g1073(.A0(new_new_n283_), .A1(new_new_n162_), .B0(new_new_n89_), .Y(new_new_n1096_));
  NA3        g1074(.A(new_new_n806_), .B(new_new_n307_), .C(new_new_n80_), .Y(new_new_n1097_));
  AOI210     g1075(.A0(new_new_n1097_), .A1(new_new_n1096_), .B0(i_11_), .Y(new_new_n1098_));
  NA2        g1076(.A(new_new_n655_), .B(new_new_n224_), .Y(new_new_n1099_));
  OAI210     g1077(.A0(new_new_n1099_), .A1(new_new_n956_), .B0(new_new_n214_), .Y(new_new_n1100_));
  NA2        g1078(.A(new_new_n168_), .B(i_5_), .Y(new_new_n1101_));
  NO2        g1079(.A(new_new_n1100_), .B(new_new_n1101_), .Y(new_new_n1102_));
  NO3        g1080(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1103_));
  OAI210     g1081(.A0(new_new_n967_), .A1(new_new_n326_), .B0(new_new_n1103_), .Y(new_new_n1104_));
  NO2        g1082(.A(new_new_n1104_), .B(new_new_n772_), .Y(new_new_n1105_));
  NO2        g1083(.A(new_new_n859_), .B(new_new_n386_), .Y(new_new_n1106_));
  NO2        g1084(.A(new_new_n1106_), .B(new_new_n41_), .Y(new_new_n1107_));
  NO4        g1085(.A(new_new_n1107_), .B(new_new_n1105_), .C(new_new_n1102_), .D(new_new_n1098_), .Y(new_new_n1108_));
  OAI210     g1086(.A0(new_new_n1095_), .A1(i_4_), .B0(new_new_n1108_), .Y(new_new_n1109_));
  NO3        g1087(.A(new_new_n1109_), .B(new_new_n1085_), .C(new_new_n1083_), .Y(new_new_n1110_));
  NA4        g1088(.A(new_new_n1110_), .B(new_new_n1065_), .C(new_new_n994_), .D(new_new_n915_), .Y(zz04));
  INV        g1089(.A(i_2_), .Y(new_new_n1114_));
  INV        g1090(.A(new_new_n761_), .Y(new_new_n1115_));
  INV        g1091(.A(new_new_n518_), .Y(new_new_n1116_));
  INV        g1092(.A(i_7_), .Y(new_new_n1117_));
endmodule


